

module b17_C_gen_AntiSAT_k_256_4 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, 
        keyinput_f65, keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, 
        keyinput_f70, keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, 
        keyinput_f75, keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, 
        keyinput_f80, keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, 
        keyinput_f85, keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, 
        keyinput_f90, keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, 
        keyinput_f95, keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, 
        keyinput_f100, keyinput_f101, keyinput_f102, keyinput_f103, 
        keyinput_f104, keyinput_f105, keyinput_f106, keyinput_f107, 
        keyinput_f108, keyinput_f109, keyinput_f110, keyinput_f111, 
        keyinput_f112, keyinput_f113, keyinput_f114, keyinput_f115, 
        keyinput_f116, keyinput_f117, keyinput_f118, keyinput_f119, 
        keyinput_f120, keyinput_f121, keyinput_f122, keyinput_f123, 
        keyinput_f124, keyinput_f125, keyinput_f126, keyinput_f127, 
        keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, 
        keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, 
        keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, 
        keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, 
        keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, 
        keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, 
        keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, 
        keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, 
        keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, 
        keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, 
        keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, 
        keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, 
        keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, keyinput_g64, 
        keyinput_g65, keyinput_g66, keyinput_g67, keyinput_g68, keyinput_g69, 
        keyinput_g70, keyinput_g71, keyinput_g72, keyinput_g73, keyinput_g74, 
        keyinput_g75, keyinput_g76, keyinput_g77, keyinput_g78, keyinput_g79, 
        keyinput_g80, keyinput_g81, keyinput_g82, keyinput_g83, keyinput_g84, 
        keyinput_g85, keyinput_g86, keyinput_g87, keyinput_g88, keyinput_g89, 
        keyinput_g90, keyinput_g91, keyinput_g92, keyinput_g93, keyinput_g94, 
        keyinput_g95, keyinput_g96, keyinput_g97, keyinput_g98, keyinput_g99, 
        keyinput_g100, keyinput_g101, keyinput_g102, keyinput_g103, 
        keyinput_g104, keyinput_g105, keyinput_g106, keyinput_g107, 
        keyinput_g108, keyinput_g109, keyinput_g110, keyinput_g111, 
        keyinput_g112, keyinput_g113, keyinput_g114, keyinput_g115, 
        keyinput_g116, keyinput_g117, keyinput_g118, keyinput_g119, 
        keyinput_g120, keyinput_g121, keyinput_g122, keyinput_g123, 
        keyinput_g124, keyinput_g125, keyinput_g126, keyinput_g127, U355, U356, 
        U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, 
        U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, 
        U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, 
        U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, 
        U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, 
        U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, 
        U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, 
        U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, 
        P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, 
        P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, 
        P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, 
        P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, 
        P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, 
        P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, 
        P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, 
        P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, 
        P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, 
        P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, 
        P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, 
        P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, 
        P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, 
        P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, 
        P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, 
        P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, 
        P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, 
        P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, 
        P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, 
        P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, 
        P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, 
        P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, 
        P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, 
        P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, 
        P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, 
        P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, 
        P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, 
        P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, 
        P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, 
        P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, 
        P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, 
        P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, 
        P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, 
        P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, 
        P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, 
        P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, 
        P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, 
        P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, 
        P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, 
        P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, 
        P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, 
        P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, 
        P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, 
        P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, 
        P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, 
        P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, 
        P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, 
        P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, 
        P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, 
        P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, 
        P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, 
        P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, 
        P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, 
        P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, 
        P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, 
        P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, 
        P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, 
        P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, 
        P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, 
        P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, 
        P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, 
        P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, 
        P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, 
        P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, 
        P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, 
        P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, 
        P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, 
        P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, 
        P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, 
        P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, 
        P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, 
        P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, 
        P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, 
        P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, 
        P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, 
        P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, 
        P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, 
        P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, 
        P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, 
        P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, 
        P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, 
        P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, 
        P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, 
        P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, 
        P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, 
        P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, 
        P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, 
        P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, 
        P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, 
        P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, 
        P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, 
        P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, 
        P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, 
        P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, 
        P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, 
        P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, 
        P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, 
        P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, 
        P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, 
        P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, 
        P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, 
        P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, 
        P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, 
        P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, 
        P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, 
        P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, 
        P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, 
        P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, 
        P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, 
        P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, 
        P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, 
        P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, 
        P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, 
        P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, 
        P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, 
        P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, 
        P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, 
        P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, 
        P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, 
        P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, 
        P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, 
        P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, 
        P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, 
        P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, 
        P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, 
        P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, 
        P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, 
        P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, 
        P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, 
        P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, 
        P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, 
        P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, 
        P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, 
        P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, 
        P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, 
        P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, 
        P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, 
        P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, 
        P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, 
        P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, 
        P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, 
        P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, 
        P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, 
        P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, 
        P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, 
        P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, 
        P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, 
        P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, 
        P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, 
        P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, 
        P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, 
        P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, 
        P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, 
        P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, 
        P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, 
        P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, 
        P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, 
        P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, 
        P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, 
        P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, 
        P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, 
        P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, 
        P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, 
        P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, 
        P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, 
        P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, 
        P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, 
        P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, 
        P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, 
        P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, 
        P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, 
        P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, 
        P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, 
        P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, 
        P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, 
        P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, 
        P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, 
        P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, 
        P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, 
        P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9810, n9811, n9812, n9813, n9814, n9815, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9832, n9833, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9940, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322;

  NAND2_X2 U11254 ( .A1(n17870), .A2(n17776), .ZN(n17815) );
  INV_X1 U11255 ( .A(n18026), .ZN(n18036) );
  NOR2_X1 U11256 ( .A1(n18021), .A2(n17993), .ZN(n17919) );
  OR2_X1 U11257 ( .A1(n10470), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17681) );
  NOR2_X1 U11258 ( .A1(n14877), .A2(n10237), .ZN(n10240) );
  NAND2_X2 U11259 ( .A1(n18804), .A2(n18802), .ZN(n18202) );
  OAI21_X2 U11260 ( .B1(n13064), .B2(n10055), .A(n13066), .ZN(n16153) );
  NAND3_X1 U11261 ( .A1(n16173), .A2(n18375), .A3(n18366), .ZN(n17382) );
  CLKBUF_X1 U11263 ( .A(n11690), .Z(n14593) );
  NAND2_X1 U11264 ( .A1(n12396), .A2(n12397), .ZN(n13034) );
  INV_X2 U11265 ( .A(n20051), .ZN(n20050) );
  CLKBUF_X2 U11266 ( .A(n10548), .Z(n17224) );
  AND2_X1 U11267 ( .A1(n10868), .A2(n13827), .ZN(n11900) );
  AND2_X1 U11268 ( .A1(n10674), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11571) );
  AND2_X1 U11269 ( .A1(n10868), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11072) );
  AND2_X1 U11270 ( .A1(n10157), .A2(n10156), .ZN(n11840) );
  BUF_X1 U11271 ( .A(n11064), .Z(n11901) );
  CLKBUF_X2 U11272 ( .A(n9822), .Z(n9922) );
  AND2_X1 U11273 ( .A1(n10674), .A2(n13827), .ZN(n11902) );
  AND3_X1 U11274 ( .A1(n20243), .A2(n12301), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n13059) );
  INV_X1 U11275 ( .A(n11300), .ZN(n10773) );
  CLKBUF_X2 U11276 ( .A(n10342), .Z(n9814) );
  BUF_X2 U11277 ( .A(n10342), .Z(n9813) );
  CLKBUF_X2 U11278 ( .A(n12610), .Z(n12967) );
  CLKBUF_X1 U11279 ( .A(n13588), .Z(n9938) );
  CLKBUF_X3 U11280 ( .A(n10356), .Z(n17331) );
  BUF_X2 U11281 ( .A(n17122), .Z(n17167) );
  INV_X1 U11282 ( .A(n17121), .ZN(n17348) );
  CLKBUF_X3 U11283 ( .A(n10380), .Z(n9821) );
  AND2_X1 U11284 ( .A1(n12239), .A2(n12243), .ZN(n13086) );
  AND3_X2 U11285 ( .A1(n12186), .A2(n12185), .A3(n12184), .ZN(n13587) );
  CLKBUF_X2 U11287 ( .A(n9942), .Z(n9944) );
  AND2_X1 U11288 ( .A1(n12095), .A2(n12087), .ZN(n12223) );
  NAND2_X2 U11289 ( .A1(n12094), .A2(n13537), .ZN(n12961) );
  BUF_X2 U11290 ( .A(n10653), .Z(n9818) );
  NAND2_X1 U11291 ( .A1(n9950), .A2(n13885), .ZN(n12986) );
  NOR2_X2 U11292 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13792) );
  AND2_X1 U11293 ( .A1(n10641), .A2(n13802), .ZN(n10653) );
  AND2_X2 U11294 ( .A1(n9951), .A2(n12087), .ZN(n12702) );
  AND2_X2 U11295 ( .A1(n12088), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12087) );
  CLKBUF_X2 U11296 ( .A(n12223), .Z(n12859) );
  INV_X1 U11298 ( .A(n13010), .ZN(n14429) );
  INV_X1 U11300 ( .A(n11400), .ZN(n14585) );
  INV_X2 U11301 ( .A(n10556), .ZN(n17341) );
  CLKBUF_X3 U11302 ( .A(n10394), .Z(n9833) );
  INV_X1 U11303 ( .A(n9938), .ZN(n14631) );
  INV_X1 U11304 ( .A(n15140), .ZN(n16276) );
  INV_X1 U11305 ( .A(n12634), .ZN(n13879) );
  INV_X1 U11306 ( .A(n12241), .ZN(n10059) );
  INV_X1 U11307 ( .A(n17815), .ZN(n18018) );
  INV_X1 U11308 ( .A(n18812), .ZN(n18802) );
  OR2_X2 U11309 ( .A1(n12220), .A2(n12219), .ZN(n20243) );
  NAND2_X1 U11310 ( .A1(n15151), .A2(n15150), .ZN(n15152) );
  NAND2_X1 U11311 ( .A1(n15089), .A2(n15088), .ZN(n15079) );
  INV_X1 U11312 ( .A(n19206), .ZN(n10206) );
  INV_X1 U11313 ( .A(n19181), .ZN(n19172) );
  INV_X1 U11314 ( .A(n16960), .ZN(n17047) );
  INV_X1 U11315 ( .A(n17756), .ZN(n17836) );
  INV_X1 U11317 ( .A(n17926), .ZN(n17946) );
  NAND2_X1 U11318 ( .A1(n10641), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9810) );
  BUF_X1 U11319 ( .A(n9942), .Z(n9943) );
  CLKBUF_X3 U11320 ( .A(n13900), .Z(n9951) );
  NAND2_X1 U11321 ( .A1(n15058), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15010) );
  OR2_X2 U11322 ( .A1(n15470), .A2(n10264), .ZN(n10261) );
  OAI21_X4 U11323 ( .B1(n16176), .B2(n17591), .A(n16175), .ZN(n17401) );
  BUF_X4 U11324 ( .A(n10803), .Z(n9959) );
  NAND2_X2 U11325 ( .A1(n15152), .A2(n9970), .ZN(n9889) );
  NAND2_X1 U11327 ( .A1(n12247), .A2(n20243), .ZN(n14462) );
  INV_X2 U11328 ( .A(n10406), .ZN(n10417) );
  AND2_X1 U11329 ( .A1(n12390), .A2(n12389), .ZN(n12414) );
  OAI21_X2 U11330 ( .B1(n10975), .B2(n10974), .A(n10985), .ZN(n14013) );
  BUF_X2 U11331 ( .A(n10436), .Z(n9812) );
  NOR2_X4 U11332 ( .A1(n17960), .A2(n17974), .ZN(n16937) );
  AND2_X1 U11333 ( .A1(n9950), .A2(n12087), .ZN(n9957) );
  NOR2_X4 U11334 ( .A1(n18202), .A2(n18817), .ZN(n18297) );
  NAND2_X1 U11335 ( .A1(n10814), .A2(n10815), .ZN(n10828) );
  INV_X2 U11336 ( .A(n14134), .ZN(n20035) );
  BUF_X4 U11338 ( .A(n10358), .Z(n17347) );
  OR2_X4 U11339 ( .A1(n11717), .A2(n19032), .ZN(n11400) );
  XNOR2_X1 U11341 ( .A(n14582), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14605) );
  NAND2_X1 U11342 ( .A1(n9848), .A2(n9847), .ZN(n14637) );
  CLKBUF_X1 U11343 ( .A(n15612), .Z(n15613) );
  CLKBUF_X1 U11344 ( .A(n15670), .Z(n15671) );
  CLKBUF_X1 U11345 ( .A(n15690), .Z(n15691) );
  NAND2_X1 U11346 ( .A1(n9879), .A2(n10136), .ZN(n15635) );
  NAND2_X1 U11347 ( .A1(n10119), .A2(n9971), .ZN(n9882) );
  AND2_X1 U11348 ( .A1(n17681), .A2(n10165), .ZN(n17666) );
  NOR2_X1 U11349 ( .A1(n17681), .A2(n16598), .ZN(n9904) );
  NAND2_X1 U11350 ( .A1(n14292), .A2(n14293), .ZN(n10119) );
  NAND2_X1 U11351 ( .A1(n10470), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17680) );
  NOR2_X1 U11352 ( .A1(n17692), .A2(n9864), .ZN(n10470) );
  NOR2_X1 U11353 ( .A1(n14448), .A2(n10049), .ZN(n10048) );
  NOR2_X1 U11354 ( .A1(n17693), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17692) );
  NOR2_X1 U11356 ( .A1(n10132), .A2(n10131), .ZN(n10130) );
  NAND2_X1 U11357 ( .A1(n9867), .A2(n9825), .ZN(n9866) );
  INV_X1 U11358 ( .A(n17723), .ZN(n9825) );
  INV_X1 U11359 ( .A(n17865), .ZN(n17791) );
  NAND2_X1 U11360 ( .A1(n10115), .A2(n9924), .ZN(n11159) );
  NAND2_X1 U11361 ( .A1(n10973), .A2(n10972), .ZN(n11165) );
  INV_X2 U11362 ( .A(n18032), .ZN(n18021) );
  AND4_X1 U11363 ( .A1(n10912), .A2(n10914), .A3(n10913), .A4(n10911), .ZN(
        n10927) );
  NOR2_X1 U11364 ( .A1(n17660), .A2(n17484), .ZN(n17478) );
  NAND2_X1 U11365 ( .A1(n10330), .A2(n11777), .ZN(n10832) );
  AOI21_X1 U11366 ( .B1(n19571), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n19356), .ZN(n10824) );
  NOR2_X1 U11367 ( .A1(n10854), .A2(n10836), .ZN(n10941) );
  NAND2_X1 U11368 ( .A1(n13357), .A2(n11786), .ZN(n13468) );
  AND2_X1 U11369 ( .A1(n13322), .A2(n11555), .ZN(n14072) );
  NAND2_X1 U11370 ( .A1(n17961), .A2(n10451), .ZN(n10452) );
  CLKBUF_X2 U11371 ( .A(n10819), .Z(n10829) );
  AND2_X1 U11372 ( .A1(n14090), .A2(n14002), .ZN(n14170) );
  NAND2_X1 U11373 ( .A1(n11731), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10803) );
  BUF_X2 U11374 ( .A(n10773), .Z(n11383) );
  NAND2_X1 U11375 ( .A1(n10730), .A2(n13781), .ZN(n11731) );
  INV_X1 U11376 ( .A(n11680), .ZN(n11668) );
  NAND2_X1 U11377 ( .A1(n14631), .A2(n14517), .ZN(n13325) );
  NAND2_X1 U11378 ( .A1(n12067), .A2(n11520), .ZN(n11680) );
  NAND2_X1 U11379 ( .A1(n14462), .A2(n14480), .ZN(n13597) );
  INV_X2 U11380 ( .A(n18397), .ZN(n10597) );
  NAND2_X1 U11381 ( .A1(n13578), .A2(n20268), .ZN(n12248) );
  INV_X2 U11382 ( .A(n13364), .ZN(n11511) );
  NOR2_X2 U11383 ( .A1(n14134), .A2(n11507), .ZN(n11409) );
  OR2_X2 U11385 ( .A1(n12238), .A2(n12237), .ZN(n12268) );
  NAND2_X1 U11386 ( .A1(n12203), .A2(n9982), .ZN(n20263) );
  INV_X2 U11387 ( .A(n10723), .ZN(n9819) );
  CLKBUF_X2 U11388 ( .A(n12808), .Z(n9945) );
  NOR3_X1 U11389 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n18825), .ZN(n10342) );
  INV_X4 U11391 ( .A(n12988), .ZN(n12753) );
  INV_X2 U11392 ( .A(n12961), .ZN(n12880) );
  INV_X1 U11393 ( .A(n12232), .ZN(n12808) );
  BUF_X1 U11394 ( .A(n10548), .Z(n17346) );
  BUF_X2 U11395 ( .A(n12855), .Z(n12993) );
  INV_X1 U11396 ( .A(n9961), .ZN(n9820) );
  CLKBUF_X2 U11397 ( .A(n10862), .Z(n9954) );
  CLKBUF_X2 U11398 ( .A(n10716), .Z(n12047) );
  CLKBUF_X2 U11399 ( .A(n10862), .Z(n9955) );
  CLKBUF_X2 U11400 ( .A(n10862), .Z(n9956) );
  OR2_X1 U11401 ( .A1(n18969), .A2(n10346), .ZN(n17121) );
  CLKBUF_X3 U11402 ( .A(n10425), .Z(n9835) );
  INV_X2 U11403 ( .A(n12848), .ZN(n9822) );
  NOR3_X1 U11404 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18969), .A3(
        n18826), .ZN(n10425) );
  BUF_X4 U11405 ( .A(n10862), .Z(n9823) );
  OR2_X1 U11408 ( .A1(n11762), .A2(n15966), .ZN(n11755) );
  AOI21_X1 U11409 ( .B1(n14637), .B2(n20188), .A(n14616), .ZN(n14617) );
  OAI211_X1 U11410 ( .C1(n11472), .C2(n15759), .A(n11471), .B(n11470), .ZN(
        n15575) );
  AND3_X1 U11411 ( .A1(n10254), .A2(n10253), .A3(n11470), .ZN(n15587) );
  OR2_X1 U11412 ( .A1(n11467), .A2(n11290), .ZN(n10254) );
  INV_X1 U11413 ( .A(n11289), .ZN(n11467) );
  NOR2_X1 U11414 ( .A1(n11289), .A2(n11284), .ZN(n11469) );
  NAND2_X1 U11415 ( .A1(n9933), .A2(n9905), .ZN(n11289) );
  NOR3_X1 U11416 ( .A1(n10291), .A2(n9851), .A3(n9850), .ZN(n9849) );
  CLKBUF_X1 U11417 ( .A(n14670), .Z(n14671) );
  INV_X1 U11418 ( .A(n15670), .ZN(n9824) );
  OAI21_X1 U11419 ( .B1(n15630), .B2(n9988), .A(n10130), .ZN(n9906) );
  NAND2_X1 U11420 ( .A1(n14726), .A2(n10279), .ZN(n14685) );
  OAI21_X1 U11421 ( .B1(n15729), .B2(n15730), .A(n9842), .ZN(n15731) );
  AOI21_X1 U11422 ( .B1(n14602), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14601), .ZN(n14603) );
  OR2_X1 U11423 ( .A1(n14874), .A2(n14787), .ZN(n14865) );
  AOI21_X1 U11424 ( .B1(n16588), .B2(n18250), .A(n9870), .ZN(n16100) );
  NAND2_X1 U11425 ( .A1(n15635), .A2(n15636), .ZN(n11271) );
  OAI21_X1 U11426 ( .B1(n11440), .B2(n14136), .A(n11439), .ZN(n11441) );
  XNOR2_X1 U11427 ( .A(n11958), .B(n11955), .ZN(n15457) );
  XNOR2_X1 U11428 ( .A(n9872), .B(n9871), .ZN(n16588) );
  NAND2_X1 U11429 ( .A1(n9882), .A2(n9880), .ZN(n9879) );
  XNOR2_X1 U11430 ( .A(n14591), .B(n14590), .ZN(n15366) );
  OR2_X1 U11431 ( .A1(n9904), .A2(n10251), .ZN(n9872) );
  NAND2_X1 U11432 ( .A1(n9904), .A2(n9871), .ZN(n11449) );
  OR2_X1 U11433 ( .A1(n15429), .A2(n15428), .ZN(n16377) );
  NAND2_X1 U11434 ( .A1(n9882), .A2(n11206), .ZN(n15719) );
  NOR2_X1 U11435 ( .A1(n15427), .A2(n11404), .ZN(n16398) );
  AND2_X1 U11436 ( .A1(n15446), .A2(n15445), .ZN(n16412) );
  NAND2_X1 U11437 ( .A1(n15136), .A2(n10048), .ZN(n10047) );
  XNOR2_X1 U11438 ( .A(n15429), .B(n14584), .ZN(n15379) );
  AOI21_X1 U11439 ( .B1(n19234), .B2(n16558), .A(n14599), .ZN(n14600) );
  AND2_X1 U11440 ( .A1(n15479), .A2(n11910), .ZN(n10323) );
  XNOR2_X1 U11441 ( .A(n14596), .B(n14595), .ZN(n19234) );
  NAND2_X1 U11442 ( .A1(n10060), .A2(n16285), .ZN(n14402) );
  NAND2_X1 U11443 ( .A1(n14232), .A2(n14309), .ZN(n14308) );
  OAI211_X1 U11444 ( .C1(n17826), .C2(n17723), .A(n9865), .B(n10329), .ZN(
        n17693) );
  OR2_X1 U11445 ( .A1(n17714), .A2(n10468), .ZN(n9864) );
  NOR2_X1 U11446 ( .A1(n15511), .A2(n15510), .ZN(n15513) );
  AND2_X1 U11447 ( .A1(n14159), .A2(n12526), .ZN(n14209) );
  NOR2_X1 U11448 ( .A1(n14446), .A2(n16253), .ZN(n14447) );
  AOI21_X1 U11449 ( .B1(n15095), .B2(n14445), .A(n14442), .ZN(n16252) );
  XNOR2_X1 U11450 ( .A(n11183), .B(n14295), .ZN(n14293) );
  NAND2_X1 U11451 ( .A1(n16498), .A2(n16497), .ZN(n11041) );
  OR2_X1 U11452 ( .A1(n11088), .A2(n16545), .ZN(n11089) );
  INV_X1 U11453 ( .A(n14445), .ZN(n16253) );
  NAND2_X1 U11454 ( .A1(n9843), .A2(n10988), .ZN(n16498) );
  CLKBUF_X1 U11455 ( .A(n15388), .Z(n15526) );
  OR2_X1 U11456 ( .A1(n14373), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16286) );
  OAI21_X1 U11457 ( .B1(n14011), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n14009), .ZN(n9901) );
  NOR2_X1 U11458 ( .A1(n15120), .A2(n14439), .ZN(n15106) );
  AND2_X1 U11459 ( .A1(n16263), .A2(n16267), .ZN(n14445) );
  AND2_X1 U11460 ( .A1(n15118), .A2(n15114), .ZN(n15103) );
  AND2_X1 U11461 ( .A1(n15104), .A2(n14441), .ZN(n16263) );
  NAND3_X1 U11462 ( .A1(n10135), .A2(n10134), .A3(n14150), .ZN(n14011) );
  AND2_X1 U11463 ( .A1(n15594), .A2(n10186), .ZN(n9905) );
  OR2_X1 U11464 ( .A1(n15216), .A2(n14531), .ZN(n15206) );
  NAND2_X1 U11465 ( .A1(n17733), .A2(n9891), .ZN(n17724) );
  NAND2_X1 U11466 ( .A1(n11159), .A2(n11036), .ZN(n10159) );
  AOI21_X1 U11467 ( .B1(n11036), .B2(n11165), .A(n14578), .ZN(n10158) );
  XNOR2_X1 U11468 ( .A(n10985), .B(n11547), .ZN(n14187) );
  XNOR2_X1 U11469 ( .A(n11159), .B(n11165), .ZN(n11174) );
  INV_X1 U11470 ( .A(n17870), .ZN(n17890) );
  AND2_X1 U11471 ( .A1(n10137), .A2(n11263), .ZN(n10136) );
  NOR2_X1 U11472 ( .A1(n10139), .A2(n9881), .ZN(n9880) );
  NAND2_X1 U11473 ( .A1(n11033), .A2(n11032), .ZN(n11036) );
  NAND2_X1 U11474 ( .A1(n9841), .A2(n9840), .ZN(n10985) );
  AND2_X1 U11475 ( .A1(n14060), .A2(n10183), .ZN(n14389) );
  AND2_X1 U11476 ( .A1(n11280), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15615) );
  NAND2_X1 U11477 ( .A1(n17821), .A2(n17932), .ZN(n17733) );
  NOR3_X2 U11478 ( .A1(n17100), .A2(n17099), .A3(n17154), .ZN(n17140) );
  NOR2_X1 U11479 ( .A1(n9852), .A2(n14007), .ZN(n13985) );
  NAND2_X1 U11480 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17919), .ZN(n17870) );
  AND2_X1 U11481 ( .A1(n10897), .A2(n10117), .ZN(n9840) );
  OR2_X1 U11482 ( .A1(n9963), .A2(n14677), .ZN(n14679) );
  NAND2_X1 U11483 ( .A1(n10067), .A2(n10066), .ZN(n14356) );
  AND2_X1 U11484 ( .A1(n10897), .A2(n10978), .ZN(n10974) );
  NAND2_X1 U11485 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17163), .ZN(n17154) );
  NOR2_X1 U11486 ( .A1(n15395), .A2(n11169), .ZN(n11280) );
  NAND2_X1 U11487 ( .A1(n13855), .A2(n13854), .ZN(n9852) );
  XNOR2_X1 U11488 ( .A(n13529), .B(n13531), .ZN(n19988) );
  AND2_X1 U11489 ( .A1(n12448), .A2(n12447), .ZN(n14007) );
  AND3_X1 U11490 ( .A1(n10463), .A2(n9875), .A3(n10247), .ZN(n17822) );
  OAI21_X1 U11491 ( .B1(n20238), .B2(n10283), .A(n12425), .ZN(n13854) );
  AOI21_X1 U11492 ( .B1(n10466), .B2(n18078), .A(n10465), .ZN(n9892) );
  AND4_X1 U11493 ( .A1(n10901), .A2(n10899), .A3(n10898), .A4(n10900), .ZN(
        n10928) );
  NAND2_X1 U11494 ( .A1(n12449), .A2(n12416), .ZN(n20238) );
  NOR2_X1 U11495 ( .A1(n13934), .A2(n11335), .ZN(n13190) );
  OAI22_X1 U11496 ( .A1(n11023), .A2(n19428), .B1(n10990), .B2(n10989), .ZN(
        n10991) );
  NAND2_X1 U11497 ( .A1(n12477), .A2(n12476), .ZN(n10068) );
  NAND2_X1 U11498 ( .A1(n10462), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9875) );
  OAI21_X2 U11499 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19008), .A(n16719), 
        .ZN(n18032) );
  AND2_X1 U11500 ( .A1(n10831), .A2(n10830), .ZN(n10861) );
  NAND2_X1 U11501 ( .A1(n17909), .A2(n13119), .ZN(n10462) );
  OAI21_X1 U11502 ( .B1(n17877), .B2(n9873), .A(n17932), .ZN(n10463) );
  NAND2_X1 U11503 ( .A1(n12414), .A2(n13920), .ZN(n12449) );
  NOR2_X1 U11504 ( .A1(n11276), .A2(n10199), .ZN(n11282) );
  OAI211_X1 U11505 ( .C1(n19632), .C2(n10826), .A(n10825), .B(n10824), .ZN(
        n10827) );
  NAND2_X1 U11506 ( .A1(n17931), .A2(n10460), .ZN(n17909) );
  NOR2_X1 U11507 ( .A1(n14262), .A2(n10832), .ZN(n19425) );
  NAND2_X1 U11508 ( .A1(n17892), .A2(n10461), .ZN(n17877) );
  NOR2_X2 U11509 ( .A1(n10832), .A2(n13472), .ZN(n10957) );
  INV_X1 U11510 ( .A(n19350), .ZN(n19347) );
  INV_X1 U11511 ( .A(n10902), .ZN(n10940) );
  INV_X1 U11512 ( .A(n19632), .ZN(n19641) );
  INV_X1 U11513 ( .A(n10903), .ZN(n19797) );
  INV_X1 U11514 ( .A(n14124), .ZN(n10956) );
  OAI21_X1 U11515 ( .B1(n13468), .B2(n13470), .A(n13469), .ZN(n11793) );
  AND2_X1 U11516 ( .A1(n10330), .A2(n10841), .ZN(n19350) );
  INV_X1 U11517 ( .A(n19571), .ZN(n10942) );
  NAND2_X1 U11518 ( .A1(n9845), .A2(n9990), .ZN(n19675) );
  AND2_X1 U11519 ( .A1(n10941), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10904) );
  AND2_X1 U11520 ( .A1(n10330), .A2(n10843), .ZN(n19488) );
  NAND2_X1 U11521 ( .A1(n9845), .A2(n10842), .ZN(n19632) );
  INV_X1 U11522 ( .A(n19517), .ZN(n10995) );
  NAND2_X1 U11523 ( .A1(n10849), .A2(n9990), .ZN(n10903) );
  NAND2_X1 U11524 ( .A1(n9845), .A2(n10848), .ZN(n10902) );
  INV_X1 U11525 ( .A(n19397), .ZN(n10998) );
  NAND2_X1 U11526 ( .A1(n9845), .A2(n10822), .ZN(n19700) );
  INV_X1 U11527 ( .A(n19464), .ZN(n10945) );
  NOR2_X1 U11528 ( .A1(n17904), .A2(n10172), .ZN(n17892) );
  AND2_X1 U11529 ( .A1(n10823), .A2(n13532), .ZN(n19571) );
  OR2_X1 U11530 ( .A1(n10854), .A2(n10853), .ZN(n14124) );
  NAND2_X2 U11531 ( .A1(n14983), .A2(n13769), .ZN(n14987) );
  NAND2_X1 U11532 ( .A1(n11770), .A2(n11769), .ZN(n11797) );
  AND2_X1 U11533 ( .A1(n13532), .A2(n13414), .ZN(n10330) );
  AND2_X1 U11534 ( .A1(n9903), .A2(n17952), .ZN(n9876) );
  AND2_X1 U11535 ( .A1(n10837), .A2(n13532), .ZN(n19397) );
  XNOR2_X1 U11536 ( .A(n10459), .B(n18263), .ZN(n18267) );
  AND2_X1 U11537 ( .A1(n10821), .A2(n13532), .ZN(n19464) );
  NAND2_X1 U11538 ( .A1(n17952), .A2(n10454), .ZN(n10459) );
  AND2_X1 U11539 ( .A1(n13586), .A2(n13585), .ZN(n13612) );
  NOR2_X1 U11540 ( .A1(n10053), .A2(n17826), .ZN(n9903) );
  NAND2_X1 U11541 ( .A1(n12413), .A2(n12412), .ZN(n13920) );
  AND2_X1 U11542 ( .A1(n11249), .A2(n11248), .ZN(n11259) );
  AND2_X1 U11543 ( .A1(n17401), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17550) );
  NAND2_X2 U11544 ( .A1(n19014), .A2(n18297), .ZN(n18225) );
  AND2_X1 U11545 ( .A1(n11231), .A2(n11230), .ZN(n19097) );
  BUF_X1 U11546 ( .A(n11765), .Z(n10813) );
  INV_X1 U11547 ( .A(n14744), .ZN(n9854) );
  NAND2_X1 U11548 ( .A1(n17953), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17952) );
  AND2_X1 U11549 ( .A1(n10840), .A2(n10822), .ZN(n10821) );
  INV_X1 U11550 ( .A(n10838), .ZN(n10840) );
  NAND2_X1 U11551 ( .A1(n13818), .A2(n13414), .ZN(n10853) );
  XNOR2_X1 U11552 ( .A(n10452), .B(n10248), .ZN(n17953) );
  CLKBUF_X1 U11553 ( .A(n13748), .Z(n20528) );
  NOR2_X2 U11554 ( .A1(n19292), .A2(n19792), .ZN(n14132) );
  NOR2_X1 U11555 ( .A1(n14027), .A2(n14026), .ZN(n14192) );
  NOR2_X2 U11556 ( .A1(n19357), .A2(n19792), .ZN(n19358) );
  INV_X1 U11557 ( .A(n19224), .ZN(n13414) );
  AND2_X1 U11558 ( .A1(n9915), .A2(n9916), .ZN(n12359) );
  NOR2_X2 U11559 ( .A1(n19362), .A2(n19792), .ZN(n19363) );
  OR2_X1 U11560 ( .A1(n11235), .A2(n11234), .ZN(n11238) );
  AOI221_X1 U11561 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16170), .C1(n20025), .C2(
        n16170), .A(n19833), .ZN(n20021) );
  AND2_X1 U11562 ( .A1(n10036), .A2(n10038), .ZN(n10035) );
  AND2_X1 U11563 ( .A1(n10794), .A2(n10808), .ZN(n10795) );
  INV_X1 U11564 ( .A(n10799), .ZN(n9886) );
  OAI21_X1 U11565 ( .B1(n17980), .B2(n9859), .A(n9856), .ZN(n17961) );
  AND2_X1 U11566 ( .A1(n16153), .A2(n20936), .ZN(n16142) );
  NAND2_X1 U11567 ( .A1(n20358), .A2(n12361), .ZN(n12364) );
  NAND2_X1 U11568 ( .A1(n11211), .A2(n11212), .ZN(n11235) );
  AOI21_X1 U11569 ( .B1(n10449), .B2(n9858), .A(n9857), .ZN(n9856) );
  INV_X1 U11570 ( .A(n10449), .ZN(n9859) );
  INV_X1 U11571 ( .A(n11299), .ZN(n9887) );
  AND2_X1 U11572 ( .A1(n12307), .A2(n12306), .ZN(n12361) );
  OR2_X1 U11573 ( .A1(n9839), .A2(n11297), .ZN(n11298) );
  NAND2_X1 U11574 ( .A1(n12395), .A2(n12394), .ZN(n20400) );
  NAND2_X1 U11575 ( .A1(n17986), .A2(n10444), .ZN(n10447) );
  NAND2_X1 U11576 ( .A1(n10586), .A2(n10583), .ZN(n10588) );
  INV_X1 U11577 ( .A(n10796), .ZN(n10810) );
  AND2_X1 U11578 ( .A1(n10790), .A2(n10789), .ZN(n10797) );
  AND3_X1 U11579 ( .A1(n11303), .A2(n11302), .A3(n11301), .ZN(n13623) );
  NAND2_X1 U11580 ( .A1(n10062), .A2(n10061), .ZN(n10064) );
  NAND2_X1 U11581 ( .A1(n10299), .A2(n12271), .ZN(n12306) );
  OR2_X1 U11582 ( .A1(n13374), .A2(n13375), .ZN(n13377) );
  AOI21_X1 U11583 ( .B1(n10783), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10784), .ZN(n10796) );
  OAI21_X1 U11584 ( .B1(n18004), .B2(n9863), .A(n9860), .ZN(n17986) );
  NAND2_X1 U11585 ( .A1(n17826), .A2(n18162), .ZN(n10247) );
  NAND2_X1 U11586 ( .A1(n10777), .A2(n10758), .ZN(n10783) );
  AOI21_X1 U11587 ( .B1(n18383), .B2(n10574), .A(n13106), .ZN(n10586) );
  AND2_X1 U11588 ( .A1(n13459), .A2(n12270), .ZN(n12271) );
  AND2_X1 U11589 ( .A1(n9861), .A2(n17988), .ZN(n9860) );
  INV_X1 U11590 ( .A(n17963), .ZN(n9857) );
  NOR2_X2 U11591 ( .A1(n17524), .A2(n16601), .ZN(n17826) );
  AND2_X1 U11592 ( .A1(n10750), .A2(n10749), .ZN(n10777) );
  INV_X1 U11593 ( .A(n10442), .ZN(n9863) );
  NAND3_X2 U11594 ( .A1(n19014), .A2(n18848), .A3(n17593), .ZN(n17642) );
  NOR2_X2 U11595 ( .A1(n16718), .A2(n10580), .ZN(n14415) );
  NAND2_X1 U11596 ( .A1(n10442), .A2(n9862), .ZN(n9861) );
  AND2_X1 U11597 ( .A1(n11519), .A2(n11518), .ZN(n11527) );
  XNOR2_X1 U11598 ( .A(n10441), .B(n18308), .ZN(n18004) );
  NAND2_X1 U11599 ( .A1(n11491), .A2(n10757), .ZN(n11300) );
  AOI21_X1 U11600 ( .B1(n13034), .B2(n12268), .A(n13033), .ZN(n13044) );
  AND3_X1 U11601 ( .A1(n10728), .A2(n10727), .A3(n11703), .ZN(n10763) );
  NAND2_X1 U11602 ( .A1(n9902), .A2(n12262), .ZN(n13448) );
  OR2_X1 U11603 ( .A1(n13415), .A2(n13993), .ZN(n13067) );
  XNOR2_X1 U11604 ( .A(n10249), .B(n10614), .ZN(n10443) );
  INV_X1 U11605 ( .A(n13848), .ZN(n11491) );
  NOR2_X1 U11606 ( .A1(n17696), .A2(n17695), .ZN(n17667) );
  INV_X1 U11607 ( .A(n11680), .ZN(n9826) );
  NAND2_X1 U11608 ( .A1(n10747), .A2(n10746), .ZN(n13838) );
  NAND2_X1 U11609 ( .A1(n10729), .A2(n11409), .ZN(n11707) );
  NAND2_X1 U11610 ( .A1(n13597), .A2(n12248), .ZN(n9902) );
  NAND2_X1 U11611 ( .A1(n10733), .A2(n14134), .ZN(n9896) );
  NAND2_X1 U11612 ( .A1(n10435), .A2(n18023), .ZN(n18015) );
  NAND2_X1 U11613 ( .A1(n10739), .A2(n20035), .ZN(n11483) );
  NAND2_X1 U11614 ( .A1(n12189), .A2(n12254), .ZN(n12206) );
  NAND2_X1 U11615 ( .A1(n9890), .A2(n18024), .ZN(n18023) );
  NAND2_X1 U11616 ( .A1(n13446), .A2(n9853), .ZN(n12251) );
  AND2_X1 U11617 ( .A1(n12240), .A2(n13078), .ZN(n12261) );
  NOR2_X1 U11618 ( .A1(n17730), .A2(n17745), .ZN(n17718) );
  NOR2_X1 U11619 ( .A1(n10585), .A2(n18379), .ZN(n13115) );
  NOR2_X1 U11620 ( .A1(n17367), .A2(n10578), .ZN(n10599) );
  BUF_X4 U11621 ( .A(n11277), .Z(n14575) );
  OR2_X1 U11622 ( .A1(n12334), .A2(n12333), .ZN(n13693) );
  CLKBUF_X3 U11623 ( .A(n14480), .Z(n14517) );
  INV_X1 U11624 ( .A(n11409), .ZN(n9846) );
  NOR2_X1 U11625 ( .A1(n11507), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11520) );
  CLKBUF_X1 U11626 ( .A(n12243), .Z(n13015) );
  AND2_X1 U11627 ( .A1(n16179), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n9890) );
  INV_X1 U11628 ( .A(n10607), .ZN(n17543) );
  NAND2_X2 U11629 ( .A1(n10129), .A2(n10127), .ZN(n13364) );
  NAND2_X2 U11630 ( .A1(n10341), .A2(n10318), .ZN(n12239) );
  NAND4_X1 U11631 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12243) );
  AND2_X2 U11632 ( .A1(n10698), .A2(n10697), .ZN(n10738) );
  NAND2_X2 U11633 ( .A1(n10126), .A2(n10122), .ZN(n19373) );
  INV_X1 U11634 ( .A(n19361), .ZN(n9827) );
  AND2_X1 U11635 ( .A1(n12183), .A2(n12182), .ZN(n12184) );
  OR2_X2 U11636 ( .A1(n16668), .A2(n16615), .ZN(n16670) );
  NAND2_X1 U11637 ( .A1(n10665), .A2(n10664), .ZN(n10723) );
  OR2_X1 U11638 ( .A1(n10884), .A2(n10883), .ZN(n13240) );
  INV_X2 U11639 ( .A(U212), .ZN(n16655) );
  NAND2_X1 U11640 ( .A1(n10704), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10711) );
  NAND2_X1 U11641 ( .A1(n9986), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10126) );
  NAND2_X1 U11642 ( .A1(n10709), .A2(n13827), .ZN(n10710) );
  NAND2_X1 U11643 ( .A1(n10147), .A2(n10146), .ZN(n11513) );
  NAND2_X1 U11644 ( .A1(n9987), .A2(n9966), .ZN(n10698) );
  OAI21_X1 U11645 ( .B1(n10121), .B2(n10128), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10127) );
  AND4_X1 U11646 ( .A1(n12193), .A2(n12192), .A3(n12191), .A4(n12190), .ZN(
        n12203) );
  AND4_X1 U11647 ( .A1(n12127), .A2(n12126), .A3(n12125), .A4(n12124), .ZN(
        n12133) );
  AND4_X1 U11648 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12132) );
  AND4_X1 U11649 ( .A1(n12106), .A2(n12105), .A3(n12104), .A4(n12103), .ZN(
        n10341) );
  AND2_X1 U11650 ( .A1(n12165), .A2(n12164), .ZN(n12166) );
  AND4_X1 U11651 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(
        n12159) );
  INV_X2 U11652 ( .A(U214), .ZN(n16668) );
  AND2_X1 U11653 ( .A1(n12142), .A2(n12141), .ZN(n12146) );
  AND4_X1 U11654 ( .A1(n12151), .A2(n12150), .A3(n12149), .A4(n12148), .ZN(
        n12157) );
  CLKBUF_X1 U11655 ( .A(n9815), .Z(n13000) );
  INV_X2 U11656 ( .A(n12434), .ZN(n12752) );
  INV_X2 U11657 ( .A(n12986), .ZN(n12610) );
  INV_X1 U11658 ( .A(n9810), .ZN(n9930) );
  INV_X2 U11659 ( .A(n18345), .ZN(n9828) );
  INV_X2 U11660 ( .A(n12988), .ZN(n9952) );
  INV_X2 U11661 ( .A(n20895), .ZN(n9829) );
  OR2_X1 U11662 ( .A1(n10556), .A2(n9895), .ZN(n9894) );
  NAND2_X2 U11663 ( .A1(n20050), .A2(n19917), .ZN(n19974) );
  NAND2_X1 U11664 ( .A1(n10458), .A2(n9874), .ZN(n9873) );
  INV_X1 U11665 ( .A(n12909), .ZN(n12998) );
  NAND2_X2 U11666 ( .A1(n18955), .A2(n18888), .ZN(n18947) );
  INV_X1 U11667 ( .A(n17166), .ZN(n17342) );
  BUF_X2 U11668 ( .A(n17122), .Z(n16071) );
  INV_X2 U11669 ( .A(n20142), .ZN(n20164) );
  INV_X2 U11670 ( .A(n12294), .ZN(n12751) );
  AND2_X1 U11671 ( .A1(n10645), .A2(n10644), .ZN(n10649) );
  BUF_X4 U11672 ( .A(n10405), .Z(n9830) );
  INV_X2 U11673 ( .A(n16704), .ZN(U215) );
  NAND2_X1 U11674 ( .A1(n9942), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12150) );
  CLKBUF_X3 U11675 ( .A(n10378), .Z(n17299) );
  INV_X1 U11676 ( .A(n12909), .ZN(n9962) );
  OR2_X1 U11677 ( .A1(n18826), .A2(n10242), .ZN(n10556) );
  INV_X2 U11678 ( .A(n20939), .ZN(n20927) );
  BUF_X4 U11679 ( .A(n10424), .Z(n9832) );
  INV_X2 U11680 ( .A(n16708), .ZN(n16710) );
  INV_X2 U11681 ( .A(n17063), .ZN(n18825) );
  OR2_X1 U11682 ( .A1(n10345), .A2(n18818), .ZN(n17166) );
  NOR2_X1 U11683 ( .A1(n10344), .A2(n18818), .ZN(n17122) );
  NAND2_X2 U11685 ( .A1(n12094), .A2(n12095), .ZN(n12988) );
  NAND2_X1 U11686 ( .A1(n13886), .A2(n9951), .ZN(n12848) );
  NAND2_X1 U11687 ( .A1(n13536), .A2(n12088), .ZN(n12232) );
  NAND2_X2 U11688 ( .A1(n12093), .A2(n13886), .ZN(n12959) );
  NAND2_X1 U11689 ( .A1(n12093), .A2(n13885), .ZN(n12909) );
  AND2_X2 U11690 ( .A1(n12093), .A2(n12087), .ZN(n12855) );
  AND3_X2 U11691 ( .A1(n9838), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10862) );
  AND2_X2 U11692 ( .A1(n11118), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10863) );
  NAND2_X1 U11693 ( .A1(n18969), .A2(n18994), .ZN(n10242) );
  AND2_X2 U11694 ( .A1(n11118), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9953) );
  NOR2_X2 U11695 ( .A1(n9855), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12095) );
  NAND2_X1 U11696 ( .A1(n18979), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n18830) );
  BUF_X1 U11697 ( .A(n13900), .Z(n9950) );
  NAND2_X1 U11698 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17992) );
  INV_X1 U11699 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9907) );
  INV_X1 U11700 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9908) );
  INV_X1 U11701 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9855) );
  AND2_X1 U11702 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13885) );
  NOR2_X2 U11703 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13900) );
  INV_X1 U11704 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12381) );
  INV_X2 U11705 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12088) );
  INV_X1 U11706 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14250) );
  AND2_X1 U11707 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11118) );
  INV_X2 U11708 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13802) );
  NOR2_X1 U11709 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10641) );
  AND2_X1 U11710 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13783) );
  INV_X1 U11711 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9838) );
  INV_X1 U11712 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10058) );
  NAND2_X1 U11713 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10345) );
  NAND2_X1 U11714 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18799) );
  INV_X2 U11715 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18969) );
  INV_X2 U11716 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18994) );
  NAND2_X1 U11717 ( .A1(n9838), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11096) );
  AOI21_X1 U11718 ( .B1(n13819), .B2(n9837), .A(n9836), .ZN(n13816) );
  AND2_X1 U11719 ( .A1(n10759), .A2(n9838), .ZN(n9836) );
  XNOR2_X1 U11720 ( .A(n9932), .B(n9838), .ZN(n9837) );
  XNOR2_X2 U11721 ( .A(n11297), .B(n9839), .ZN(n11299) );
  OAI21_X2 U11722 ( .B1(n9960), .B2(n14030), .A(n10807), .ZN(n9839) );
  NAND2_X1 U11723 ( .A1(n9841), .A2(n10925), .ZN(n9923) );
  NAND2_X1 U11724 ( .A1(n10927), .A2(n10928), .ZN(n9841) );
  NAND2_X2 U11725 ( .A1(n9842), .A2(n11089), .ZN(n15717) );
  NAND2_X1 U11726 ( .A1(n15728), .A2(n15730), .ZN(n9842) );
  NAND2_X1 U11727 ( .A1(n9844), .A2(n10986), .ZN(n9843) );
  OAI22_X1 U11728 ( .A1(n14013), .A2(n14012), .B1(n14030), .B2(n10984), .ZN(
        n9844) );
  AND2_X2 U11729 ( .A1(n10813), .A2(n10840), .ZN(n9845) );
  NAND2_X2 U11730 ( .A1(n9846), .A2(n10762), .ZN(n11703) );
  INV_X2 U11731 ( .A(n11513), .ZN(n11507) );
  OAI21_X1 U11732 ( .B1(n10291), .B2(n9851), .A(n9850), .ZN(n9847) );
  INV_X1 U11733 ( .A(n9849), .ZN(n9848) );
  INV_X1 U11734 ( .A(n14430), .ZN(n9850) );
  INV_X1 U11735 ( .A(n10291), .ZN(n14659) );
  INV_X1 U11736 ( .A(n14427), .ZN(n9851) );
  OAI21_X1 U11737 ( .B1(n13855), .B2(n13854), .A(n9852), .ZN(n14173) );
  XNOR2_X1 U11738 ( .A(n14008), .B(n9852), .ZN(n20187) );
  NAND2_X1 U11739 ( .A1(n9853), .A2(n16165), .ZN(n13753) );
  NAND2_X2 U11740 ( .A1(n9853), .A2(n20243), .ZN(n14378) );
  NAND2_X2 U11741 ( .A1(n13309), .A2(n9853), .ZN(n13069) );
  OAI21_X2 U11742 ( .B1(n9898), .B2(n9853), .A(n13696), .ZN(n13862) );
  NOR2_X2 U11743 ( .A1(n20178), .A2(n9853), .ZN(n13682) );
  NOR2_X2 U11744 ( .A1(n20276), .A2(n9853), .ZN(n20797) );
  INV_X2 U11745 ( .A(n12268), .ZN(n9853) );
  AND2_X2 U11746 ( .A1(n14209), .A2(n14233), .ZN(n14232) );
  NOR2_X2 U11747 ( .A1(n14161), .A2(n14160), .ZN(n14159) );
  NAND2_X2 U11748 ( .A1(n12284), .A2(n12283), .ZN(n12391) );
  NAND2_X2 U11749 ( .A1(n12364), .A2(n12276), .ZN(n12284) );
  XNOR2_X2 U11750 ( .A(n10064), .B(n12272), .ZN(n20358) );
  INV_X1 U11751 ( .A(n12784), .ZN(n14743) );
  NOR2_X2 U11752 ( .A1(n14685), .A2(n14686), .ZN(n14670) );
  AND2_X2 U11753 ( .A1(n12784), .A2(n9854), .ZN(n14726) );
  AND2_X2 U11754 ( .A1(n10052), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12094) );
  INV_X1 U11755 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10052) );
  INV_X1 U11756 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U11757 ( .A1(n17979), .A2(n10449), .ZN(n17962) );
  NAND2_X1 U11758 ( .A1(n17980), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17979) );
  INV_X1 U11759 ( .A(n18005), .ZN(n9862) );
  NAND2_X1 U11760 ( .A1(n18003), .A2(n10442), .ZN(n17987) );
  NAND2_X1 U11761 ( .A1(n18004), .A2(n18005), .ZN(n18003) );
  AND2_X1 U11762 ( .A1(n9866), .A2(n17826), .ZN(n17714) );
  NAND2_X1 U11763 ( .A1(n9866), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9865) );
  NOR2_X1 U11764 ( .A1(n17734), .A2(n18091), .ZN(n9867) );
  AND2_X1 U11766 ( .A1(n9828), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n9870) );
  INV_X1 U11767 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9871) );
  NOR2_X1 U11768 ( .A1(n17877), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17858) );
  INV_X1 U11769 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n9874) );
  NAND3_X1 U11770 ( .A1(n9903), .A2(n18263), .A3(n17952), .ZN(n17904) );
  NAND3_X1 U11771 ( .A1(n9878), .A2(n10975), .A3(n11169), .ZN(n10135) );
  AND2_X1 U11772 ( .A1(n9877), .A2(n10925), .ZN(n10975) );
  NAND2_X1 U11773 ( .A1(n10927), .A2(n10928), .ZN(n9877) );
  INV_X1 U11774 ( .A(n10974), .ZN(n9878) );
  NAND4_X1 U11775 ( .A1(n10861), .A2(n10860), .A3(n10858), .A4(n10859), .ZN(
        n10897) );
  INV_X1 U11776 ( .A(n11206), .ZN(n9881) );
  NAND2_X1 U11777 ( .A1(n10800), .A2(n10799), .ZN(n9888) );
  OAI211_X2 U11778 ( .C1(n10800), .C2(n9887), .A(n9885), .B(n9883), .ZN(n11765) );
  NAND2_X1 U11779 ( .A1(n10800), .A2(n9884), .ZN(n9883) );
  NOR2_X1 U11780 ( .A1(n11299), .A2(n9886), .ZN(n9884) );
  NAND2_X1 U11781 ( .A1(n9886), .A2(n11299), .ZN(n9885) );
  OAI21_X1 U11782 ( .B1(n9888), .B2(n11299), .A(n11298), .ZN(n13624) );
  NAND2_X2 U11783 ( .A1(n13873), .A2(n13874), .ZN(n14340) );
  OAI211_X2 U11784 ( .C1(n15152), .C2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10042), .B(n9889), .ZN(n13873) );
  NAND2_X1 U11785 ( .A1(n13861), .A2(n13860), .ZN(n15150) );
  XNOR2_X1 U11786 ( .A(n13867), .B(n20232), .ZN(n15151) );
  INV_X1 U11787 ( .A(n16179), .ZN(n18031) );
  XNOR2_X1 U11788 ( .A(n9812), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18024) );
  NAND3_X1 U11789 ( .A1(n10387), .A2(n10389), .A3(n10388), .ZN(n10436) );
  NOR2_X2 U11790 ( .A1(n17724), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17723) );
  INV_X1 U11791 ( .A(n9892), .ZN(n9891) );
  NAND2_X1 U11792 ( .A1(n17822), .A2(n18145), .ZN(n17821) );
  OAI211_X1 U11793 ( .C1(n16059), .C2(n17344), .A(n9894), .B(n9893), .ZN(
        n10431) );
  NAND2_X1 U11794 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n9893) );
  INV_X1 U11795 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U11796 ( .A1(n11483), .A2(n9896), .ZN(n11695) );
  OAI211_X2 U11797 ( .C1(n9897), .C2(n11707), .A(n11483), .B(n9896), .ZN(
        n10759) );
  NAND3_X1 U11798 ( .A1(n11277), .A2(n10738), .A3(n13364), .ZN(n9897) );
  INV_X2 U11799 ( .A(n11508), .ZN(n11277) );
  INV_X1 U11800 ( .A(n10731), .ZN(n10729) );
  NAND2_X1 U11801 ( .A1(n10452), .A2(n10453), .ZN(n10454) );
  OAI21_X2 U11802 ( .B1(n12371), .B2(n9898), .A(n12366), .ZN(n12388) );
  XNOR2_X2 U11803 ( .A(n9920), .B(n9898), .ZN(n13913) );
  OAI21_X4 U11804 ( .B1(n13748), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12365), 
        .ZN(n9898) );
  NAND2_X1 U11805 ( .A1(n9899), .A2(n11158), .ZN(n16500) );
  NAND2_X1 U11806 ( .A1(n14189), .A2(n14190), .ZN(n9899) );
  NAND2_X1 U11807 ( .A1(n9901), .A2(n9900), .ZN(n14189) );
  NAND2_X1 U11808 ( .A1(n14011), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9900) );
  NAND2_X2 U11809 ( .A1(n20268), .A2(n12268), .ZN(n14480) );
  INV_X1 U11810 ( .A(n9906), .ZN(n9933) );
  AND2_X2 U11811 ( .A1(n9908), .A2(n9907), .ZN(n13886) );
  AND2_X2 U11812 ( .A1(n12381), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12093) );
  NAND2_X1 U11813 ( .A1(n20184), .A2(n9909), .ZN(n16297) );
  INV_X1 U11814 ( .A(n10302), .ZN(n9909) );
  AND2_X2 U11815 ( .A1(n14346), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10302) );
  NAND2_X2 U11816 ( .A1(n14405), .A2(n10303), .ZN(n15136) );
  NAND2_X2 U11817 ( .A1(n14402), .A2(n14401), .ZN(n14405) );
  INV_X2 U11818 ( .A(n10803), .ZN(n11402) );
  NAND2_X1 U11819 ( .A1(n11402), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10790) );
  INV_X1 U11820 ( .A(n9942), .ZN(n12850) );
  AND2_X2 U11821 ( .A1(n9950), .A2(n12094), .ZN(n9942) );
  AND2_X2 U11822 ( .A1(n14329), .A2(n11366), .ZN(n15413) );
  INV_X1 U11823 ( .A(n9933), .ZN(n15601) );
  OAI22_X1 U11824 ( .A1(n14013), .A2(n14012), .B1(n10984), .B2(n14030), .ZN(
        n9910) );
  AND2_X1 U11825 ( .A1(n16534), .A2(n16502), .ZN(n9911) );
  AND2_X1 U11826 ( .A1(n19337), .A2(n16533), .ZN(n9912) );
  AND2_X1 U11827 ( .A1(n16503), .A2(n16532), .ZN(n9913) );
  NOR3_X1 U11828 ( .A1(n9911), .A2(n9912), .A3(n9913), .ZN(n16470) );
  INV_X2 U11829 ( .A(n14038), .ZN(n11819) );
  OR2_X2 U11830 ( .A1(n12986), .A2(n12140), .ZN(n12141) );
  NAND2_X1 U11831 ( .A1(n10119), .A2(n9971), .ZN(n9914) );
  XNOR2_X1 U11832 ( .A(n10291), .B(n14427), .ZN(n14649) );
  OR2_X1 U11833 ( .A1(n13592), .A2(n12245), .ZN(n12258) );
  OAI22_X1 U11834 ( .A1(n13705), .A2(n19347), .B1(n11003), .B2(n10950), .ZN(
        n10951) );
  AND4_X2 U11835 ( .A1(n12146), .A2(n12145), .A3(n9985), .A4(n12144), .ZN(
        n12158) );
  OR2_X2 U11836 ( .A1(n15431), .A2(n15430), .ZN(n15495) );
  AOI21_X2 U11837 ( .B1(n17393), .B2(n17098), .A(n17147), .ZN(n17137) );
  NOR2_X2 U11838 ( .A1(n16935), .A2(n17295), .ZN(n17258) );
  NOR2_X2 U11839 ( .A1(n17362), .A2(n17361), .ZN(n17366) );
  INV_X1 U11840 ( .A(n18809), .ZN(n18817) );
  NAND2_X2 U11841 ( .A1(n18820), .A2(n13151), .ZN(n18812) );
  NOR2_X2 U11842 ( .A1(n15450), .A2(n11980), .ZN(n12003) );
  NOR2_X2 U11843 ( .A1(n14072), .A2(n10014), .ZN(n13435) );
  NOR2_X2 U11844 ( .A1(n13632), .A2(n10148), .ZN(n14043) );
  NOR2_X2 U11845 ( .A1(n15404), .A2(n15405), .ZN(n15389) );
  NAND2_X1 U11846 ( .A1(n10041), .A2(n9918), .ZN(n9915) );
  OR2_X1 U11847 ( .A1(n9917), .A2(n12376), .ZN(n9916) );
  INV_X1 U11848 ( .A(n12339), .ZN(n9917) );
  AND2_X1 U11849 ( .A1(n12336), .A2(n12339), .ZN(n9918) );
  NAND2_X1 U11850 ( .A1(n15012), .A2(n15030), .ZN(n9919) );
  NAND2_X1 U11851 ( .A1(n12366), .A2(n12360), .ZN(n9920) );
  AND2_X1 U11852 ( .A1(n15089), .A2(n9921), .ZN(n15066) );
  AND2_X1 U11853 ( .A1(n15088), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9921) );
  AOI21_X2 U11854 ( .B1(n15051), .B2(n15190), .A(n14546), .ZN(n15012) );
  NAND2_X1 U11855 ( .A1(n12366), .A2(n12360), .ZN(n12371) );
  AND2_X1 U11856 ( .A1(n10897), .A2(n10116), .ZN(n10115) );
  NAND2_X1 U11857 ( .A1(n15457), .A2(n15456), .ZN(n15455) );
  INV_X1 U11858 ( .A(n11777), .ZN(n13818) );
  NAND2_X1 U11859 ( .A1(n10928), .A2(n10927), .ZN(n9924) );
  OR2_X2 U11860 ( .A1(n13592), .A2(n12245), .ZN(n9925) );
  NAND2_X1 U11861 ( .A1(n12206), .A2(n12205), .ZN(n9926) );
  NAND2_X1 U11862 ( .A1(n12206), .A2(n12205), .ZN(n12250) );
  INV_X1 U11863 ( .A(n13780), .ZN(n9927) );
  NAND2_X1 U11864 ( .A1(n11520), .A2(n11508), .ZN(n11661) );
  INV_X1 U11865 ( .A(n9810), .ZN(n9928) );
  INV_X1 U11866 ( .A(n9810), .ZN(n9929) );
  INV_X1 U11867 ( .A(n9810), .ZN(n9931) );
  INV_X1 U11868 ( .A(n10738), .ZN(n19384) );
  AND4_X1 U11869 ( .A1(n10751), .A2(n11511), .A3(n19373), .A4(n10738), .ZN(
        n11702) );
  OR2_X2 U11870 ( .A1(n13359), .A2(n13358), .ZN(n13357) );
  NOR2_X2 U11871 ( .A1(n12007), .A2(n12004), .ZN(n15441) );
  NOR2_X2 U11872 ( .A1(n15449), .A2(n15451), .ZN(n15450) );
  INV_X1 U11873 ( .A(n10738), .ZN(n10722) );
  NOR2_X1 U11874 ( .A1(n10699), .A2(n10751), .ZN(n10739) );
  INV_X1 U11875 ( .A(n13108), .ZN(n10579) );
  AOI21_X2 U11876 ( .B1(n10584), .B2(n15992), .A(n10588), .ZN(n18819) );
  AND2_X2 U11877 ( .A1(n10722), .A2(n11508), .ZN(n12066) );
  NOR2_X1 U11878 ( .A1(n9926), .A2(n12222), .ZN(n9934) );
  INV_X1 U11879 ( .A(n15040), .ZN(n9935) );
  NAND2_X2 U11880 ( .A1(n15058), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9936) );
  CLKBUF_X1 U11881 ( .A(n13866), .Z(n9937) );
  NOR2_X1 U11882 ( .A1(n12250), .A2(n12222), .ZN(n13309) );
  NAND2_X2 U11883 ( .A1(n13618), .A2(n11798), .ZN(n13617) );
  AOI21_X2 U11884 ( .B1(n11795), .B2(n11796), .A(n11794), .ZN(n13618) );
  NAND2_X2 U11885 ( .A1(n13536), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12516) );
  INV_X1 U11887 ( .A(n12294), .ZN(n9940) );
  MUX2_X2 U11889 ( .A(n12204), .B(n12221), .S(n20263), .Z(n12205) );
  NAND2_X2 U11890 ( .A1(n12252), .A2(n12188), .ZN(n12254) );
  OR2_X2 U11891 ( .A1(n14308), .A2(n14900), .ZN(n9979) );
  NOR2_X1 U11892 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10346), .ZN(
        n10380) );
  AND2_X1 U11893 ( .A1(n12095), .A2(n12087), .ZN(n9946) );
  AND2_X1 U11894 ( .A1(n12095), .A2(n12087), .ZN(n9947) );
  OAI211_X2 U11895 ( .C1(n9959), .C2(n13367), .A(n10782), .B(n10781), .ZN(
        n10815) );
  AOI21_X2 U11896 ( .B1(n10302), .B2(n16296), .A(n10000), .ZN(n10301) );
  NOR2_X2 U11897 ( .A1(n13942), .A2(n11804), .ZN(n13943) );
  NOR2_X2 U11898 ( .A1(n14755), .A2(n14757), .ZN(n12784) );
  XNOR2_X2 U11899 ( .A(n11911), .B(n11910), .ZN(n15470) );
  INV_X1 U11900 ( .A(n11680), .ZN(n9948) );
  INV_X1 U11901 ( .A(n11668), .ZN(n9949) );
  OAI21_X2 U11902 ( .B1(n13562), .B2(n13872), .A(n13561), .ZN(n13563) );
  XNOR2_X2 U11903 ( .A(n14346), .B(n14521), .ZN(n20183) );
  NAND2_X2 U11904 ( .A1(n14340), .A2(n14339), .ZN(n14346) );
  AND2_X1 U11905 ( .A1(n9951), .A2(n12087), .ZN(n9958) );
  BUF_X1 U11906 ( .A(n10803), .Z(n9960) );
  INV_X2 U11907 ( .A(n12909), .ZN(n9961) );
  NAND2_X1 U11908 ( .A1(n11693), .A2(n10324), .ZN(n10749) );
  INV_X1 U11909 ( .A(n12475), .ZN(n12477) );
  AOI21_X1 U11910 ( .B1(n11402), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10737), .ZN(n10792) );
  OR2_X1 U11911 ( .A1(n11300), .A2(n10734), .ZN(n10735) );
  NAND2_X1 U11912 ( .A1(n10756), .A2(n10755), .ZN(n10779) );
  NAND2_X1 U11913 ( .A1(n10754), .A2(n9819), .ZN(n10755) );
  NAND2_X1 U11914 ( .A1(n10238), .A2(n14861), .ZN(n10237) );
  AND2_X1 U11915 ( .A1(n14404), .A2(n14435), .ZN(n10303) );
  INV_X1 U11916 ( .A(n14434), .ZN(n14435) );
  INV_X1 U11917 ( .A(n12376), .ZN(n10040) );
  INV_X1 U11918 ( .A(n13059), .ZN(n13052) );
  NAND2_X1 U11919 ( .A1(n11267), .A2(n11283), .ZN(n11266) );
  NOR2_X1 U11920 ( .A1(n9984), .A2(n10194), .ZN(n10193) );
  INV_X1 U11921 ( .A(n11189), .ZN(n10194) );
  NOR2_X1 U11922 ( .A1(n11141), .A2(n11140), .ZN(n11155) );
  NAND2_X1 U11923 ( .A1(n11400), .A2(n14250), .ZN(n10768) );
  NAND2_X1 U11924 ( .A1(n9819), .A2(n19361), .ZN(n10731) );
  INV_X1 U11925 ( .A(n15480), .ZN(n10267) );
  NOR2_X1 U11926 ( .A1(n11031), .A2(n11030), .ZN(n11551) );
  AND2_X1 U11927 ( .A1(n14194), .A2(n14102), .ZN(n10144) );
  INV_X1 U11928 ( .A(n15602), .ZN(n10186) );
  OR2_X1 U11929 ( .A1(n10200), .A2(n11285), .ZN(n15593) );
  INV_X1 U11930 ( .A(n11043), .ZN(n10089) );
  NAND2_X1 U11931 ( .A1(n13838), .A2(n10748), .ZN(n11693) );
  AND4_X1 U11932 ( .A1(n10578), .A2(n15993), .A3(n10577), .A4(n10576), .ZN(
        n10587) );
  NOR3_X1 U11933 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n18830), .ZN(n10394) );
  AOI21_X1 U11934 ( .B1(n18848), .B2(n18375), .A(n18827), .ZN(n16176) );
  OAI211_X1 U11935 ( .C1(n10577), .C2(n18383), .A(n10573), .B(n10572), .ZN(
        n13106) );
  NOR2_X1 U11936 ( .A1(n18379), .A2(n10569), .ZN(n10575) );
  NAND2_X1 U11937 ( .A1(n14670), .A2(n10289), .ZN(n10291) );
  NOR2_X1 U11938 ( .A1(n14660), .A2(n10290), .ZN(n10289) );
  INV_X1 U11939 ( .A(n14672), .ZN(n10290) );
  AND2_X1 U11940 ( .A1(n14169), .A2(n14168), .ZN(n14167) );
  AND2_X1 U11941 ( .A1(n15334), .A2(n14523), .ZN(n16334) );
  NOR2_X1 U11942 ( .A1(n12163), .A2(n10316), .ZN(n12186) );
  NAND2_X1 U11943 ( .A1(n12378), .A2(n20932), .ZN(n10041) );
  NAND2_X1 U11944 ( .A1(n12378), .A2(n10037), .ZN(n10036) );
  NOR2_X1 U11945 ( .A1(n10040), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U11946 ( .A1(n13206), .A2(n9977), .ZN(n15353) );
  NAND2_X1 U11947 ( .A1(n14573), .A2(n16407), .ZN(n16405) );
  AND2_X1 U11948 ( .A1(n11197), .A2(n11324), .ZN(n11202) );
  NOR2_X1 U11949 ( .A1(n15353), .A2(n16381), .ZN(n15352) );
  NOR2_X2 U11950 ( .A1(n10180), .A2(n10179), .ZN(n15429) );
  INV_X1 U11951 ( .A(n15426), .ZN(n10179) );
  NOR2_X1 U11952 ( .A1(n16392), .A2(n11169), .ZN(n11468) );
  XNOR2_X1 U11953 ( .A(n15496), .B(n14592), .ZN(n15374) );
  NAND2_X1 U11954 ( .A1(n10151), .A2(n13930), .ZN(n10150) );
  INV_X1 U11955 ( .A(n13198), .ZN(n10151) );
  AND2_X1 U11956 ( .A1(n11504), .A2(n13362), .ZN(n11753) );
  NAND2_X1 U11957 ( .A1(n18379), .A2(n10587), .ZN(n13108) );
  AND2_X1 U11958 ( .A1(n16759), .A2(n10084), .ZN(n16752) );
  NOR2_X1 U11959 ( .A1(n16740), .A2(n16763), .ZN(n16591) );
  NOR2_X1 U11960 ( .A1(n10309), .A2(n15808), .ZN(n10308) );
  INV_X1 U11961 ( .A(n15744), .ZN(n10310) );
  NOR2_X1 U11962 ( .A1(n10058), .A2(n20932), .ZN(n10063) );
  AOI22_X1 U11963 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10659) );
  NOR2_X1 U11964 ( .A1(n12381), .A2(n20932), .ZN(n10297) );
  AOI22_X1 U11965 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10863), .B1(
        n10652), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10670) );
  AND4_X1 U11966 ( .A1(n11056), .A2(n11055), .A3(n11054), .A4(n11053), .ZN(
        n11083) );
  AND4_X1 U11967 ( .A1(n11080), .A2(n11079), .A3(n11078), .A4(n11077), .ZN(
        n11081) );
  NAND2_X1 U11968 ( .A1(n10753), .A2(n13364), .ZN(n11712) );
  AOI22_X1 U11969 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9954), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10655) );
  OR2_X1 U11970 ( .A1(n10249), .A2(n17535), .ZN(n10445) );
  INV_X1 U11971 ( .A(n12387), .ZN(n10282) );
  NAND2_X1 U11972 ( .A1(n14815), .A2(n10285), .ZN(n14755) );
  AND2_X1 U11973 ( .A1(n10286), .A2(n14853), .ZN(n10285) );
  OR2_X1 U11974 ( .A1(n13015), .A2(n20929), .ZN(n13010) );
  CLKBUF_X1 U11975 ( .A(n12716), .Z(n13741) );
  NOR2_X1 U11976 ( .A1(n14788), .A2(n10011), .ZN(n10238) );
  INV_X1 U11977 ( .A(n12501), .ZN(n10066) );
  INV_X1 U11978 ( .A(n10068), .ZN(n10067) );
  NAND2_X1 U11979 ( .A1(n10068), .A2(n12501), .ZN(n14357) );
  INV_X1 U11980 ( .A(n14510), .ZN(n14504) );
  NAND2_X1 U11981 ( .A1(n14467), .A2(n14517), .ZN(n14510) );
  NOR2_X1 U11982 ( .A1(n20268), .A2(n20263), .ZN(n13881) );
  NAND2_X1 U11983 ( .A1(n20527), .A2(n20932), .ZN(n12413) );
  AND2_X1 U11985 ( .A1(n11979), .A2(n10331), .ZN(n11980) );
  AND2_X1 U11986 ( .A1(n10269), .A2(n15484), .ZN(n10268) );
  NOR2_X1 U11987 ( .A1(n10971), .A2(n10970), .ZN(n11550) );
  NOR2_X1 U11988 ( .A1(n15705), .A2(n10220), .ZN(n10219) );
  NOR2_X1 U11989 ( .A1(n16472), .A2(n10223), .ZN(n10222) );
  INV_X1 U11990 ( .A(n13168), .ZN(n10214) );
  NAND2_X1 U11991 ( .A1(n10802), .A2(n10801), .ZN(n11297) );
  NAND2_X1 U11992 ( .A1(n13223), .A2(n10175), .ZN(n10180) );
  AND2_X1 U11993 ( .A1(n10177), .A2(n10176), .ZN(n10175) );
  INV_X1 U11994 ( .A(n11403), .ZN(n10176) );
  OR2_X1 U11995 ( .A1(n14573), .A2(n11169), .ZN(n11286) );
  INV_X1 U11996 ( .A(n11274), .ZN(n10133) );
  NOR2_X1 U11997 ( .A1(n9988), .A2(n15629), .ZN(n10132) );
  OR2_X1 U11998 ( .A1(n10273), .A2(n10274), .ZN(n10272) );
  NOR2_X1 U11999 ( .A1(n11264), .A2(n10275), .ZN(n10274) );
  NAND2_X1 U12000 ( .A1(n10272), .A2(n10138), .ZN(n10137) );
  INV_X1 U12001 ( .A(n15642), .ZN(n10138) );
  NAND2_X1 U12002 ( .A1(n15568), .A2(n10026), .ZN(n14283) );
  INV_X1 U12003 ( .A(n15690), .ZN(n11093) );
  AND2_X1 U12004 ( .A1(n14178), .A2(n14213), .ZN(n10185) );
  OR2_X1 U12005 ( .A1(n13727), .A2(n10166), .ZN(n13934) );
  NAND2_X1 U12006 ( .A1(n10167), .A2(n13936), .ZN(n10166) );
  INV_X1 U12007 ( .A(n10168), .ZN(n10167) );
  NAND2_X1 U12008 ( .A1(n10171), .A2(n13722), .ZN(n10170) );
  INV_X1 U12009 ( .A(n13713), .ZN(n10171) );
  NAND2_X1 U12010 ( .A1(n11085), .A2(n14578), .ZN(n11088) );
  INV_X1 U12011 ( .A(n11044), .ZN(n11085) );
  AND2_X1 U12012 ( .A1(n11494), .A2(n13364), .ZN(n10727) );
  OAI21_X1 U12013 ( .B1(n10726), .B2(n10725), .A(n10724), .ZN(n10728) );
  OR2_X1 U12014 ( .A1(n10738), .A2(n14134), .ZN(n10726) );
  OAI21_X1 U12015 ( .B1(n11159), .B2(n11165), .A(n11036), .ZN(n10160) );
  NOR2_X1 U12016 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  NAND2_X1 U12017 ( .A1(n10763), .A2(n10729), .ZN(n13781) );
  INV_X1 U12018 ( .A(n10763), .ZN(n13814) );
  OAI211_X1 U12019 ( .C1(n10742), .C2(n10741), .A(n20035), .B(n10740), .ZN(
        n11711) );
  AND2_X1 U12020 ( .A1(n10839), .A2(n13532), .ZN(n19517) );
  AOI21_X1 U12021 ( .B1(n10652), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10644) );
  NAND2_X1 U12022 ( .A1(n10863), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10645) );
  NOR2_X1 U12023 ( .A1(n10345), .A2(n18830), .ZN(n10424) );
  NOR2_X1 U12024 ( .A1(n16775), .A2(n10071), .ZN(n10070) );
  INV_X1 U12025 ( .A(n17829), .ZN(n10069) );
  INV_X1 U12026 ( .A(n10454), .ZN(n10053) );
  AOI21_X1 U12027 ( .B1(n17524), .B2(n16601), .A(n17826), .ZN(n10453) );
  INV_X1 U12028 ( .A(n17528), .ZN(n10609) );
  NAND2_X1 U12029 ( .A1(n18014), .A2(n10438), .ZN(n10441) );
  OR2_X1 U12030 ( .A1(n18329), .A2(n10437), .ZN(n10438) );
  NAND2_X1 U12031 ( .A1(n9812), .A2(n17543), .ZN(n10440) );
  XNOR2_X1 U12032 ( .A(n9812), .B(n17543), .ZN(n10437) );
  NOR2_X1 U12033 ( .A1(n10345), .A2(n18825), .ZN(n10406) );
  NOR2_X2 U12034 ( .A1(n10533), .A2(n10532), .ZN(n10585) );
  OR2_X1 U12035 ( .A1(n13458), .A2(n13581), .ZN(n14623) );
  NAND2_X1 U12036 ( .A1(n14831), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13752) );
  INV_X1 U12037 ( .A(n13686), .ZN(n12385) );
  NOR2_X1 U12038 ( .A1(n12268), .A2(n20243), .ZN(n13588) );
  AND2_X1 U12039 ( .A1(n12950), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12951) );
  NAND2_X1 U12040 ( .A1(n12899), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12949) );
  NOR2_X1 U12041 ( .A1(n10280), .A2(n14703), .ZN(n10279) );
  INV_X1 U12042 ( .A(n10008), .ZN(n10280) );
  NAND2_X1 U12043 ( .A1(n10232), .A2(n14683), .ZN(n10231) );
  INV_X1 U12044 ( .A(n10233), .ZN(n10232) );
  NOR3_X1 U12045 ( .A1(n14741), .A2(n10234), .A3(n10233), .ZN(n14700) );
  NOR2_X1 U12046 ( .A1(n14741), .A2(n14733), .ZN(n14735) );
  AND2_X1 U12047 ( .A1(n14089), .A2(n14001), .ZN(n14002) );
  NAND2_X1 U12048 ( .A1(n13563), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13864) );
  OAI211_X1 U12049 ( .C1(n13052), .C2(n12788), .A(n12338), .B(n12337), .ZN(
        n12376) );
  INV_X1 U12050 ( .A(n12336), .ZN(n10039) );
  INV_X1 U12051 ( .A(n12306), .ZN(n10298) );
  NAND2_X1 U12052 ( .A1(n20932), .A2(n20242), .ZN(n20406) );
  INV_X1 U12053 ( .A(n16153), .ZN(n14625) );
  AND2_X1 U12054 ( .A1(n13913), .A2(n13562), .ZN(n20718) );
  AND2_X1 U12055 ( .A1(n13914), .A2(n13920), .ZN(n20719) );
  NAND2_X1 U12056 ( .A1(n20932), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10056) );
  NOR2_X1 U12057 ( .A1(n16405), .A2(n11293), .ZN(n11475) );
  NAND2_X1 U12058 ( .A1(n13206), .A2(n10216), .ZN(n15356) );
  OAI22_X1 U12059 ( .A1(n15381), .A2(n10025), .B1(n10206), .B2(n16424), .ZN(
        n16422) );
  OAI21_X1 U12060 ( .B1(n11282), .B2(n10029), .A(n10198), .ZN(n10201) );
  NAND2_X1 U12061 ( .A1(n11282), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U12062 ( .A1(n15397), .A2(n19206), .ZN(n15381) );
  NAND2_X1 U12063 ( .A1(n10205), .A2(n15619), .ZN(n10207) );
  INV_X1 U12064 ( .A(n15381), .ZN(n10205) );
  NAND2_X1 U12065 ( .A1(n11249), .A2(n10196), .ZN(n11246) );
  AND2_X1 U12066 ( .A1(n13739), .A2(n10190), .ZN(n10189) );
  NAND2_X1 U12067 ( .A1(n11213), .A2(n11283), .ZN(n11211) );
  NAND2_X1 U12068 ( .A1(n10193), .A2(n11186), .ZN(n10192) );
  INV_X1 U12069 ( .A(n13205), .ZN(n19206) );
  AND2_X1 U12070 ( .A1(n11428), .A2(n11128), .ZN(n13828) );
  AND2_X1 U12071 ( .A1(n11356), .A2(n11355), .ZN(n14218) );
  NOR2_X1 U12072 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10157) );
  NOR2_X1 U12073 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10156) );
  NOR2_X1 U12074 ( .A1(n10762), .A2(n10731), .ZN(n10732) );
  NAND2_X1 U12075 ( .A1(n12046), .A2(n12062), .ZN(n10260) );
  NOR2_X1 U12076 ( .A1(n10257), .A2(n12062), .ZN(n10256) );
  INV_X1 U12077 ( .A(n15430), .ZN(n10257) );
  OR2_X1 U12078 ( .A1(n15465), .A2(n15472), .ZN(n10264) );
  OR2_X1 U12079 ( .A1(n15470), .A2(n15472), .ZN(n10266) );
  AND2_X1 U12080 ( .A1(n10141), .A2(n13319), .ZN(n10140) );
  OR2_X1 U12081 ( .A1(n10144), .A2(n10142), .ZN(n10141) );
  INV_X1 U12082 ( .A(n11552), .ZN(n10142) );
  NAND2_X1 U12083 ( .A1(n14192), .A2(n10144), .ZN(n14100) );
  INV_X1 U12084 ( .A(n11405), .ZN(n13332) );
  NAND2_X1 U12085 ( .A1(n13210), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13217) );
  NAND2_X1 U12086 ( .A1(n13163), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13214) );
  NAND2_X1 U12087 ( .A1(n13223), .A2(n10177), .ZN(n15446) );
  NOR2_X1 U12088 ( .A1(n10114), .A2(n15808), .ZN(n10113) );
  NAND2_X1 U12089 ( .A1(n15413), .A2(n10181), .ZN(n15403) );
  AND2_X1 U12090 ( .A1(n10182), .A2(n9972), .ZN(n10181) );
  INV_X1 U12091 ( .A(n15401), .ZN(n10182) );
  NAND2_X1 U12092 ( .A1(n10149), .A2(n16509), .ZN(n10148) );
  INV_X1 U12093 ( .A(n10150), .ZN(n10149) );
  XNOR2_X1 U12094 ( .A(n11088), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15730) );
  NAND2_X1 U12095 ( .A1(n13702), .A2(n13728), .ZN(n13727) );
  INV_X1 U12096 ( .A(n10751), .ZN(n10746) );
  AND2_X1 U12097 ( .A1(n19988), .A2(n20017), .ZN(n19578) );
  AND2_X1 U12098 ( .A1(n19998), .A2(n20007), .ZN(n19639) );
  INV_X1 U12099 ( .A(n19759), .ZN(n19640) );
  INV_X1 U12100 ( .A(n19758), .ZN(n19756) );
  OR2_X1 U12101 ( .A1(n19988), .A2(n20017), .ZN(n19789) );
  OR2_X1 U12102 ( .A1(n19988), .A2(n19342), .ZN(n19759) );
  INV_X1 U12103 ( .A(n19788), .ZN(n19838) );
  INV_X1 U12104 ( .A(n19833), .ZN(n19792) );
  OAI21_X1 U12105 ( .B1(n10595), .B2(n10594), .A(n10593), .ZN(n18793) );
  INV_X1 U12106 ( .A(n17803), .ZN(n17792) );
  NAND2_X1 U12107 ( .A1(n10450), .A2(n10609), .ZN(n16601) );
  AOI21_X2 U12108 ( .B1(n10585), .B2(n18819), .A(n14415), .ZN(n18820) );
  XNOR2_X1 U12109 ( .A(n10437), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18016) );
  INV_X1 U12110 ( .A(n18793), .ZN(n16172) );
  INV_X2 U12111 ( .A(n19014), .ZN(n18375) );
  AOI211_X1 U12112 ( .C1(n9814), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n10540), .B(n10539), .ZN(n10541) );
  AND2_X1 U12113 ( .A1(n14615), .A2(n13747), .ZN(n20084) );
  OR2_X1 U12114 ( .A1(n20189), .A2(n13567), .ZN(n15131) );
  AND2_X1 U12115 ( .A1(n16131), .A2(n13585), .ZN(n20189) );
  XNOR2_X1 U12116 ( .A(n10044), .B(n15006), .ZN(n15167) );
  NAND2_X1 U12117 ( .A1(n10046), .A2(n10045), .ZN(n10044) );
  NAND2_X1 U12118 ( .A1(n15004), .A2(n10012), .ZN(n10045) );
  NAND2_X1 U12119 ( .A1(n15005), .A2(n15140), .ZN(n10046) );
  NAND2_X1 U12120 ( .A1(n10054), .A2(n9997), .ZN(n15216) );
  INV_X1 U12121 ( .A(n15232), .ZN(n10054) );
  OR2_X1 U12122 ( .A1(n20363), .A2(n20628), .ZN(n20403) );
  OR2_X1 U12123 ( .A1(n20497), .A2(n20628), .ZN(n20525) );
  INV_X1 U12124 ( .A(n13838), .ZN(n20027) );
  NAND2_X1 U12125 ( .A1(n16503), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10109) );
  OAI21_X1 U12126 ( .B1(n15578), .B2(n10105), .A(n15581), .ZN(n10104) );
  NAND2_X1 U12127 ( .A1(n16503), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10105) );
  NAND2_X1 U12128 ( .A1(n15588), .A2(n11292), .ZN(n11296) );
  NAND2_X1 U12129 ( .A1(n20004), .A2(n19833), .ZN(n14136) );
  OR2_X1 U12130 ( .A1(n13253), .A2(n19356), .ZN(n19333) );
  AND2_X1 U12131 ( .A1(n11733), .A2(n11732), .ZN(n11751) );
  OR2_X1 U12132 ( .A1(n15379), .A2(n15976), .ZN(n11732) );
  INV_X1 U12133 ( .A(n15976), .ZN(n16565) );
  INV_X1 U12134 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20012) );
  NAND2_X1 U12135 ( .A1(n13833), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15988) );
  INV_X1 U12136 ( .A(n16755), .ZN(n10075) );
  OR2_X1 U12137 ( .A1(n16769), .A2(n18950), .ZN(n10074) );
  XNOR2_X1 U12138 ( .A(n16752), .B(n16751), .ZN(n10077) );
  NAND2_X1 U12139 ( .A1(n12093), .A2(n12094), .ZN(n12294) );
  NAND2_X1 U12140 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12018) );
  NAND2_X1 U12141 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12011) );
  NAND2_X1 U12142 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U12143 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11972) );
  NAND2_X1 U12144 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11965) );
  AOI21_X1 U12145 ( .B1(n10652), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n10099), .ZN(n10098) );
  NAND2_X1 U12146 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10095) );
  INV_X1 U12147 ( .A(n19829), .ZN(n11010) );
  INV_X1 U12148 ( .A(n19700), .ZN(n10993) );
  AND4_X1 U12149 ( .A1(n11068), .A2(n11067), .A3(n11066), .A4(n11065), .ZN(
        n11082) );
  OR2_X1 U12150 ( .A1(n10476), .A2(n10477), .ZN(n10472) );
  INV_X1 U12151 ( .A(n20268), .ZN(n12247) );
  AOI21_X1 U12153 ( .B1(n10300), .B2(n10063), .A(n12257), .ZN(n10061) );
  NAND2_X1 U12154 ( .A1(n9925), .A2(n10063), .ZN(n10062) );
  NOR2_X1 U12155 ( .A1(n10762), .A2(n19032), .ZN(n10757) );
  CLKBUF_X1 U12156 ( .A(n9818), .Z(n12028) );
  NAND2_X1 U12157 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12034) );
  NAND2_X1 U12158 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12027) );
  INV_X1 U12159 ( .A(n11089), .ZN(n10102) );
  INV_X1 U12160 ( .A(n11159), .ZN(n10161) );
  AOI22_X1 U12161 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n10956), .B1(
        n19797), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10960) );
  NAND2_X1 U12162 ( .A1(n19373), .A2(n19384), .ZN(n10162) );
  NAND2_X1 U12163 ( .A1(n10722), .A2(n10721), .ZN(n10752) );
  NAND2_X1 U12164 ( .A1(n10250), .A2(n17540), .ZN(n10249) );
  INV_X1 U12165 ( .A(n10440), .ZN(n10250) );
  NOR2_X1 U12166 ( .A1(n10585), .A2(n10597), .ZN(n10576) );
  AND2_X1 U12167 ( .A1(n10059), .A2(n20243), .ZN(n13029) );
  NAND2_X1 U12168 ( .A1(n10059), .A2(n12239), .ZN(n13078) );
  INV_X1 U12169 ( .A(n12253), .ZN(n13084) );
  NOR2_X1 U12170 ( .A1(n10010), .A2(n10287), .ZN(n10286) );
  INV_X1 U12171 ( .A(n10288), .ZN(n10287) );
  NOR2_X1 U12172 ( .A1(n12643), .A2(n16230), .ZN(n12721) );
  AND2_X1 U12173 ( .A1(n14883), .A2(n14796), .ZN(n10288) );
  NAND2_X1 U12174 ( .A1(n10278), .A2(n10277), .ZN(n14812) );
  INV_X1 U12175 ( .A(n14810), .ZN(n10277) );
  INV_X1 U12176 ( .A(n14308), .ZN(n10278) );
  XNOR2_X1 U12177 ( .A(n14356), .B(n12504), .ZN(n14366) );
  INV_X1 U12178 ( .A(n14698), .ZN(n10234) );
  OR2_X1 U12179 ( .A1(n10235), .A2(n14733), .ZN(n10233) );
  INV_X1 U12180 ( .A(n14713), .ZN(n10235) );
  NAND2_X1 U12181 ( .A1(n15106), .A2(n14440), .ZN(n15095) );
  INV_X1 U12182 ( .A(n14374), .ZN(n14379) );
  OR2_X1 U12183 ( .A1(n12411), .A2(n12410), .ZN(n14349) );
  NAND2_X1 U12184 ( .A1(n12168), .A2(n12167), .ZN(n12169) );
  INV_X1 U12185 ( .A(n20263), .ZN(n13578) );
  NAND2_X1 U12186 ( .A1(n10296), .A2(n10294), .ZN(n12307) );
  NAND2_X1 U12187 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  OR2_X1 U12188 ( .A1(n10295), .A2(n10297), .ZN(n10292) );
  INV_X1 U12189 ( .A(n12396), .ZN(n14376) );
  NAND2_X1 U12190 ( .A1(n13751), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12397) );
  OR2_X1 U12191 ( .A1(n12301), .A2(n20932), .ZN(n12396) );
  INV_X1 U12192 ( .A(n12302), .ZN(n13869) );
  OAI211_X1 U12193 ( .C1(n20245), .C2(n13566), .A(n12282), .B(n12281), .ZN(
        n12283) );
  OR2_X1 U12194 ( .A1(n12280), .A2(n10052), .ZN(n12282) );
  AOI22_X1 U12195 ( .A1(n9962), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12212) );
  OAI21_X1 U12196 ( .B1(n13906), .B2(n16368), .A(n20914), .ZN(n20242) );
  INV_X1 U12197 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20585) );
  OR2_X1 U12198 ( .A1(n10896), .A2(n10895), .ZN(n11099) );
  NOR2_X1 U12199 ( .A1(n16410), .A2(n10217), .ZN(n10216) );
  INV_X1 U12200 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10217) );
  NAND2_X1 U12201 ( .A1(n11249), .A2(n10195), .ZN(n11267) );
  NOR2_X1 U12202 ( .A1(n10197), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10195) );
  NOR2_X1 U12203 ( .A1(n11161), .A2(n9984), .ZN(n11190) );
  OAI21_X1 U12204 ( .B1(n11111), .B2(n14575), .A(n11139), .ZN(n11140) );
  NAND2_X1 U12205 ( .A1(n14575), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11139) );
  OR2_X1 U12206 ( .A1(n11568), .A2(n11567), .ZN(n11799) );
  AOI21_X1 U12207 ( .B1(n10863), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n10032), .ZN(n12057) );
  NAND2_X1 U12208 ( .A1(n10153), .A2(n15502), .ZN(n10152) );
  INV_X1 U12209 ( .A(n15510), .ZN(n10153) );
  NAND2_X1 U12210 ( .A1(n15455), .A2(n11961), .ZN(n11979) );
  INV_X1 U12211 ( .A(n15465), .ZN(n10265) );
  NOR2_X1 U12212 ( .A1(n11861), .A2(n14041), .ZN(n10269) );
  NOR2_X1 U12213 ( .A1(n10204), .A2(n10203), .ZN(n10202) );
  NAND2_X1 U12214 ( .A1(n13213), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13215) );
  NOR2_X1 U12215 ( .A1(n10178), .A2(n15444), .ZN(n10177) );
  INV_X1 U12216 ( .A(n13224), .ZN(n10178) );
  AND2_X1 U12217 ( .A1(n15389), .A2(n15390), .ZN(n15388) );
  OR2_X1 U12218 ( .A1(n16110), .A2(n11169), .ZN(n11269) );
  NAND2_X1 U12219 ( .A1(n10307), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10306) );
  NOR2_X1 U12220 ( .A1(n15853), .A2(n15662), .ZN(n10307) );
  INV_X1 U12221 ( .A(n15559), .ZN(n10145) );
  OAI21_X1 U12222 ( .B1(n15728), .B2(n10102), .A(n10100), .ZN(n15690) );
  INV_X1 U12223 ( .A(n10101), .ZN(n10100) );
  OAI21_X1 U12224 ( .B1(n15730), .B2(n10102), .A(n10304), .ZN(n10101) );
  AND2_X1 U12225 ( .A1(n15913), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10304) );
  INV_X1 U12226 ( .A(n13941), .ZN(n11335) );
  NAND2_X1 U12227 ( .A1(n10169), .A2(n13735), .ZN(n10168) );
  INV_X1 U12228 ( .A(n10170), .ZN(n10169) );
  NAND2_X1 U12229 ( .A1(n10155), .A2(n13404), .ZN(n10154) );
  INV_X1 U12230 ( .A(n14071), .ZN(n10155) );
  AND2_X1 U12231 ( .A1(n10978), .A2(n10925), .ZN(n10117) );
  NAND2_X1 U12232 ( .A1(n11507), .A2(n14134), .ZN(n10762) );
  OR2_X1 U12233 ( .A1(n11135), .A2(n14575), .ZN(n11525) );
  AOI22_X1 U12234 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10718) );
  XNOR2_X1 U12235 ( .A(n10797), .B(n10810), .ZN(n10811) );
  NAND2_X1 U12236 ( .A1(n10658), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10665) );
  AOI22_X1 U12237 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9953), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10680) );
  AOI21_X1 U12238 ( .B1(n10652), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n10124), .ZN(n10123) );
  NAND2_X1 U12239 ( .A1(n10125), .A2(n13827), .ZN(n10124) );
  OR2_X1 U12240 ( .A1(n10854), .A2(n10852), .ZN(n19829) );
  NAND3_X1 U12241 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18986), .A3(
        n18994), .ZN(n10346) );
  NAND2_X1 U12242 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18969), .ZN(
        n10344) );
  NOR2_X1 U12243 ( .A1(n10344), .A2(n18825), .ZN(n10405) );
  NOR2_X1 U12244 ( .A1(n17531), .A2(n10445), .ZN(n10450) );
  NAND2_X1 U12245 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18799), .ZN(
        n18818) );
  NOR2_X1 U12246 ( .A1(n10523), .A2(n10522), .ZN(n10578) );
  NOR2_X1 U12247 ( .A1(n10554), .A2(n10553), .ZN(n15993) );
  OR2_X1 U12248 ( .A1(n20934), .A2(n13743), .ZN(n14831) );
  NAND2_X1 U12249 ( .A1(n13953), .A2(n13952), .ZN(n13959) );
  AND2_X1 U12250 ( .A1(n12764), .A2(n12763), .ZN(n14853) );
  AND3_X1 U12251 ( .A1(n12525), .A2(n12524), .A3(n12523), .ZN(n14207) );
  INV_X1 U12252 ( .A(n12370), .ZN(n10284) );
  AOI21_X1 U12253 ( .B1(n12370), .B2(n10283), .A(n10282), .ZN(n10281) );
  NAND2_X1 U12254 ( .A1(n13913), .A2(n12640), .ZN(n12375) );
  AND2_X1 U12255 ( .A1(n12898), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12899) );
  OR2_X1 U12256 ( .A1(n15017), .A2(n12982), .ZN(n12927) );
  AND2_X1 U12257 ( .A1(n12873), .A2(n12872), .ZN(n14711) );
  OR2_X1 U12258 ( .A1(n15035), .A2(n12982), .ZN(n12873) );
  OR2_X1 U12259 ( .A1(n12785), .A2(n15061), .ZN(n12786) );
  OR2_X1 U12260 ( .A1(n12786), .A2(n14746), .ZN(n12843) );
  CLKBUF_X1 U12261 ( .A(n14755), .Z(n14756) );
  AND2_X1 U12262 ( .A1(n12679), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12659) );
  NAND2_X1 U12263 ( .A1(n12626), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12643) );
  NAND2_X1 U12264 ( .A1(n14815), .A2(n10288), .ZN(n14886) );
  AND2_X1 U12265 ( .A1(n14815), .A2(n14796), .ZN(n14884) );
  INV_X1 U12266 ( .A(n12590), .ZN(n12623) );
  AND2_X1 U12267 ( .A1(n12560), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12561) );
  NAND2_X1 U12268 ( .A1(n12527), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12556) );
  INV_X1 U12269 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20073) );
  NAND2_X1 U12270 ( .A1(n12505), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12522) );
  AOI21_X1 U12271 ( .B1(n14357), .B2(n12640), .A(n12498), .ZN(n14092) );
  CLKBUF_X1 U12272 ( .A(n13986), .Z(n13987) );
  NAND2_X1 U12273 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12418) );
  NOR2_X1 U12274 ( .A1(n12418), .A2(n12417), .ZN(n12466) );
  INV_X1 U12275 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12417) );
  NAND2_X1 U12276 ( .A1(n10276), .A2(n12387), .ZN(n13855) );
  AND2_X1 U12277 ( .A1(n15014), .A2(n9976), .ZN(n14552) );
  OR2_X1 U12278 ( .A1(n14856), .A2(n14498), .ZN(n14741) );
  NAND2_X1 U12279 ( .A1(n10240), .A2(n10239), .ZN(n14856) );
  INV_X1 U12280 ( .A(n14854), .ZN(n10239) );
  INV_X1 U12281 ( .A(n10240), .ZN(n14863) );
  INV_X1 U12282 ( .A(n10238), .ZN(n10236) );
  NOR2_X1 U12283 ( .A1(n14877), .A2(n14788), .ZN(n14868) );
  OR2_X1 U12284 ( .A1(n14882), .A2(n14875), .ZN(n14877) );
  NAND2_X1 U12285 ( .A1(n14801), .A2(n14880), .ZN(n14882) );
  NOR2_X1 U12286 ( .A1(n14893), .A2(n14817), .ZN(n14819) );
  OR2_X1 U12287 ( .A1(n14901), .A2(n14891), .ZN(n14893) );
  NAND2_X1 U12288 ( .A1(n10228), .A2(n10227), .ZN(n14901) );
  INV_X1 U12289 ( .A(n14904), .ZN(n10227) );
  INV_X1 U12290 ( .A(n14903), .ZN(n10228) );
  NAND2_X1 U12291 ( .A1(n10226), .A2(n10224), .ZN(n14903) );
  NOR2_X1 U12292 ( .A1(n9965), .A2(n10225), .ZN(n10224) );
  INV_X1 U12293 ( .A(n14315), .ZN(n10225) );
  NOR2_X1 U12294 ( .A1(n14229), .A2(n9965), .ZN(n14316) );
  NAND2_X1 U12295 ( .A1(n10226), .A2(n10229), .ZN(n14239) );
  AND2_X1 U12296 ( .A1(n14000), .A2(n13999), .ZN(n14001) );
  NAND2_X1 U12297 ( .A1(n10043), .A2(n14520), .ZN(n10042) );
  INV_X1 U12298 ( .A(n13868), .ZN(n10043) );
  AND4_X1 U12299 ( .A1(n13953), .A2(n13957), .A3(n13952), .A4(n10241), .ZN(
        n14090) );
  INV_X1 U12300 ( .A(n13972), .ZN(n10241) );
  OR2_X1 U12301 ( .A1(n13958), .A2(n13959), .ZN(n13973) );
  XNOR2_X1 U12302 ( .A(n13864), .B(n13862), .ZN(n13697) );
  INV_X1 U12303 ( .A(n14523), .ZN(n14539) );
  AND2_X1 U12304 ( .A1(n13612), .A2(n13611), .ZN(n20221) );
  NAND4_X1 U12305 ( .A1(n13881), .A2(n9938), .A3(n13086), .A4(n10059), .ZN(
        n13595) );
  NAND2_X1 U12306 ( .A1(n13599), .A2(n13598), .ZN(n13949) );
  NOR2_X1 U12307 ( .A1(n13587), .A2(n12187), .ZN(n12188) );
  OR2_X1 U12308 ( .A1(n20238), .A2(n13914), .ZN(n20629) );
  INV_X1 U12309 ( .A(n13587), .ZN(n12301) );
  INV_X1 U12310 ( .A(n20276), .ZN(n20289) );
  AND2_X1 U12311 ( .A1(n10188), .A2(n10187), .ZN(n11111) );
  NAND2_X1 U12312 ( .A1(n11505), .A2(n11418), .ZN(n10187) );
  NAND2_X1 U12313 ( .A1(n11541), .A2(n20026), .ZN(n10188) );
  NAND2_X1 U12314 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  INV_X1 U12315 ( .A(n16403), .ZN(n10208) );
  INV_X1 U12316 ( .A(n16402), .ZN(n10209) );
  NAND2_X1 U12317 ( .A1(n13206), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15354) );
  OR2_X1 U12318 ( .A1(n13226), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16404) );
  OR2_X1 U12319 ( .A1(n11275), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10199) );
  OAI21_X1 U12320 ( .B1(n19206), .B2(n16103), .A(n16102), .ZN(n15398) );
  INV_X1 U12321 ( .A(n10193), .ZN(n10191) );
  OR2_X1 U12322 ( .A1(n11161), .A2(n11160), .ZN(n11180) );
  NOR2_X1 U12323 ( .A1(n10780), .A2(n10335), .ZN(n10781) );
  AND2_X1 U12324 ( .A1(n13846), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10765) );
  NAND2_X1 U12325 ( .A1(n10120), .A2(n13827), .ZN(n10129) );
  INV_X1 U12326 ( .A(n10667), .ZN(n10121) );
  CLKBUF_X1 U12327 ( .A(n15404), .Z(n15540) );
  NAND2_X1 U12328 ( .A1(n15568), .A2(n14201), .ZN(n15558) );
  NOR2_X1 U12329 ( .A1(n15793), .A2(n11388), .ZN(n10311) );
  NAND2_X1 U12330 ( .A1(n13208), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13209) );
  AND2_X1 U12331 ( .A1(n9973), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10218) );
  NAND2_X1 U12332 ( .A1(n13213), .A2(n9973), .ZN(n13216) );
  NAND2_X1 U12333 ( .A1(n13165), .A2(n9968), .ZN(n13174) );
  AND2_X1 U12334 ( .A1(n9968), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10221) );
  NAND2_X1 U12335 ( .A1(n13165), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13172) );
  NAND2_X1 U12336 ( .A1(n13167), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13171) );
  NOR2_X1 U12337 ( .A1(n16507), .A2(n10215), .ZN(n10212) );
  NOR2_X1 U12338 ( .A1(n10213), .A2(n16507), .ZN(n10211) );
  NOR2_X1 U12339 ( .A1(n14015), .A2(n13168), .ZN(n13170) );
  NAND2_X1 U12340 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13168) );
  NOR2_X1 U12341 ( .A1(n15578), .A2(n15759), .ZN(n10106) );
  AND2_X1 U12342 ( .A1(n15593), .A2(n11288), .ZN(n11470) );
  XNOR2_X1 U12343 ( .A(n11286), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15594) );
  AND2_X1 U12344 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15807), .ZN(
        n15794) );
  INV_X1 U12345 ( .A(n15616), .ZN(n10131) );
  NAND2_X1 U12346 ( .A1(n11382), .A2(n11381), .ZN(n15459) );
  INV_X1 U12347 ( .A(n15403), .ZN(n11382) );
  NAND2_X1 U12348 ( .A1(n9824), .A2(n10305), .ZN(n15612) );
  NOR2_X1 U12349 ( .A1(n10306), .A2(n15820), .ZN(n10305) );
  NAND2_X1 U12350 ( .A1(n15413), .A2(n9972), .ZN(n15477) );
  INV_X1 U12351 ( .A(n10272), .ZN(n10139) );
  CLKBUF_X1 U12352 ( .A(n14283), .Z(n15416) );
  AND2_X1 U12353 ( .A1(n15694), .A2(n15693), .ZN(n15683) );
  AND2_X1 U12354 ( .A1(n10185), .A2(n10184), .ZN(n10183) );
  INV_X1 U12355 ( .A(n14218), .ZN(n10184) );
  OAI21_X1 U12356 ( .B1(n15700), .B2(n15701), .A(n15652), .ZN(n15694) );
  NAND2_X1 U12357 ( .A1(n14060), .A2(n10185), .ZN(n14217) );
  INV_X1 U12358 ( .A(n16454), .ZN(n10163) );
  AND2_X1 U12359 ( .A1(n14060), .A2(n14178), .ZN(n14212) );
  AND2_X1 U12360 ( .A1(n11720), .A2(n16542), .ZN(n15914) );
  AND3_X1 U12361 ( .A1(n11585), .A2(n11584), .A3(n11583), .ZN(n13436) );
  AND3_X1 U12362 ( .A1(n11321), .A2(n11320), .A3(n11319), .ZN(n13713) );
  CLKBUF_X1 U12363 ( .A(n15970), .Z(n15971) );
  AND3_X1 U12364 ( .A1(n11312), .A2(n11311), .A3(n11310), .ZN(n13701) );
  NAND2_X1 U12365 ( .A1(n13625), .A2(n13636), .ZN(n13700) );
  AND3_X1 U12366 ( .A1(n11544), .A2(n11543), .A3(n11542), .ZN(n14026) );
  AND2_X1 U12367 ( .A1(n11701), .A2(n11700), .ZN(n13784) );
  AND2_X1 U12368 ( .A1(n11533), .A2(n11532), .ZN(n13343) );
  NAND2_X1 U12369 ( .A1(n13344), .A2(n13343), .ZN(n13342) );
  NAND2_X1 U12370 ( .A1(n11481), .A2(n11430), .ZN(n13833) );
  INV_X1 U12371 ( .A(n19675), .ZN(n10992) );
  AND2_X1 U12372 ( .A1(n19998), .A2(n19986), .ZN(n19984) );
  INV_X1 U12373 ( .A(n19789), .ZN(n19668) );
  NAND2_X2 U12374 ( .A1(n10651), .A2(n10650), .ZN(n19361) );
  INV_X1 U12375 ( .A(n19389), .ZN(n19379) );
  INV_X1 U12376 ( .A(n19388), .ZN(n19377) );
  OR2_X1 U12377 ( .A1(n19998), .A2(n20007), .ZN(n19788) );
  INV_X1 U12378 ( .A(n10733), .ZN(n13848) );
  NAND2_X1 U12379 ( .A1(n16174), .A2(n18375), .ZN(n10580) );
  OR3_X1 U12380 ( .A1(n18848), .A2(n14415), .A3(n18827), .ZN(n18792) );
  NOR2_X1 U12381 ( .A1(n16771), .A2(n17047), .ZN(n16761) );
  OR2_X1 U12382 ( .A1(n16761), .A2(n16762), .ZN(n16759) );
  OAI22_X1 U12383 ( .A1(n16784), .A2(n10082), .B1(n10084), .B2(n16772), .ZN(
        n16771) );
  NAND2_X1 U12384 ( .A1(n17672), .A2(n10083), .ZN(n10082) );
  INV_X1 U12385 ( .A(n17684), .ZN(n10083) );
  OR2_X1 U12386 ( .A1(n16784), .A2(n17684), .ZN(n10085) );
  AND2_X1 U12387 ( .A1(n16827), .A2(n10084), .ZN(n16816) );
  OR2_X1 U12388 ( .A1(n16829), .A2(n17752), .ZN(n16827) );
  NAND2_X1 U12389 ( .A1(n10079), .A2(n10078), .ZN(n10080) );
  AOI21_X1 U12390 ( .B1(n16960), .B2(n17781), .A(n17773), .ZN(n10078) );
  NAND2_X1 U12391 ( .A1(n16848), .A2(n10084), .ZN(n10079) );
  OR2_X1 U12392 ( .A1(n16848), .A2(n17781), .ZN(n10081) );
  NAND2_X1 U12393 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17366), .ZN(n17324) );
  NAND2_X1 U12394 ( .A1(n17667), .A2(n9975), .ZN(n16740) );
  NAND2_X1 U12395 ( .A1(n17680), .A2(n17826), .ZN(n10165) );
  NAND4_X1 U12396 ( .A1(n10069), .A2(n16937), .A3(n10602), .A4(n10327), .ZN(
        n10603) );
  INV_X1 U12397 ( .A(n10603), .ZN(n16889) );
  NAND2_X1 U12398 ( .A1(n16937), .A2(n10327), .ZN(n17866) );
  NAND2_X1 U12399 ( .A1(n10086), .A2(n9998), .ZN(n17960) );
  INV_X1 U12400 ( .A(n17992), .ZN(n10086) );
  NOR2_X1 U12401 ( .A1(n18844), .A2(n18856), .ZN(n10601) );
  INV_X1 U12402 ( .A(n11449), .ZN(n11446) );
  NOR2_X1 U12403 ( .A1(n18043), .A2(n13128), .ZN(n16589) );
  NOR2_X1 U12404 ( .A1(n17854), .A2(n18147), .ZN(n18168) );
  NOR2_X1 U12405 ( .A1(n18200), .A2(n9874), .ZN(n17849) );
  NAND2_X1 U12406 ( .A1(n10174), .A2(n10173), .ZN(n10172) );
  NOR2_X1 U12407 ( .A1(n9876), .A2(n18263), .ZN(n18227) );
  INV_X1 U12408 ( .A(n17826), .ZN(n17932) );
  INV_X1 U12409 ( .A(n10453), .ZN(n10248) );
  XNOR2_X1 U12410 ( .A(n10450), .B(n17970), .ZN(n17963) );
  XNOR2_X1 U12411 ( .A(n10447), .B(n10446), .ZN(n17980) );
  INV_X1 U12412 ( .A(n10448), .ZN(n10446) );
  NAND2_X1 U12413 ( .A1(n18015), .A2(n18016), .ZN(n18014) );
  INV_X1 U12414 ( .A(n18820), .ZN(n18816) );
  NOR2_X2 U12415 ( .A1(n13151), .A2(n18816), .ZN(n18827) );
  INV_X1 U12416 ( .A(n10578), .ZN(n18383) );
  INV_X1 U12417 ( .A(n10585), .ZN(n18392) );
  AOI22_X1 U12418 ( .A1(n18797), .A2(n18790), .B1(n18795), .B2(n18791), .ZN(
        n18844) );
  NOR2_X2 U12419 ( .A1(n10493), .A2(n10492), .ZN(n19014) );
  OR2_X1 U12420 ( .A1(n13316), .A2(n14634), .ZN(n13324) );
  INV_X1 U12421 ( .A(n14378), .ZN(n20930) );
  INV_X1 U12422 ( .A(n14839), .ZN(n20075) );
  INV_X1 U12423 ( .A(n20104), .ZN(n20127) );
  AND2_X1 U12424 ( .A1(n13761), .A2(n13760), .ZN(n20126) );
  AND2_X1 U12425 ( .A1(n14897), .A2(n12187), .ZN(n14906) );
  INV_X1 U12426 ( .A(n14906), .ZN(n14898) );
  INV_X1 U12427 ( .A(n14957), .ZN(n14966) );
  INV_X1 U12428 ( .A(n14983), .ZN(n14965) );
  NAND2_X1 U12429 ( .A1(n13439), .A2(n13585), .ZN(n13083) );
  OR2_X1 U12430 ( .A1(n14965), .A2(n13769), .ZN(n14986) );
  BUF_X1 U12431 ( .A(n16167), .Z(n20163) );
  INV_X1 U12432 ( .A(n13652), .ZN(n20179) );
  OR2_X1 U12433 ( .A1(n13744), .A2(n14557), .ZN(n13745) );
  INV_X1 U12434 ( .A(n15131), .ZN(n20182) );
  XNOR2_X1 U12435 ( .A(n14519), .B(n14518), .ZN(n14636) );
  NAND2_X1 U12436 ( .A1(n15014), .A2(n14457), .ZN(n10065) );
  AND2_X1 U12437 ( .A1(n15197), .A2(n14537), .ZN(n15180) );
  NAND2_X1 U12438 ( .A1(n15248), .A2(n14530), .ZN(n15232) );
  NOR2_X1 U12439 ( .A1(n14542), .A2(n16303), .ZN(n15260) );
  NAND2_X1 U12440 ( .A1(n16297), .A2(n16296), .ZN(n16295) );
  OAI21_X1 U12441 ( .B1(n14523), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n15330), .ZN(n20212) );
  INV_X1 U12442 ( .A(n20225), .ZN(n20205) );
  OR2_X1 U12443 ( .A1(n13612), .A2(n10057), .ZN(n15330) );
  INV_X1 U12444 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20690) );
  NAND2_X1 U12445 ( .A1(n10041), .A2(n9994), .ZN(n10034) );
  NAND2_X1 U12446 ( .A1(n10039), .A2(n12376), .ZN(n10038) );
  AND2_X2 U12447 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13537) );
  AND2_X1 U12448 ( .A1(n13463), .A2(n13455), .ZN(n20918) );
  OR2_X1 U12449 ( .A1(n20363), .A2(n20454), .ZN(n20394) );
  OAI21_X1 U12450 ( .B1(n20423), .B2(n20407), .A(n20730), .ZN(n20425) );
  INV_X1 U12451 ( .A(n20441), .ZN(n20450) );
  OAI211_X1 U12452 ( .C1(n20550), .C2(n20664), .A(n20589), .B(n20534), .ZN(
        n20552) );
  INV_X1 U12453 ( .A(n20525), .ZN(n20551) );
  OAI211_X1 U12454 ( .C1(n20592), .C2(n20591), .A(n20590), .B(n20589), .ZN(
        n20617) );
  OAI211_X1 U12455 ( .C1(n20681), .C2(n20664), .A(n20730), .B(n20663), .ZN(
        n20683) );
  NOR2_X2 U12456 ( .A1(n20629), .A2(n20628), .ZN(n20682) );
  INV_X1 U12457 ( .A(n20782), .ZN(n20724) );
  INV_X1 U12458 ( .A(n20783), .ZN(n20725) );
  INV_X1 U12459 ( .A(n20803), .ZN(n20742) );
  INV_X1 U12460 ( .A(n20809), .ZN(n20747) );
  INV_X1 U12461 ( .A(n20810), .ZN(n20748) );
  INV_X1 U12462 ( .A(n20816), .ZN(n20753) );
  INV_X1 U12463 ( .A(n20817), .ZN(n20754) );
  INV_X1 U12464 ( .A(n20832), .ZN(n20764) );
  OAI211_X1 U12465 ( .C1(n20770), .C2(n20731), .A(n20730), .B(n20729), .ZN(
        n20773) );
  INV_X1 U12466 ( .A(n20732), .ZN(n20772) );
  AND2_X1 U12467 ( .A1(n20719), .A2(n20241), .ZN(n20843) );
  INV_X1 U12468 ( .A(n20614), .ZN(n20840) );
  NAND2_X1 U12469 ( .A1(n13065), .A2(n10056), .ZN(n10055) );
  INV_X1 U12470 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20849) );
  NAND2_X1 U12471 ( .A1(n15429), .A2(n14584), .ZN(n14591) );
  NAND2_X1 U12472 ( .A1(n16378), .A2(n19223), .ZN(n16385) );
  OR2_X1 U12473 ( .A1(n16379), .A2(n19217), .ZN(n16384) );
  OAI22_X1 U12474 ( .A1(n16402), .A2(n10024), .B1(n10206), .B2(n16394), .ZN(
        n16393) );
  AND2_X1 U12475 ( .A1(n10210), .A2(n10206), .ZN(n16395) );
  NAND2_X1 U12476 ( .A1(n11294), .A2(n10339), .ZN(n16392) );
  NOR2_X1 U12477 ( .A1(n15357), .A2(n19206), .ZN(n16402) );
  INV_X1 U12478 ( .A(n10210), .ZN(n16401) );
  NAND2_X1 U12479 ( .A1(n11283), .A2(n16404), .ZN(n14573) );
  AND2_X1 U12480 ( .A1(n10207), .A2(n10206), .ZN(n16423) );
  INV_X1 U12481 ( .A(n10207), .ZN(n15380) );
  NAND2_X1 U12482 ( .A1(n11202), .A2(n13739), .ZN(n11203) );
  OR2_X1 U12483 ( .A1(n15358), .A2(n13182), .ZN(n19168) );
  INV_X1 U12484 ( .A(n19199), .ZN(n19220) );
  OR2_X1 U12485 ( .A1(n20043), .A2(n13186), .ZN(n19217) );
  NOR2_X1 U12486 ( .A1(n10206), .A2(n19895), .ZN(n19228) );
  INV_X1 U12487 ( .A(n19155), .ZN(n19229) );
  INV_X1 U12488 ( .A(n19202), .ZN(n19223) );
  AND2_X1 U12489 ( .A1(n11801), .A2(n10271), .ZN(n10270) );
  INV_X1 U12490 ( .A(n13721), .ZN(n10271) );
  OR2_X1 U12491 ( .A1(n11595), .A2(n11594), .ZN(n13733) );
  CLKBUF_X1 U12492 ( .A(n13731), .Z(n13732) );
  OR2_X1 U12493 ( .A1(n11782), .A2(n13386), .ZN(n19342) );
  NAND2_X1 U12494 ( .A1(n15496), .A2(n14592), .ZN(n14596) );
  INV_X1 U12495 ( .A(n10259), .ZN(n10258) );
  OAI22_X1 U12496 ( .A1(n15430), .A2(n10260), .B1(n12046), .B2(n12062), .ZN(
        n10259) );
  AND2_X1 U12497 ( .A1(n10263), .A2(n10266), .ZN(n15463) );
  INV_X1 U12498 ( .A(n10323), .ZN(n10263) );
  INV_X1 U12499 ( .A(n10266), .ZN(n15471) );
  AND2_X1 U12500 ( .A1(n19250), .A2(n12067), .ZN(n16430) );
  NAND2_X1 U12501 ( .A1(n14100), .A2(n11552), .ZN(n13320) );
  NOR2_X1 U12502 ( .A1(n14193), .A2(n10143), .ZN(n14101) );
  INV_X1 U12503 ( .A(n14194), .ZN(n10143) );
  AND2_X1 U12504 ( .A1(n19257), .A2(n15552), .ZN(n19252) );
  INV_X1 U12505 ( .A(n19250), .ZN(n19284) );
  CLKBUF_X1 U12507 ( .A(n13515), .Z(n20047) );
  INV_X1 U12508 ( .A(n13329), .ZN(n13305) );
  XNOR2_X1 U12509 ( .A(n13176), .B(n13175), .ZN(n14608) );
  INV_X1 U12510 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16507) );
  NAND2_X1 U12511 ( .A1(n13253), .A2(n11433), .ZN(n16506) );
  AND2_X1 U12512 ( .A1(n16506), .A2(n13411), .ZN(n16496) );
  INV_X1 U12513 ( .A(n16496), .ZN(n19341) );
  INV_X1 U12514 ( .A(n19333), .ZN(n16502) );
  NAND2_X1 U12515 ( .A1(n10112), .A2(n10111), .ZN(n15743) );
  NAND2_X1 U12516 ( .A1(n10103), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10111) );
  NAND2_X1 U12517 ( .A1(n15577), .A2(n10106), .ZN(n10112) );
  INV_X1 U12518 ( .A(n15578), .ZN(n10103) );
  OR2_X1 U12519 ( .A1(n15803), .A2(n11748), .ZN(n15799) );
  OR2_X1 U12520 ( .A1(n15872), .A2(n11744), .ZN(n15838) );
  NOR2_X1 U12521 ( .A1(n13632), .A2(n10150), .ZN(n16508) );
  NAND2_X1 U12522 ( .A1(n15643), .A2(n16454), .ZN(n10164) );
  NAND2_X1 U12523 ( .A1(n11217), .A2(n15721), .ZN(n16455) );
  NAND2_X1 U12524 ( .A1(n15719), .A2(n15642), .ZN(n11217) );
  CLKBUF_X1 U12525 ( .A(n15728), .Z(n15729) );
  CLKBUF_X1 U12526 ( .A(n15973), .Z(n15974) );
  NOR2_X2 U12527 ( .A1(n11754), .A2(n20030), .ZN(n16566) );
  NAND2_X1 U12528 ( .A1(n11753), .A2(n11731), .ZN(n15976) );
  INV_X1 U12529 ( .A(n19342), .ZN(n20017) );
  INV_X1 U12530 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20011) );
  INV_X1 U12531 ( .A(n19986), .ZN(n20007) );
  INV_X1 U12532 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20002) );
  XNOR2_X1 U12533 ( .A(n13468), .B(n13471), .ZN(n19998) );
  XNOR2_X1 U12534 ( .A(n13469), .B(n13470), .ZN(n13471) );
  CLKBUF_X1 U12535 ( .A(n13530), .Z(n13531) );
  CLKBUF_X1 U12536 ( .A(n11483), .Z(n11484) );
  OAI21_X1 U12537 ( .B1(n19496), .B2(n19495), .A(n19494), .ZN(n19514) );
  AND2_X1 U12538 ( .A1(n19578), .A2(n19984), .ZN(n19513) );
  OR3_X1 U12539 ( .A1(n19549), .A2(n19792), .A3(n19548), .ZN(n19568) );
  INV_X1 U12540 ( .A(n19591), .ZN(n19595) );
  OAI21_X1 U12541 ( .B1(n19623), .B2(n19603), .A(n19833), .ZN(n19626) );
  AND2_X1 U12542 ( .A1(n19578), .A2(n19838), .ZN(n19624) );
  AND2_X1 U12543 ( .A1(n19668), .A2(n19639), .ZN(n19655) );
  OAI21_X1 U12544 ( .B1(n19676), .B2(n19691), .A(n19833), .ZN(n19694) );
  AND2_X1 U12545 ( .A1(n19640), .A2(n19639), .ZN(n19693) );
  OR2_X1 U12546 ( .A1(n14127), .A2(n14126), .ZN(n19747) );
  INV_X1 U12547 ( .A(n19779), .ZN(n19784) );
  OAI21_X1 U12548 ( .B1(n19800), .B2(n19796), .A(n19795), .ZN(n19824) );
  NOR2_X1 U12549 ( .A1(n19759), .A2(n19758), .ZN(n19821) );
  INV_X1 U12550 ( .A(n19890), .ZN(n19822) );
  INV_X1 U12551 ( .A(n19763), .ZN(n19840) );
  INV_X1 U12552 ( .A(n19809), .ZN(n19865) );
  INV_X1 U12553 ( .A(n19780), .ZN(n19868) );
  INV_X1 U12554 ( .A(n19776), .ZN(n19871) );
  NOR2_X1 U12555 ( .A1(n19789), .A2(n19788), .ZN(n19875) );
  INV_X1 U12556 ( .A(n19819), .ZN(n19874) );
  NAND2_X1 U12557 ( .A1(n17593), .A2(n18792), .ZN(n19026) );
  NOR2_X2 U12558 ( .A1(n18848), .A2(n10579), .ZN(n16718) );
  INV_X1 U12559 ( .A(n10601), .ZN(n16719) );
  INV_X1 U12560 ( .A(n10085), .ZN(n16783) );
  AND2_X1 U12561 ( .A1(n10080), .A2(n16960), .ZN(n16829) );
  AND2_X1 U12562 ( .A1(n10081), .A2(n16960), .ZN(n16838) );
  NOR2_X1 U12563 ( .A1(n18915), .A2(n16916), .ZN(n16897) );
  NOR2_X1 U12564 ( .A1(n17084), .A2(n13154), .ZN(n16931) );
  NOR2_X2 U12565 ( .A1(n19028), .A2(n18850), .ZN(n17067) );
  INV_X1 U12566 ( .A(n17094), .ZN(n17079) );
  NAND4_X1 U12567 ( .A1(n18345), .A2(n19026), .A3(n18866), .A4(n18854), .ZN(
        n17094) );
  INV_X1 U12568 ( .A(n17078), .ZN(n17090) );
  NOR2_X1 U12569 ( .A1(n17192), .A2(n17193), .ZN(n17164) );
  NOR2_X1 U12570 ( .A1(n18402), .A2(n17217), .ZN(n17204) );
  NAND2_X1 U12571 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17311), .ZN(n17295) );
  NOR2_X1 U12572 ( .A1(n17297), .A2(n17322), .ZN(n17311) );
  NAND2_X1 U12573 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17339), .ZN(n17322) );
  NOR2_X2 U12574 ( .A1(n16980), .A2(n17324), .ZN(n17339) );
  NOR2_X2 U12575 ( .A1(n10513), .A2(n10512), .ZN(n17367) );
  NOR2_X1 U12576 ( .A1(n17617), .A2(n17426), .ZN(n17420) );
  NAND2_X1 U12577 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17429), .ZN(n17426) );
  NOR3_X1 U12578 ( .A1(n18402), .A2(n17477), .A3(n17597), .ZN(n17469) );
  INV_X1 U12579 ( .A(n17451), .ZN(n17475) );
  AND2_X1 U12580 ( .A1(n18402), .A2(n17401), .ZN(n17513) );
  INV_X1 U12581 ( .A(n16600), .ZN(n17524) );
  NOR2_X1 U12582 ( .A1(n10423), .A2(n10422), .ZN(n17528) );
  INV_X1 U12583 ( .A(n10611), .ZN(n17531) );
  AOI211_X1 U12584 ( .C1(n9832), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n10386), .B(n10385), .ZN(n10387) );
  INV_X1 U12585 ( .A(n17513), .ZN(n17549) );
  INV_X1 U12586 ( .A(n17539), .ZN(n17547) );
  CLKBUF_X1 U12587 ( .A(n17567), .Z(n17587) );
  CLKBUF_X1 U12588 ( .A(n19011), .Z(n17588) );
  CLKBUF_X1 U12589 ( .A(n17640), .Z(n17658) );
  CLKBUF_X1 U12590 ( .A(n17654), .Z(n17657) );
  NAND2_X1 U12591 ( .A1(n17667), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17663) );
  NAND2_X1 U12592 ( .A1(n9967), .A2(n10326), .ZN(n17730) );
  NAND2_X1 U12593 ( .A1(n17792), .A2(n9974), .ZN(n17778) );
  AOI21_X1 U12594 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17750), .A(
        n18738), .ZN(n17865) );
  NAND2_X1 U12595 ( .A1(n16889), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17803) );
  NOR2_X2 U12596 ( .A1(n17524), .A2(n18035), .ZN(n17926) );
  AND3_X1 U12597 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17978) );
  INV_X1 U12598 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17994) );
  CLKBUF_X1 U12599 ( .A(n18384), .Z(n18738) );
  XNOR2_X1 U12600 ( .A(n10246), .B(n16164), .ZN(n16161) );
  NAND2_X1 U12601 ( .A1(n11449), .A2(n11445), .ZN(n10246) );
  NOR2_X1 U12602 ( .A1(n17680), .A2(n16597), .ZN(n10251) );
  INV_X1 U12603 ( .A(n17681), .ZN(n16599) );
  NAND2_X1 U12604 ( .A1(n19017), .A2(n14414), .ZN(n18804) );
  AOI21_X1 U12605 ( .B1(n14419), .B2(n13116), .A(n18856), .ZN(n18326) );
  NOR2_X1 U12606 ( .A1(n18225), .A2(n18344), .ZN(n18339) );
  INV_X1 U12607 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18368) );
  INV_X1 U12608 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18367) );
  INV_X1 U12609 ( .A(n18992), .ZN(n18995) );
  CLKBUF_X1 U12611 ( .A(n16699), .Z(n16704) );
  NAND2_X1 U12612 ( .A1(n15167), .A2(n20189), .ZN(n15007) );
  AOI21_X1 U12613 ( .B1(n15369), .B2(n15368), .A(n19895), .ZN(n15370) );
  NAND2_X1 U12614 ( .A1(n15577), .A2(n10108), .ZN(n10107) );
  INV_X1 U12615 ( .A(n10104), .ZN(n10110) );
  NOR2_X1 U12616 ( .A1(n15578), .A2(n10109), .ZN(n10108) );
  INV_X1 U12617 ( .A(n11441), .ZN(n11442) );
  NAND2_X1 U12618 ( .A1(n10076), .A2(n10072), .ZN(P3_U2641) );
  NOR2_X1 U12619 ( .A1(n16756), .A2(n10073), .ZN(n10072) );
  NAND2_X1 U12620 ( .A1(n10077), .A2(n17069), .ZN(n10076) );
  NAND2_X1 U12621 ( .A1(n10245), .A2(n10243), .ZN(P3_U2832) );
  NOR3_X1 U12622 ( .A1(n16159), .A2(n10244), .A3(n16160), .ZN(n10243) );
  NAND2_X1 U12623 ( .A1(n16161), .A2(n18250), .ZN(n10245) );
  AOI21_X1 U12624 ( .B1(n16163), .B2(n16162), .A(n16164), .ZN(n10244) );
  AND2_X1 U12625 ( .A1(n9955), .A2(n13827), .ZN(n11064) );
  NAND2_X1 U12626 ( .A1(n12268), .A2(n20243), .ZN(n13993) );
  NAND2_X1 U12628 ( .A1(n10161), .A2(n11034), .ZN(n11044) );
  AND2_X2 U12629 ( .A1(n12047), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10886) );
  AND2_X1 U12630 ( .A1(n10652), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11021) );
  OR3_X1 U12631 ( .A1(n14741), .A2(n10234), .A3(n10231), .ZN(n9963) );
  NAND2_X1 U12632 ( .A1(n14726), .A2(n10008), .ZN(n14701) );
  NAND2_X1 U12633 ( .A1(n11819), .A2(n10268), .ZN(n15478) );
  NAND2_X1 U12634 ( .A1(n11095), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15606) );
  NAND2_X1 U12635 ( .A1(n11095), .A2(n10113), .ZN(n15582) );
  OR2_X1 U12636 ( .A1(n15670), .A2(n15853), .ZN(n9964) );
  AND2_X1 U12637 ( .A1(n15568), .A2(n10023), .ZN(n14282) );
  OR2_X1 U12639 ( .A1(n14228), .A2(n14238), .ZN(n9965) );
  AND2_X1 U12640 ( .A1(n10691), .A2(n10690), .ZN(n9966) );
  AND2_X1 U12641 ( .A1(n17792), .A2(n10013), .ZN(n9967) );
  AND2_X1 U12642 ( .A1(n10222), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9968) );
  XNOR2_X1 U12643 ( .A(n11979), .B(n10331), .ZN(n15449) );
  NOR2_X1 U12644 ( .A1(n17664), .A2(n10030), .ZN(n9969) );
  AND2_X1 U12645 ( .A1(n13868), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9970) );
  AND2_X1 U12646 ( .A1(n11184), .A2(n10009), .ZN(n9971) );
  INV_X1 U12647 ( .A(n11169), .ZN(n14578) );
  AND2_X1 U12648 ( .A1(n15414), .A2(n15475), .ZN(n9972) );
  AND2_X1 U12649 ( .A1(n10219), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9973) );
  AND2_X1 U12650 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9974) );
  AND2_X1 U12651 ( .A1(n10070), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9975) );
  OR2_X1 U12652 ( .A1(n10939), .A2(n10938), .ZN(n11108) );
  AND2_X1 U12653 ( .A1(n14457), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9976) );
  OR2_X1 U12654 ( .A1(n14072), .A2(n10154), .ZN(n13403) );
  AND2_X1 U12655 ( .A1(n10216), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9977) );
  NAND2_X1 U12656 ( .A1(n15136), .A2(n14436), .ZN(n15094) );
  OR2_X1 U12657 ( .A1(n11238), .A2(n11219), .ZN(n9978) );
  AND2_X2 U12658 ( .A1(n12047), .A2(n13827), .ZN(n10929) );
  INV_X2 U12659 ( .A(n11513), .ZN(n13179) );
  NAND2_X1 U12660 ( .A1(n10119), .A2(n11184), .ZN(n15732) );
  NOR2_X1 U12662 ( .A1(n15670), .A2(n10306), .ZN(n15624) );
  AND2_X1 U12663 ( .A1(n14815), .A2(n10286), .ZN(n14852) );
  NOR2_X1 U12664 ( .A1(n15606), .A2(n15793), .ZN(n15591) );
  NAND2_X1 U12665 ( .A1(n15630), .A2(n15629), .ZN(n15631) );
  NOR2_X1 U12666 ( .A1(n18870), .A2(n18021), .ZN(n17750) );
  AND2_X1 U12667 ( .A1(n13827), .A2(n10652), .ZN(n9980) );
  AND2_X1 U12668 ( .A1(n15717), .A2(n15913), .ZN(n9981) );
  AND4_X1 U12669 ( .A1(n12202), .A2(n12201), .A3(n12200), .A4(n12199), .ZN(
        n9982) );
  AND2_X1 U12670 ( .A1(n9824), .A2(n10307), .ZN(n9983) );
  OR2_X1 U12671 ( .A1(n11179), .A2(n11160), .ZN(n9984) );
  OR2_X1 U12672 ( .A1(n12232), .A2(n12143), .ZN(n9985) );
  OAI21_X1 U12673 ( .B1(n9925), .B2(n10300), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12280) );
  AND4_X1 U12674 ( .A1(n10681), .A2(n10680), .A3(n10679), .A4(n10678), .ZN(
        n9986) );
  AND3_X1 U12675 ( .A1(n10689), .A2(n13827), .A3(n10688), .ZN(n9987) );
  AND2_X1 U12676 ( .A1(n11044), .A2(n10160), .ZN(n11178) );
  OR2_X1 U12677 ( .A1(n15615), .A2(n10133), .ZN(n9988) );
  NAND2_X1 U12678 ( .A1(n15631), .A2(n11274), .ZN(n15614) );
  NAND2_X1 U12679 ( .A1(n14405), .A2(n14404), .ZN(n14433) );
  AND2_X2 U12680 ( .A1(n9931), .A2(n13827), .ZN(n11558) );
  AND2_X1 U12681 ( .A1(n16296), .A2(n20185), .ZN(n9989) );
  AND2_X1 U12682 ( .A1(n11777), .A2(n13414), .ZN(n9990) );
  NAND2_X1 U12683 ( .A1(n11781), .A2(n11780), .ZN(n11782) );
  NOR2_X1 U12684 ( .A1(n11161), .A2(n10191), .ZN(n9991) );
  NAND2_X1 U12685 ( .A1(n15152), .A2(n13868), .ZN(n14338) );
  INV_X1 U12686 ( .A(n10200), .ZN(n16418) );
  NAND2_X1 U12687 ( .A1(n10201), .A2(n11283), .ZN(n10200) );
  NOR2_X1 U12688 ( .A1(n15459), .A2(n15458), .ZN(n13223) );
  INV_X1 U12689 ( .A(n14228), .ZN(n10229) );
  OR2_X1 U12690 ( .A1(n15511), .A2(n10152), .ZN(n9992) );
  AND2_X1 U12691 ( .A1(n10643), .A2(n10642), .ZN(n9993) );
  AND2_X1 U12692 ( .A1(n12336), .A2(n10040), .ZN(n9994) );
  INV_X1 U12693 ( .A(n17540), .ZN(n10439) );
  INV_X1 U12694 ( .A(n15612), .ZN(n11095) );
  AND3_X1 U12695 ( .A1(n10717), .A2(n10718), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9995) );
  AND3_X1 U12696 ( .A1(n10712), .A2(n10713), .A3(n13827), .ZN(n9996) );
  BUF_X1 U12697 ( .A(n10762), .Z(n11505) );
  NAND2_X1 U12698 ( .A1(n16338), .A2(n14544), .ZN(n9997) );
  INV_X1 U12699 ( .A(n13472), .ZN(n14262) );
  AND2_X1 U12700 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9998) );
  AND2_X1 U12701 ( .A1(n14450), .A2(n14449), .ZN(n9999) );
  INV_X1 U12702 ( .A(n10832), .ZN(n10087) );
  AND2_X1 U12703 ( .A1(n14355), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10000) );
  AND2_X1 U12704 ( .A1(n12268), .A2(n12241), .ZN(n14375) );
  NAND2_X1 U12705 ( .A1(n13223), .A2(n13224), .ZN(n13222) );
  OR2_X1 U12706 ( .A1(n12232), .A2(n12904), .ZN(n10001) );
  AND2_X2 U12707 ( .A1(n9818), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11069) );
  AND2_X1 U12708 ( .A1(n10683), .A2(n10096), .ZN(n10002) );
  INV_X1 U12709 ( .A(n17535), .ZN(n10614) );
  NOR2_X1 U12710 ( .A1(n10412), .A2(n10411), .ZN(n17535) );
  NAND2_X1 U12711 ( .A1(n14453), .A2(n16276), .ZN(n15057) );
  OR2_X1 U12712 ( .A1(n11276), .A2(n11275), .ZN(n10003) );
  AND2_X1 U12713 ( .A1(n11470), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10004) );
  AND2_X1 U12714 ( .A1(n10085), .A2(n10084), .ZN(n10005) );
  INV_X1 U12715 ( .A(n12260), .ZN(n10295) );
  INV_X1 U12717 ( .A(n13179), .ZN(n19356) );
  OAI22_X1 U12718 ( .A1(n14608), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19032), 
        .B2(n14588), .ZN(n13205) );
  INV_X1 U12719 ( .A(n12640), .ZN(n10283) );
  NAND2_X1 U12720 ( .A1(n11819), .A2(n11818), .ZN(n14039) );
  OR2_X1 U12721 ( .A1(n13632), .A2(n13198), .ZN(n10006) );
  AND2_X1 U12722 ( .A1(n13191), .A2(n14061), .ZN(n14060) );
  AND2_X1 U12723 ( .A1(n11819), .A2(n10269), .ZN(n14279) );
  NOR2_X1 U12724 ( .A1(n13217), .A2(n15663), .ZN(n13208) );
  NOR2_X1 U12725 ( .A1(n13214), .A2(n16445), .ZN(n13213) );
  NOR2_X1 U12726 ( .A1(n13727), .A2(n13713), .ZN(n13712) );
  NOR2_X1 U12727 ( .A1(n13171), .A2(n16485), .ZN(n13165) );
  NOR2_X1 U12728 ( .A1(n13166), .A2(n16494), .ZN(n13167) );
  AND2_X1 U12729 ( .A1(n13165), .A2(n10221), .ZN(n13163) );
  AND2_X1 U12730 ( .A1(n13213), .A2(n10219), .ZN(n13212) );
  AND3_X1 U12731 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10214), .A3(
        n10211), .ZN(n10007) );
  AND2_X1 U12732 ( .A1(n14711), .A2(n14728), .ZN(n10008) );
  AND2_X1 U12733 ( .A1(n15735), .A2(n15968), .ZN(n10009) );
  OR2_X1 U12734 ( .A1(n10338), .A2(n14872), .ZN(n10010) );
  OR2_X1 U12735 ( .A1(n14772), .A2(n14775), .ZN(n10011) );
  NOR2_X1 U12736 ( .A1(n14877), .A2(n10236), .ZN(n14773) );
  AND2_X1 U12737 ( .A1(n13165), .A2(n10222), .ZN(n13164) );
  INV_X1 U12738 ( .A(n15721), .ZN(n10275) );
  INV_X1 U12739 ( .A(n14436), .ZN(n10049) );
  NAND2_X1 U12740 ( .A1(n10050), .A2(n10301), .ZN(n16290) );
  NAND2_X1 U12741 ( .A1(n10051), .A2(n14365), .ZN(n16284) );
  AND2_X1 U12742 ( .A1(n15413), .A2(n15414), .ZN(n15412) );
  AOI21_X1 U12743 ( .B1(n10838), .B2(n11791), .A(n11790), .ZN(n13469) );
  AND2_X1 U12744 ( .A1(n14043), .A2(n14044), .ZN(n14042) );
  AND2_X1 U12745 ( .A1(n13190), .A2(n13189), .ZN(n13191) );
  AND2_X1 U12746 ( .A1(n16276), .A2(n15003), .ZN(n10012) );
  NAND2_X1 U12747 ( .A1(n14389), .A2(n14388), .ZN(n14330) );
  AND2_X1 U12748 ( .A1(n9974), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10013) );
  INV_X2 U12749 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20932) );
  OR2_X1 U12750 ( .A1(n10154), .A2(n13436), .ZN(n10014) );
  NOR2_X1 U12751 ( .A1(n14741), .A2(n10233), .ZN(n14697) );
  NOR2_X1 U12752 ( .A1(n15644), .A2(n10163), .ZN(n10015) );
  AND2_X1 U12753 ( .A1(n10268), .A2(n10267), .ZN(n10016) );
  AND2_X1 U12754 ( .A1(n10270), .A2(n13733), .ZN(n10017) );
  INV_X1 U12755 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10213) );
  AND2_X1 U12756 ( .A1(n11134), .A2(n19356), .ZN(n16503) );
  INV_X1 U12757 ( .A(n16503), .ZN(n19332) );
  INV_X1 U12758 ( .A(n14224), .ZN(n14214) );
  NAND2_X1 U12759 ( .A1(n13617), .A2(n11801), .ZN(n13716) );
  NOR2_X1 U12760 ( .A1(n13727), .A2(n10168), .ZN(n13734) );
  NOR2_X1 U12761 ( .A1(n13727), .A2(n10170), .ZN(n10018) );
  NOR2_X1 U12762 ( .A1(n13700), .A2(n13701), .ZN(n13702) );
  NOR2_X1 U12763 ( .A1(n20527), .A2(n20247), .ZN(n10019) );
  AND2_X1 U12764 ( .A1(n17667), .A2(n10070), .ZN(n10020) );
  NOR2_X1 U12765 ( .A1(n14072), .A2(n14071), .ZN(n13402) );
  AND2_X1 U12766 ( .A1(n13213), .A2(n10218), .ZN(n13210) );
  NAND3_X1 U12767 ( .A1(n16937), .A2(n10327), .A3(n10069), .ZN(n10021) );
  INV_X1 U12768 ( .A(n17047), .ZN(n10084) );
  AND2_X1 U12769 ( .A1(n13208), .A2(n10202), .ZN(n10022) );
  AND2_X1 U12770 ( .A1(n11753), .A2(n11697), .ZN(n16558) );
  INV_X1 U12771 ( .A(n16558), .ZN(n16544) );
  AND2_X1 U12772 ( .A1(n10145), .A2(n14201), .ZN(n10023) );
  AND2_X1 U12773 ( .A1(n14819), .A2(n14802), .ZN(n14801) );
  NOR2_X1 U12774 ( .A1(n13207), .A2(n15608), .ZN(n13206) );
  OR2_X1 U12775 ( .A1(n16394), .A2(n16403), .ZN(n10024) );
  OR2_X1 U12776 ( .A1(n16424), .A2(n15382), .ZN(n10025) );
  AND2_X1 U12777 ( .A1(n13435), .A2(n13499), .ZN(n13498) );
  AND2_X1 U12778 ( .A1(n10023), .A2(n14284), .ZN(n10026) );
  INV_X1 U12779 ( .A(n10197), .ZN(n10196) );
  NAND2_X1 U12780 ( .A1(n11248), .A2(n15491), .ZN(n10197) );
  AND2_X1 U12781 ( .A1(n10202), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10027) );
  AND2_X1 U12782 ( .A1(n13617), .A2(n10270), .ZN(n10028) );
  XNOR2_X1 U12783 ( .A(n13949), .B(n13951), .ZN(n13948) );
  AND2_X1 U12784 ( .A1(n14575), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10029) );
  AND2_X2 U12785 ( .A1(n13537), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13536) );
  NAND2_X1 U12786 ( .A1(n14170), .A2(n14167), .ZN(n14229) );
  INV_X1 U12787 ( .A(n14229), .ZN(n10226) );
  OR2_X1 U12788 ( .A1(n16601), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10030) );
  NOR3_X2 U12789 ( .A1(n18860), .A2(n18636), .A3(n18496), .ZN(n10031) );
  INV_X1 U12790 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10071) );
  INV_X1 U12791 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10204) );
  AND2_X1 U12792 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10032) );
  INV_X1 U12793 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10173) );
  INV_X1 U12794 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10174) );
  INV_X1 U12795 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10220) );
  INV_X1 U12796 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10203) );
  INV_X1 U12797 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10215) );
  INV_X1 U12798 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10223) );
  INV_X1 U12799 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n10190) );
  NAND2_X2 U12800 ( .A1(n19027), .A2(n18859), .ZN(n18345) );
  OAI21_X2 U12801 ( .B1(n15988), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11432), 
        .ZN(n19833) );
  AOI22_X2 U12802 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19389), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19388), .ZN(n19879) );
  NOR3_X2 U12803 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18860), .A3(
        n18588), .ZN(n18558) );
  INV_X1 U12804 ( .A(n10311), .ZN(n10114) );
  NAND2_X1 U12805 ( .A1(n10310), .A2(n10311), .ZN(n10309) );
  AOI22_X2 U12806 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19389), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19388), .ZN(n19827) );
  NOR2_X2 U12807 ( .A1(n14135), .A2(n14136), .ZN(n19388) );
  NOR3_X2 U12808 ( .A1(n18860), .A2(n18660), .A3(n18635), .ZN(n18628) );
  NOR2_X2 U12809 ( .A1(n14137), .A2(n14136), .ZN(n19389) );
  OAI21_X4 U12810 ( .B1(n12076), .B2(n12075), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14137) );
  NOR2_X1 U12811 ( .A1(n19373), .A2(n19390), .ZN(n10033) );
  NAND2_X2 U12812 ( .A1(n10035), .A2(n10034), .ZN(n13562) );
  NAND2_X2 U12813 ( .A1(n10047), .A2(n14447), .ZN(n15089) );
  NAND2_X1 U12814 ( .A1(n16290), .A2(n14364), .ZN(n10051) );
  NAND2_X1 U12815 ( .A1(n9989), .A2(n20183), .ZN(n10050) );
  NAND2_X2 U12816 ( .A1(n15010), .A2(n15057), .ZN(n15051) );
  NAND2_X2 U12817 ( .A1(n14454), .A2(n15140), .ZN(n15058) );
  NOR2_X2 U12818 ( .A1(n15206), .A2(n14535), .ZN(n15197) );
  INV_X2 U12819 ( .A(n20222), .ZN(n10057) );
  INV_X2 U12820 ( .A(n20243), .ZN(n13751) );
  NOR2_X2 U12821 ( .A1(n10059), .A2(n12239), .ZN(n12252) );
  INV_X1 U12822 ( .A(n12239), .ZN(n13604) );
  NAND2_X1 U12823 ( .A1(n16284), .A2(n16286), .ZN(n10060) );
  NAND2_X1 U12824 ( .A1(n9925), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12272) );
  NAND2_X1 U12825 ( .A1(n14989), .A2(n10065), .ZN(n14990) );
  NAND2_X1 U12826 ( .A1(n15104), .A2(n14437), .ZN(n15120) );
  NAND2_X1 U12827 ( .A1(n9936), .A2(n15140), .ZN(n15030) );
  NAND3_X1 U12828 ( .A1(n12414), .A2(n13920), .A3(n12450), .ZN(n12475) );
  NAND3_X1 U12829 ( .A1(n16758), .A2(n10075), .A3(n10074), .ZN(n10073) );
  INV_X1 U12830 ( .A(n10081), .ZN(n16847) );
  INV_X1 U12831 ( .A(n10080), .ZN(n16837) );
  NAND3_X1 U12832 ( .A1(n10087), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A3(
        n13472), .ZN(n10830) );
  NAND3_X1 U12833 ( .A1(n10087), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A3(
        n13472), .ZN(n10898) );
  NAND2_X1 U12834 ( .A1(n14291), .A2(n11043), .ZN(n10091) );
  OAI211_X1 U12835 ( .C1(n14291), .C2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10090), .B(n10088), .ZN(n15970) );
  NAND2_X1 U12836 ( .A1(n10089), .A2(n16543), .ZN(n10088) );
  NAND3_X1 U12837 ( .A1(n14291), .A2(n11043), .A3(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U12838 ( .A1(n10091), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11087) );
  NAND2_X1 U12839 ( .A1(n9953), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10092) );
  INV_X1 U12840 ( .A(n10686), .ZN(n10094) );
  NAND2_X1 U12841 ( .A1(n10092), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10099) );
  OAI21_X2 U12842 ( .B1(n10097), .B2(n10094), .A(n10093), .ZN(n10721) );
  NAND4_X1 U12843 ( .A1(n10095), .A2(n10682), .A3(n10002), .A4(n10684), .ZN(
        n10093) );
  AOI21_X1 U12844 ( .B1(n9953), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10096) );
  NAND3_X1 U12845 ( .A1(n10687), .A2(n10685), .A3(n10098), .ZN(n10097) );
  OAI211_X1 U12846 ( .C1(n15754), .C2(n19333), .A(n10110), .B(n10107), .ZN(
        P2_U2985) );
  AND2_X1 U12847 ( .A1(n10118), .A2(n10978), .ZN(n10116) );
  NOR2_X1 U12848 ( .A1(n10926), .A2(n11547), .ZN(n10118) );
  NAND2_X1 U12849 ( .A1(n10957), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10899) );
  NAND4_X1 U12850 ( .A1(n10670), .A2(n10672), .A3(n10673), .A4(n10671), .ZN(
        n10120) );
  NAND4_X1 U12851 ( .A1(n19361), .A2(n19373), .A3(n13364), .A4(n10723), .ZN(
        n10745) );
  NAND4_X1 U12852 ( .A1(n10676), .A2(n10677), .A3(n10675), .A4(n10123), .ZN(
        n10122) );
  NAND2_X1 U12853 ( .A1(n9953), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10125) );
  NAND3_X1 U12854 ( .A1(n10666), .A2(n10668), .A3(n10669), .ZN(n10128) );
  NAND3_X1 U12855 ( .A1(n9923), .A2(n10974), .A3(n11169), .ZN(n10134) );
  OAI21_X1 U12856 ( .B1(n14192), .B2(n10142), .A(n10140), .ZN(n13322) );
  NOR2_X2 U12857 ( .A1(n14283), .A2(n15417), .ZN(n15541) );
  NAND3_X1 U12858 ( .A1(n9995), .A2(n10719), .A3(n10720), .ZN(n10146) );
  NAND3_X1 U12859 ( .A1(n9996), .A2(n10714), .A3(n10715), .ZN(n10147) );
  NOR3_X4 U12860 ( .A1(n15511), .A2(n10152), .A3(n15497), .ZN(n15496) );
  AND2_X2 U12861 ( .A1(n13783), .A2(n13802), .ZN(n10716) );
  NAND3_X1 U12862 ( .A1(n11044), .A2(n10158), .A3(n10159), .ZN(n11182) );
  OAI21_X1 U12863 ( .B1(n13364), .B2(n19373), .A(n10162), .ZN(n10741) );
  NAND2_X1 U12864 ( .A1(n15643), .A2(n10015), .ZN(n16439) );
  XNOR2_X1 U12865 ( .A(n10164), .B(n15912), .ZN(n16446) );
  OAI21_X2 U12866 ( .B1(n15711), .B2(n15648), .A(n15650), .ZN(n15700) );
  NOR2_X2 U12867 ( .A1(n17666), .A2(n17665), .ZN(n17664) );
  INV_X1 U12868 ( .A(n10180), .ZN(n15427) );
  OR2_X2 U12869 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18826) );
  INV_X2 U12870 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18986) );
  INV_X2 U12871 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18979) );
  NAND2_X1 U12872 ( .A1(n11202), .A2(n10189), .ZN(n11213) );
  NOR2_X2 U12873 ( .A1(n11161), .A2(n10192), .ZN(n11197) );
  NAND2_X1 U12874 ( .A1(n13208), .A2(n10027), .ZN(n13207) );
  NAND4_X1 U12875 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10214), .A3(
        n10212), .A4(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13166) );
  NAND3_X1 U12876 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10214), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13169) );
  NAND2_X1 U12877 ( .A1(n13763), .A2(n10230), .ZN(n13951) );
  NAND3_X1 U12878 ( .A1(n12246), .A2(n14467), .A3(n21099), .ZN(n10230) );
  NOR2_X2 U12879 ( .A1(n14630), .A2(n14517), .ZN(n14500) );
  NOR2_X2 U12880 ( .A1(n10252), .A2(n18969), .ZN(n10356) );
  NAND3_X1 U12881 ( .A1(n18979), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n18994), .ZN(n10252) );
  NAND3_X1 U12882 ( .A1(n10253), .A2(n10254), .A3(n10004), .ZN(n15588) );
  INV_X1 U12883 ( .A(n11469), .ZN(n10253) );
  NAND2_X1 U12884 ( .A1(n15431), .A2(n10256), .ZN(n10255) );
  OAI211_X1 U12885 ( .C1(n15431), .C2(n10260), .A(n10258), .B(n10255), .ZN(
        n14621) );
  NAND2_X1 U12886 ( .A1(n15431), .A2(n15430), .ZN(n15432) );
  OAI21_X1 U12887 ( .B1(n14621), .B2(n15493), .A(n14620), .ZN(P2_U2857) );
  NOR2_X2 U12888 ( .A1(n15464), .A2(n11934), .ZN(n11958) );
  NAND2_X1 U12889 ( .A1(n10261), .A2(n10262), .ZN(n15464) );
  NAND2_X1 U12890 ( .A1(n10323), .A2(n10265), .ZN(n10262) );
  AND2_X2 U12891 ( .A1(n11819), .A2(n10016), .ZN(n11911) );
  NOR2_X1 U12892 ( .A1(n15601), .A2(n15602), .ZN(n15592) );
  NAND2_X1 U12893 ( .A1(n13617), .A2(n10017), .ZN(n13731) );
  NOR2_X1 U12894 ( .A1(n15659), .A2(n10275), .ZN(n10273) );
  NAND2_X1 U12895 ( .A1(n13773), .A2(n10276), .ZN(n15148) );
  NAND2_X1 U12896 ( .A1(n12386), .A2(n12385), .ZN(n10276) );
  AND2_X1 U12897 ( .A1(n14726), .A2(n14728), .ZN(n14710) );
  OAI21_X1 U12898 ( .B1(n13914), .B2(n10284), .A(n10281), .ZN(n13772) );
  XNOR2_X2 U12899 ( .A(n12389), .B(n12388), .ZN(n13914) );
  NAND2_X1 U12900 ( .A1(n14670), .A2(n14672), .ZN(n14658) );
  NAND3_X1 U12901 ( .A1(n12256), .A2(n12255), .A3(n12267), .ZN(n10300) );
  NAND4_X1 U12902 ( .A1(n12256), .A2(n12255), .A3(n12267), .A4(n12260), .ZN(
        n10293) );
  NAND2_X1 U12903 ( .A1(n12258), .A2(n10297), .ZN(n10296) );
  INV_X1 U12904 ( .A(n12266), .ZN(n10299) );
  XNOR2_X2 U12905 ( .A(n12307), .B(n10298), .ZN(n12378) );
  NAND2_X1 U12906 ( .A1(n20183), .A2(n20185), .ZN(n20184) );
  NAND2_X1 U12907 ( .A1(n15022), .A2(n9919), .ZN(n15014) );
  NAND3_X1 U12908 ( .A1(n15022), .A2(n14455), .A3(n14456), .ZN(n14989) );
  NOR2_X2 U12909 ( .A1(n14989), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14553) );
  NAND3_X1 U12910 ( .A1(n15057), .A2(n9936), .A3(n15221), .ZN(n15031) );
  AND3_X4 U12911 ( .A1(n14250), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10652) );
  AND2_X2 U12912 ( .A1(n11095), .A2(n10308), .ZN(n15578) );
  OAI21_X1 U12913 ( .B1(n14572), .B2(n14571), .A(n10340), .ZN(n14581) );
  NAND2_X1 U12914 ( .A1(n20297), .A2(n12364), .ZN(n13748) );
  NAND2_X1 U12915 ( .A1(n10001), .A2(n12166), .ZN(n12170) );
  AND2_X1 U12916 ( .A1(n12003), .A2(n12002), .ZN(n12004) );
  AOI211_X1 U12917 ( .C1(n19224), .C2(n19223), .A(n19222), .B(n19221), .ZN(
        n19232) );
  NAND2_X1 U12918 ( .A1(n19224), .A2(n11791), .ZN(n11781) );
  AOI22_X1 U12919 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12348), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12215) );
  INV_X1 U12920 ( .A(n10776), .ZN(n10782) );
  CLKBUF_X1 U12921 ( .A(n13535), .Z(n20655) );
  NAND2_X1 U12922 ( .A1(n10663), .A2(n13827), .ZN(n10664) );
  NAND2_X1 U12923 ( .A1(n15973), .A2(n11087), .ZN(n15728) );
  NAND2_X1 U12924 ( .A1(n11037), .A2(n11036), .ZN(n11038) );
  AND4_X1 U12925 ( .A1(n10847), .A2(n10846), .A3(n10845), .A4(n10844), .ZN(
        n10859) );
  AND2_X1 U12926 ( .A1(n10692), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10696) );
  AND2_X1 U12927 ( .A1(n12243), .A2(n13587), .ZN(n12240) );
  INV_X1 U12928 ( .A(n14649), .ZN(n14847) );
  XNOR2_X1 U12929 ( .A(n14460), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14618) );
  NAND2_X1 U12930 ( .A1(n14459), .A2(n14458), .ZN(n14460) );
  OAI21_X1 U12931 ( .B1(n12284), .B2(n12283), .A(n12391), .ZN(n13535) );
  NOR2_X1 U12932 ( .A1(n19373), .A2(n19390), .ZN(n19860) );
  MUX2_X1 U12933 ( .A(n12066), .B(n11490), .S(n19373), .Z(n10753) );
  INV_X1 U12934 ( .A(n12388), .ZN(n12390) );
  AND3_X1 U12935 ( .A1(n18994), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n17063), .ZN(n10312) );
  AND3_X1 U12936 ( .A1(n20658), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10313) );
  INV_X1 U12937 ( .A(n14897), .ZN(n14905) );
  OR2_X1 U12938 ( .A1(n14583), .A2(n14597), .ZN(n10314) );
  INV_X1 U12939 ( .A(n16552), .ZN(n16563) );
  OR2_X1 U12940 ( .A1(n18036), .A2(n13134), .ZN(n10315) );
  AND2_X1 U12941 ( .A1(n10863), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11020) );
  INV_X1 U12942 ( .A(n11741), .ZN(n11092) );
  AND2_X1 U12943 ( .A1(n9940), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10316) );
  AND2_X1 U12944 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10317) );
  INV_X1 U12945 ( .A(n11290), .ZN(n11284) );
  AND4_X1 U12946 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n10318) );
  AND4_X1 U12947 ( .A1(n11009), .A2(n11008), .A3(n11007), .A4(n11006), .ZN(
        n10319) );
  AND4_X1 U12948 ( .A1(n10955), .A2(n10954), .A3(n10953), .A4(n10952), .ZN(
        n10320) );
  AND4_X1 U12949 ( .A1(n10961), .A2(n10960), .A3(n10959), .A4(n10958), .ZN(
        n10321) );
  AND2_X1 U12950 ( .A1(n16384), .A2(n16383), .ZN(n10322) );
  AND2_X1 U12951 ( .A1(n13848), .A2(n13332), .ZN(n10324) );
  OR2_X1 U12952 ( .A1(n10634), .A2(n13128), .ZN(n10325) );
  AND2_X1 U12953 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10326) );
  AND3_X1 U12954 ( .A1(n17894), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10327) );
  NOR2_X2 U12955 ( .A1(n9978), .A2(n11222), .ZN(n11223) );
  AND4_X1 U12956 ( .A1(n11014), .A2(n11013), .A3(n11012), .A4(n11011), .ZN(
        n10328) );
  OR2_X1 U12957 ( .A1(n17932), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10329) );
  INV_X1 U12958 ( .A(n11959), .ZN(n11955) );
  AND2_X1 U12959 ( .A1(n11978), .A2(n12000), .ZN(n10331) );
  INV_X1 U12960 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11094) );
  AND3_X1 U12961 ( .A1(n11465), .A2(n11464), .A3(n10315), .ZN(n10332) );
  AND3_X1 U12962 ( .A1(n10636), .A2(n10635), .A3(n10325), .ZN(n10333) );
  OR2_X1 U12963 ( .A1(n15410), .A2(n15665), .ZN(n10334) );
  AND3_X1 U12964 ( .A1(n10779), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10778), 
        .ZN(n10335) );
  OR3_X1 U12965 ( .A1(n15770), .A2(n15744), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10336) );
  INV_X1 U12966 ( .A(n12294), .ZN(n12797) );
  AND3_X1 U12967 ( .A1(n10640), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10639), .ZN(n10337) );
  NAND2_X1 U12968 ( .A1(n10463), .A2(n10462), .ZN(n10466) );
  OR2_X1 U12969 ( .A1(n12719), .A2(n14767), .ZN(n10338) );
  NAND2_X1 U12970 ( .A1(n16405), .A2(n11293), .ZN(n10339) );
  AND2_X1 U12971 ( .A1(n14570), .A2(n15574), .ZN(n10340) );
  INV_X1 U12972 ( .A(n12702), .ZN(n12907) );
  INV_X1 U12973 ( .A(n12293), .ZN(n12434) );
  INV_X1 U12974 ( .A(n19488), .ZN(n11003) );
  INV_X1 U12975 ( .A(n13034), .ZN(n13037) );
  NOR2_X1 U12976 ( .A1(n13037), .A2(n13071), .ZN(n13048) );
  OR2_X1 U12977 ( .A1(n12261), .A2(n14378), .ZN(n12264) );
  NOR2_X1 U12978 ( .A1(n11036), .A2(n11165), .ZN(n11034) );
  NAND2_X1 U12979 ( .A1(n12066), .A2(n10723), .ZN(n10724) );
  AND2_X1 U12980 ( .A1(n10456), .A2(n10455), .ZN(n10457) );
  OR2_X1 U12981 ( .A1(n12463), .A2(n12462), .ZN(n14359) );
  OR2_X1 U12982 ( .A1(n12300), .A2(n12299), .ZN(n12302) );
  OR2_X1 U12983 ( .A1(n12440), .A2(n12439), .ZN(n14348) );
  OR2_X1 U12984 ( .A1(n12354), .A2(n12353), .ZN(n13692) );
  NAND2_X1 U12985 ( .A1(n11960), .A2(n11955), .ZN(n11961) );
  AOI22_X1 U12986 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10639) );
  OR2_X1 U12987 ( .A1(n12491), .A2(n12490), .ZN(n14368) );
  OR2_X1 U12988 ( .A1(n12988), .A2(n12147), .ZN(n12151) );
  AOI22_X1 U12989 ( .A1(n9931), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10716), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10703) );
  AND2_X1 U12990 ( .A1(n16405), .A2(n14578), .ZN(n11290) );
  AOI22_X1 U12991 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19350), .B1(
        n19488), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10911) );
  AND2_X1 U12992 ( .A1(n11126), .A2(n11097), .ZN(n11105) );
  OR2_X1 U12993 ( .A1(n17963), .A2(n18284), .ZN(n10451) );
  INV_X1 U12994 ( .A(n14207), .ZN(n12526) );
  AOI22_X1 U12995 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12348), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12234) );
  OR2_X1 U12996 ( .A1(n12321), .A2(n12320), .ZN(n14374) );
  OR2_X1 U12997 ( .A1(n11407), .A2(n11101), .ZN(n11126) );
  INV_X1 U12998 ( .A(n11933), .ZN(n11910) );
  INV_X1 U12999 ( .A(n15386), .ZN(n11381) );
  INV_X1 U13000 ( .A(n10925), .ZN(n10926) );
  OAI21_X1 U13001 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18979), .A(
        n10472), .ZN(n10473) );
  NOR2_X1 U13002 ( .A1(n17367), .A2(n18366), .ZN(n10577) );
  NOR2_X1 U13003 ( .A1(n18826), .A2(n10344), .ZN(n10548) );
  AND2_X1 U13004 ( .A1(n13059), .A2(n14375), .ZN(n13055) );
  NOR2_X1 U13005 ( .A1(n12843), .A2(n15044), .ZN(n12844) );
  INV_X1 U13006 ( .A(n14500), .ZN(n14514) );
  AND3_X1 U13007 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A3(n12623), .ZN(n12626) );
  INV_X1 U13008 ( .A(n12522), .ZN(n12527) );
  AND2_X1 U13009 ( .A1(n20929), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14428) );
  INV_X1 U13010 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13020) );
  INV_X1 U13011 ( .A(n20691), .ZN(n20778) );
  NAND2_X1 U13012 ( .A1(n15352), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13176) );
  OR2_X1 U13013 ( .A1(n14598), .A2(n14606), .ZN(n14599) );
  AND2_X1 U13014 ( .A1(n11088), .A2(n11086), .ZN(n15972) );
  AND2_X1 U13015 ( .A1(n19988), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19574) );
  AOI21_X1 U13016 ( .B1(n18636), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10471), .ZN(n10477) );
  INV_X1 U13017 ( .A(n11450), .ZN(n11451) );
  NAND2_X1 U13018 ( .A1(n10587), .A2(n10586), .ZN(n13151) );
  NOR2_X1 U13019 ( .A1(n12739), .A2(n16192), .ZN(n12740) );
  NOR2_X1 U13020 ( .A1(n12696), .A2(n12697), .ZN(n12679) );
  INV_X1 U13021 ( .A(n16242), .ZN(n16246) );
  INV_X1 U13022 ( .A(n20133), .ZN(n20115) );
  INV_X1 U13023 ( .A(n14719), .ZN(n20112) );
  AND2_X1 U13024 ( .A1(n13761), .A2(n13757), .ZN(n14839) );
  INV_X1 U13025 ( .A(n13958), .ZN(n13957) );
  OR2_X1 U13026 ( .A1(n12718), .A2(n14768), .ZN(n14767) );
  NAND2_X1 U13027 ( .A1(n12659), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12739) );
  NAND2_X1 U13028 ( .A1(n12721), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12696) );
  NOR2_X1 U13029 ( .A1(n12556), .A2(n20073), .ZN(n12560) );
  AND3_X1 U13030 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(n12466), .ZN(n12492) );
  OR3_X1 U13031 ( .A1(n15211), .A2(n15190), .A3(n14546), .ZN(n15172) );
  OAI21_X1 U13032 ( .B1(n15292), .B2(n15293), .A(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16303) );
  INV_X1 U13033 ( .A(n20221), .ZN(n20196) );
  NOR2_X1 U13034 ( .A1(n20664), .A2(n14625), .ZN(n13550) );
  AND2_X1 U13035 ( .A1(n13921), .A2(n20790), .ZN(n20787) );
  INV_X1 U13036 ( .A(n13562), .ZN(n20240) );
  AND2_X1 U13037 ( .A1(n20722), .A2(n20292), .ZN(n20589) );
  INV_X1 U13038 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20658) );
  NOR2_X1 U13039 ( .A1(n20584), .A2(n20406), .ZN(n20730) );
  AOI21_X1 U13040 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20690), .A(n20406), 
        .ZN(n20789) );
  NAND2_X1 U13041 ( .A1(n13205), .A2(n10334), .ZN(n16102) );
  NAND2_X1 U13042 ( .A1(n9991), .A2(n11508), .ZN(n11283) );
  NAND2_X1 U13043 ( .A1(n11155), .A2(n11154), .ZN(n11161) );
  INV_X1 U13044 ( .A(n11505), .ZN(n20026) );
  AND2_X1 U13045 ( .A1(n11557), .A2(n11556), .ZN(n14071) );
  OR2_X1 U13046 ( .A1(n19998), .A2(n19986), .ZN(n19758) );
  NAND2_X1 U13047 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19833), .ZN(n19390) );
  INV_X1 U13048 ( .A(n18225), .ZN(n18790) );
  INV_X1 U13049 ( .A(n16750), .ZN(n16751) );
  OAI21_X1 U13050 ( .B1(n16855), .B2(n17047), .A(n16891), .ZN(n16848) );
  INV_X1 U13051 ( .A(n17067), .ZN(n17084) );
  NOR2_X1 U13052 ( .A1(n10400), .A2(n10399), .ZN(n10607) );
  AOI21_X1 U13053 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n11448), .A(
        n11447), .ZN(n11456) );
  NOR2_X1 U13054 ( .A1(n10632), .A2(n17933), .ZN(n17854) );
  INV_X1 U13055 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18636) );
  NOR2_X1 U13056 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18365), .ZN(n18662) );
  NAND2_X1 U13057 ( .A1(n12740), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12785) );
  AND2_X1 U13058 ( .A1(n14839), .A2(n14777), .ZN(n16242) );
  INV_X1 U13059 ( .A(n14809), .ZN(n20106) );
  AND2_X1 U13060 ( .A1(n14831), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20133) );
  OR2_X1 U13061 ( .A1(n14623), .A2(n16153), .ZN(n13992) );
  INV_X1 U13062 ( .A(n14948), .ZN(n14967) );
  AND2_X1 U13063 ( .A1(n13421), .A2(n13420), .ZN(n20144) );
  OR2_X1 U13064 ( .A1(n14886), .A2(n14872), .ZN(n14874) );
  NAND2_X1 U13065 ( .A1(n12561), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12590) );
  AND2_X1 U13066 ( .A1(n12492), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12505) );
  INV_X1 U13067 ( .A(n20193), .ZN(n16270) );
  INV_X1 U13068 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14554) );
  NOR2_X1 U13069 ( .A1(n15239), .A2(n14451), .ZN(n15236) );
  NAND2_X1 U13070 ( .A1(n16334), .A2(n20196), .ZN(n16338) );
  AND2_X1 U13071 ( .A1(n13612), .A2(n13593), .ZN(n20215) );
  INV_X1 U13072 ( .A(n13550), .ZN(n20914) );
  INV_X1 U13073 ( .A(n20308), .ZN(n20321) );
  NAND2_X1 U13074 ( .A1(n20239), .A2(n20238), .ZN(n20363) );
  OR2_X1 U13075 ( .A1(n20361), .A2(n20787), .ZN(n20367) );
  INV_X1 U13076 ( .A(n20403), .ZN(n20424) );
  OR2_X1 U13077 ( .A1(n13913), .A2(n20240), .ZN(n20526) );
  OR2_X1 U13078 ( .A1(n13913), .A2(n13562), .ZN(n20688) );
  NAND2_X1 U13079 ( .A1(n13913), .A2(n20240), .ZN(n20628) );
  INV_X1 U13080 ( .A(n20526), .ZN(n20651) );
  NOR2_X2 U13081 ( .A1(n20629), .A2(n20688), .ZN(n20616) );
  INV_X1 U13082 ( .A(n20629), .ZN(n20579) );
  INV_X1 U13083 ( .A(n20406), .ZN(n20292) );
  AND2_X1 U13084 ( .A1(n20719), .A2(n20651), .ZN(n20714) );
  INV_X1 U13085 ( .A(n20802), .ZN(n20741) );
  INV_X1 U13086 ( .A(n20830), .ZN(n20763) );
  INV_X1 U13087 ( .A(n20669), .ZN(n20796) );
  INV_X1 U13088 ( .A(n20678), .ZN(n20823) );
  AND2_X1 U13089 ( .A1(n20292), .A2(n20291), .ZN(n20839) );
  NOR2_X1 U13090 ( .A1(n15368), .A2(n15369), .ZN(n15367) );
  NAND2_X1 U13091 ( .A1(n16385), .A2(n10322), .ZN(n16386) );
  NAND2_X1 U13092 ( .A1(n11282), .A2(n11386), .ZN(n13226) );
  AND2_X1 U13093 ( .A1(n20043), .A2(n13185), .ZN(n19199) );
  NOR2_X1 U13094 ( .A1(n19206), .A2(n14252), .ZN(n14265) );
  INV_X1 U13095 ( .A(n13943), .ZN(n14057) );
  INV_X1 U13096 ( .A(n15493), .ZN(n15481) );
  INV_X1 U13097 ( .A(n19257), .ZN(n19286) );
  INV_X1 U13098 ( .A(n15552), .ZN(n19285) );
  INV_X1 U13099 ( .A(n13308), .ZN(n13297) );
  INV_X1 U13100 ( .A(n14137), .ZN(n14135) );
  OR2_X1 U13101 ( .A1(n15916), .A2(n11743), .ZN(n15872) );
  NOR2_X1 U13102 ( .A1(n15936), .A2(n15915), .ZN(n16468) );
  NAND2_X1 U13103 ( .A1(n13338), .A2(n15888), .ZN(n15889) );
  NAND2_X1 U13104 ( .A1(n13357), .A2(n13360), .ZN(n19986) );
  OAI21_X1 U13105 ( .B1(n19353), .B2(n19352), .A(n19351), .ZN(n19393) );
  INV_X1 U13106 ( .A(n19424), .ZN(n19413) );
  INV_X1 U13107 ( .A(n19416), .ZN(n19450) );
  INV_X1 U13108 ( .A(n19479), .ZN(n19483) );
  AND2_X1 U13109 ( .A1(n19578), .A2(n19756), .ZN(n19567) );
  AND2_X1 U13110 ( .A1(n19988), .A2(n19342), .ZN(n19543) );
  NAND2_X1 U13111 ( .A1(n19607), .A2(n19606), .ZN(n19625) );
  INV_X1 U13112 ( .A(n19650), .ZN(n19664) );
  INV_X1 U13113 ( .A(n19729), .ZN(n19721) );
  INV_X1 U13114 ( .A(n19750), .ZN(n19742) );
  INV_X1 U13115 ( .A(n19848), .ZN(n19764) );
  OAI21_X1 U13116 ( .B1(n19800), .B2(n19799), .A(n19798), .ZN(n19823) );
  INV_X1 U13117 ( .A(n19343), .ZN(n19832) );
  INV_X1 U13118 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19032) );
  NOR2_X1 U13119 ( .A1(n10503), .A2(n10502), .ZN(n16174) );
  INV_X1 U13120 ( .A(n16793), .ZN(n16780) );
  INV_X1 U13121 ( .A(n17056), .ZN(n17091) );
  NOR2_X1 U13122 ( .A1(n17067), .A2(n17079), .ZN(n16923) );
  NOR2_X2 U13123 ( .A1(n18963), .A2(n17079), .ZN(n17043) );
  NAND2_X1 U13124 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17232), .ZN(n17217) );
  NAND2_X1 U13125 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17420), .ZN(n17417) );
  NAND2_X1 U13126 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17435), .ZN(n17434) );
  NOR2_X1 U13127 ( .A1(n17601), .A2(n17465), .ZN(n17460) );
  NAND2_X1 U13128 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17478), .ZN(n17477) );
  NOR2_X1 U13129 ( .A1(n17548), .A2(n17482), .ZN(n17521) );
  INV_X1 U13130 ( .A(n18808), .ZN(n16178) );
  INV_X1 U13131 ( .A(n17536), .ZN(n17546) );
  INV_X1 U13132 ( .A(n17590), .ZN(n17554) );
  INV_X1 U13133 ( .A(n16712), .ZN(n17593) );
  NAND2_X1 U13134 ( .A1(n18227), .A2(n18184), .ZN(n18200) );
  INV_X1 U13135 ( .A(n17854), .ZN(n18224) );
  NAND2_X1 U13136 ( .A1(n17849), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18170) );
  INV_X1 U13137 ( .A(n18330), .ZN(n18334) );
  NOR2_X1 U13138 ( .A1(n13112), .A2(n13107), .ZN(n18791) );
  INV_X1 U13139 ( .A(n18662), .ZN(n18707) );
  NAND3_X1 U13140 ( .A1(n10543), .A2(n10542), .A3(n10541), .ZN(n18379) );
  INV_X1 U13141 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18972) );
  NAND2_X1 U13142 ( .A1(n13324), .A2(n13475), .ZN(n20934) );
  INV_X1 U13143 ( .A(n20126), .ZN(n20080) );
  OR2_X1 U13144 ( .A1(n14615), .A2(n13746), .ZN(n14809) );
  INV_X1 U13145 ( .A(n20084), .ZN(n20140) );
  NAND2_X1 U13146 ( .A1(n14649), .A2(n13085), .ZN(n13104) );
  OR2_X1 U13147 ( .A1(n14859), .A2(n14771), .ZN(n15082) );
  NAND2_X2 U13148 ( .A1(n13083), .A2(n13082), .ZN(n14983) );
  NOR2_X1 U13149 ( .A1(n20144), .A2(n20164), .ZN(n16167) );
  INV_X1 U13150 ( .A(n20144), .ZN(n20166) );
  OAI21_X1 U13151 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n16238) );
  INV_X1 U13152 ( .A(n20189), .ZN(n20056) );
  NAND2_X1 U13153 ( .A1(n15131), .A2(n13684), .ZN(n20193) );
  NAND2_X1 U13154 ( .A1(n13612), .A2(n13596), .ZN(n20225) );
  INV_X1 U13155 ( .A(n20215), .ZN(n16326) );
  OR2_X1 U13156 ( .A1(n20363), .A2(n20526), .ZN(n20308) );
  OR2_X1 U13157 ( .A1(n20363), .A2(n20688), .ZN(n20352) );
  OR2_X1 U13158 ( .A1(n20497), .A2(n20526), .ZN(n20441) );
  OR2_X1 U13159 ( .A1(n20497), .A2(n20688), .ZN(n20484) );
  OR2_X1 U13160 ( .A1(n20497), .A2(n20454), .ZN(n20518) );
  NAND2_X1 U13161 ( .A1(n20579), .A2(n20651), .ZN(n20578) );
  AOI22_X1 U13162 ( .A1(n20587), .A2(n20591), .B1(n20584), .B2(n20583), .ZN(
        n20620) );
  NAND2_X1 U13163 ( .A1(n20579), .A2(n20718), .ZN(n20649) );
  AOI22_X1 U13164 ( .A1(n20662), .A2(n20659), .B1(n20657), .B2(n20656), .ZN(
        n20687) );
  NAND2_X1 U13165 ( .A1(n20719), .A2(n20689), .ZN(n20732) );
  NAND2_X1 U13166 ( .A1(n20719), .A2(n20718), .ZN(n20847) );
  OR2_X1 U13167 ( .A1(n13252), .A2(n16580), .ZN(n20043) );
  OR2_X1 U13168 ( .A1(n20043), .A2(n13847), .ZN(n19214) );
  INV_X1 U13169 ( .A(n15366), .ZN(n15425) );
  AND2_X1 U13170 ( .A1(n12065), .A2(n13362), .ZN(n19250) );
  AND2_X1 U13171 ( .A1(n15534), .A2(n13323), .ZN(n19291) );
  NOR2_X1 U13172 ( .A1(n19293), .A2(n20047), .ZN(n19312) );
  INV_X1 U13173 ( .A(n19293), .ZN(n19326) );
  OR2_X1 U13174 ( .A1(n11762), .A2(n19332), .ZN(n11763) );
  INV_X1 U13175 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16494) );
  OAI21_X1 U13176 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15584), .A(
        n15583), .ZN(n15778) );
  INV_X1 U13177 ( .A(n16566), .ZN(n15966) );
  INV_X1 U13178 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20020) );
  NAND2_X1 U13179 ( .A1(n19639), .A2(n19543), .ZN(n19424) );
  NAND2_X1 U13180 ( .A1(n19543), .A2(n19984), .ZN(n19479) );
  INV_X1 U13181 ( .A(n19513), .ZN(n19491) );
  NAND2_X1 U13182 ( .A1(n19543), .A2(n19756), .ZN(n19537) );
  INV_X1 U13183 ( .A(n19567), .ZN(n19564) );
  NAND2_X1 U13184 ( .A1(n19838), .A2(n19543), .ZN(n19591) );
  INV_X1 U13185 ( .A(n19624), .ZN(n19618) );
  AND2_X1 U13186 ( .A1(n19638), .A2(n19637), .ZN(n19650) );
  INV_X1 U13187 ( .A(n19655), .ZN(n19667) );
  NAND2_X1 U13188 ( .A1(n19668), .A2(n19984), .ZN(n19729) );
  NAND2_X1 U13189 ( .A1(n19640), .A2(n19984), .ZN(n19750) );
  NAND2_X1 U13190 ( .A1(n19668), .A2(n19756), .ZN(n19779) );
  INV_X1 U13191 ( .A(n19821), .ZN(n19818) );
  INV_X1 U13192 ( .A(n19875), .ZN(n19889) );
  OR2_X1 U13193 ( .A1(n16174), .A2(n19026), .ZN(n19028) );
  NOR3_X1 U13194 ( .A1(n16746), .A2(n16745), .A3(n16744), .ZN(n16747) );
  INV_X1 U13195 ( .A(n17043), .ZN(n17080) );
  INV_X1 U13196 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17374) );
  AND2_X1 U13197 ( .A1(n18402), .A2(n17397), .ZN(n17394) );
  NAND2_X1 U13198 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17550), .ZN(n17548) );
  NOR2_X1 U13199 ( .A1(n19011), .A2(n17554), .ZN(n17567) );
  NAND2_X1 U13200 ( .A1(n17593), .A2(n17553), .ZN(n17590) );
  INV_X1 U13201 ( .A(n17943), .ZN(n17901) );
  INV_X1 U13202 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17974) );
  INV_X1 U13203 ( .A(n18326), .ZN(n18344) );
  INV_X1 U13204 ( .A(n18250), .ZN(n18271) );
  INV_X1 U13205 ( .A(n18339), .ZN(n18352) );
  INV_X1 U13206 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18963) );
  INV_X1 U13207 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18886) );
  AND2_X1 U13208 ( .A1(n13096), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20236)
         );
  NAND2_X1 U13209 ( .A1(n13104), .A2(n13103), .ZN(P1_U2874) );
  NAND2_X1 U13210 ( .A1(n11466), .A2(n10332), .ZN(P3_U2799) );
  NOR2_X2 U13211 ( .A1(n18986), .A2(n18979), .ZN(n17063) );
  AOI22_X1 U13212 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U13213 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9832), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10354) );
  INV_X1 U13214 ( .A(n10406), .ZN(n16059) );
  INV_X1 U13215 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17364) );
  NOR2_X2 U13216 ( .A1(n18826), .A2(n10345), .ZN(n10358) );
  AOI22_X1 U13217 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10343) );
  OAI21_X1 U13218 ( .B1(n16059), .B2(n17364), .A(n10343), .ZN(n10352) );
  NOR2_X2 U13219 ( .A1(n18830), .A2(n10344), .ZN(n10378) );
  AOI22_X1 U13220 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13221 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10349) );
  BUF_X4 U13222 ( .A(n10312), .Z(n17325) );
  AOI22_X1 U13223 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13224 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10347) );
  NAND4_X1 U13225 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n10351) );
  AOI211_X1 U13226 ( .C1(n17167), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n10352), .B(n10351), .ZN(n10353) );
  NAND3_X1 U13227 ( .A1(n10355), .A2(n10354), .A3(n10353), .ZN(n16600) );
  AOI22_X1 U13228 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U13229 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10366) );
  INV_X1 U13230 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17372) );
  AOI22_X1 U13231 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10357) );
  OAI21_X1 U13232 ( .B1(n16059), .B2(n17372), .A(n10357), .ZN(n10364) );
  AOI22_X1 U13233 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13234 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U13235 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13236 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10359) );
  NAND4_X1 U13237 ( .A1(n10362), .A2(n10361), .A3(n10360), .A4(n10359), .ZN(
        n10363) );
  AOI211_X1 U13238 ( .C1(n9835), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n10364), .B(n10363), .ZN(n10365) );
  NAND3_X1 U13239 ( .A1(n10367), .A2(n10366), .A3(n10365), .ZN(n10611) );
  AOI22_X1 U13240 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9832), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13241 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10376) );
  INV_X1 U13242 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17379) );
  AOI22_X1 U13243 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10368) );
  OAI21_X1 U13244 ( .B1(n16059), .B2(n17379), .A(n10368), .ZN(n10374) );
  AOI22_X1 U13245 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10372) );
  AOI22_X1 U13246 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13247 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13248 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10312), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10369) );
  NAND4_X1 U13249 ( .A1(n10372), .A2(n10371), .A3(n10370), .A4(n10369), .ZN(
        n10373) );
  AOI211_X1 U13250 ( .C1(n9830), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n10374), .B(n10373), .ZN(n10375) );
  NAND3_X1 U13251 ( .A1(n10377), .A2(n10376), .A3(n10375), .ZN(n17540) );
  AOI22_X1 U13252 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13253 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10388) );
  INV_X1 U13254 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U13255 ( .A1(n10378), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10358), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10379) );
  OAI21_X1 U13256 ( .B1(n16059), .B2(n17389), .A(n10379), .ZN(n10386) );
  AOI22_X1 U13257 ( .A1(n10425), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10356), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U13258 ( .A1(n10405), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10312), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U13259 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13260 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10381) );
  NAND4_X1 U13261 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10385) );
  AOI22_X1 U13262 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U13263 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9821), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10392) );
  AOI22_X1 U13264 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13265 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10312), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10390) );
  NAND4_X1 U13266 ( .A1(n10393), .A2(n10392), .A3(n10391), .A4(n10390), .ZN(
        n10400) );
  AOI22_X1 U13267 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10406), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U13268 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13269 ( .A1(n9814), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U13270 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10395) );
  NAND4_X1 U13271 ( .A1(n10398), .A2(n10397), .A3(n10396), .A4(n10395), .ZN(
        n10399) );
  AOI22_X1 U13272 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10404) );
  AOI22_X1 U13273 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10403) );
  INV_X2 U13274 ( .A(n17166), .ZN(n17113) );
  AOI22_X1 U13275 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U13276 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10401) );
  NAND4_X1 U13277 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n10412) );
  AOI22_X1 U13278 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U13279 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U13280 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9832), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U13281 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10407) );
  NAND4_X1 U13282 ( .A1(n10410), .A2(n10409), .A3(n10408), .A4(n10407), .ZN(
        n10411) );
  AOI22_X1 U13283 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U13284 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13285 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13286 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10413) );
  NAND4_X1 U13287 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10423) );
  INV_X4 U13288 ( .A(n10417), .ZN(n17340) );
  AOI22_X1 U13289 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10421) );
  AOI22_X1 U13290 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9832), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10420) );
  AOI22_X1 U13291 ( .A1(n9814), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10419) );
  AOI22_X1 U13292 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10418) );
  NAND4_X1 U13293 ( .A1(n10421), .A2(n10420), .A3(n10419), .A4(n10418), .ZN(
        n10422) );
  INV_X1 U13294 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18973) );
  OR2_X1 U13295 ( .A1(n9812), .A2(n18973), .ZN(n10435) );
  AOI22_X1 U13296 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13297 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10433) );
  INV_X1 U13298 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17344) );
  AOI22_X1 U13299 ( .A1(n10425), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10424), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13300 ( .A1(n10548), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13301 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10312), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13302 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10426) );
  NAND4_X1 U13303 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10430) );
  AOI211_X1 U13304 ( .C1(n9830), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n10431), .B(n10430), .ZN(n10432) );
  NAND3_X1 U13305 ( .A1(n10434), .A2(n10433), .A3(n10432), .ZN(n16179) );
  INV_X1 U13306 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18991) );
  INV_X1 U13307 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18329) );
  INV_X1 U13308 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18308) );
  XOR2_X1 U13309 ( .A(n10440), .B(n10439), .Z(n18005) );
  NAND2_X1 U13310 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n10441), .ZN(
        n10442) );
  XOR2_X1 U13311 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n10443), .Z(
        n17988) );
  NAND2_X1 U13312 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n10443), .ZN(
        n10444) );
  XNOR2_X1 U13313 ( .A(n10445), .B(n10611), .ZN(n10448) );
  NAND2_X1 U13314 ( .A1(n10448), .A2(n10447), .ZN(n10449) );
  XNOR2_X1 U13315 ( .A(n10609), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17970) );
  INV_X1 U13316 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18284) );
  INV_X1 U13317 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18263) );
  INV_X1 U13318 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10461) );
  INV_X1 U13319 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10456) );
  INV_X1 U13320 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10455) );
  INV_X1 U13321 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18190) );
  AND2_X1 U13322 ( .A1(n10457), .A2(n18190), .ZN(n10458) );
  NAND2_X1 U13323 ( .A1(n18267), .A2(n17932), .ZN(n17931) );
  NAND2_X1 U13324 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n10459), .ZN(
        n10460) );
  NAND2_X1 U13325 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18230) );
  NOR2_X1 U13326 ( .A1(n18230), .A2(n10461), .ZN(n18214) );
  INV_X1 U13327 ( .A(n18214), .ZN(n18201) );
  NOR2_X1 U13328 ( .A1(n18201), .A2(n10456), .ZN(n18184) );
  NAND2_X1 U13329 ( .A1(n18184), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18191) );
  OR2_X1 U13330 ( .A1(n18190), .A2(n18191), .ZN(n18172) );
  NOR2_X1 U13331 ( .A1(n10455), .A2(n18172), .ZN(n13119) );
  INV_X1 U13332 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18162) );
  INV_X1 U13333 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18145) );
  NAND2_X1 U13334 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18102) );
  INV_X1 U13335 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17814) );
  NOR2_X1 U13336 ( .A1(n18102), .A2(n17814), .ZN(n17770) );
  INV_X1 U13337 ( .A(n17770), .ZN(n17783) );
  INV_X1 U13338 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17801) );
  INV_X1 U13339 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18098) );
  NOR2_X1 U13340 ( .A1(n17801), .A2(n18098), .ZN(n18120) );
  NAND2_X1 U13341 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18120), .ZN(
        n18105) );
  NOR2_X1 U13342 ( .A1(n17783), .A2(n18105), .ZN(n18107) );
  INV_X1 U13343 ( .A(n18107), .ZN(n18097) );
  INV_X1 U13344 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18114) );
  NOR2_X1 U13345 ( .A1(n18097), .A2(n18114), .ZN(n18037) );
  NAND2_X1 U13346 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18037), .ZN(
        n18064) );
  INV_X1 U13347 ( .A(n18064), .ZN(n18078) );
  NOR2_X1 U13348 ( .A1(n17826), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17809) );
  NAND2_X1 U13349 ( .A1(n17809), .A2(n17801), .ZN(n10464) );
  NOR2_X1 U13350 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n10464), .ZN(
        n17768) );
  INV_X1 U13351 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18116) );
  NAND2_X1 U13352 ( .A1(n17768), .A2(n18116), .ZN(n17753) );
  NOR3_X1 U13353 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17753), .ZN(n10465) );
  INV_X1 U13354 ( .A(n18102), .ZN(n18143) );
  NAND2_X1 U13355 ( .A1(n18143), .A2(n10466), .ZN(n17766) );
  NAND2_X1 U13356 ( .A1(n17733), .A2(n17766), .ZN(n17767) );
  NOR2_X1 U13357 ( .A1(n18105), .A2(n18114), .ZN(n13120) );
  AND2_X1 U13358 ( .A1(n13120), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10467) );
  NAND2_X1 U13359 ( .A1(n17767), .A2(n10467), .ZN(n17734) );
  INV_X1 U13360 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18091) );
  INV_X1 U13361 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18069) );
  NAND2_X1 U13362 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18042) );
  AND2_X1 U13363 ( .A1(n17826), .A2(n18042), .ZN(n10468) );
  NAND2_X1 U13364 ( .A1(n17826), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16597) );
  NOR2_X1 U13365 ( .A1(n17680), .A2(n16597), .ZN(n10469) );
  NAND2_X1 U13366 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n10469), .ZN(
        n11445) );
  INV_X1 U13367 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17661) );
  NAND2_X1 U13368 ( .A1(n17932), .A2(n17661), .ZN(n16598) );
  INV_X1 U13369 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18363) );
  OAI22_X1 U13370 ( .A1(n18979), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18367), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10476) );
  OAI22_X1 U13371 ( .A1(n18986), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18636), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U13372 ( .A1(n18368), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10591) );
  NOR2_X1 U13373 ( .A1(n10592), .A2(n10591), .ZN(n10471) );
  OAI22_X1 U13374 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18363), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n10473), .ZN(n10478) );
  NOR2_X1 U13375 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18363), .ZN(
        n10474) );
  NAND2_X1 U13376 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10473), .ZN(
        n10479) );
  AOI22_X1 U13377 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n10478), .B1(
        n10474), .B2(n10479), .ZN(n10483) );
  OAI21_X1 U13378 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18368), .A(
        n10591), .ZN(n10590) );
  NOR2_X1 U13379 ( .A1(n10592), .A2(n10590), .ZN(n10482) );
  OAI21_X1 U13380 ( .B1(n10477), .B2(n10476), .A(n10483), .ZN(n10475) );
  AOI21_X1 U13381 ( .B1(n10477), .B2(n10476), .A(n10475), .ZN(n10589) );
  AOI21_X1 U13382 ( .B1(n10479), .B2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n10478), .ZN(n10480) );
  AOI21_X1 U13383 ( .B1(n18363), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n10480), .ZN(n10593) );
  INV_X1 U13384 ( .A(n10593), .ZN(n10481) );
  AOI211_X2 U13385 ( .C1(n10483), .C2(n10482), .A(n10589), .B(n10481), .ZN(
        n18797) );
  AOI22_X1 U13386 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13387 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13388 ( .A1(n17113), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13389 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10484) );
  NAND4_X1 U13390 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10493) );
  AOI22_X1 U13391 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10491) );
  AOI22_X1 U13392 ( .A1(n9814), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13393 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13394 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10488) );
  NAND4_X1 U13395 ( .A1(n10491), .A2(n10490), .A3(n10489), .A4(n10488), .ZN(
        n10492) );
  AOI22_X1 U13396 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9833), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13397 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13398 ( .A1(n17113), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U13399 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10494) );
  NAND4_X1 U13400 ( .A1(n10497), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        n10503) );
  AOI22_X1 U13401 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U13402 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13403 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13404 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10498) );
  NAND4_X1 U13405 ( .A1(n10501), .A2(n10500), .A3(n10499), .A4(n10498), .ZN(
        n10502) );
  INV_X2 U13406 ( .A(n16174), .ZN(n18366) );
  NAND2_X1 U13407 ( .A1(n19014), .A2(n18366), .ZN(n10566) );
  NAND2_X1 U13408 ( .A1(n10580), .A2(n10566), .ZN(n19025) );
  INV_X1 U13409 ( .A(n19025), .ZN(n19017) );
  AOI22_X1 U13410 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17299), .ZN(n10507) );
  AOI22_X1 U13411 ( .A1(n17340), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17325), .ZN(n10506) );
  INV_X2 U13412 ( .A(n17121), .ZN(n17326) );
  AOI22_X1 U13413 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17326), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10505) );
  AOI22_X1 U13414 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9821), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10504) );
  NAND4_X1 U13415 ( .A1(n10507), .A2(n10506), .A3(n10505), .A4(n10504), .ZN(
        n10513) );
  AOI22_X1 U13416 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n9813), .ZN(n10511) );
  AOI22_X1 U13417 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13418 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9832), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13419 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17347), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n9833), .ZN(n10508) );
  NAND4_X1 U13420 ( .A1(n10511), .A2(n10510), .A3(n10509), .A4(n10508), .ZN(
        n10512) );
  AOI22_X1 U13421 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10517) );
  AOI22_X1 U13422 ( .A1(n17340), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U13423 ( .A1(n17113), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13424 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10514) );
  NAND4_X1 U13425 ( .A1(n10517), .A2(n10516), .A3(n10515), .A4(n10514), .ZN(
        n10523) );
  AOI22_X1 U13426 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13427 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13428 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9813), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13429 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10518) );
  NAND4_X1 U13430 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10522) );
  AOI22_X1 U13431 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13432 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13433 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13434 ( .A1(n17113), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10524) );
  NAND4_X1 U13435 ( .A1(n10527), .A2(n10526), .A3(n10525), .A4(n10524), .ZN(
        n10533) );
  AOI22_X1 U13436 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13437 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13438 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13439 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9813), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10528) );
  NAND4_X1 U13440 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10532) );
  AOI22_X1 U13441 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13442 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10542) );
  INV_X1 U13443 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U13444 ( .A1(n17340), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10534) );
  OAI21_X1 U13445 ( .B1(n10556), .B2(n17387), .A(n10534), .ZN(n10540) );
  AOI22_X1 U13446 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10538) );
  AOI22_X1 U13447 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9832), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13448 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13449 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10535) );
  NAND4_X1 U13450 ( .A1(n10538), .A2(n10537), .A3(n10536), .A4(n10535), .ZN(
        n10539) );
  AOI22_X1 U13451 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13452 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13453 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13454 ( .A1(n17113), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10544) );
  NAND4_X1 U13455 ( .A1(n10547), .A2(n10546), .A3(n10545), .A4(n10544), .ZN(
        n10554) );
  AOI22_X1 U13456 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9813), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U13457 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U13458 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U13459 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10549) );
  NAND4_X1 U13460 ( .A1(n10552), .A2(n10551), .A3(n10550), .A4(n10549), .ZN(
        n10553) );
  AOI22_X1 U13461 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13462 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10564) );
  INV_X1 U13463 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U13464 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10555) );
  OAI21_X1 U13465 ( .B1(n10556), .B2(n17369), .A(n10555), .ZN(n10562) );
  AOI22_X1 U13466 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9833), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13467 ( .A1(n17347), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13468 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13469 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10557) );
  NAND4_X1 U13470 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n10561) );
  AOI211_X1 U13471 ( .C1(n9835), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n10562), .B(n10561), .ZN(n10563) );
  NAND3_X1 U13472 ( .A1(n10565), .A2(n10564), .A3(n10563), .ZN(n18397) );
  NOR2_X1 U13473 ( .A1(n15993), .A2(n18397), .ZN(n10584) );
  AND3_X1 U13474 ( .A1(n10599), .A2(n13115), .A3(n10584), .ZN(n14414) );
  NOR2_X2 U13475 ( .A1(n18383), .A2(n18379), .ZN(n15992) );
  NAND2_X1 U13476 ( .A1(n10597), .A2(n15993), .ZN(n10569) );
  NAND2_X1 U13477 ( .A1(n10597), .A2(n18392), .ZN(n18808) );
  NOR2_X1 U13478 ( .A1(n17367), .A2(n16178), .ZN(n16177) );
  NOR2_X1 U13479 ( .A1(n10566), .A2(n16177), .ZN(n13105) );
  INV_X1 U13480 ( .A(n13105), .ZN(n10567) );
  OAI21_X1 U13481 ( .B1(n13115), .B2(n10575), .A(n10567), .ZN(n10574) );
  INV_X1 U13482 ( .A(n10576), .ZN(n10571) );
  INV_X1 U13483 ( .A(n18379), .ZN(n13109) );
  NAND2_X1 U13484 ( .A1(n13109), .A2(n10580), .ZN(n10596) );
  AOI21_X1 U13485 ( .B1(n13109), .B2(n16174), .A(n16178), .ZN(n10568) );
  AOI21_X1 U13486 ( .B1(n10569), .B2(n10571), .A(n10568), .ZN(n10570) );
  AOI21_X1 U13487 ( .B1(n10571), .B2(n10596), .A(n10570), .ZN(n10573) );
  INV_X1 U13488 ( .A(n15993), .ZN(n18387) );
  OAI21_X1 U13489 ( .B1(n17367), .B2(n10576), .A(n18387), .ZN(n10572) );
  INV_X1 U13490 ( .A(n10599), .ZN(n10582) );
  AND4_X2 U13491 ( .A1(n18366), .A2(n10599), .A3(n10585), .A4(n10575), .ZN(
        n18848) );
  INV_X1 U13492 ( .A(n14415), .ZN(n10581) );
  NAND3_X1 U13493 ( .A1(n10582), .A2(n18375), .A3(n10581), .ZN(n10583) );
  AOI21_X4 U13494 ( .B1(n15992), .B2(n18820), .A(n10588), .ZN(n18809) );
  INV_X1 U13495 ( .A(n10589), .ZN(n10594) );
  NOR2_X1 U13496 ( .A1(n10594), .A2(n10590), .ZN(n13113) );
  XNOR2_X1 U13497 ( .A(n10592), .B(n10591), .ZN(n10595) );
  NOR2_X1 U13498 ( .A1(n13113), .A2(n18793), .ZN(n18795) );
  NOR2_X1 U13499 ( .A1(n19014), .A2(n18379), .ZN(n13111) );
  NAND2_X1 U13500 ( .A1(n13111), .A2(n18397), .ZN(n13112) );
  INV_X1 U13501 ( .A(n10596), .ZN(n10600) );
  NOR2_X1 U13502 ( .A1(n10597), .A2(n18392), .ZN(n15991) );
  OAI21_X1 U13503 ( .B1(n15991), .B2(n18387), .A(n18808), .ZN(n10598) );
  NAND3_X1 U13504 ( .A1(n10600), .A2(n10599), .A3(n10598), .ZN(n13107) );
  NAND2_X1 U13505 ( .A1(n18972), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18862) );
  INV_X1 U13506 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18354) );
  NOR2_X1 U13507 ( .A1(n18862), .A2(n18354), .ZN(n19009) );
  INV_X1 U13508 ( .A(n19009), .ZN(n18856) );
  NAND2_X2 U13509 ( .A1(n10601), .A2(n18375), .ZN(n18035) );
  NAND2_X1 U13510 ( .A1(n16161), .A2(n17926), .ZN(n10637) );
  NAND2_X1 U13511 ( .A1(n18972), .A2(n18963), .ZN(n18967) );
  NAND2_X1 U13512 ( .A1(n18354), .A2(n18963), .ZN(n16714) );
  AND2_X1 U13513 ( .A1(n18967), .A2(n16714), .ZN(n19008) );
  INV_X1 U13514 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19013) );
  NOR2_X1 U13515 ( .A1(n18972), .A2(n19013), .ZN(n17993) );
  INV_X1 U13516 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16754) );
  INV_X1 U13517 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16763) );
  NAND2_X1 U13518 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17936) );
  INV_X1 U13519 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17918) );
  NOR2_X1 U13520 ( .A1(n17936), .A2(n17918), .ZN(n17894) );
  INV_X1 U13521 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17882) );
  INV_X1 U13522 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17868) );
  NOR2_X1 U13523 ( .A1(n17882), .A2(n17868), .ZN(n17867) );
  NAND2_X1 U13524 ( .A1(n17867), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17829) );
  NAND2_X1 U13525 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17830) );
  INV_X1 U13526 ( .A(n17830), .ZN(n10602) );
  INV_X1 U13527 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17777) );
  INV_X1 U13528 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17745) );
  NAND3_X1 U13529 ( .A1(n17718), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17696) );
  INV_X1 U13530 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17695) );
  INV_X1 U13531 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16775) );
  XNOR2_X1 U13532 ( .A(n16754), .B(n16591), .ZN(n16750) );
  NOR2_X1 U13533 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18967), .ZN(n19027) );
  INV_X1 U13534 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18859) );
  INV_X1 U13535 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18950) );
  NOR2_X1 U13536 ( .A1(n18345), .A2(n18950), .ZN(n16160) );
  NAND2_X1 U13537 ( .A1(n18859), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18870) );
  INV_X1 U13538 ( .A(n17750), .ZN(n17776) );
  NOR2_X1 U13539 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17776), .ZN(
        n16592) );
  INV_X1 U13540 ( .A(n18870), .ZN(n17862) );
  NOR2_X1 U13541 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18963), .ZN(
        n18988) );
  NOR2_X1 U13542 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19018) );
  AOI21_X1 U13543 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n19018), .ZN(n18867) );
  NOR2_X1 U13544 ( .A1(n18988), .A2(n18867), .ZN(n18365) );
  NAND3_X1 U13545 ( .A1(n18354), .A2(n18963), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18611) );
  NOR2_X1 U13546 ( .A1(n18707), .A2(n18611), .ZN(n18384) );
  NAND2_X1 U13547 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n10020), .ZN(
        n10605) );
  AOI22_X1 U13548 ( .A1(n17862), .A2(n16740), .B1(n18738), .B2(n10605), .ZN(
        n10604) );
  NAND2_X1 U13549 ( .A1(n10604), .A2(n18032), .ZN(n16584) );
  NOR2_X1 U13550 ( .A1(n16592), .A2(n16584), .ZN(n11458) );
  OR2_X1 U13551 ( .A1(n10605), .A2(n17865), .ZN(n11460) );
  AOI22_X1 U13552 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n11458), .B1(
        n11460), .B2(n16754), .ZN(n10606) );
  AOI211_X1 U13553 ( .C1(n17890), .C2(n16750), .A(n16160), .B(n10606), .ZN(
        n10636) );
  NOR2_X2 U13554 ( .A1(n18170), .A2(n10455), .ZN(n18169) );
  INV_X1 U13555 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18083) );
  NOR2_X1 U13556 ( .A1(n18064), .A2(n18083), .ZN(n17712) );
  INV_X1 U13557 ( .A(n17712), .ZN(n18068) );
  NOR2_X1 U13558 ( .A1(n18068), .A2(n18042), .ZN(n17683) );
  NAND2_X1 U13559 ( .A1(n18169), .A2(n17683), .ZN(n18043) );
  NAND2_X1 U13560 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16094) );
  OR2_X1 U13561 ( .A1(n16094), .A2(n9871), .ZN(n13128) );
  NOR2_X2 U13562 ( .A1(n16600), .A2(n18035), .ZN(n17943) );
  NAND2_X1 U13563 ( .A1(n9812), .A2(n16179), .ZN(n10618) );
  NAND2_X1 U13564 ( .A1(n10607), .A2(n10618), .ZN(n10616) );
  NAND2_X1 U13565 ( .A1(n17540), .A2(n10616), .ZN(n10613) );
  NOR2_X1 U13566 ( .A1(n17535), .A2(n10613), .ZN(n10610) );
  NAND2_X1 U13567 ( .A1(n10610), .A2(n10611), .ZN(n17966) );
  NOR2_X1 U13568 ( .A1(n17528), .A2(n17966), .ZN(n10608) );
  NAND2_X1 U13569 ( .A1(n10608), .A2(n16600), .ZN(n10627) );
  XNOR2_X1 U13570 ( .A(n16600), .B(n10608), .ZN(n17948) );
  INV_X1 U13571 ( .A(n17966), .ZN(n17968) );
  XOR2_X1 U13572 ( .A(n10609), .B(n17968), .Z(n10626) );
  XOR2_X1 U13573 ( .A(n10611), .B(n10610), .Z(n10612) );
  NAND2_X1 U13574 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n10612), .ZN(
        n10625) );
  XOR2_X1 U13575 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n10612), .Z(
        n17977) );
  XNOR2_X1 U13576 ( .A(n10614), .B(n10613), .ZN(n10615) );
  NAND2_X1 U13577 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n10615), .ZN(
        n10624) );
  XOR2_X1 U13578 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n10615), .Z(
        n17991) );
  XOR2_X1 U13579 ( .A(n17540), .B(n10616), .Z(n10617) );
  NAND2_X1 U13580 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n10617), .ZN(
        n10623) );
  XOR2_X1 U13581 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n10617), .Z(
        n18002) );
  XNOR2_X1 U13582 ( .A(n17543), .B(n10618), .ZN(n10621) );
  OR2_X1 U13583 ( .A1(n18329), .A2(n10621), .ZN(n10622) );
  AOI21_X1 U13584 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n9812), .A(
        n16179), .ZN(n10620) );
  NOR2_X1 U13585 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n9812), .ZN(
        n10619) );
  AOI221_X1 U13586 ( .B1(n16179), .B2(n9812), .C1(n10620), .C2(n18991), .A(
        n10619), .ZN(n18013) );
  XOR2_X1 U13587 ( .A(n18329), .B(n10621), .Z(n18012) );
  NAND2_X1 U13588 ( .A1(n18013), .A2(n18012), .ZN(n18011) );
  NAND2_X1 U13589 ( .A1(n10622), .A2(n18011), .ZN(n18001) );
  NAND2_X1 U13590 ( .A1(n18002), .A2(n18001), .ZN(n18000) );
  NAND2_X1 U13591 ( .A1(n10623), .A2(n18000), .ZN(n17990) );
  NAND2_X1 U13592 ( .A1(n17991), .A2(n17990), .ZN(n17989) );
  NAND2_X1 U13593 ( .A1(n10624), .A2(n17989), .ZN(n17976) );
  NAND2_X1 U13594 ( .A1(n17977), .A2(n17976), .ZN(n17975) );
  NAND2_X1 U13595 ( .A1(n10625), .A2(n17975), .ZN(n17967) );
  AOI222_X1 U13596 ( .A1(n10626), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n10626), .B2(n17967), .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(
        n17967), .ZN(n17949) );
  NAND2_X1 U13597 ( .A1(n17948), .A2(n17949), .ZN(n17947) );
  NAND2_X1 U13598 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17947), .ZN(
        n10630) );
  NOR2_X1 U13599 ( .A1(n10627), .A2(n10630), .ZN(n10632) );
  INV_X1 U13600 ( .A(n10627), .ZN(n10631) );
  NOR2_X1 U13601 ( .A1(n17948), .A2(n17949), .ZN(n10629) );
  NOR2_X1 U13602 ( .A1(n10631), .A2(n10630), .ZN(n10628) );
  AOI211_X1 U13603 ( .C1(n10631), .C2(n10630), .A(n10629), .B(n10628), .ZN(
        n17934) );
  NOR2_X1 U13604 ( .A1(n17934), .A2(n18263), .ZN(n17933) );
  INV_X1 U13605 ( .A(n13119), .ZN(n18147) );
  NAND2_X1 U13606 ( .A1(n17683), .A2(n18168), .ZN(n18045) );
  NOR2_X1 U13607 ( .A1(n13128), .A2(n18045), .ZN(n16585) );
  NOR2_X2 U13608 ( .A1(n18375), .A2(n16719), .ZN(n18026) );
  OAI22_X1 U13609 ( .A1(n16589), .A2(n17901), .B1(n16585), .B2(n18036), .ZN(
        n10633) );
  NAND2_X1 U13610 ( .A1(n10633), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10635) );
  AOI22_X1 U13611 ( .A1(n17943), .A2(n18227), .B1(n18026), .B2(n18224), .ZN(
        n17930) );
  INV_X1 U13612 ( .A(n17930), .ZN(n17900) );
  NAND2_X1 U13613 ( .A1(n17900), .A2(n13119), .ZN(n17756) );
  INV_X1 U13614 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16164) );
  NAND3_X1 U13615 ( .A1(n17683), .A2(n17836), .A3(n16164), .ZN(n10634) );
  NAND2_X1 U13616 ( .A1(n10637), .A2(n10333), .ZN(P3_U2800) );
  NOR2_X2 U13617 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10638) );
  AND2_X4 U13618 ( .A1(n10638), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10868) );
  AOI22_X1 U13619 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10640) );
  AND2_X4 U13620 ( .A1(n13792), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10674) );
  AOI22_X1 U13621 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10643) );
  AOI22_X1 U13622 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9954), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U13623 ( .A1(n10337), .A2(n9993), .ZN(n10651) );
  AOI22_X1 U13624 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13625 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9955), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U13626 ( .A1(n9931), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10646) );
  NAND4_X1 U13627 ( .A1(n10649), .A2(n10648), .A3(n10647), .A4(n10646), .ZN(
        n10650) );
  AOI22_X1 U13628 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13629 ( .A1(n9928), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13630 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10654) );
  NAND4_X1 U13631 ( .A1(n10657), .A2(n10656), .A3(n10655), .A4(n10654), .ZN(
        n10658) );
  AOI22_X1 U13632 ( .A1(n9929), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13633 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10661) );
  AOI22_X1 U13634 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10660) );
  NAND4_X1 U13635 ( .A1(n10662), .A2(n10661), .A3(n10660), .A4(n10659), .ZN(
        n10663) );
  AOI22_X1 U13636 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9953), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10669) );
  AOI22_X1 U13637 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13638 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9955), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13639 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13640 ( .A1(n9928), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13641 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13642 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13643 ( .A1(n9931), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13644 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U13645 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13646 ( .A1(n9929), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13647 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13648 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10678) );
  NAND4_X1 U13649 ( .A1(n9827), .A2(n9819), .A3(n13364), .A4(n19373), .ZN(
        n10699) );
  AOI22_X1 U13650 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13651 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9956), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13652 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13653 ( .A1(n9931), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10687) );
  AOI22_X1 U13654 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9956), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U13655 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10685) );
  AOI22_X1 U13656 ( .A1(n9928), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13657 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13658 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U13659 ( .A1(n9817), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13660 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13661 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13662 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13663 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10693) );
  NAND4_X1 U13664 ( .A1(n10696), .A2(n10695), .A3(n10694), .A4(n10693), .ZN(
        n10697) );
  AOI22_X1 U13665 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10863), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13666 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13667 ( .A1(n9956), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10700) );
  NAND4_X1 U13668 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(
        n10704) );
  AOI22_X1 U13669 ( .A1(n9929), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U13670 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13671 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9954), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13672 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9953), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10705) );
  NAND4_X1 U13673 ( .A1(n10708), .A2(n10707), .A3(n10706), .A4(n10705), .ZN(
        n10709) );
  NOR2_X2 U13674 ( .A1(n10745), .A2(n10752), .ZN(n10733) );
  AOI22_X1 U13675 ( .A1(n9929), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13676 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13677 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13678 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9953), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13679 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9955), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10717) );
  AOI22_X1 U13680 ( .A1(n9929), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13681 ( .A1(n9818), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10719) );
  INV_X2 U13682 ( .A(n10721), .ZN(n11508) );
  NAND2_X1 U13683 ( .A1(n10759), .A2(n11513), .ZN(n10730) );
  NAND2_X1 U13684 ( .A1(n10721), .A2(n9819), .ZN(n10725) );
  INV_X1 U13685 ( .A(n19373), .ZN(n11494) );
  INV_X1 U13686 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14394) );
  NAND2_X1 U13687 ( .A1(n11702), .A2(n10732), .ZN(n11717) );
  NAND2_X1 U13688 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10736) );
  INV_X1 U13689 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10734) );
  OAI211_X1 U13690 ( .C1(n11400), .C2(n14273), .A(n10736), .B(n10735), .ZN(
        n10737) );
  INV_X1 U13691 ( .A(n11702), .ZN(n10754) );
  NOR2_X1 U13692 ( .A1(n12066), .A2(n13179), .ZN(n11704) );
  NAND2_X1 U13693 ( .A1(n10754), .A2(n11704), .ZN(n10778) );
  NAND2_X1 U13694 ( .A1(n10778), .A2(n20035), .ZN(n10743) );
  OAI211_X1 U13695 ( .C1(n12066), .C2(n9819), .A(n19361), .B(n10751), .ZN(
        n10742) );
  INV_X1 U13696 ( .A(n10739), .ZN(n10740) );
  NAND2_X1 U13697 ( .A1(n10743), .A2(n11711), .ZN(n10744) );
  NAND2_X1 U13698 ( .A1(n10744), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10750) );
  INV_X1 U13699 ( .A(n10745), .ZN(n10747) );
  AND2_X1 U13700 ( .A1(n13179), .A2(n19361), .ZN(n10748) );
  NAND2_X1 U13701 ( .A1(n14134), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11405) );
  NAND2_X1 U13702 ( .A1(n10752), .A2(n10751), .ZN(n11490) );
  NAND2_X1 U13703 ( .A1(n11712), .A2(n10723), .ZN(n10756) );
  NAND2_X1 U13704 ( .A1(n10779), .A2(n10757), .ZN(n10758) );
  NAND2_X1 U13705 ( .A1(n10783), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10761) );
  NOR2_X1 U13706 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U13707 ( .A1(n10759), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13846), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10760) );
  NAND2_X1 U13708 ( .A1(n10761), .A2(n10760), .ZN(n10791) );
  XNOR2_X1 U13709 ( .A(n10792), .B(n10791), .ZN(n10819) );
  NAND2_X1 U13710 ( .A1(n10768), .A2(n20026), .ZN(n10764) );
  NAND2_X1 U13711 ( .A1(n10764), .A2(n13814), .ZN(n10767) );
  AND2_X1 U13712 ( .A1(n10729), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10766) );
  AOI21_X1 U13713 ( .B1(n10767), .B2(n10766), .A(n10765), .ZN(n10770) );
  NAND2_X1 U13714 ( .A1(n10783), .A2(n10768), .ZN(n10769) );
  NAND2_X1 U13715 ( .A1(n10770), .A2(n10769), .ZN(n10814) );
  INV_X1 U13716 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13367) );
  INV_X1 U13717 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11136) );
  INV_X1 U13718 ( .A(n13846), .ZN(n10772) );
  NAND2_X1 U13719 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10771) );
  AND2_X1 U13720 ( .A1(n10772), .A2(n10771), .ZN(n10775) );
  NAND2_X1 U13721 ( .A1(n10773), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10774) );
  OAI211_X1 U13722 ( .C1(n11400), .C2(n11136), .A(n10775), .B(n10774), .ZN(
        n10776) );
  INV_X1 U13723 ( .A(n10777), .ZN(n10780) );
  NAND2_X1 U13724 ( .A1(n10819), .A2(n10828), .ZN(n10809) );
  INV_X1 U13725 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n14396) );
  OAI21_X1 U13726 ( .B1(n20002), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n14396), 
        .ZN(n10784) );
  INV_X1 U13727 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10787) );
  NAND2_X1 U13728 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10786) );
  NAND2_X1 U13729 ( .A1(n10773), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10785) );
  OAI211_X1 U13730 ( .C1(n11400), .C2(n10787), .A(n10786), .B(n10785), .ZN(
        n10788) );
  INV_X1 U13731 ( .A(n10788), .ZN(n10789) );
  NAND2_X1 U13732 ( .A1(n10796), .A2(n10797), .ZN(n10794) );
  INV_X1 U13733 ( .A(n10791), .ZN(n10793) );
  NAND2_X1 U13734 ( .A1(n10793), .A2(n10792), .ZN(n10808) );
  NAND2_X1 U13735 ( .A1(n10809), .A2(n10795), .ZN(n10800) );
  INV_X1 U13736 ( .A(n10797), .ZN(n10798) );
  NAND2_X1 U13737 ( .A1(n10810), .A2(n10798), .ZN(n10799) );
  NAND2_X1 U13738 ( .A1(n10783), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10802) );
  NAND2_X1 U13739 ( .A1(n13846), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10801) );
  INV_X1 U13740 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14030) );
  INV_X1 U13741 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n14148) );
  NAND2_X1 U13742 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10805) );
  NAND2_X1 U13743 ( .A1(n10773), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10804) );
  OAI211_X1 U13744 ( .C1(n11400), .C2(n14148), .A(n10805), .B(n10804), .ZN(
        n10806) );
  INV_X1 U13745 ( .A(n10806), .ZN(n10807) );
  NAND2_X1 U13746 ( .A1(n10809), .A2(n10808), .ZN(n10812) );
  XNOR2_X2 U13747 ( .A(n10812), .B(n10811), .ZN(n10838) );
  INV_X1 U13748 ( .A(n10814), .ZN(n10817) );
  INV_X1 U13749 ( .A(n10815), .ZN(n10816) );
  NAND2_X1 U13750 ( .A1(n10817), .A2(n10816), .ZN(n10818) );
  AND2_X2 U13751 ( .A1(n10818), .A2(n10828), .ZN(n19224) );
  INV_X1 U13752 ( .A(n10829), .ZN(n10820) );
  NAND2_X1 U13753 ( .A1(n19224), .A2(n10820), .ZN(n10836) );
  INV_X1 U13754 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U13755 ( .A1(n19224), .A2(n10829), .ZN(n10852) );
  INV_X1 U13756 ( .A(n10852), .ZN(n10822) );
  INV_X2 U13757 ( .A(n11765), .ZN(n13532) );
  NAND2_X1 U13758 ( .A1(n19464), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10825) );
  AND2_X1 U13759 ( .A1(n10822), .A2(n10838), .ZN(n10823) );
  INV_X1 U13760 ( .A(n10827), .ZN(n10831) );
  XNOR2_X2 U13761 ( .A(n10829), .B(n10828), .ZN(n11777) );
  INV_X1 U13762 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10834) );
  NAND2_X1 U13763 ( .A1(n10838), .A2(n11765), .ZN(n10854) );
  INV_X1 U13764 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10833) );
  OAI22_X1 U13765 ( .A1(n10834), .A2(n19829), .B1(n19675), .B2(n10833), .ZN(
        n10835) );
  AOI21_X1 U13766 ( .B1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n10957), .A(
        n10835), .ZN(n10860) );
  INV_X1 U13767 ( .A(n10836), .ZN(n10842) );
  AND2_X1 U13768 ( .A1(n10840), .A2(n10842), .ZN(n10837) );
  AND2_X1 U13769 ( .A1(n10838), .A2(n10842), .ZN(n10839) );
  AOI22_X1 U13770 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19397), .B1(
        n19517), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10847) );
  AND2_X1 U13771 ( .A1(n10840), .A2(n13818), .ZN(n10841) );
  NAND2_X1 U13772 ( .A1(n19350), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10846) );
  NAND2_X1 U13773 ( .A1(n10941), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10845) );
  AND2_X1 U13774 ( .A1(n10838), .A2(n13818), .ZN(n10843) );
  NAND2_X1 U13775 ( .A1(n19488), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10844) );
  INV_X1 U13776 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10851) );
  INV_X1 U13777 ( .A(n10853), .ZN(n10848) );
  INV_X1 U13778 ( .A(n10854), .ZN(n10849) );
  INV_X1 U13779 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10850) );
  OAI22_X1 U13780 ( .A1(n10851), .A2(n10902), .B1(n10903), .B2(n10850), .ZN(
        n10857) );
  INV_X1 U13781 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10855) );
  INV_X1 U13782 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n19732) );
  OAI22_X1 U13783 ( .A1(n10855), .A2(n19700), .B1(n14124), .B2(n19732), .ZN(
        n10856) );
  NOR2_X1 U13784 ( .A1(n10857), .A2(n10856), .ZN(n10858) );
  AOI22_X1 U13785 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11064), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13786 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n11021), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10866) );
  AND2_X2 U13787 ( .A1(n9931), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11057) );
  INV_X1 U13788 ( .A(n10863), .ZN(n13787) );
  AND2_X2 U13789 ( .A1(n9953), .A2(n13827), .ZN(n13809) );
  AOI22_X1 U13790 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13791 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9980), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10864) );
  NAND4_X1 U13792 ( .A1(n10867), .A2(n10866), .A3(n10865), .A4(n10864), .ZN(
        n10874) );
  AOI22_X1 U13793 ( .A1(n10929), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n11840), .ZN(n10872) );
  AOI22_X1 U13794 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11558), .B1(
        n11069), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10871) );
  AND2_X2 U13795 ( .A1(n9954), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11022) );
  AOI22_X1 U13796 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n11022), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10870) );
  AOI22_X1 U13797 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11020), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10869) );
  NAND4_X1 U13798 ( .A1(n10872), .A2(n10871), .A3(n10870), .A4(n10869), .ZN(
        n10873) );
  NOR2_X1 U13799 ( .A1(n10874), .A2(n10873), .ZN(n11135) );
  AOI22_X1 U13800 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11558), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13801 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11840), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13802 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U13803 ( .A1(n11064), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10875) );
  NAND4_X1 U13804 ( .A1(n10878), .A2(n10877), .A3(n10876), .A4(n10875), .ZN(
        n10884) );
  AOI22_X1 U13805 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11021), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10882) );
  AOI22_X1 U13806 ( .A1(n13809), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13807 ( .A1(n10929), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13808 ( .A1(n11022), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10879) );
  NAND4_X1 U13809 ( .A1(n10882), .A2(n10881), .A3(n10880), .A4(n10879), .ZN(
        n10883) );
  NAND2_X1 U13810 ( .A1(n19356), .A2(n13240), .ZN(n10885) );
  OR2_X1 U13811 ( .A1(n11135), .A2(n10885), .ZN(n10979) );
  AOI22_X1 U13812 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n9980), .B1(
        n11020), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U13813 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n11021), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10889) );
  AOI22_X1 U13814 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10888) );
  AOI22_X1 U13815 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10887) );
  NAND4_X1 U13816 ( .A1(n10890), .A2(n10889), .A3(n10888), .A4(n10887), .ZN(
        n10896) );
  AOI22_X1 U13817 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13818 ( .A1(n11558), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11064), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13819 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n11022), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13820 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n11840), .ZN(n10891) );
  NAND4_X1 U13821 ( .A1(n10894), .A2(n10893), .A3(n10892), .A4(n10891), .ZN(
        n10895) );
  INV_X1 U13822 ( .A(n11099), .ZN(n11529) );
  NAND2_X1 U13823 ( .A1(n10979), .A2(n11529), .ZN(n10978) );
  AOI22_X1 U13824 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19641), .B1(
        n10992), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10901) );
  AOI22_X1 U13825 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n11010), .B1(
        n10956), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10900) );
  AOI22_X1 U13826 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10993), .B1(
        n10940), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10914) );
  AOI21_X1 U13827 ( .B1(n19797), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n10904), .ZN(n10913) );
  INV_X1 U13828 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10906) );
  INV_X1 U13829 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10905) );
  OAI22_X1 U13830 ( .A1(n10906), .A2(n10998), .B1(n10945), .B2(n10905), .ZN(
        n10910) );
  INV_X1 U13831 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10908) );
  INV_X1 U13832 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10907) );
  OAI22_X1 U13833 ( .A1(n10908), .A2(n10942), .B1(n10995), .B2(n10907), .ZN(
        n10909) );
  NOR2_X1 U13834 ( .A1(n10910), .A2(n10909), .ZN(n10912) );
  AOI22_X1 U13835 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n9980), .B1(
        n11020), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U13836 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n11021), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U13837 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13838 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11901), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10915) );
  NAND4_X1 U13839 ( .A1(n10918), .A2(n10917), .A3(n10916), .A4(n10915), .ZN(
        n10924) );
  AOI22_X1 U13840 ( .A1(n11558), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13841 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11022), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U13842 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U13843 ( .A1(n11571), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n11840), .ZN(n10919) );
  NAND4_X1 U13844 ( .A1(n10922), .A2(n10921), .A3(n10920), .A4(n10919), .ZN(
        n10923) );
  NOR2_X1 U13845 ( .A1(n10924), .A2(n10923), .ZN(n11541) );
  NAND2_X1 U13846 ( .A1(n11541), .A2(n19356), .ZN(n10925) );
  AOI22_X1 U13847 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n9980), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U13848 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11020), .B1(
        n11021), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10932) );
  AOI22_X1 U13849 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U13850 ( .A1(n11558), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10930) );
  NAND4_X1 U13851 ( .A1(n10933), .A2(n10932), .A3(n10931), .A4(n10930), .ZN(
        n10939) );
  AOI22_X1 U13852 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n11840), .ZN(n10937) );
  AOI22_X1 U13853 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11022), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U13854 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U13855 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11900), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10934) );
  NAND4_X1 U13856 ( .A1(n10937), .A2(n10936), .A3(n10935), .A4(n10934), .ZN(
        n10938) );
  AOI22_X1 U13857 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n10940), .B1(
        n10941), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U13858 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n10992), .B1(
        n10993), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10954) );
  INV_X1 U13859 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10944) );
  INV_X1 U13860 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10943) );
  OAI22_X1 U13861 ( .A1(n10944), .A2(n10942), .B1(n10998), .B2(n10943), .ZN(
        n10949) );
  INV_X1 U13862 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10947) );
  INV_X1 U13863 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10946) );
  OAI22_X1 U13864 ( .A1(n10947), .A2(n10945), .B1(n10995), .B2(n10946), .ZN(
        n10948) );
  NOR2_X1 U13865 ( .A1(n10949), .A2(n10948), .ZN(n10953) );
  INV_X1 U13866 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13705) );
  INV_X1 U13867 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10950) );
  INV_X1 U13868 ( .A(n10951), .ZN(n10952) );
  AOI22_X1 U13869 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n11010), .B1(
        n19641), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10961) );
  NAND2_X1 U13870 ( .A1(n19425), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10959) );
  NAND2_X1 U13871 ( .A1(n10957), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10958) );
  NAND2_X1 U13872 ( .A1(n10320), .A2(n10321), .ZN(n10973) );
  AOI22_X1 U13873 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11558), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U13874 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11840), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U13875 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U13876 ( .A1(n11064), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10962) );
  NAND4_X1 U13877 ( .A1(n10965), .A2(n10964), .A3(n10963), .A4(n10962), .ZN(
        n10971) );
  AOI22_X1 U13878 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11021), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U13879 ( .A1(n13809), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10968) );
  AOI22_X1 U13880 ( .A1(n10929), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U13881 ( .A1(n11022), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10966) );
  NAND4_X1 U13882 ( .A1(n10969), .A2(n10968), .A3(n10967), .A4(n10966), .ZN(
        n10970) );
  NAND2_X1 U13883 ( .A1(n11550), .A2(n19356), .ZN(n10972) );
  INV_X1 U13884 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16570) );
  NAND2_X1 U13885 ( .A1(n11174), .A2(n16570), .ZN(n16497) );
  OR3_X1 U13886 ( .A1(n13240), .A2(n13367), .A3(n11135), .ZN(n10977) );
  NOR2_X1 U13887 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13240), .ZN(
        n10976) );
  XOR2_X1 U13888 ( .A(n11135), .B(n10976), .Z(n13373) );
  NAND2_X1 U13889 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13373), .ZN(
        n13372) );
  NAND2_X1 U13890 ( .A1(n10977), .A2(n13372), .ZN(n10980) );
  XOR2_X1 U13891 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10980), .Z(
        n13341) );
  OAI21_X1 U13892 ( .B1(n10979), .B2(n11529), .A(n10978), .ZN(n13339) );
  NAND2_X1 U13893 ( .A1(n13341), .A2(n13339), .ZN(n10982) );
  NAND2_X1 U13894 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10980), .ZN(
        n10981) );
  NAND2_X1 U13895 ( .A1(n10982), .A2(n10981), .ZN(n10983) );
  XNOR2_X1 U13896 ( .A(n10983), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14012) );
  INV_X1 U13897 ( .A(n10983), .ZN(n10984) );
  INV_X1 U13898 ( .A(n11108), .ZN(n11547) );
  INV_X1 U13899 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16556) );
  NAND2_X1 U13900 ( .A1(n14187), .A2(n16556), .ZN(n10986) );
  INV_X1 U13901 ( .A(n14187), .ZN(n10987) );
  NAND2_X1 U13902 ( .A1(n10987), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10988) );
  INV_X1 U13903 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11023) );
  INV_X1 U13904 ( .A(n19425), .ZN(n19428) );
  INV_X1 U13905 ( .A(n10957), .ZN(n10990) );
  INV_X1 U13906 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10989) );
  INV_X1 U13907 ( .A(n10991), .ZN(n11015) );
  AOI22_X1 U13908 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10941), .B1(
        n10992), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U13909 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10993), .B1(
        n19641), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11008) );
  INV_X1 U13910 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10996) );
  INV_X1 U13911 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10994) );
  OAI22_X1 U13912 ( .A1(n10996), .A2(n10942), .B1(n10995), .B2(n10994), .ZN(
        n11001) );
  INV_X1 U13913 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10999) );
  INV_X1 U13914 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10997) );
  OAI22_X1 U13915 ( .A1(n10999), .A2(n10998), .B1(n10945), .B2(n10997), .ZN(
        n11000) );
  NOR2_X1 U13916 ( .A1(n11001), .A2(n11000), .ZN(n11007) );
  INV_X1 U13917 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11004) );
  INV_X1 U13918 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11002) );
  OAI22_X1 U13919 ( .A1(n11004), .A2(n19347), .B1(n11003), .B2(n11002), .ZN(
        n11005) );
  INV_X1 U13920 ( .A(n11005), .ZN(n11006) );
  NAND2_X1 U13921 ( .A1(n10940), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11014) );
  NAND2_X1 U13922 ( .A1(n19797), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11013) );
  NAND2_X1 U13923 ( .A1(n11010), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11012) );
  NAND2_X1 U13924 ( .A1(n10956), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11011) );
  NAND3_X1 U13925 ( .A1(n11015), .A2(n10319), .A3(n10328), .ZN(n11033) );
  AOI22_X1 U13926 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11558), .B1(
        n11057), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U13927 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n11840), .ZN(n11018) );
  AOI22_X1 U13928 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11072), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U13929 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11901), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11016) );
  NAND4_X1 U13930 ( .A1(n11019), .A2(n11018), .A3(n11017), .A4(n11016), .ZN(
        n11031) );
  AOI22_X1 U13931 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11020), .B1(
        n11021), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U13932 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n9980), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U13933 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11027) );
  INV_X1 U13934 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11024) );
  INV_X1 U13935 ( .A(n11022), .ZN(n11050) );
  INV_X1 U13936 ( .A(n11902), .ZN(n11052) );
  OAI22_X1 U13937 ( .A1(n11024), .A2(n11050), .B1(n11052), .B2(n11023), .ZN(
        n11025) );
  INV_X1 U13938 ( .A(n11025), .ZN(n11026) );
  NAND4_X1 U13939 ( .A1(n11029), .A2(n11028), .A3(n11027), .A4(n11026), .ZN(
        n11030) );
  NAND2_X1 U13940 ( .A1(n11551), .A2(n19356), .ZN(n11032) );
  INV_X1 U13941 ( .A(n11174), .ZN(n11035) );
  NAND2_X1 U13942 ( .A1(n11035), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11040) );
  NAND3_X1 U13943 ( .A1(n11041), .A2(n11178), .A3(n11040), .ZN(n11039) );
  INV_X1 U13944 ( .A(n11040), .ZN(n11037) );
  OAI211_X1 U13945 ( .C1(n11041), .C2(n11178), .A(n11039), .B(n11038), .ZN(
        n14290) );
  NAND2_X1 U13946 ( .A1(n14290), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14291) );
  NAND2_X1 U13947 ( .A1(n11041), .A2(n11040), .ZN(n11042) );
  NAND2_X1 U13948 ( .A1(n11042), .A2(n11178), .ZN(n11043) );
  INV_X1 U13949 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16543) );
  NAND2_X1 U13950 ( .A1(n11021), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11048) );
  NAND2_X1 U13951 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11047) );
  NAND2_X1 U13952 ( .A1(n9980), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11046) );
  NAND2_X1 U13953 ( .A1(n13809), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11045) );
  AND4_X1 U13954 ( .A1(n11048), .A2(n11047), .A3(n11046), .A4(n11045), .ZN(
        n11084) );
  NAND2_X1 U13955 ( .A1(n10929), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11056) );
  NAND2_X1 U13956 ( .A1(n10886), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11055) );
  INV_X1 U13957 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11049) );
  OR2_X1 U13958 ( .A1(n11050), .A2(n11049), .ZN(n11054) );
  INV_X1 U13959 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11051) );
  OR2_X1 U13960 ( .A1(n11052), .A2(n11051), .ZN(n11053) );
  INV_X1 U13961 ( .A(n11057), .ZN(n11059) );
  INV_X1 U13962 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11058) );
  OR2_X1 U13963 ( .A1(n11059), .A2(n11058), .ZN(n11068) );
  INV_X1 U13964 ( .A(n11558), .ZN(n11061) );
  INV_X1 U13965 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11060) );
  OR2_X1 U13966 ( .A1(n11061), .A2(n11060), .ZN(n11067) );
  INV_X1 U13967 ( .A(n11900), .ZN(n11063) );
  INV_X1 U13968 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11062) );
  OR2_X1 U13969 ( .A1(n11063), .A2(n11062), .ZN(n11066) );
  NAND2_X1 U13970 ( .A1(n11901), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11065) );
  INV_X1 U13971 ( .A(n11069), .ZN(n11071) );
  INV_X1 U13972 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11070) );
  OR2_X1 U13973 ( .A1(n11071), .A2(n11070), .ZN(n11080) );
  NAND2_X1 U13974 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11840), .ZN(
        n11079) );
  INV_X1 U13975 ( .A(n11072), .ZN(n11074) );
  INV_X1 U13976 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11073) );
  OR2_X1 U13977 ( .A1(n11074), .A2(n11073), .ZN(n11078) );
  INV_X1 U13978 ( .A(n11571), .ZN(n11076) );
  INV_X1 U13979 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11075) );
  OR2_X1 U13980 ( .A1(n11076), .A2(n11075), .ZN(n11077) );
  NAND4_X1 U13981 ( .A1(n11084), .A2(n11083), .A3(n11082), .A4(n11081), .ZN(
        n11185) );
  INV_X1 U13982 ( .A(n11185), .ZN(n11169) );
  NAND2_X1 U13983 ( .A1(n11044), .A2(n11169), .ZN(n11086) );
  NAND2_X1 U13984 ( .A1(n15970), .A2(n15972), .ZN(n15973) );
  INV_X1 U13985 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16545) );
  NAND2_X1 U13986 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16535) );
  INV_X1 U13987 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15962) );
  NOR2_X1 U13988 ( .A1(n16535), .A2(n15962), .ZN(n15917) );
  AND2_X1 U13989 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11090) );
  AND2_X1 U13990 ( .A1(n15917), .A2(n11090), .ZN(n15913) );
  INV_X1 U13991 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11243) );
  NAND3_X1 U13992 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15873) );
  INV_X1 U13993 ( .A(n15873), .ZN(n11091) );
  NAND2_X1 U13994 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n11091), .ZN(
        n11741) );
  NAND2_X1 U13995 ( .A1(n11093), .A2(n11092), .ZN(n15670) );
  NAND2_X1 U13996 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15853) );
  INV_X1 U13997 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15808) );
  INV_X1 U13998 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15793) );
  INV_X1 U13999 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15771) );
  NOR2_X2 U14000 ( .A1(n15582), .A2(n15771), .ZN(n15577) );
  XNOR2_X1 U14001 ( .A(n15577), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15766) );
  NAND2_X1 U14002 ( .A1(n20011), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11097) );
  NAND2_X1 U14003 ( .A1(n11097), .A2(n11096), .ZN(n11407) );
  NAND2_X1 U14004 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20020), .ZN(
        n11101) );
  NAND2_X1 U14005 ( .A1(n13802), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11106) );
  OAI21_X1 U14006 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13802), .A(
        n11106), .ZN(n11098) );
  XNOR2_X1 U14007 ( .A(n11105), .B(n11098), .ZN(n11123) );
  INV_X1 U14008 ( .A(n11123), .ZN(n11408) );
  MUX2_X1 U14009 ( .A(n11099), .B(n11408), .S(n11505), .Z(n11138) );
  INV_X1 U14010 ( .A(n11138), .ZN(n11103) );
  OAI21_X1 U14011 ( .B1(n9932), .B2(n20020), .A(n11101), .ZN(n11410) );
  INV_X1 U14012 ( .A(n11410), .ZN(n11100) );
  MUX2_X1 U14013 ( .A(n13240), .B(n11100), .S(n11505), .Z(n11147) );
  NAND2_X1 U14014 ( .A1(n11407), .A2(n11101), .ZN(n11125) );
  NAND2_X1 U14015 ( .A1(n11147), .A2(n11125), .ZN(n11102) );
  NAND2_X1 U14016 ( .A1(n11103), .A2(n11102), .ZN(n11112) );
  NAND2_X1 U14017 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20002), .ZN(
        n11104) );
  NAND2_X1 U14018 ( .A1(n11105), .A2(n11104), .ZN(n11107) );
  NAND2_X1 U14019 ( .A1(n11107), .A2(n11106), .ZN(n11110) );
  XNOR2_X1 U14020 ( .A(n13827), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11109) );
  OAI22_X1 U14021 ( .A1(n11110), .A2(n11109), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13827), .ZN(n11114) );
  NAND2_X1 U14022 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11119), .ZN(
        n11115) );
  OR2_X1 U14023 ( .A1(n11114), .A2(n11115), .ZN(n11419) );
  MUX2_X1 U14024 ( .A(n11108), .B(n11419), .S(n11505), .Z(n11422) );
  XNOR2_X1 U14025 ( .A(n11110), .B(n11109), .ZN(n11418) );
  NAND3_X1 U14026 ( .A1(n11112), .A2(n11422), .A3(n11111), .ZN(n11117) );
  INV_X1 U14027 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16171) );
  AND2_X1 U14028 ( .A1(n16171), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11113) );
  OR2_X1 U14029 ( .A1(n11114), .A2(n11113), .ZN(n11116) );
  NAND2_X1 U14030 ( .A1(n11116), .A2(n11115), .ZN(n11428) );
  NAND2_X1 U14031 ( .A1(n11117), .A2(n11428), .ZN(n20023) );
  AND2_X1 U14032 ( .A1(n14134), .A2(n19356), .ZN(n13197) );
  NAND2_X1 U14033 ( .A1(n20027), .A2(n13197), .ZN(n20030) );
  NAND2_X1 U14034 ( .A1(n9927), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11120) );
  INV_X1 U14035 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11119) );
  NAND2_X1 U14036 ( .A1(n11120), .A2(n11119), .ZN(n16089) );
  INV_X1 U14037 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n11121) );
  OAI21_X1 U14038 ( .B1(n11022), .B2(n16089), .A(n11121), .ZN(n11122) );
  NAND2_X1 U14039 ( .A1(n11122), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16572) );
  INV_X1 U14040 ( .A(n11419), .ZN(n11124) );
  OR3_X1 U14041 ( .A1(n11124), .A2(n11123), .A3(n11418), .ZN(n11129) );
  AND2_X1 U14042 ( .A1(n11126), .A2(n11125), .ZN(n11411) );
  INV_X1 U14043 ( .A(n11129), .ZN(n11127) );
  NAND2_X1 U14044 ( .A1(n11411), .A2(n11127), .ZN(n11128) );
  OAI211_X1 U14045 ( .C1(n11410), .C2(n11129), .A(n13828), .B(n14396), .ZN(
        n11130) );
  AND2_X1 U14046 ( .A1(n16572), .A2(n11130), .ZN(n20025) );
  INV_X1 U14047 ( .A(n20025), .ZN(n11131) );
  NAND3_X1 U14048 ( .A1(n20027), .A2(n13179), .A3(n11131), .ZN(n11132) );
  OAI21_X1 U14049 ( .B1(n20023), .B2(n20030), .A(n11132), .ZN(n11500) );
  NAND2_X1 U14050 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14396), .ZN(n19898) );
  INV_X1 U14051 ( .A(n19898), .ZN(n11133) );
  NAND2_X1 U14052 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11133), .ZN(n16580) );
  INV_X1 U14053 ( .A(n16580), .ZN(n13362) );
  AND2_X1 U14054 ( .A1(n14134), .A2(n13362), .ZN(n13178) );
  NAND2_X1 U14055 ( .A1(n11500), .A2(n13178), .ZN(n13253) );
  INV_X1 U14056 ( .A(n13253), .ZN(n11134) );
  INV_X1 U14057 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14273) );
  NAND3_X1 U14058 ( .A1(n11277), .A2(n14273), .A3(n11136), .ZN(n11137) );
  NAND2_X1 U14059 ( .A1(n11525), .A2(n11137), .ZN(n11151) );
  MUX2_X1 U14060 ( .A(n11138), .B(n10787), .S(n14575), .Z(n11150) );
  NAND2_X1 U14061 ( .A1(n11151), .A2(n11150), .ZN(n11141) );
  INV_X1 U14062 ( .A(n11155), .ZN(n11143) );
  NAND2_X1 U14063 ( .A1(n11141), .A2(n11140), .ZN(n11142) );
  NAND2_X1 U14064 ( .A1(n11143), .A2(n11142), .ZN(n14150) );
  INV_X1 U14065 ( .A(n11151), .ZN(n11146) );
  AND2_X1 U14066 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11144) );
  NAND2_X1 U14067 ( .A1(n14575), .A2(n11144), .ZN(n11145) );
  NAND2_X1 U14068 ( .A1(n11146), .A2(n11145), .ZN(n14271) );
  MUX2_X1 U14069 ( .A(n11147), .B(P2_EBX_REG_0__SCAN_IN), .S(n14575), .Z(
        n19216) );
  NAND2_X1 U14070 ( .A1(n19216), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13368) );
  OAI21_X1 U14071 ( .B1(n14271), .B2(n14394), .A(n13368), .ZN(n11149) );
  NAND2_X1 U14072 ( .A1(n14271), .A2(n14394), .ZN(n11148) );
  AND2_X1 U14073 ( .A1(n11149), .A2(n11148), .ZN(n13345) );
  XNOR2_X1 U14074 ( .A(n11151), .B(n11150), .ZN(n14260) );
  XNOR2_X1 U14075 ( .A(n14260), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13346) );
  NAND2_X1 U14076 ( .A1(n13345), .A2(n13346), .ZN(n13388) );
  INV_X1 U14077 ( .A(n14260), .ZN(n11152) );
  NAND2_X1 U14078 ( .A1(n11152), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11153) );
  NAND2_X1 U14079 ( .A1(n13388), .A2(n11153), .ZN(n14009) );
  INV_X1 U14080 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19196) );
  MUX2_X1 U14081 ( .A(n11422), .B(n19196), .S(n14575), .Z(n11154) );
  OR2_X1 U14082 ( .A1(n11155), .A2(n11154), .ZN(n11156) );
  NAND2_X1 U14083 ( .A1(n11161), .A2(n11156), .ZN(n19197) );
  XNOR2_X1 U14084 ( .A(n19197), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14190) );
  INV_X1 U14085 ( .A(n19197), .ZN(n11157) );
  NAND2_X1 U14086 ( .A1(n11157), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11158) );
  MUX2_X1 U14087 ( .A(n11550), .B(P2_EBX_REG_5__SCAN_IN), .S(n14575), .Z(
        n11160) );
  NAND2_X1 U14088 ( .A1(n11161), .A2(n11160), .ZN(n11162) );
  NAND2_X1 U14089 ( .A1(n11180), .A2(n11162), .ZN(n14109) );
  AND2_X1 U14090 ( .A1(n14109), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11166) );
  INV_X1 U14091 ( .A(n11166), .ZN(n11164) );
  NOR2_X1 U14092 ( .A1(n14578), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11167) );
  INV_X1 U14093 ( .A(n11167), .ZN(n11163) );
  MUX2_X1 U14094 ( .A(n11164), .B(n11163), .S(n11165), .Z(n11173) );
  MUX2_X1 U14095 ( .A(n11167), .B(n11166), .S(n11165), .Z(n11168) );
  NAND2_X1 U14096 ( .A1(n11159), .A2(n11168), .ZN(n11172) );
  OAI21_X1 U14097 ( .B1(n11169), .B2(n16570), .A(n14109), .ZN(n11170) );
  OAI21_X1 U14098 ( .B1(n14109), .B2(n16570), .A(n11170), .ZN(n11171) );
  OAI211_X1 U14099 ( .C1(n11159), .C2(n11173), .A(n11172), .B(n11171), .ZN(
        n16501) );
  NAND2_X1 U14100 ( .A1(n16500), .A2(n16501), .ZN(n11177) );
  OAI21_X1 U14101 ( .B1(n11174), .B2(n14578), .A(n14109), .ZN(n11175) );
  NAND2_X1 U14102 ( .A1(n11175), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11176) );
  NAND2_X1 U14103 ( .A1(n11177), .A2(n11176), .ZN(n14292) );
  MUX2_X1 U14104 ( .A(n11551), .B(P2_EBX_REG_6__SCAN_IN), .S(n14575), .Z(
        n11179) );
  AND2_X1 U14105 ( .A1(n11180), .A2(n11179), .ZN(n11181) );
  OR2_X1 U14106 ( .A1(n11181), .A2(n11190), .ZN(n19183) );
  NAND2_X1 U14107 ( .A1(n11182), .A2(n19183), .ZN(n11183) );
  INV_X1 U14108 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14295) );
  NAND2_X1 U14109 ( .A1(n11183), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11184) );
  INV_X1 U14110 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11315) );
  MUX2_X1 U14111 ( .A(n11185), .B(n11315), .S(n14575), .Z(n11189) );
  NAND2_X1 U14112 ( .A1(n14575), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11186) );
  INV_X1 U14113 ( .A(n11197), .ZN(n11188) );
  OR2_X1 U14114 ( .A1(n9991), .A2(n11186), .ZN(n11187) );
  NAND2_X1 U14115 ( .A1(n11188), .A2(n11187), .ZN(n19170) );
  NOR2_X1 U14116 ( .A1(n19170), .A2(n11169), .ZN(n11194) );
  NAND2_X1 U14117 ( .A1(n11194), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15735) );
  NOR2_X1 U14118 ( .A1(n11190), .A2(n11189), .ZN(n11191) );
  OR2_X1 U14119 ( .A1(n9991), .A2(n11191), .ZN(n11196) );
  INV_X1 U14120 ( .A(n11196), .ZN(n14068) );
  NAND2_X1 U14121 ( .A1(n14068), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15968) );
  NAND2_X1 U14122 ( .A1(n14575), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11192) );
  INV_X1 U14123 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11324) );
  MUX2_X1 U14124 ( .A(n11192), .B(P2_EBX_REG_10__SCAN_IN), .S(n11202), .Z(
        n11193) );
  NAND2_X1 U14125 ( .A1(n11193), .A2(n11283), .ZN(n19156) );
  OR2_X1 U14126 ( .A1(n19156), .A2(n11169), .ZN(n11209) );
  INV_X1 U14127 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15946) );
  NAND2_X1 U14128 ( .A1(n11209), .A2(n15946), .ZN(n16464) );
  INV_X1 U14129 ( .A(n11194), .ZN(n11195) );
  NAND2_X1 U14130 ( .A1(n11195), .A2(n16545), .ZN(n15734) );
  NAND2_X1 U14131 ( .A1(n11196), .A2(n16543), .ZN(n15967) );
  AND2_X1 U14132 ( .A1(n15734), .A2(n15967), .ZN(n15938) );
  NAND2_X1 U14133 ( .A1(n14575), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11198) );
  MUX2_X1 U14134 ( .A(n11198), .B(n11277), .S(n11197), .Z(n11200) );
  INV_X1 U14135 ( .A(n11202), .ZN(n11199) );
  NAND2_X1 U14136 ( .A1(n11200), .A2(n11199), .ZN(n14120) );
  OR2_X1 U14137 ( .A1(n14120), .A2(n11169), .ZN(n11201) );
  NAND2_X1 U14138 ( .A1(n11201), .A2(n15962), .ZN(n15939) );
  INV_X1 U14139 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13739) );
  AND3_X1 U14140 ( .A1(n11277), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n11203), .ZN(
        n11204) );
  OR2_X1 U14141 ( .A1(n11211), .A2(n11204), .ZN(n14088) );
  OR2_X1 U14142 ( .A1(n14088), .A2(n11169), .ZN(n11205) );
  INV_X1 U14143 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U14144 ( .A1(n11205), .A2(n11332), .ZN(n16462) );
  AND4_X1 U14145 ( .A1(n16464), .A2(n15938), .A3(n15939), .A4(n16462), .ZN(
        n11206) );
  NAND2_X1 U14146 ( .A1(n14578), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11207) );
  OR2_X1 U14147 ( .A1(n14088), .A2(n11207), .ZN(n16461) );
  NAND2_X1 U14148 ( .A1(n14578), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11208) );
  OR2_X1 U14149 ( .A1(n14120), .A2(n11208), .ZN(n15940) );
  OR2_X1 U14150 ( .A1(n15946), .A2(n11209), .ZN(n15941) );
  NAND2_X1 U14151 ( .A1(n15940), .A2(n15941), .ZN(n16463) );
  INV_X1 U14152 ( .A(n16463), .ZN(n11210) );
  AND2_X1 U14153 ( .A1(n16461), .A2(n11210), .ZN(n15718) );
  NAND2_X1 U14154 ( .A1(n14575), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11212) );
  INV_X1 U14155 ( .A(n11212), .ZN(n11214) );
  NAND2_X1 U14156 ( .A1(n11214), .A2(n11213), .ZN(n11215) );
  NAND2_X1 U14157 ( .A1(n11235), .A2(n11215), .ZN(n19144) );
  INV_X1 U14158 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15929) );
  OR3_X1 U14159 ( .A1(n19144), .A2(n11169), .A3(n15929), .ZN(n15720) );
  AND2_X1 U14160 ( .A1(n15718), .A2(n15720), .ZN(n15642) );
  OR2_X1 U14161 ( .A1(n19144), .A2(n11169), .ZN(n11216) );
  NAND2_X1 U14162 ( .A1(n11216), .A2(n15929), .ZN(n15721) );
  AND2_X1 U14163 ( .A1(n14575), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11234) );
  INV_X1 U14164 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11343) );
  INV_X1 U14165 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n14065) );
  NAND2_X1 U14166 ( .A1(n11343), .A2(n14065), .ZN(n11218) );
  AND2_X1 U14167 ( .A1(n14575), .A2(n11218), .ZN(n11219) );
  INV_X1 U14168 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11349) );
  INV_X1 U14169 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11220) );
  NAND2_X1 U14170 ( .A1(n11349), .A2(n11220), .ZN(n11221) );
  AND2_X1 U14171 ( .A1(n14575), .A2(n11221), .ZN(n11222) );
  NAND2_X1 U14172 ( .A1(n14575), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11224) );
  AND2_X2 U14173 ( .A1(n11223), .A2(n11224), .ZN(n11249) );
  NOR2_X1 U14174 ( .A1(n11223), .A2(n11224), .ZN(n11225) );
  OR2_X1 U14175 ( .A1(n11249), .A2(n11225), .ZN(n19082) );
  NOR2_X1 U14176 ( .A1(n19082), .A2(n11169), .ZN(n11251) );
  INV_X1 U14177 ( .A(n11251), .ZN(n11226) );
  INV_X1 U14178 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15876) );
  NAND2_X1 U14179 ( .A1(n11226), .A2(n15876), .ZN(n15692) );
  NAND2_X1 U14180 ( .A1(n14575), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11227) );
  MUX2_X1 U14181 ( .A(P2_EBX_REG_16__SCAN_IN), .B(n11227), .S(n9978), .Z(
        n11228) );
  NAND2_X1 U14182 ( .A1(n11228), .A2(n11283), .ZN(n19109) );
  NOR2_X1 U14183 ( .A1(n19109), .A2(n11169), .ZN(n11229) );
  INV_X1 U14184 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15909) );
  XNOR2_X1 U14185 ( .A(n11229), .B(n15909), .ZN(n15710) );
  INV_X1 U14186 ( .A(n11223), .ZN(n11231) );
  OAI211_X1 U14187 ( .C1(n9978), .C2(P2_EBX_REG_16__SCAN_IN), .A(
        P2_EBX_REG_17__SCAN_IN), .B(n14575), .ZN(n11230) );
  INV_X1 U14188 ( .A(n19097), .ZN(n11232) );
  INV_X1 U14189 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15898) );
  OAI21_X1 U14190 ( .B1(n11232), .B2(n11169), .A(n15898), .ZN(n15652) );
  OR2_X1 U14191 ( .A1(n11238), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11240) );
  NAND3_X1 U14192 ( .A1(n11240), .A2(n14575), .A3(P2_EBX_REG_15__SCAN_IN), 
        .ZN(n11233) );
  AND2_X1 U14193 ( .A1(n11233), .A2(n9978), .ZN(n11257) );
  INV_X1 U14194 ( .A(n11257), .ZN(n19126) );
  INV_X1 U14195 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16513) );
  OAI21_X1 U14196 ( .B1(n19126), .B2(n11169), .A(n16513), .ZN(n16437) );
  INV_X1 U14197 ( .A(n15853), .ZN(n11721) );
  XNOR2_X1 U14198 ( .A(n11235), .B(n11234), .ZN(n11252) );
  INV_X1 U14199 ( .A(n11252), .ZN(n13187) );
  NAND2_X1 U14200 ( .A1(n13187), .A2(n14578), .ZN(n11236) );
  INV_X1 U14201 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11338) );
  NAND2_X1 U14202 ( .A1(n11236), .A2(n11338), .ZN(n16454) );
  AND4_X1 U14203 ( .A1(n16437), .A2(n11721), .A3(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n16454), .ZN(n11237) );
  AND2_X1 U14204 ( .A1(n15652), .A2(n11237), .ZN(n11245) );
  NAND2_X1 U14205 ( .A1(n14575), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11239) );
  MUX2_X1 U14206 ( .A(n11277), .B(n11239), .S(n11238), .Z(n11241) );
  NAND2_X1 U14207 ( .A1(n11241), .A2(n11240), .ZN(n19136) );
  INV_X1 U14208 ( .A(n19136), .ZN(n11242) );
  NAND2_X1 U14209 ( .A1(n11242), .A2(n14578), .ZN(n11244) );
  NAND2_X1 U14210 ( .A1(n11244), .A2(n11243), .ZN(n15911) );
  NAND4_X1 U14211 ( .A1(n15692), .A2(n15710), .A3(n11245), .A4(n15911), .ZN(
        n11264) );
  NAND2_X1 U14212 ( .A1(n14575), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11248) );
  INV_X1 U14213 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15491) );
  AND3_X1 U14214 ( .A1(n11246), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n14575), .ZN(
        n11247) );
  NOR2_X1 U14215 ( .A1(n11266), .A2(n11247), .ZN(n15411) );
  NAND3_X1 U14216 ( .A1(n15411), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n14578), .ZN(n11262) );
  NOR2_X1 U14217 ( .A1(n11249), .A2(n11248), .ZN(n11250) );
  OR2_X1 U14218 ( .A1(n11259), .A2(n11250), .ZN(n19073) );
  NOR2_X1 U14219 ( .A1(n19073), .A2(n11169), .ZN(n15653) );
  NAND2_X1 U14220 ( .A1(n15653), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15680) );
  NAND2_X1 U14221 ( .A1(n11251), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15693) );
  OR3_X1 U14222 ( .A1(n11252), .A2(n11169), .A3(n11338), .ZN(n16453) );
  AND2_X1 U14223 ( .A1(n14578), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11253) );
  NAND2_X1 U14224 ( .A1(n19097), .A2(n11253), .ZN(n15651) );
  AND4_X1 U14225 ( .A1(n15680), .A2(n15693), .A3(n16453), .A4(n15651), .ZN(
        n11261) );
  NAND2_X1 U14226 ( .A1(n14578), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11254) );
  NOR2_X1 U14227 ( .A1(n19109), .A2(n11254), .ZN(n15649) );
  NAND2_X1 U14228 ( .A1(n14578), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11255) );
  OR2_X1 U14229 ( .A1(n19136), .A2(n11255), .ZN(n16438) );
  AND2_X1 U14230 ( .A1(n14578), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11256) );
  NAND2_X1 U14231 ( .A1(n11257), .A2(n11256), .ZN(n16436) );
  NAND2_X1 U14232 ( .A1(n16438), .A2(n16436), .ZN(n15645) );
  NOR2_X1 U14233 ( .A1(n15649), .A2(n15645), .ZN(n11260) );
  AND2_X1 U14234 ( .A1(n14575), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11258) );
  XNOR2_X1 U14235 ( .A(n11259), .B(n11258), .ZN(n19062) );
  NAND2_X1 U14236 ( .A1(n19062), .A2(n14578), .ZN(n15656) );
  INV_X1 U14237 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15655) );
  OR2_X1 U14238 ( .A1(n15656), .A2(n15655), .ZN(n15658) );
  AND4_X1 U14239 ( .A1(n11262), .A2(n11261), .A3(n11260), .A4(n15658), .ZN(
        n11263) );
  NAND2_X1 U14240 ( .A1(n15411), .A2(n14578), .ZN(n15659) );
  NAND2_X1 U14241 ( .A1(n14575), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11265) );
  NAND2_X1 U14242 ( .A1(n11266), .A2(n11265), .ZN(n11276) );
  NAND3_X1 U14243 ( .A1(n11267), .A2(n14575), .A3(P2_EBX_REG_22__SCAN_IN), 
        .ZN(n11268) );
  NAND2_X1 U14244 ( .A1(n11276), .A2(n11268), .ZN(n16110) );
  NAND2_X1 U14245 ( .A1(n11269), .A2(n11094), .ZN(n15636) );
  INV_X1 U14246 ( .A(n11269), .ZN(n11270) );
  NAND2_X1 U14247 ( .A1(n11270), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15637) );
  NAND2_X1 U14248 ( .A1(n11271), .A2(n15637), .ZN(n15630) );
  AND2_X1 U14249 ( .A1(n14575), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11275) );
  INV_X1 U14250 ( .A(n11275), .ZN(n11272) );
  XNOR2_X1 U14251 ( .A(n11276), .B(n11272), .ZN(n15396) );
  NAND2_X1 U14252 ( .A1(n15396), .A2(n14578), .ZN(n11273) );
  XNOR2_X1 U14253 ( .A(n11273), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15629) );
  INV_X1 U14254 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15820) );
  OR2_X1 U14255 ( .A1(n11273), .A2(n15820), .ZN(n11274) );
  NAND3_X1 U14256 ( .A1(n10003), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n11277), 
        .ZN(n11278) );
  NAND2_X1 U14257 ( .A1(n11278), .A2(n11283), .ZN(n11279) );
  OR2_X1 U14258 ( .A1(n11279), .A2(n11282), .ZN(n15395) );
  INV_X1 U14259 ( .A(n11280), .ZN(n11281) );
  NAND2_X1 U14260 ( .A1(n11281), .A2(n15808), .ZN(n15616) );
  AOI21_X1 U14261 ( .B1(n16418), .B2(n14578), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15602) );
  INV_X1 U14262 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n11386) );
  NAND2_X1 U14263 ( .A1(n14575), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16407) );
  NAND2_X1 U14264 ( .A1(n14578), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11285) );
  INV_X1 U14265 ( .A(n11286), .ZN(n11287) );
  NAND2_X1 U14266 ( .A1(n11287), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11288) );
  INV_X1 U14267 ( .A(n11470), .ZN(n11291) );
  OAI21_X1 U14268 ( .B1(n11467), .B2(n11291), .A(n11290), .ZN(n11292) );
  AND2_X1 U14269 ( .A1(n14575), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11293) );
  INV_X1 U14270 ( .A(n11475), .ZN(n11294) );
  XOR2_X1 U14271 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n11468), .Z(
        n11295) );
  XNOR2_X1 U14272 ( .A(n11296), .B(n11295), .ZN(n15762) );
  OR2_X1 U14273 ( .A1(n9959), .A2(n16556), .ZN(n11303) );
  AOI22_X1 U14274 ( .A1(n11383), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11302) );
  NAND2_X1 U14275 ( .A1(n14585), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11301) );
  OR2_X1 U14276 ( .A1(n9960), .A2(n16570), .ZN(n11309) );
  INV_X1 U14277 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n11306) );
  NAND2_X1 U14278 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11305) );
  NAND2_X1 U14279 ( .A1(n11383), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11304) );
  OAI211_X1 U14280 ( .C1(n11400), .C2(n11306), .A(n11305), .B(n11304), .ZN(
        n11307) );
  INV_X1 U14281 ( .A(n11307), .ZN(n11308) );
  NAND2_X1 U14282 ( .A1(n11309), .A2(n11308), .ZN(n13636) );
  OR2_X1 U14283 ( .A1(n9960), .A2(n14295), .ZN(n11312) );
  AOI22_X1 U14284 ( .A1(n11383), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11311) );
  NAND2_X1 U14285 ( .A1(n14585), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11310) );
  OR2_X1 U14286 ( .A1(n9959), .A2(n16543), .ZN(n11318) );
  NAND2_X1 U14287 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11314) );
  NAND2_X1 U14288 ( .A1(n11383), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11313) );
  OAI211_X1 U14289 ( .C1(n11400), .C2(n11315), .A(n11314), .B(n11313), .ZN(
        n11316) );
  INV_X1 U14290 ( .A(n11316), .ZN(n11317) );
  NAND2_X1 U14291 ( .A1(n11318), .A2(n11317), .ZN(n13728) );
  OR2_X1 U14292 ( .A1(n9959), .A2(n16545), .ZN(n11321) );
  AOI22_X1 U14293 ( .A1(n11383), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11320) );
  NAND2_X1 U14294 ( .A1(n14585), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11319) );
  OR2_X1 U14295 ( .A1(n9959), .A2(n15962), .ZN(n11327) );
  NAND2_X1 U14296 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11323) );
  NAND2_X1 U14297 ( .A1(n11383), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11322) );
  OAI211_X1 U14298 ( .C1(n11400), .C2(n11324), .A(n11323), .B(n11322), .ZN(
        n11325) );
  INV_X1 U14299 ( .A(n11325), .ZN(n11326) );
  NAND2_X1 U14300 ( .A1(n11327), .A2(n11326), .ZN(n13722) );
  AOI22_X1 U14301 ( .A1(n11383), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11329) );
  NAND2_X1 U14302 ( .A1(n14585), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11328) );
  OAI211_X1 U14303 ( .C1(n9959), .C2(n15946), .A(n11329), .B(n11328), .ZN(
        n13735) );
  AOI22_X1 U14304 ( .A1(n11383), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11331) );
  NAND2_X1 U14305 ( .A1(n14585), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11330) );
  OAI211_X1 U14306 ( .C1(n9960), .C2(n11332), .A(n11331), .B(n11330), .ZN(
        n13936) );
  AOI22_X1 U14307 ( .A1(n11383), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11334) );
  NAND2_X1 U14308 ( .A1(n14585), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11333) );
  OAI211_X1 U14309 ( .C1(n9959), .C2(n15929), .A(n11334), .B(n11333), .ZN(
        n13941) );
  AOI22_X1 U14310 ( .A1(n11383), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11337) );
  NAND2_X1 U14311 ( .A1(n14585), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11336) );
  OAI211_X1 U14312 ( .C1(n9960), .C2(n11338), .A(n11337), .B(n11336), .ZN(
        n13189) );
  AOI22_X1 U14313 ( .A1(n11383), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11340) );
  NAND2_X1 U14314 ( .A1(n14585), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11339) );
  OAI211_X1 U14315 ( .C1(n9960), .C2(n11243), .A(n11340), .B(n11339), .ZN(
        n14061) );
  OR2_X1 U14316 ( .A1(n9959), .A2(n16513), .ZN(n11346) );
  NAND2_X1 U14317 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U14318 ( .A1(n11383), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11341) );
  OAI211_X1 U14319 ( .C1(n11400), .C2(n11343), .A(n11342), .B(n11341), .ZN(
        n11344) );
  INV_X1 U14320 ( .A(n11344), .ZN(n11345) );
  NAND2_X1 U14321 ( .A1(n11346), .A2(n11345), .ZN(n14178) );
  OR2_X1 U14322 ( .A1(n9960), .A2(n15909), .ZN(n11352) );
  NAND2_X1 U14323 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11348) );
  NAND2_X1 U14324 ( .A1(n11383), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11347) );
  OAI211_X1 U14325 ( .C1(n11400), .C2(n11349), .A(n11348), .B(n11347), .ZN(
        n11350) );
  INV_X1 U14326 ( .A(n11350), .ZN(n11351) );
  NAND2_X1 U14327 ( .A1(n11352), .A2(n11351), .ZN(n14213) );
  OR2_X1 U14328 ( .A1(n9959), .A2(n15898), .ZN(n11356) );
  AOI22_X1 U14329 ( .A1(n11383), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11354) );
  NAND2_X1 U14330 ( .A1(n14585), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11353) );
  AND2_X1 U14331 ( .A1(n11354), .A2(n11353), .ZN(n11355) );
  AOI22_X1 U14332 ( .A1(n11383), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11358) );
  NAND2_X1 U14333 ( .A1(n14585), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11357) );
  OAI211_X1 U14334 ( .C1(n9959), .C2(n15876), .A(n11358), .B(n11357), .ZN(
        n14388) );
  INV_X1 U14335 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11361) );
  NAND2_X1 U14336 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11360) );
  NAND2_X1 U14337 ( .A1(n11383), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11359) );
  OAI211_X1 U14338 ( .C1(n11400), .C2(n11361), .A(n11360), .B(n11359), .ZN(
        n11362) );
  AOI21_X1 U14339 ( .B1(n11402), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11362), .ZN(n14331) );
  NOR2_X2 U14340 ( .A1(n14330), .A2(n14331), .ZN(n14329) );
  NAND2_X1 U14341 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11364) );
  INV_X1 U14342 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19952) );
  OR2_X1 U14343 ( .A1(n11300), .A2(n19952), .ZN(n11363) );
  OAI211_X1 U14344 ( .C1(n11400), .C2(n15491), .A(n11364), .B(n11363), .ZN(
        n11365) );
  AOI21_X1 U14345 ( .B1(n11402), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11365), .ZN(n15487) );
  INV_X1 U14346 ( .A(n15487), .ZN(n11366) );
  INV_X1 U14347 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15662) );
  OR2_X1 U14348 ( .A1(n9960), .A2(n15662), .ZN(n11370) );
  AOI22_X1 U14349 ( .A1(n11383), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11368) );
  NAND2_X1 U14350 ( .A1(n14585), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11367) );
  AND2_X1 U14351 ( .A1(n11368), .A2(n11367), .ZN(n11369) );
  NAND2_X1 U14352 ( .A1(n11370), .A2(n11369), .ZN(n15414) );
  AOI22_X1 U14353 ( .A1(n11383), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11372) );
  NAND2_X1 U14354 ( .A1(n14585), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11371) );
  OAI211_X1 U14355 ( .C1(n9959), .C2(n11094), .A(n11372), .B(n11371), .ZN(
        n15475) );
  INV_X1 U14356 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11375) );
  NAND2_X1 U14357 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11374) );
  INV_X1 U14358 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19958) );
  OR2_X1 U14359 ( .A1(n11300), .A2(n19958), .ZN(n11373) );
  OAI211_X1 U14360 ( .C1(n11400), .C2(n11375), .A(n11374), .B(n11373), .ZN(
        n11376) );
  AOI21_X1 U14361 ( .B1(n11402), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11376), .ZN(n15401) );
  INV_X1 U14362 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11379) );
  NAND2_X1 U14363 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11378) );
  INV_X1 U14364 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19960) );
  OR2_X1 U14365 ( .A1(n11300), .A2(n19960), .ZN(n11377) );
  OAI211_X1 U14366 ( .C1(n11400), .C2(n11379), .A(n11378), .B(n11377), .ZN(
        n11380) );
  AOI21_X1 U14367 ( .B1(n11402), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11380), .ZN(n15386) );
  NAND2_X1 U14368 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11385) );
  NAND2_X1 U14369 ( .A1(n11383), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11384) );
  OAI211_X1 U14370 ( .C1(n11400), .C2(n11386), .A(n11385), .B(n11384), .ZN(
        n11387) );
  AOI21_X1 U14371 ( .B1(n11402), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11387), .ZN(n15458) );
  INV_X1 U14372 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11388) );
  OR2_X1 U14373 ( .A1(n9959), .A2(n11388), .ZN(n11392) );
  AOI22_X1 U14374 ( .A1(n11383), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11390) );
  NAND2_X1 U14375 ( .A1(n14585), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11389) );
  AND2_X1 U14376 ( .A1(n11390), .A2(n11389), .ZN(n11391) );
  NAND2_X1 U14377 ( .A1(n11392), .A2(n11391), .ZN(n13224) );
  INV_X1 U14378 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n11395) );
  NAND2_X1 U14379 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11394) );
  NAND2_X1 U14380 ( .A1(n10773), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11393) );
  OAI211_X1 U14381 ( .C1(n11400), .C2(n11395), .A(n11394), .B(n11393), .ZN(
        n11396) );
  AOI21_X1 U14382 ( .B1(n11402), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11396), .ZN(n15444) );
  INV_X1 U14383 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n11399) );
  NAND2_X1 U14384 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11398) );
  INV_X1 U14385 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19968) );
  OR2_X1 U14386 ( .A1(n11300), .A2(n19968), .ZN(n11397) );
  OAI211_X1 U14387 ( .C1(n11400), .C2(n11399), .A(n11398), .B(n11397), .ZN(
        n11401) );
  AOI21_X1 U14388 ( .B1(n11402), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11401), .ZN(n11403) );
  AND2_X1 U14389 ( .A1(n15446), .A2(n11403), .ZN(n11404) );
  INV_X1 U14390 ( .A(n16398), .ZN(n11440) );
  NOR2_X2 U14391 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19990) );
  INV_X1 U14392 ( .A(n19990), .ZN(n19599) );
  INV_X1 U14393 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19629) );
  NOR2_X1 U14394 ( .A1(n19599), .A2(n19629), .ZN(n20004) );
  NAND2_X1 U14395 ( .A1(n13179), .A2(n11405), .ZN(n11406) );
  MUX2_X1 U14396 ( .A(n11406), .B(n11505), .S(n11408), .Z(n11417) );
  OAI21_X1 U14397 ( .B1(n11410), .B2(n11407), .A(n20026), .ZN(n11415) );
  NAND2_X1 U14398 ( .A1(n11409), .A2(n11408), .ZN(n11414) );
  NAND2_X1 U14399 ( .A1(n11513), .A2(n11410), .ZN(n11412) );
  NAND3_X1 U14400 ( .A1(n11412), .A2(n20035), .A3(n11411), .ZN(n11413) );
  NAND3_X1 U14401 ( .A1(n11415), .A2(n11414), .A3(n11413), .ZN(n11416) );
  NAND2_X1 U14402 ( .A1(n11417), .A2(n11416), .ZN(n11421) );
  INV_X1 U14403 ( .A(n11418), .ZN(n11423) );
  NAND3_X1 U14404 ( .A1(n11421), .A2(n11423), .A3(n11419), .ZN(n11420) );
  NAND2_X1 U14405 ( .A1(n11420), .A2(n20026), .ZN(n11426) );
  INV_X1 U14406 ( .A(n11421), .ZN(n11424) );
  NAND3_X1 U14407 ( .A1(n11424), .A2(n11423), .A3(n11422), .ZN(n11425) );
  NAND3_X1 U14408 ( .A1(n11426), .A2(n11425), .A3(n11428), .ZN(n11427) );
  MUX2_X1 U14409 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11427), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11481) );
  INV_X1 U14410 ( .A(n11428), .ZN(n11429) );
  NAND2_X1 U14411 ( .A1(n11429), .A2(n13332), .ZN(n11430) );
  OAI21_X1 U14412 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n19032), .ZN(n20038) );
  INV_X1 U14413 ( .A(n20038), .ZN(n11431) );
  NAND2_X1 U14414 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n13851) );
  NAND2_X1 U14415 ( .A1(n11431), .A2(n13851), .ZN(n11432) );
  NOR2_X1 U14416 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19033) );
  OR2_X1 U14417 ( .A1(n19990), .A2(n19033), .ZN(n20016) );
  NAND2_X1 U14418 ( .A1(n20016), .A2(n19032), .ZN(n11433) );
  INV_X1 U14419 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11437) );
  NAND2_X1 U14420 ( .A1(n19032), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11766) );
  NAND2_X1 U14421 ( .A1(n19629), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11434) );
  NAND2_X1 U14422 ( .A1(n11766), .A2(n11434), .ZN(n13411) );
  INV_X1 U14423 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14015) );
  INV_X1 U14424 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16485) );
  INV_X1 U14425 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16472) );
  INV_X1 U14426 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16459) );
  INV_X1 U14427 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16445) );
  INV_X1 U14428 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15705) );
  INV_X1 U14429 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n13211) );
  INV_X1 U14430 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15663) );
  INV_X1 U14431 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15608) );
  INV_X1 U14432 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16410) );
  INV_X1 U14433 ( .A(n15353), .ZN(n11435) );
  AOI21_X1 U14434 ( .B1(n11437), .B2(n15356), .A(n11435), .ZN(n16394) );
  NAND2_X1 U14435 ( .A1(n16496), .A2(n16394), .ZN(n11436) );
  AND2_X1 U14436 ( .A1(n13846), .A2(n19990), .ZN(n19328) );
  NAND2_X1 U14437 ( .A1(n19328), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15758) );
  OAI211_X1 U14438 ( .C1(n16506), .C2(n11437), .A(n11436), .B(n15758), .ZN(
        n11438) );
  INV_X1 U14439 ( .A(n11438), .ZN(n11439) );
  OAI21_X1 U14440 ( .B1(n15762), .B2(n19333), .A(n11442), .ZN(n11443) );
  INV_X1 U14441 ( .A(n11443), .ZN(n11444) );
  OAI21_X1 U14442 ( .B1(n15766), .B2(n19332), .A(n11444), .ZN(P2_U2986) );
  NAND2_X1 U14443 ( .A1(n17826), .A2(n11445), .ZN(n11448) );
  AOI21_X1 U14444 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11446), .A(
        n17826), .ZN(n11447) );
  NAND2_X1 U14445 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17826), .ZN(
        n11455) );
  NAND2_X1 U14446 ( .A1(n11449), .A2(n11448), .ZN(n11453) );
  INV_X1 U14447 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18974) );
  NAND2_X1 U14448 ( .A1(n18974), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11452) );
  OAI22_X1 U14449 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17826), .B1(
        n11455), .B2(n16164), .ZN(n11450) );
  AOI21_X1 U14450 ( .B1(n11453), .B2(n11452), .A(n11451), .ZN(n11454) );
  AOI21_X1 U14451 ( .B1(n11456), .B2(n11455), .A(n11454), .ZN(n13117) );
  NAND2_X1 U14452 ( .A1(n13117), .A2(n17926), .ZN(n11466) );
  NAND2_X1 U14453 ( .A1(n16591), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11457) );
  INV_X1 U14454 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16749) );
  XNOR2_X2 U14455 ( .A(n11457), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16960) );
  INV_X1 U14456 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18948) );
  NOR2_X1 U14457 ( .A1(n18948), .A2(n18345), .ZN(n13130) );
  XNOR2_X1 U14458 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11459) );
  OAI22_X1 U14459 ( .A1(n11460), .A2(n11459), .B1(n11458), .B2(n16749), .ZN(
        n11461) );
  AOI211_X1 U14460 ( .C1(n17890), .C2(n16960), .A(n13130), .B(n11461), .ZN(
        n11465) );
  NAND2_X1 U14461 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16589), .ZN(
        n11462) );
  XOR2_X1 U14462 ( .A(n11462), .B(n18974), .Z(n13136) );
  NAND2_X1 U14463 ( .A1(n13136), .A2(n17943), .ZN(n11464) );
  NAND2_X1 U14464 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16585), .ZN(
        n11463) );
  NOR2_X1 U14465 ( .A1(n16094), .A2(n18045), .ZN(n16605) );
  NOR3_X1 U14466 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n9871), .A3(
        n16164), .ZN(n13132) );
  AOI22_X1 U14467 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n11463), .B1(
        n16605), .B2(n13132), .ZN(n13134) );
  AOI21_X1 U14468 ( .B1(n11467), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11468), .ZN(n11472) );
  INV_X1 U14469 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15759) );
  OAI21_X1 U14470 ( .B1(n11469), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11468), .ZN(n11471) );
  NAND2_X1 U14471 ( .A1(n14575), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11474) );
  XNOR2_X1 U14472 ( .A(n11475), .B(n11474), .ZN(n16379) );
  INV_X1 U14473 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11728) );
  OAI21_X1 U14474 ( .B1(n16379), .B2(n11169), .A(n11728), .ZN(n15573) );
  NAND2_X1 U14475 ( .A1(n15575), .A2(n15573), .ZN(n14572) );
  INV_X1 U14476 ( .A(n16379), .ZN(n11473) );
  NAND3_X1 U14477 ( .A1(n11473), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14578), .ZN(n15574) );
  NAND2_X1 U14478 ( .A1(n14572), .A2(n15574), .ZN(n11480) );
  NAND2_X1 U14479 ( .A1(n11475), .A2(n11474), .ZN(n14574) );
  NAND2_X1 U14480 ( .A1(n14575), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11476) );
  XNOR2_X1 U14481 ( .A(n14574), .B(n11476), .ZN(n15376) );
  AOI21_X1 U14482 ( .B1(n15376), .B2(n14578), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14571) );
  INV_X1 U14483 ( .A(n14571), .ZN(n11478) );
  AND2_X1 U14484 ( .A1(n14578), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11477) );
  NAND2_X1 U14485 ( .A1(n15376), .A2(n11477), .ZN(n14570) );
  NAND2_X1 U14486 ( .A1(n11478), .A2(n14570), .ZN(n11479) );
  XNOR2_X1 U14487 ( .A(n11480), .B(n11479), .ZN(n11761) );
  NAND2_X1 U14488 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20046) );
  INV_X1 U14489 ( .A(n20046), .ZN(n20040) );
  INV_X1 U14490 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19900) );
  NAND2_X1 U14491 ( .A1(n19900), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20051) );
  NAND2_X2 U14492 ( .A1(n20050), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19972) );
  OR2_X1 U14493 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19910) );
  NAND3_X1 U14494 ( .A1(n19900), .A2(n19972), .A3(n19910), .ZN(n19906) );
  NOR2_X1 U14495 ( .A1(n20040), .A2(n19906), .ZN(n13250) );
  NAND2_X1 U14496 ( .A1(n9827), .A2(n13250), .ZN(n11503) );
  NAND2_X1 U14497 ( .A1(n13833), .A2(n13179), .ZN(n13794) );
  AOI21_X1 U14498 ( .B1(n11481), .B2(n20035), .A(n19373), .ZN(n11482) );
  NAND2_X1 U14499 ( .A1(n13794), .A2(n11482), .ZN(n11502) );
  OAI21_X1 U14500 ( .B1(n12066), .B2(n19373), .A(n19361), .ZN(n11485) );
  NAND2_X1 U14501 ( .A1(n11484), .A2(n11485), .ZN(n11489) );
  NAND2_X1 U14502 ( .A1(n11494), .A2(n19356), .ZN(n11698) );
  NAND2_X1 U14503 ( .A1(n11698), .A2(n20035), .ZN(n11486) );
  NAND2_X1 U14504 ( .A1(n11486), .A2(n13364), .ZN(n11487) );
  AOI21_X1 U14505 ( .B1(n11487), .B2(n19361), .A(n10729), .ZN(n11488) );
  AND2_X1 U14506 ( .A1(n11489), .A2(n11488), .ZN(n11701) );
  NAND3_X1 U14507 ( .A1(n11491), .A2(n13828), .A3(n13250), .ZN(n11493) );
  NAND2_X1 U14508 ( .A1(n11490), .A2(n13364), .ZN(n11492) );
  NAND2_X1 U14509 ( .A1(n11492), .A2(n13197), .ZN(n11713) );
  OAI211_X1 U14510 ( .C1(n11490), .C2(n11494), .A(n11493), .B(n11713), .ZN(
        n11495) );
  INV_X1 U14511 ( .A(n11495), .ZN(n11496) );
  AND2_X1 U14512 ( .A1(n11701), .A2(n11496), .ZN(n13799) );
  MUX2_X1 U14513 ( .A(n11491), .B(n9827), .S(n19356), .Z(n11497) );
  NAND3_X1 U14514 ( .A1(n11497), .A2(n13828), .A3(n20046), .ZN(n11498) );
  NAND2_X1 U14515 ( .A1(n13799), .A2(n11498), .ZN(n11499) );
  NOR2_X1 U14516 ( .A1(n11500), .A2(n11499), .ZN(n11501) );
  OAI211_X1 U14517 ( .C1(n11503), .C2(n13794), .A(n11502), .B(n11501), .ZN(
        n11504) );
  NOR2_X1 U14518 ( .A1(n13838), .A2(n11505), .ZN(n11506) );
  NAND2_X1 U14519 ( .A1(n11753), .A2(n11506), .ZN(n16552) );
  INV_X1 U14520 ( .A(n13240), .ZN(n13239) );
  NOR2_X1 U14521 ( .A1(n13364), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11517) );
  AND2_X1 U14522 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11509) );
  NOR2_X1 U14523 ( .A1(n11517), .A2(n11509), .ZN(n11510) );
  NAND2_X1 U14524 ( .A1(n12066), .A2(n11538), .ZN(n11530) );
  OAI211_X1 U14525 ( .C1(n13239), .C2(n11661), .A(n11510), .B(n11530), .ZN(
        n13238) );
  AND2_X1 U14526 ( .A1(n14575), .A2(n13364), .ZN(n12067) );
  NAND2_X1 U14527 ( .A1(n9826), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11516) );
  NAND2_X1 U14528 ( .A1(n11511), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11512) );
  OAI211_X1 U14529 ( .C1(n11513), .C2(n13367), .A(n11512), .B(n20012), .ZN(
        n11514) );
  INV_X1 U14530 ( .A(n11514), .ZN(n11515) );
  NAND2_X1 U14531 ( .A1(n11516), .A2(n11515), .ZN(n13237) );
  NAND2_X1 U14532 ( .A1(n13238), .A2(n13237), .ZN(n11526) );
  NAND2_X1 U14533 ( .A1(n9826), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14534 ( .A1(n11690), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11538), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11518) );
  XNOR2_X1 U14535 ( .A(n11526), .B(n11527), .ZN(n13374) );
  INV_X1 U14536 ( .A(n11520), .ZN(n11524) );
  INV_X1 U14537 ( .A(n12066), .ZN(n11521) );
  NAND2_X1 U14538 ( .A1(n11521), .A2(n13364), .ZN(n11522) );
  MUX2_X1 U14539 ( .A(n11522), .B(n20011), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11523) );
  OAI21_X1 U14540 ( .B1(n11525), .B2(n11524), .A(n11523), .ZN(n13375) );
  NAND2_X1 U14541 ( .A1(n11527), .A2(n11526), .ZN(n11528) );
  NAND2_X1 U14542 ( .A1(n13377), .A2(n11528), .ZN(n11535) );
  OR2_X1 U14543 ( .A1(n11661), .A2(n11529), .ZN(n11531) );
  OAI211_X1 U14544 ( .C1(n20012), .C2(n20002), .A(n11531), .B(n11530), .ZN(
        n11534) );
  XNOR2_X1 U14545 ( .A(n11535), .B(n11534), .ZN(n13344) );
  NAND2_X1 U14546 ( .A1(n9948), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14547 ( .A1(n14593), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11538), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11532) );
  INV_X1 U14548 ( .A(n11534), .ZN(n11536) );
  NAND2_X1 U14549 ( .A1(n11536), .A2(n11535), .ZN(n11537) );
  NAND2_X1 U14550 ( .A1(n13342), .A2(n11537), .ZN(n14027) );
  NAND2_X1 U14551 ( .A1(n11668), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14552 ( .A1(n11538), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11540) );
  NAND2_X1 U14553 ( .A1(n14593), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11539) );
  AND2_X1 U14554 ( .A1(n11540), .A2(n11539), .ZN(n11543) );
  OR2_X1 U14555 ( .A1(n11661), .A2(n11541), .ZN(n11542) );
  NAND2_X1 U14556 ( .A1(n9948), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14557 ( .A1(n14593), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11538), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11545) );
  OAI211_X1 U14558 ( .C1(n11661), .C2(n11547), .A(n11546), .B(n11545), .ZN(
        n14194) );
  NAND2_X1 U14559 ( .A1(n9948), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14560 ( .A1(n14593), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11538), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11548) );
  OAI211_X1 U14561 ( .C1(n11661), .C2(n11550), .A(n11549), .B(n11548), .ZN(
        n14102) );
  OR2_X1 U14562 ( .A1(n11661), .A2(n11551), .ZN(n11552) );
  NAND2_X1 U14563 ( .A1(n11668), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14564 ( .A1(n14593), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11538), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11553) );
  NAND2_X1 U14565 ( .A1(n11554), .A2(n11553), .ZN(n13319) );
  OR2_X1 U14566 ( .A1(n11661), .A2(n11169), .ZN(n11555) );
  NAND2_X1 U14567 ( .A1(n11668), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14568 ( .A1(n14593), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11538), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14569 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11558), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14570 ( .A1(n11900), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11840), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14571 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U14572 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11559) );
  NAND4_X1 U14573 ( .A1(n11562), .A2(n11561), .A3(n11560), .A4(n11559), .ZN(
        n11568) );
  AOI22_X1 U14574 ( .A1(n11021), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14575 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14576 ( .A1(n10929), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14577 ( .A1(n11901), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11022), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11563) );
  NAND4_X1 U14578 ( .A1(n11566), .A2(n11565), .A3(n11564), .A4(n11563), .ZN(
        n11567) );
  INV_X1 U14579 ( .A(n11799), .ZN(n13714) );
  NAND2_X1 U14580 ( .A1(n11668), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14581 ( .A1(n14593), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11538), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11569) );
  OAI211_X1 U14582 ( .C1(n11661), .C2(n13714), .A(n11570), .B(n11569), .ZN(
        n13404) );
  NAND2_X1 U14583 ( .A1(n11668), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14584 ( .A1(n14593), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11538), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14585 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11558), .B1(
        n11057), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14586 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n11840), .ZN(n11574) );
  AOI22_X1 U14587 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11571), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14588 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11901), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11572) );
  NAND4_X1 U14589 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11582) );
  INV_X1 U14590 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14591 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11020), .B1(
        n11021), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14592 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n13809), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14593 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14594 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n11022), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11577) );
  NAND4_X1 U14595 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n11581) );
  NOR2_X1 U14596 ( .A1(n11582), .A2(n11581), .ZN(n13721) );
  OR2_X1 U14597 ( .A1(n11661), .A2(n13721), .ZN(n11583) );
  AOI22_X1 U14598 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11021), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14599 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11020), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14600 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14601 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11586) );
  NAND4_X1 U14602 ( .A1(n11589), .A2(n11588), .A3(n11587), .A4(n11586), .ZN(
        n11595) );
  AOI22_X1 U14603 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n11840), .ZN(n11593) );
  AOI22_X1 U14604 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n11022), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U14605 ( .A1(n11558), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11901), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U14606 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11900), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11590) );
  NAND4_X1 U14607 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n11594) );
  INV_X1 U14608 ( .A(n13733), .ZN(n11598) );
  NAND2_X1 U14609 ( .A1(n11668), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14610 ( .A1(n14593), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11596) );
  OAI211_X1 U14611 ( .C1(n11661), .C2(n11598), .A(n11597), .B(n11596), .ZN(
        n13499) );
  AOI22_X1 U14612 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11558), .B1(
        n11057), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14613 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n11840), .ZN(n11601) );
  AOI22_X1 U14614 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11571), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14615 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11901), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11599) );
  NAND4_X1 U14616 ( .A1(n11602), .A2(n11601), .A3(n11600), .A4(n11599), .ZN(
        n11608) );
  AOI22_X1 U14617 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11020), .B1(
        n11021), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U14618 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n13809), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14619 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14620 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n11022), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11603) );
  NAND4_X1 U14621 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11607) );
  NOR2_X1 U14622 ( .A1(n11608), .A2(n11607), .ZN(n13933) );
  NAND2_X1 U14623 ( .A1(n9948), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14624 ( .A1(n14593), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11609) );
  OAI211_X1 U14625 ( .C1(n11661), .C2(n13933), .A(n11610), .B(n11609), .ZN(
        n13628) );
  AND2_X2 U14626 ( .A1(n13498), .A2(n13628), .ZN(n13634) );
  AOI22_X1 U14627 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11021), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14628 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11020), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14629 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14630 ( .A1(n11558), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11022), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11611) );
  NAND4_X1 U14631 ( .A1(n11614), .A2(n11613), .A3(n11612), .A4(n11611), .ZN(
        n11620) );
  AOI22_X1 U14632 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11901), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14633 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14634 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14635 ( .A1(n11571), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n11840), .ZN(n11615) );
  NAND4_X1 U14636 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(
        n11619) );
  OR2_X1 U14637 ( .A1(n11620), .A2(n11619), .ZN(n13944) );
  INV_X1 U14638 ( .A(n13944), .ZN(n11804) );
  NAND2_X1 U14639 ( .A1(n11668), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14640 ( .A1(n14593), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11621) );
  OAI211_X1 U14641 ( .C1(n11661), .C2(n11804), .A(n11622), .B(n11621), .ZN(
        n13633) );
  NAND2_X1 U14643 ( .A1(n11668), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14644 ( .A1(n14593), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14645 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11558), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14646 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11840), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14647 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14648 ( .A1(n11064), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11623) );
  NAND4_X1 U14649 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11632) );
  AOI22_X1 U14650 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11021), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14651 ( .A1(n13809), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14652 ( .A1(n10929), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U14653 ( .A1(n11022), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11627) );
  NAND4_X1 U14654 ( .A1(n11630), .A2(n11629), .A3(n11628), .A4(n11627), .ZN(
        n11631) );
  OR2_X1 U14655 ( .A1(n11632), .A2(n11631), .ZN(n11806) );
  INV_X1 U14656 ( .A(n11806), .ZN(n14056) );
  OR2_X1 U14657 ( .A1(n11661), .A2(n14056), .ZN(n11633) );
  AND3_X1 U14658 ( .A1(n11635), .A2(n11634), .A3(n11633), .ZN(n13198) );
  AOI22_X1 U14659 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11020), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14660 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11021), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14661 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14662 ( .A1(n11558), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11022), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11636) );
  NAND4_X1 U14663 ( .A1(n11639), .A2(n11638), .A3(n11637), .A4(n11636), .ZN(
        n11645) );
  AOI22_X1 U14664 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n11840), .ZN(n11643) );
  AOI22_X1 U14665 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11901), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14666 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14667 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11571), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11640) );
  NAND4_X1 U14668 ( .A1(n11643), .A2(n11642), .A3(n11641), .A4(n11640), .ZN(
        n11644) );
  OR2_X1 U14669 ( .A1(n11645), .A2(n11644), .ZN(n11805) );
  INV_X1 U14670 ( .A(n11805), .ZN(n14055) );
  NAND2_X1 U14671 ( .A1(n11668), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14672 ( .A1(n14593), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11646) );
  OAI211_X1 U14673 ( .C1(n11661), .C2(n14055), .A(n11647), .B(n11646), .ZN(
        n13930) );
  AOI22_X1 U14674 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11558), .B1(
        n11057), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14675 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n11840), .ZN(n11650) );
  AOI22_X1 U14676 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n11571), .B1(
        n11072), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14677 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11901), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11648) );
  NAND4_X1 U14678 ( .A1(n11651), .A2(n11650), .A3(n11649), .A4(n11648), .ZN(
        n11657) );
  AOI22_X1 U14679 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11020), .B1(
        n11021), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14680 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n9980), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14681 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14682 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n11022), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11652) );
  NAND4_X1 U14683 ( .A1(n11655), .A2(n11654), .A3(n11653), .A4(n11652), .ZN(
        n11656) );
  OR2_X1 U14684 ( .A1(n11657), .A2(n11656), .ZN(n14176) );
  INV_X1 U14685 ( .A(n14176), .ZN(n11660) );
  NAND2_X1 U14686 ( .A1(n9948), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14687 ( .A1(n14593), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11658) );
  OAI211_X1 U14688 ( .C1(n11661), .C2(n11660), .A(n11659), .B(n11658), .ZN(
        n16509) );
  NAND2_X1 U14689 ( .A1(n11668), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14690 ( .A1(n14593), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11662) );
  NAND2_X1 U14691 ( .A1(n11663), .A2(n11662), .ZN(n14044) );
  NAND2_X1 U14692 ( .A1(n11668), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14693 ( .A1(n14593), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U14694 ( .A1(n11665), .A2(n11664), .ZN(n15566) );
  AND2_X2 U14695 ( .A1(n14042), .A2(n15566), .ZN(n15568) );
  NAND2_X1 U14696 ( .A1(n9948), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14697 ( .A1(n14593), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14698 ( .A1(n11667), .A2(n11666), .ZN(n14201) );
  NAND2_X1 U14699 ( .A1(n11668), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14700 ( .A1(n11690), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11669) );
  AND2_X1 U14701 ( .A1(n11670), .A2(n11669), .ZN(n15559) );
  NAND2_X1 U14702 ( .A1(n11668), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14703 ( .A1(n11690), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11671) );
  NAND2_X1 U14704 ( .A1(n11672), .A2(n11671), .ZN(n14284) );
  NAND2_X1 U14705 ( .A1(n9948), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14706 ( .A1(n11690), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11673) );
  AND2_X1 U14707 ( .A1(n11674), .A2(n11673), .ZN(n15417) );
  NAND2_X1 U14708 ( .A1(n11668), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14709 ( .A1(n11690), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11675) );
  NAND2_X1 U14710 ( .A1(n11676), .A2(n11675), .ZN(n15542) );
  NAND2_X1 U14711 ( .A1(n15541), .A2(n15542), .ZN(n15404) );
  NAND2_X1 U14712 ( .A1(n11668), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14713 ( .A1(n11690), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11677) );
  AND2_X1 U14714 ( .A1(n11678), .A2(n11677), .ZN(n15405) );
  AOI22_X1 U14715 ( .A1(n11690), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11679) );
  OAI21_X1 U14716 ( .B1(n9949), .B2(n19960), .A(n11679), .ZN(n15390) );
  NAND2_X1 U14717 ( .A1(n9948), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14718 ( .A1(n11690), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11681) );
  NAND2_X1 U14719 ( .A1(n11682), .A2(n11681), .ZN(n15525) );
  NAND2_X1 U14720 ( .A1(n15388), .A2(n15525), .ZN(n13227) );
  NAND2_X1 U14721 ( .A1(n9948), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14722 ( .A1(n14593), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11683) );
  AND2_X1 U14723 ( .A1(n11684), .A2(n11683), .ZN(n13228) );
  OR2_X2 U14724 ( .A1(n13227), .A2(n13228), .ZN(n15511) );
  NAND2_X1 U14725 ( .A1(n9948), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14726 ( .A1(n11690), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11685) );
  AND2_X1 U14727 ( .A1(n11686), .A2(n11685), .ZN(n15510) );
  NAND2_X1 U14728 ( .A1(n9948), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14729 ( .A1(n11690), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11687) );
  NAND2_X1 U14730 ( .A1(n11688), .A2(n11687), .ZN(n15502) );
  AOI222_X1 U14731 ( .A1(n9948), .A2(P2_REIP_REG_29__SCAN_IN), .B1(n14593), 
        .B2(P2_EAX_REG_29__SCAN_IN), .C1(n11538), .C2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15497) );
  NAND2_X1 U14732 ( .A1(n9948), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14733 ( .A1(n11690), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11538), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11691) );
  NAND2_X1 U14734 ( .A1(n11692), .A2(n11691), .ZN(n14592) );
  INV_X1 U14735 ( .A(n11693), .ZN(n11694) );
  NAND2_X1 U14736 ( .A1(n10763), .A2(n11694), .ZN(n13785) );
  NAND2_X1 U14737 ( .A1(n11695), .A2(n13179), .ZN(n11696) );
  NAND2_X1 U14738 ( .A1(n13785), .A2(n11696), .ZN(n11697) );
  NAND2_X1 U14739 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15781) );
  INV_X1 U14740 ( .A(n15781), .ZN(n11722) );
  NOR2_X1 U14741 ( .A1(n11094), .A2(n15820), .ZN(n15819) );
  NAND2_X1 U14742 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11734) );
  NOR2_X1 U14743 ( .A1(n14394), .A2(n13367), .ZN(n13366) );
  NOR2_X1 U14744 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13366), .ZN(
        n11736) );
  INV_X1 U14745 ( .A(n11698), .ZN(n11699) );
  AND2_X1 U14746 ( .A1(n11713), .A2(n11699), .ZN(n11700) );
  NAND2_X1 U14747 ( .A1(n11753), .A2(n13784), .ZN(n13338) );
  INV_X1 U14748 ( .A(n13366), .ZN(n11735) );
  OAI21_X1 U14749 ( .B1(n11704), .B2(n11702), .A(n11703), .ZN(n11705) );
  NAND2_X1 U14750 ( .A1(n11705), .A2(n10729), .ZN(n11710) );
  OAI22_X1 U14751 ( .A1(n11703), .A2(n19373), .B1(n20035), .B2(n19361), .ZN(
        n11706) );
  INV_X1 U14752 ( .A(n11706), .ZN(n11709) );
  INV_X1 U14753 ( .A(n11707), .ZN(n11708) );
  NAND2_X1 U14754 ( .A1(n11708), .A2(n11702), .ZN(n12064) );
  AND4_X1 U14755 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n12064), .ZN(
        n11716) );
  NAND2_X1 U14756 ( .A1(n11712), .A2(n13179), .ZN(n13815) );
  NAND2_X1 U14757 ( .A1(n13815), .A2(n11713), .ZN(n11714) );
  NAND2_X1 U14758 ( .A1(n11714), .A2(n10723), .ZN(n11715) );
  AND2_X1 U14759 ( .A1(n11716), .A2(n11715), .ZN(n13817) );
  NAND2_X1 U14760 ( .A1(n13817), .A2(n11717), .ZN(n11718) );
  NAND2_X1 U14761 ( .A1(n11753), .A2(n11718), .ZN(n15888) );
  INV_X1 U14762 ( .A(n15888), .ZN(n11737) );
  NAND2_X1 U14763 ( .A1(n11737), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11719) );
  OAI22_X1 U14764 ( .A1(n11736), .A2(n13338), .B1(n11735), .B2(n11719), .ZN(
        n14029) );
  NAND2_X1 U14765 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14029), .ZN(
        n16554) );
  NOR2_X1 U14766 ( .A1(n11734), .A2(n16554), .ZN(n14296) );
  NAND2_X1 U14767 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14296), .ZN(
        n16541) );
  INV_X1 U14768 ( .A(n16541), .ZN(n11720) );
  NOR2_X1 U14769 ( .A1(n16543), .A2(n16545), .ZN(n16542) );
  NAND3_X1 U14770 ( .A1(n15913), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15914), .ZN(n16512) );
  NOR2_X1 U14771 ( .A1(n16512), .A2(n11741), .ZN(n15861) );
  NAND2_X1 U14772 ( .A1(n15861), .A2(n11721), .ZN(n15840) );
  NOR2_X1 U14773 ( .A1(n15662), .A2(n15840), .ZN(n15831) );
  AND2_X1 U14774 ( .A1(n15819), .A2(n15831), .ZN(n15807) );
  NAND2_X1 U14775 ( .A1(n11722), .A2(n15794), .ZN(n15770) );
  AND2_X1 U14776 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15745) );
  NAND2_X1 U14777 ( .A1(n15745), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15744) );
  INV_X2 U14778 ( .A(n19328), .ZN(n19181) );
  INV_X1 U14779 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n11723) );
  NOR2_X1 U14780 ( .A1(n19181), .A2(n11723), .ZN(n11757) );
  INV_X1 U14781 ( .A(n11757), .ZN(n11724) );
  OAI211_X1 U14782 ( .C1(n15374), .C2(n16544), .A(n10336), .B(n11724), .ZN(
        n11725) );
  INV_X1 U14783 ( .A(n11725), .ZN(n11733) );
  AOI22_X1 U14784 ( .A1(n11383), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11727) );
  NAND2_X1 U14785 ( .A1(n14585), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11726) );
  OAI211_X1 U14786 ( .C1(n9960), .C2(n11728), .A(n11727), .B(n11726), .ZN(
        n15426) );
  INV_X1 U14787 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14597) );
  AOI22_X1 U14788 ( .A1(n11383), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11730) );
  NAND2_X1 U14789 ( .A1(n14585), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11729) );
  OAI211_X1 U14790 ( .C1(n9959), .C2(n14597), .A(n11730), .B(n11729), .ZN(
        n14584) );
  INV_X1 U14791 ( .A(n15889), .ZN(n15944) );
  INV_X1 U14792 ( .A(n11734), .ZN(n16555) );
  NOR2_X1 U14793 ( .A1(n11753), .A2(n19328), .ZN(n13370) );
  AOI21_X1 U14794 ( .B1(n11735), .B2(n11737), .A(n13370), .ZN(n13352) );
  INV_X1 U14795 ( .A(n13338), .ZN(n15885) );
  NAND2_X1 U14796 ( .A1(n15885), .A2(n11736), .ZN(n13347) );
  INV_X1 U14797 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U14798 ( .A1(n11737), .A2(n13351), .ZN(n13337) );
  NAND3_X1 U14799 ( .A1(n13352), .A2(n13347), .A3(n13337), .ZN(n14031) );
  AOI21_X1 U14800 ( .B1(n14030), .B2(n15889), .A(n14031), .ZN(n16571) );
  OAI21_X1 U14801 ( .B1(n15944), .B2(n16555), .A(n16571), .ZN(n14294) );
  AND2_X1 U14802 ( .A1(n15889), .A2(n14295), .ZN(n11738) );
  NOR2_X1 U14803 ( .A1(n14294), .A2(n11738), .ZN(n16546) );
  INV_X1 U14804 ( .A(n16542), .ZN(n11739) );
  NAND2_X1 U14805 ( .A1(n15889), .A2(n11739), .ZN(n11740) );
  NAND2_X1 U14806 ( .A1(n16546), .A2(n11740), .ZN(n15916) );
  NAND3_X1 U14807 ( .A1(n15913), .A2(n11092), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11742) );
  AND2_X1 U14808 ( .A1(n15889), .A2(n11742), .ZN(n11743) );
  AND2_X1 U14809 ( .A1(n15889), .A2(n15853), .ZN(n11744) );
  AND2_X1 U14810 ( .A1(n15889), .A2(n15662), .ZN(n11745) );
  NOR2_X1 U14811 ( .A1(n15838), .A2(n11745), .ZN(n15828) );
  INV_X1 U14812 ( .A(n15819), .ZN(n11746) );
  NAND2_X1 U14813 ( .A1(n15889), .A2(n11746), .ZN(n11747) );
  NAND2_X1 U14814 ( .A1(n15828), .A2(n11747), .ZN(n15803) );
  AND2_X1 U14815 ( .A1(n15889), .A2(n15808), .ZN(n11748) );
  AND2_X1 U14816 ( .A1(n15889), .A2(n15781), .ZN(n11749) );
  NOR2_X1 U14817 ( .A1(n15799), .A2(n11749), .ZN(n15772) );
  NAND2_X1 U14818 ( .A1(n15889), .A2(n15744), .ZN(n11750) );
  AND2_X1 U14819 ( .A1(n15772), .A2(n11750), .ZN(n14583) );
  NAND2_X1 U14820 ( .A1(n11751), .A2(n10314), .ZN(n11752) );
  AOI21_X1 U14821 ( .B1(n11761), .B2(n16563), .A(n11752), .ZN(n11756) );
  XNOR2_X1 U14822 ( .A(n15578), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11762) );
  INV_X1 U14823 ( .A(n11753), .ZN(n11754) );
  NAND2_X1 U14824 ( .A1(n11756), .A2(n11755), .ZN(P2_U3016) );
  INV_X1 U14825 ( .A(n14136), .ZN(n19337) );
  INV_X1 U14826 ( .A(n16506), .ZN(n19329) );
  AOI21_X1 U14827 ( .B1(n19329), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n11757), .ZN(n11759) );
  INV_X1 U14828 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16381) );
  XOR2_X1 U14829 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n15352), .Z(
        n15368) );
  NAND2_X1 U14830 ( .A1(n16496), .A2(n15368), .ZN(n11758) );
  OAI211_X1 U14831 ( .C1(n15379), .C2(n14136), .A(n11759), .B(n11758), .ZN(
        n11760) );
  AOI21_X1 U14832 ( .B1(n11761), .B2(n16502), .A(n11760), .ZN(n11764) );
  NAND2_X1 U14833 ( .A1(n11764), .A2(n11763), .ZN(P2_U2984) );
  INV_X1 U14834 ( .A(n11766), .ZN(n11791) );
  NAND2_X1 U14835 ( .A1(n11765), .A2(n11791), .ZN(n11770) );
  OAI21_X1 U14836 ( .B1(n19384), .B2(n19032), .A(n20012), .ZN(n11788) );
  AND2_X1 U14837 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19698) );
  NAND2_X1 U14838 ( .A1(n19698), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19345) );
  NAND2_X1 U14839 ( .A1(n19345), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11767) );
  NOR3_X1 U14840 ( .A1(n20002), .A2(n20011), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19577) );
  NAND2_X1 U14841 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19577), .ZN(
        n19602) );
  NAND2_X1 U14842 ( .A1(n11767), .A2(n19602), .ZN(n11768) );
  AND2_X1 U14843 ( .A1(n11768), .A2(n19990), .ZN(n14128) );
  AOI21_X1 U14844 ( .B1(n11788), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14128), .ZN(n11769) );
  INV_X1 U14845 ( .A(n11797), .ZN(n11774) );
  AND2_X1 U14846 ( .A1(n19384), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11771) );
  NAND2_X1 U14847 ( .A1(n11771), .A2(n13179), .ZN(n13616) );
  INV_X1 U14848 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11772) );
  NOR2_X1 U14849 ( .A1(n13616), .A2(n11772), .ZN(n11775) );
  INV_X1 U14850 ( .A(n11775), .ZN(n11773) );
  NAND2_X1 U14851 ( .A1(n11774), .A2(n11773), .ZN(n11776) );
  NAND2_X1 U14852 ( .A1(n11797), .A2(n11775), .ZN(n13619) );
  NAND2_X1 U14853 ( .A1(n11776), .A2(n13619), .ZN(n13529) );
  INV_X1 U14854 ( .A(n13529), .ZN(n11796) );
  NAND2_X1 U14855 ( .A1(n11777), .A2(n11791), .ZN(n11779) );
  NAND2_X1 U14856 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20011), .ZN(
        n19634) );
  NAND2_X1 U14857 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20020), .ZN(
        n19670) );
  NAND2_X1 U14858 ( .A1(n19634), .A2(n19670), .ZN(n14121) );
  AND2_X1 U14859 ( .A1(n19990), .A2(n14121), .ZN(n19669) );
  AOI21_X1 U14860 ( .B1(n11788), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19669), .ZN(n11778) );
  NAND2_X1 U14861 ( .A1(n11779), .A2(n11778), .ZN(n13358) );
  AOI22_X1 U14862 ( .A1(n11788), .A2(n9932), .B1(n19990), .B2(n20020), .ZN(
        n11780) );
  NOR2_X1 U14863 ( .A1(n13616), .A2(n11576), .ZN(n11783) );
  XNOR2_X1 U14864 ( .A(n11782), .B(n11783), .ZN(n13359) );
  INV_X1 U14865 ( .A(n11782), .ZN(n11785) );
  INV_X1 U14866 ( .A(n11783), .ZN(n11784) );
  NAND2_X1 U14867 ( .A1(n11785), .A2(n11784), .ZN(n11786) );
  INV_X1 U14868 ( .A(n13616), .ZN(n12000) );
  NAND2_X1 U14869 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13470) );
  INV_X1 U14870 ( .A(n19698), .ZN(n19454) );
  NAND2_X1 U14871 ( .A1(n19454), .A2(n20002), .ZN(n11787) );
  NAND2_X1 U14872 ( .A1(n19345), .A2(n11787), .ZN(n14122) );
  NAND2_X1 U14873 ( .A1(n11788), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11789) );
  OAI21_X1 U14874 ( .B1(n19599), .B2(n14122), .A(n11789), .ZN(n11790) );
  NAND2_X1 U14875 ( .A1(n13468), .A2(n13470), .ZN(n11792) );
  NAND2_X1 U14876 ( .A1(n11793), .A2(n11792), .ZN(n13530) );
  INV_X1 U14877 ( .A(n13530), .ZN(n11795) );
  AND2_X1 U14878 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10738), .ZN(
        n11794) );
  NAND2_X1 U14879 ( .A1(n11797), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11798) );
  AND2_X1 U14880 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13707) );
  NAND4_X1 U14881 ( .A1(n11799), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .A4(n13707), .ZN(n11800) );
  NOR2_X1 U14882 ( .A1(n13616), .A2(n11800), .ZN(n11801) );
  INV_X1 U14883 ( .A(n13731), .ZN(n11803) );
  INV_X1 U14884 ( .A(n13933), .ZN(n11802) );
  NAND2_X1 U14885 ( .A1(n11803), .A2(n11802), .ZN(n13942) );
  AND2_X1 U14886 ( .A1(n11806), .A2(n11805), .ZN(n14054) );
  AND2_X1 U14887 ( .A1(n14176), .A2(n14054), .ZN(n11807) );
  NAND2_X1 U14888 ( .A1(n13943), .A2(n11807), .ZN(n14038) );
  AOI22_X1 U14889 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11558), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U14890 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11840), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U14891 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U14892 ( .A1(n11901), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11808) );
  NAND4_X1 U14893 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11817) );
  AOI22_X1 U14894 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11021), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U14895 ( .A1(n13809), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14896 ( .A1(n10929), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U14897 ( .A1(n11022), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11812) );
  NAND4_X1 U14898 ( .A1(n11815), .A2(n11814), .A3(n11813), .A4(n11812), .ZN(
        n11816) );
  NOR2_X1 U14899 ( .A1(n11817), .A2(n11816), .ZN(n14041) );
  INV_X1 U14900 ( .A(n14041), .ZN(n11818) );
  AOI22_X1 U14901 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11558), .B1(
        n11057), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U14902 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n11840), .ZN(n11822) );
  AOI22_X1 U14903 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n11072), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U14904 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11901), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11820) );
  NAND4_X1 U14905 ( .A1(n11823), .A2(n11822), .A3(n11821), .A4(n11820), .ZN(
        n11829) );
  AOI22_X1 U14906 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11021), .B1(
        n11020), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U14907 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n9980), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U14908 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14909 ( .A1(n11022), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11824) );
  NAND4_X1 U14910 ( .A1(n11827), .A2(n11826), .A3(n11825), .A4(n11824), .ZN(
        n11828) );
  OR2_X1 U14911 ( .A1(n11829), .A2(n11828), .ZN(n14278) );
  AOI22_X1 U14912 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11558), .B1(
        n11057), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U14913 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n11840), .ZN(n11832) );
  AOI22_X1 U14914 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n11072), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U14915 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11901), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11830) );
  NAND4_X1 U14916 ( .A1(n11833), .A2(n11832), .A3(n11831), .A4(n11830), .ZN(
        n11839) );
  AOI22_X1 U14917 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11021), .B1(
        n11020), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14918 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n9980), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U14919 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U14920 ( .A1(n11022), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11834) );
  NAND4_X1 U14921 ( .A1(n11837), .A2(n11836), .A3(n11835), .A4(n11834), .ZN(
        n11838) );
  OR2_X1 U14922 ( .A1(n11839), .A2(n11838), .ZN(n14199) );
  AOI22_X1 U14923 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11558), .B1(
        n11057), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14924 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n11840), .ZN(n11843) );
  AOI22_X1 U14925 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11072), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U14926 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n11901), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11841) );
  NAND4_X1 U14927 ( .A1(n11844), .A2(n11843), .A3(n11842), .A4(n11841), .ZN(
        n11850) );
  AOI22_X1 U14928 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11021), .B1(
        n11020), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14929 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n9980), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14930 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14931 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11022), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11845) );
  NAND4_X1 U14932 ( .A1(n11848), .A2(n11847), .A3(n11846), .A4(n11845), .ZN(
        n11849) );
  OR2_X1 U14933 ( .A1(n11850), .A2(n11849), .ZN(n14200) );
  AOI22_X1 U14934 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11021), .B1(
        n11020), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14935 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n9980), .B1(
        n13809), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U14936 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U14937 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11022), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11851) );
  NAND4_X1 U14938 ( .A1(n11854), .A2(n11853), .A3(n11852), .A4(n11851), .ZN(
        n11860) );
  AOI22_X1 U14939 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11558), .B1(
        n11057), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U14940 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n11840), .ZN(n11857) );
  AOI22_X1 U14941 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11072), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U14942 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11901), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11855) );
  NAND4_X1 U14943 ( .A1(n11858), .A2(n11857), .A3(n11856), .A4(n11855), .ZN(
        n11859) );
  OR2_X1 U14944 ( .A1(n11860), .A2(n11859), .ZN(n14281) );
  NAND4_X1 U14945 ( .A1(n14278), .A2(n14199), .A3(n14200), .A4(n14281), .ZN(
        n11861) );
  AOI22_X1 U14946 ( .A1(n11020), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11021), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U14947 ( .A1(n13809), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U14948 ( .A1(n10929), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U14949 ( .A1(n11022), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11862) );
  NAND4_X1 U14950 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n11871) );
  AOI22_X1 U14951 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11840), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14952 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11558), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U14953 ( .A1(n11901), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14954 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11866) );
  NAND4_X1 U14955 ( .A1(n11869), .A2(n11868), .A3(n11867), .A4(n11866), .ZN(
        n11870) );
  OR2_X1 U14956 ( .A1(n11871), .A2(n11870), .ZN(n15484) );
  AOI22_X1 U14957 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n11840), .ZN(n11875) );
  AOI22_X1 U14958 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11558), .B1(
        n11057), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14959 ( .A1(n11901), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U14960 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11072), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11872) );
  NAND4_X1 U14961 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11881) );
  AOI22_X1 U14962 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11021), .B1(
        n11020), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U14963 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n13809), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14964 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14965 ( .A1(n11022), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11876) );
  NAND4_X1 U14966 ( .A1(n11879), .A2(n11878), .A3(n11877), .A4(n11876), .ZN(
        n11880) );
  NOR2_X1 U14967 ( .A1(n11881), .A2(n11880), .ZN(n15480) );
  AOI22_X1 U14968 ( .A1(n9931), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U14969 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11882) );
  AND2_X1 U14970 ( .A1(n11883), .A2(n11882), .ZN(n11886) );
  XNOR2_X1 U14971 ( .A(n13802), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12053) );
  AOI22_X1 U14972 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12047), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U14973 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9953), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11884) );
  NAND4_X1 U14974 ( .A1(n11886), .A2(n12053), .A3(n11885), .A4(n11884), .ZN(
        n11895) );
  AOI22_X1 U14975 ( .A1(n9928), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9818), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11893) );
  NAND2_X1 U14976 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11890) );
  NAND2_X1 U14977 ( .A1(n9953), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11889) );
  NAND2_X1 U14978 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11888) );
  NAND2_X1 U14979 ( .A1(n9956), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11887) );
  AND4_X1 U14980 ( .A1(n11890), .A2(n11889), .A3(n11888), .A4(n11887), .ZN(
        n11892) );
  AOI22_X1 U14981 ( .A1(n10674), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11891) );
  INV_X1 U14982 ( .A(n12053), .ZN(n12050) );
  NAND4_X1 U14983 ( .A1(n11893), .A2(n11892), .A3(n11891), .A4(n12050), .ZN(
        n11894) );
  NAND2_X1 U14984 ( .A1(n11895), .A2(n11894), .ZN(n11932) );
  NOR2_X1 U14985 ( .A1(n19356), .A2(n11932), .ZN(n11909) );
  AOI22_X1 U14986 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n11021), .B1(
        n11020), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U14987 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n13809), .B1(
        n9980), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U14988 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10929), .B1(
        n10886), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U14989 ( .A1(n11558), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11022), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11896) );
  NAND4_X1 U14990 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n11908) );
  AOI22_X1 U14991 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11901), .B1(
        n11900), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U14992 ( .A1(n11057), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11902), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U14993 ( .A1(n11069), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11571), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U14994 ( .A1(n11072), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n11840), .ZN(n11903) );
  NAND4_X1 U14995 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n11903), .ZN(
        n11907) );
  OR2_X1 U14996 ( .A1(n11908), .A2(n11907), .ZN(n11913) );
  XNOR2_X1 U14997 ( .A(n11909), .B(n11913), .ZN(n11933) );
  INV_X1 U14998 ( .A(n11932), .ZN(n11912) );
  NAND2_X1 U14999 ( .A1(n19356), .A2(n11912), .ZN(n15472) );
  BUF_X1 U15000 ( .A(n11911), .Z(n15479) );
  NAND2_X1 U15001 ( .A1(n11913), .A2(n11912), .ZN(n11936) );
  NAND2_X1 U15002 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11917) );
  NAND2_X1 U15003 ( .A1(n10863), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11916) );
  NAND2_X1 U15004 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11915) );
  NAND2_X1 U15005 ( .A1(n9954), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11914) );
  AND4_X1 U15006 ( .A1(n11917), .A2(n11916), .A3(n11915), .A4(n11914), .ZN(
        n11920) );
  AOI22_X1 U15007 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U15008 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11918) );
  NAND4_X1 U15009 ( .A1(n11920), .A2(n11919), .A3(n11918), .A4(n12050), .ZN(
        n11929) );
  NAND2_X1 U15010 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11924) );
  NAND2_X1 U15011 ( .A1(n9953), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11923) );
  NAND2_X1 U15012 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11922) );
  NAND2_X1 U15013 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11921) );
  AND4_X1 U15014 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .ZN(
        n11927) );
  AOI22_X1 U15015 ( .A1(n9929), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U15016 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11925) );
  NAND4_X1 U15017 ( .A1(n11927), .A2(n12053), .A3(n11926), .A4(n11925), .ZN(
        n11928) );
  NAND2_X1 U15018 ( .A1(n11929), .A2(n11928), .ZN(n11935) );
  XOR2_X1 U15019 ( .A(n11936), .B(n11935), .Z(n11930) );
  NAND2_X1 U15020 ( .A1(n11930), .A2(n12000), .ZN(n15465) );
  INV_X1 U15021 ( .A(n11935), .ZN(n11931) );
  NAND2_X1 U15022 ( .A1(n19356), .A2(n11931), .ZN(n15467) );
  NOR3_X1 U15023 ( .A1(n11933), .A2(n11932), .A3(n15467), .ZN(n11934) );
  NOR2_X1 U15024 ( .A1(n11936), .A2(n11935), .ZN(n11954) );
  NAND2_X1 U15025 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U15026 ( .A1(n10863), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11940) );
  NAND2_X1 U15027 ( .A1(n10716), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n11939) );
  NAND2_X1 U15028 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11938) );
  AND4_X1 U15029 ( .A1(n11941), .A2(n11940), .A3(n11939), .A4(n11938), .ZN(
        n11944) );
  AOI22_X1 U15030 ( .A1(n9931), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U15031 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11942) );
  NAND4_X1 U15032 ( .A1(n11944), .A2(n11943), .A3(n11942), .A4(n12050), .ZN(
        n11953) );
  NAND2_X1 U15033 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11948) );
  NAND2_X1 U15034 ( .A1(n9953), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11947) );
  NAND2_X1 U15035 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11946) );
  NAND2_X1 U15036 ( .A1(n9955), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11945) );
  AND4_X1 U15037 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n11951) );
  AOI22_X1 U15038 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15039 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11949) );
  NAND4_X1 U15040 ( .A1(n11951), .A2(n12053), .A3(n11950), .A4(n11949), .ZN(
        n11952) );
  AND2_X1 U15041 ( .A1(n11953), .A2(n11952), .ZN(n11956) );
  NAND2_X1 U15042 ( .A1(n11954), .A2(n11956), .ZN(n11997) );
  OAI211_X1 U15043 ( .C1(n11954), .C2(n11956), .A(n11997), .B(n12000), .ZN(
        n11959) );
  INV_X1 U15044 ( .A(n11956), .ZN(n11957) );
  NOR2_X1 U15045 ( .A1(n13179), .A2(n11957), .ZN(n15456) );
  INV_X1 U15046 ( .A(n11958), .ZN(n11960) );
  NAND2_X1 U15047 ( .A1(n10863), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11964) );
  NAND2_X1 U15048 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11963) );
  NAND2_X1 U15049 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11962) );
  AND4_X1 U15050 ( .A1(n11965), .A2(n11964), .A3(n11963), .A4(n11962), .ZN(
        n11968) );
  AOI22_X1 U15051 ( .A1(n9928), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U15052 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11966) );
  NAND4_X1 U15053 ( .A1(n11968), .A2(n11967), .A3(n11966), .A4(n12050), .ZN(
        n11977) );
  NAND2_X1 U15054 ( .A1(n9953), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11971) );
  NAND2_X1 U15055 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11970) );
  NAND2_X1 U15056 ( .A1(n9956), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11969) );
  AND4_X1 U15057 ( .A1(n11972), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11975) );
  AOI22_X1 U15058 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15059 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11973) );
  NAND4_X1 U15060 ( .A1(n11975), .A2(n12053), .A3(n11974), .A4(n11973), .ZN(
        n11976) );
  AND2_X1 U15061 ( .A1(n11977), .A2(n11976), .ZN(n11998) );
  XNOR2_X1 U15062 ( .A(n11997), .B(n11998), .ZN(n11978) );
  NAND2_X1 U15063 ( .A1(n19356), .A2(n11998), .ZN(n15451) );
  NAND2_X1 U15064 ( .A1(n9953), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11983) );
  NAND2_X1 U15065 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11982) );
  NAND2_X1 U15066 ( .A1(n9955), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11981) );
  AND4_X1 U15067 ( .A1(n11984), .A2(n11983), .A3(n11982), .A4(n11981), .ZN(
        n11987) );
  AOI22_X1 U15068 ( .A1(n9928), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U15069 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11985) );
  NAND4_X1 U15070 ( .A1(n11987), .A2(n11986), .A3(n11985), .A4(n12050), .ZN(
        n11996) );
  NAND2_X1 U15071 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11991) );
  NAND2_X1 U15072 ( .A1(n10863), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11990) );
  NAND2_X1 U15073 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11989) );
  NAND2_X1 U15074 ( .A1(n9954), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11988) );
  AND4_X1 U15075 ( .A1(n11991), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(
        n11994) );
  AOI22_X1 U15076 ( .A1(n9931), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15077 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11992) );
  NAND4_X1 U15078 ( .A1(n11994), .A2(n12053), .A3(n11993), .A4(n11992), .ZN(
        n11995) );
  AND2_X1 U15079 ( .A1(n11996), .A2(n11995), .ZN(n12005) );
  INV_X1 U15080 ( .A(n11997), .ZN(n11999) );
  AND2_X1 U15081 ( .A1(n11999), .A2(n11998), .ZN(n12001) );
  NAND2_X1 U15082 ( .A1(n12001), .A2(n12005), .ZN(n15435) );
  OAI211_X1 U15083 ( .C1(n12005), .C2(n12001), .A(n12000), .B(n15435), .ZN(
        n12002) );
  NOR2_X1 U15084 ( .A1(n12003), .A2(n12002), .ZN(n12007) );
  INV_X1 U15085 ( .A(n12005), .ZN(n12006) );
  NOR2_X1 U15086 ( .A1(n13179), .A2(n12006), .ZN(n15443) );
  NAND2_X1 U15087 ( .A1(n15441), .A2(n15443), .ZN(n15442) );
  INV_X1 U15088 ( .A(n12007), .ZN(n15436) );
  NAND2_X1 U15089 ( .A1(n9953), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12010) );
  NAND2_X1 U15090 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12009) );
  NAND2_X1 U15091 ( .A1(n9956), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12008) );
  AND4_X1 U15092 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        n12014) );
  AOI22_X1 U15093 ( .A1(n9929), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15094 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12012) );
  NAND4_X1 U15095 ( .A1(n12014), .A2(n12013), .A3(n12012), .A4(n12050), .ZN(
        n12023) );
  NAND2_X1 U15096 ( .A1(n10863), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12017) );
  NAND2_X1 U15097 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12016) );
  NAND2_X1 U15098 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12015) );
  AND4_X1 U15099 ( .A1(n12018), .A2(n12017), .A3(n12016), .A4(n12015), .ZN(
        n12021) );
  AOI22_X1 U15100 ( .A1(n9928), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15101 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12019) );
  NAND4_X1 U15102 ( .A1(n12021), .A2(n12053), .A3(n12020), .A4(n12019), .ZN(
        n12022) );
  NAND2_X1 U15103 ( .A1(n12023), .A2(n12022), .ZN(n12041) );
  AOI21_X2 U15104 ( .B1(n15442), .B2(n15436), .A(n12041), .ZN(n15431) );
  NAND2_X1 U15105 ( .A1(n9953), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12026) );
  NAND2_X1 U15106 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12025) );
  NAND2_X1 U15107 ( .A1(n9954), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12024) );
  AND4_X1 U15108 ( .A1(n12027), .A2(n12026), .A3(n12025), .A4(n12024), .ZN(
        n12031) );
  AOI22_X1 U15109 ( .A1(n9931), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15110 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12029) );
  NAND4_X1 U15111 ( .A1(n12031), .A2(n12030), .A3(n12029), .A4(n12050), .ZN(
        n12040) );
  NAND2_X1 U15112 ( .A1(n10863), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12035) );
  NAND2_X1 U15113 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12033) );
  NAND2_X1 U15114 ( .A1(n10674), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12032) );
  AND4_X1 U15115 ( .A1(n12035), .A2(n12034), .A3(n12033), .A4(n12032), .ZN(
        n12038) );
  AOI22_X1 U15116 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15117 ( .A1(n9929), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12036) );
  NAND4_X1 U15118 ( .A1(n12038), .A2(n12053), .A3(n12037), .A4(n12036), .ZN(
        n12039) );
  NAND2_X1 U15119 ( .A1(n12040), .A2(n12039), .ZN(n12044) );
  INV_X1 U15120 ( .A(n12041), .ZN(n15437) );
  NAND2_X1 U15121 ( .A1(n13179), .A2(n15437), .ZN(n12042) );
  OR2_X1 U15122 ( .A1(n15435), .A2(n12042), .ZN(n12043) );
  NOR2_X1 U15123 ( .A1(n12043), .A2(n12044), .ZN(n12045) );
  AOI21_X1 U15124 ( .B1(n12044), .B2(n12043), .A(n12045), .ZN(n15430) );
  INV_X1 U15125 ( .A(n12045), .ZN(n12046) );
  AOI22_X1 U15126 ( .A1(n10652), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9953), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15127 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9823), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12048) );
  NAND2_X1 U15128 ( .A1(n12049), .A2(n12048), .ZN(n12061) );
  AOI22_X1 U15129 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U15130 ( .A1(n9930), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12051) );
  NAND3_X1 U15131 ( .A1(n12052), .A2(n12051), .A3(n12050), .ZN(n12060) );
  AOI22_X1 U15132 ( .A1(n9931), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9955), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15133 ( .A1(n12028), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10868), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12054) );
  NAND3_X1 U15134 ( .A1(n12055), .A2(n12054), .A3(n12053), .ZN(n12059) );
  AOI22_X1 U15135 ( .A1(n12047), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10674), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12056) );
  NAND2_X1 U15136 ( .A1(n12057), .A2(n12056), .ZN(n12058) );
  OAI22_X1 U15137 ( .A1(n12061), .A2(n12060), .B1(n12059), .B2(n12058), .ZN(
        n12062) );
  NAND2_X1 U15138 ( .A1(n11695), .A2(n13828), .ZN(n13252) );
  NAND2_X1 U15139 ( .A1(n11703), .A2(n20046), .ZN(n13249) );
  NOR2_X1 U15140 ( .A1(n13252), .A2(n13249), .ZN(n12063) );
  AOI21_X1 U15141 ( .B1(n13833), .B2(n13784), .A(n12063), .ZN(n13800) );
  NAND2_X1 U15142 ( .A1(n13800), .A2(n12064), .ZN(n12065) );
  NAND2_X1 U15143 ( .A1(n19250), .A2(n12066), .ZN(n19257) );
  NOR4_X1 U15144 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12071) );
  NOR4_X1 U15145 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12070) );
  NOR4_X1 U15146 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12069) );
  NOR4_X1 U15147 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12068) );
  NAND4_X1 U15148 ( .A1(n12071), .A2(n12070), .A3(n12069), .A4(n12068), .ZN(
        n12076) );
  NOR4_X1 U15149 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12074) );
  NOR4_X1 U15150 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12073) );
  NOR4_X1 U15151 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12072) );
  INV_X1 U15152 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19921) );
  NAND4_X1 U15153 ( .A1(n12074), .A2(n12073), .A3(n12072), .A4(n19921), .ZN(
        n12075) );
  MUX2_X1 U15154 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n14137), .Z(n13929) );
  NAND2_X1 U15155 ( .A1(n19250), .A2(n11511), .ZN(n15552) );
  INV_X1 U15156 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12077) );
  OAI22_X1 U15157 ( .A1(n15374), .A2(n15552), .B1(n19250), .B2(n12077), .ZN(
        n12078) );
  AOI21_X1 U15158 ( .B1(n16430), .B2(n13929), .A(n12078), .ZN(n12081) );
  NOR2_X1 U15159 ( .A1(n11511), .A2(n19384), .ZN(n12079) );
  NAND2_X1 U15160 ( .A1(n19250), .A2(n12079), .ZN(n13323) );
  NOR2_X2 U15161 ( .A1(n13323), .A2(n14135), .ZN(n19233) );
  NOR2_X2 U15162 ( .A1(n13323), .A2(n14137), .ZN(n19235) );
  AOI22_X1 U15163 ( .A1(n19233), .A2(BUF2_REG_30__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12080) );
  AND2_X1 U15164 ( .A1(n12081), .A2(n12080), .ZN(n12082) );
  OAI21_X1 U15165 ( .B1(n14621), .B2(n19257), .A(n12082), .ZN(P2_U2889) );
  INV_X1 U15166 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12085) );
  NAND2_X1 U15167 ( .A1(n12855), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12084) );
  NAND2_X1 U15168 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12083) );
  OAI211_X1 U15169 ( .C1(n12516), .C2(n12085), .A(n12084), .B(n12083), .ZN(
        n12086) );
  INV_X1 U15170 ( .A(n12086), .ZN(n12092) );
  AOI22_X1 U15171 ( .A1(n12880), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12091) );
  INV_X4 U15172 ( .A(n12959), .ZN(n12997) );
  AOI22_X1 U15173 ( .A1(n9962), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12090) );
  NAND2_X1 U15174 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12089) );
  NAND4_X1 U15175 ( .A1(n12092), .A2(n12091), .A3(n12090), .A4(n12089), .ZN(
        n12101) );
  AOI22_X1 U15176 ( .A1(n9822), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12099) );
  AND2_X2 U15177 ( .A1(n12095), .A2(n13885), .ZN(n12293) );
  AOI22_X1 U15178 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12098) );
  AND2_X2 U15179 ( .A1(n12095), .A2(n13886), .ZN(n12315) );
  AOI22_X1 U15180 ( .A1(n12797), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12097) );
  AND2_X2 U15181 ( .A1(n13886), .A2(n13537), .ZN(n12348) );
  AOI22_X1 U15182 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12348), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12096) );
  NAND4_X1 U15183 ( .A1(n12099), .A2(n12098), .A3(n12097), .A4(n12096), .ZN(
        n12100) );
  OR2_X2 U15184 ( .A1(n12101), .A2(n12100), .ZN(n20268) );
  AOI22_X1 U15185 ( .A1(n12797), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15186 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15187 ( .A1(n9944), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12104) );
  INV_X1 U15188 ( .A(n12348), .ZN(n12102) );
  AOI22_X1 U15189 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12348), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12103) );
  INV_X1 U15190 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12960) );
  NAND2_X1 U15191 ( .A1(n12855), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12108) );
  NAND2_X1 U15192 ( .A1(n9946), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12107) );
  OAI211_X1 U15193 ( .C1(n12516), .C2(n12960), .A(n12108), .B(n12107), .ZN(
        n12109) );
  INV_X1 U15194 ( .A(n12109), .ZN(n12113) );
  AOI22_X1 U15195 ( .A1(n12880), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15196 ( .A1(n12998), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12111) );
  NAND2_X1 U15197 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12110) );
  NAND2_X1 U15198 ( .A1(n12998), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12117) );
  NAND2_X1 U15199 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12116) );
  NAND2_X1 U15200 ( .A1(n12177), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12115) );
  NAND2_X1 U15201 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12114) );
  NAND4_X1 U15202 ( .A1(n12117), .A2(n12116), .A3(n12115), .A4(n12114), .ZN(
        n12119) );
  INV_X1 U15203 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12989) );
  NOR2_X1 U15204 ( .A1(n12232), .A2(n12989), .ZN(n12118) );
  NOR2_X1 U15205 ( .A1(n12119), .A2(n12118), .ZN(n12135) );
  INV_X1 U15206 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12122) );
  NAND2_X1 U15207 ( .A1(n12855), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12121) );
  NAND2_X1 U15208 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12120) );
  OAI211_X1 U15209 ( .C1(n12516), .C2(n12122), .A(n12121), .B(n12120), .ZN(
        n12123) );
  INV_X1 U15210 ( .A(n12123), .ZN(n12134) );
  NAND2_X1 U15211 ( .A1(n12880), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12127) );
  NAND2_X1 U15212 ( .A1(n9942), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12126) );
  NAND2_X1 U15213 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12125) );
  NAND2_X1 U15214 ( .A1(n9822), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12124) );
  NAND2_X1 U15215 ( .A1(n9940), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12131) );
  NAND2_X1 U15216 ( .A1(n12293), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12130) );
  NAND2_X1 U15217 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12129) );
  NAND2_X1 U15218 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12128) );
  NAND2_X1 U15219 ( .A1(n12247), .A2(n13086), .ZN(n12189) );
  NAND2_X1 U15220 ( .A1(n9940), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12139) );
  NAND2_X1 U15221 ( .A1(n12293), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12138) );
  NAND2_X1 U15222 ( .A1(n9822), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12137) );
  NAND2_X1 U15223 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12136) );
  NAND2_X1 U15224 ( .A1(n12998), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12142) );
  INV_X1 U15225 ( .A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12140) );
  NAND2_X1 U15226 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12145) );
  INV_X1 U15227 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12143) );
  NAND2_X1 U15228 ( .A1(n12880), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12144) );
  INV_X1 U15229 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12147) );
  NAND2_X1 U15230 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12149) );
  NAND2_X1 U15231 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12148) );
  INV_X1 U15232 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12154) );
  NAND2_X1 U15233 ( .A1(n12855), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12153) );
  NAND2_X1 U15234 ( .A1(n9946), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12152) );
  OAI211_X1 U15235 ( .C1(n12516), .C2(n12154), .A(n12153), .B(n12152), .ZN(
        n12155) );
  INV_X1 U15236 ( .A(n12155), .ZN(n12156) );
  NAND4_X4 U15237 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12241) );
  NAND2_X1 U15238 ( .A1(n9944), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12162) );
  NAND2_X1 U15239 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12161) );
  NAND2_X1 U15240 ( .A1(n12293), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12160) );
  NAND3_X1 U15241 ( .A1(n12162), .A2(n12161), .A3(n12160), .ZN(n12163) );
  INV_X1 U15242 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12904) );
  NAND2_X1 U15243 ( .A1(n9962), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12165) );
  NAND2_X1 U15244 ( .A1(n9958), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12164) );
  NAND2_X1 U15245 ( .A1(n12880), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12168) );
  NAND2_X1 U15246 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12167) );
  NOR2_X1 U15247 ( .A1(n12170), .A2(n12169), .ZN(n12185) );
  INV_X1 U15248 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12173) );
  NAND2_X1 U15249 ( .A1(n12855), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12172) );
  NAND2_X1 U15250 ( .A1(n9947), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12171) );
  OAI211_X1 U15251 ( .C1(n12516), .C2(n12173), .A(n12172), .B(n12171), .ZN(
        n12174) );
  INV_X1 U15252 ( .A(n12174), .ZN(n12183) );
  NAND2_X1 U15253 ( .A1(n9822), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12176) );
  NAND2_X1 U15254 ( .A1(n12610), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12175) );
  NAND2_X1 U15255 ( .A1(n12176), .A2(n12175), .ZN(n12181) );
  INV_X1 U15256 ( .A(n12988), .ZN(n12177) );
  NAND2_X1 U15257 ( .A1(n12177), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12179) );
  NAND2_X1 U15258 ( .A1(n12348), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12178) );
  NAND2_X1 U15259 ( .A1(n12179), .A2(n12178), .ZN(n12180) );
  NOR2_X1 U15260 ( .A1(n12181), .A2(n12180), .ZN(n12182) );
  INV_X1 U15261 ( .A(n12243), .ZN(n12187) );
  NAND2_X1 U15262 ( .A1(n12241), .A2(n12239), .ZN(n12204) );
  AND2_X2 U15263 ( .A1(n13587), .A2(n12241), .ZN(n12221) );
  AOI22_X1 U15264 ( .A1(n12797), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15265 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12348), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15266 ( .A1(n9822), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15267 ( .A1(n9944), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12190) );
  INV_X1 U15268 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12196) );
  NAND2_X1 U15269 ( .A1(n12855), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12195) );
  NAND2_X1 U15270 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12194) );
  OAI211_X1 U15271 ( .C1(n12516), .C2(n12196), .A(n12195), .B(n12194), .ZN(
        n12197) );
  INV_X1 U15272 ( .A(n12197), .ZN(n12202) );
  AOI22_X1 U15273 ( .A1(n12880), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9958), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U15274 ( .A1(n12998), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12200) );
  NAND2_X1 U15275 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12199) );
  INV_X1 U15276 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12209) );
  NAND2_X1 U15277 ( .A1(n12855), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12208) );
  NAND2_X1 U15278 ( .A1(n12223), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12207) );
  OAI211_X1 U15279 ( .C1(n12516), .C2(n12209), .A(n12208), .B(n12207), .ZN(
        n12210) );
  INV_X1 U15280 ( .A(n12210), .ZN(n12214) );
  INV_X4 U15281 ( .A(n12961), .ZN(n12915) );
  AOI22_X1 U15282 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9958), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12213) );
  NAND2_X1 U15283 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12211) );
  NAND4_X1 U15284 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n12220) );
  AOI22_X1 U15285 ( .A1(n9943), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15286 ( .A1(n12797), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15287 ( .A1(n9822), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12216) );
  NAND4_X1 U15288 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12219) );
  NAND2_X1 U15289 ( .A1(n13751), .A2(n12221), .ZN(n12222) );
  AOI22_X1 U15290 ( .A1(n12880), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9958), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15291 ( .A1(n9962), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15292 ( .A1(n12797), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12223), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15293 ( .A1(n9943), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12224) );
  NAND4_X1 U15294 ( .A1(n12227), .A2(n12226), .A3(n12225), .A4(n12224), .ZN(
        n12238) );
  AOI22_X1 U15295 ( .A1(n9822), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12236) );
  INV_X1 U15296 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12230) );
  NAND2_X1 U15297 ( .A1(n12855), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12229) );
  NAND2_X1 U15298 ( .A1(n12315), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12228) );
  OAI211_X1 U15299 ( .C1(n12516), .C2(n12230), .A(n12229), .B(n12228), .ZN(
        n12231) );
  INV_X1 U15300 ( .A(n12231), .ZN(n12235) );
  NAND2_X1 U15301 ( .A1(n12808), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12233) );
  NAND4_X1 U15302 ( .A1(n12236), .A2(n12235), .A3(n12234), .A4(n12233), .ZN(
        n12237) );
  NOR2_X1 U15303 ( .A1(n12248), .A2(n12241), .ZN(n12242) );
  NAND2_X1 U15304 ( .A1(n12261), .A2(n12242), .ZN(n13415) );
  NAND2_X1 U15305 ( .A1(n13069), .A2(n13067), .ZN(n13592) );
  INV_X1 U15306 ( .A(n12248), .ZN(n13016) );
  NAND4_X1 U15307 ( .A1(n13016), .A2(n13029), .A3(n13078), .A4(n13587), .ZN(
        n14622) );
  INV_X1 U15308 ( .A(n14622), .ZN(n12244) );
  NAND2_X1 U15309 ( .A1(n12244), .A2(n13015), .ZN(n13310) );
  XNOR2_X1 U15310 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n13416) );
  OAI21_X1 U15311 ( .B1(n13310), .B2(n13416), .A(n13595), .ZN(n12245) );
  INV_X1 U15312 ( .A(n14480), .ZN(n12246) );
  NAND2_X1 U15313 ( .A1(n12221), .A2(n12246), .ZN(n13603) );
  OAI21_X1 U15314 ( .B1(n13587), .B2(n14378), .A(n13603), .ZN(n12249) );
  NAND2_X1 U15315 ( .A1(n20243), .A2(n20263), .ZN(n12262) );
  NOR2_X2 U15316 ( .A1(n12249), .A2(n13448), .ZN(n12256) );
  INV_X1 U15317 ( .A(n13881), .ZN(n13446) );
  OAI21_X1 U15318 ( .B1(n9926), .B2(n12251), .A(n13751), .ZN(n12255) );
  NAND2_X1 U15319 ( .A1(n12261), .A2(n13084), .ZN(n13442) );
  NAND2_X1 U15320 ( .A1(n13442), .A2(n12254), .ZN(n12267) );
  NOR2_X1 U15321 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13553) );
  NAND2_X1 U15322 ( .A1(n13553), .A2(n20932), .ZN(n13566) );
  NAND2_X1 U15323 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12278) );
  OAI21_X1 U15324 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n12278), .ZN(n20582) );
  NAND2_X1 U15325 ( .A1(n20849), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16150) );
  NAND2_X1 U15326 ( .A1(n16150), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12273) );
  OAI21_X1 U15327 ( .B1(n13566), .B2(n20582), .A(n12273), .ZN(n12257) );
  INV_X1 U15328 ( .A(n16150), .ZN(n12259) );
  MUX2_X1 U15329 ( .A(n12259), .B(n13566), .S(n20690), .Z(n12260) );
  AND2_X1 U15330 ( .A1(n13084), .A2(n20268), .ZN(n12265) );
  AND3_X1 U15331 ( .A1(n12262), .A2(n13553), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12263) );
  OAI211_X1 U15332 ( .C1(n12265), .C2(n13325), .A(n12264), .B(n12263), .ZN(
        n12266) );
  NAND2_X1 U15333 ( .A1(n9926), .A2(n9938), .ZN(n13607) );
  AND2_X1 U15334 ( .A1(n13607), .A2(n13603), .ZN(n13459) );
  NAND2_X1 U15335 ( .A1(n12267), .A2(n20243), .ZN(n12269) );
  NAND2_X1 U15336 ( .A1(n12269), .A2(n12268), .ZN(n12270) );
  INV_X1 U15337 ( .A(n12272), .ZN(n12275) );
  NAND2_X1 U15338 ( .A1(n12273), .A2(n10058), .ZN(n12274) );
  NAND2_X1 U15339 ( .A1(n12275), .A2(n12274), .ZN(n12276) );
  INV_X1 U15340 ( .A(n12278), .ZN(n12277) );
  NAND2_X1 U15341 ( .A1(n12277), .A2(n13020), .ZN(n20621) );
  NAND2_X1 U15342 ( .A1(n12278), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12279) );
  AND2_X1 U15343 ( .A1(n20621), .A2(n12279), .ZN(n20245) );
  NAND2_X1 U15344 ( .A1(n16150), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12281) );
  INV_X1 U15345 ( .A(n12516), .ZN(n12634) );
  INV_X1 U15346 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12287) );
  NAND2_X1 U15347 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12286) );
  NAND2_X1 U15348 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12285) );
  OAI211_X1 U15349 ( .C1(n13879), .C2(n12287), .A(n12286), .B(n12285), .ZN(
        n12288) );
  INV_X1 U15350 ( .A(n12288), .ZN(n12292) );
  AOI22_X1 U15351 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15352 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12290) );
  NAND2_X1 U15353 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12289) );
  NAND4_X1 U15354 ( .A1(n12292), .A2(n12291), .A3(n12290), .A4(n12289), .ZN(
        n12300) );
  AOI22_X1 U15355 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12298) );
  INV_X1 U15356 ( .A(n12315), .ZN(n12956) );
  INV_X2 U15357 ( .A(n12956), .ZN(n12999) );
  AOI22_X1 U15358 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15359 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15360 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12348), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12295) );
  NAND4_X1 U15361 ( .A1(n12298), .A2(n12297), .A3(n12296), .A4(n12295), .ZN(
        n12299) );
  OAI22_X2 U15362 ( .A1(n13535), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13869), 
        .B2(n12396), .ZN(n12305) );
  INV_X1 U15363 ( .A(n12397), .ZN(n12303) );
  AOI22_X1 U15364 ( .A1(n12303), .A2(n12302), .B1(n13059), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12304) );
  XNOR2_X2 U15365 ( .A(n12305), .B(n12304), .ZN(n12389) );
  INV_X1 U15366 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12985) );
  NAND2_X1 U15367 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12309) );
  NAND2_X1 U15368 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12308) );
  OAI211_X1 U15369 ( .C1(n13879), .C2(n12985), .A(n12309), .B(n12308), .ZN(
        n12310) );
  INV_X1 U15370 ( .A(n12310), .ZN(n12314) );
  AOI22_X1 U15371 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15372 ( .A1(n12997), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12312) );
  NAND2_X1 U15373 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12311) );
  NAND4_X1 U15374 ( .A1(n12314), .A2(n12313), .A3(n12312), .A4(n12311), .ZN(
        n12321) );
  AOI22_X1 U15375 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U15376 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15377 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15378 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12316) );
  NAND4_X1 U15379 ( .A1(n12319), .A2(n12318), .A3(n12317), .A4(n12316), .ZN(
        n12320) );
  INV_X1 U15380 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12788) );
  NAND2_X1 U15381 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12323) );
  NAND2_X1 U15382 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12322) );
  OAI211_X1 U15383 ( .C1(n13879), .C2(n12788), .A(n12323), .B(n12322), .ZN(
        n12324) );
  INV_X1 U15384 ( .A(n12324), .ZN(n12328) );
  AOI22_X1 U15385 ( .A1(n12702), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15386 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12348), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12326) );
  NAND2_X1 U15387 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12325) );
  NAND4_X1 U15388 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n12325), .ZN(
        n12334) );
  AOI22_X1 U15389 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U15390 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15391 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15392 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9822), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12329) );
  NAND4_X1 U15393 ( .A1(n12332), .A2(n12331), .A3(n12330), .A4(n12329), .ZN(
        n12333) );
  XNOR2_X1 U15394 ( .A(n14379), .B(n13693), .ZN(n12335) );
  NAND2_X1 U15395 ( .A1(n12335), .A2(n14376), .ZN(n12336) );
  AOI21_X1 U15396 ( .B1(n13587), .B2(n14374), .A(n20932), .ZN(n12338) );
  NAND2_X1 U15397 ( .A1(n13751), .A2(n13693), .ZN(n12337) );
  NAND2_X1 U15398 ( .A1(n14376), .A2(n14374), .ZN(n12339) );
  INV_X1 U15399 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12342) );
  NAND2_X1 U15400 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12341) );
  NAND2_X1 U15401 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12340) );
  OAI211_X1 U15402 ( .C1(n13879), .C2(n12342), .A(n12341), .B(n12340), .ZN(
        n12343) );
  INV_X1 U15403 ( .A(n12343), .ZN(n12347) );
  AOI22_X1 U15404 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9958), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15405 ( .A1(n12997), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12345) );
  NAND2_X1 U15406 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12344) );
  NAND4_X1 U15407 ( .A1(n12347), .A2(n12346), .A3(n12345), .A4(n12344), .ZN(
        n12354) );
  AOI22_X1 U15408 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15409 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15410 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15411 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12348), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12349) );
  NAND4_X1 U15412 ( .A1(n12352), .A2(n12351), .A3(n12350), .A4(n12349), .ZN(
        n12353) );
  INV_X1 U15413 ( .A(n13692), .ZN(n12357) );
  NAND2_X1 U15414 ( .A1(n13059), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12356) );
  NAND2_X1 U15415 ( .A1(n14376), .A2(n14379), .ZN(n12355) );
  OAI211_X1 U15416 ( .C1(n12397), .C2(n12357), .A(n12356), .B(n12355), .ZN(
        n12358) );
  OR2_X2 U15417 ( .A1(n12359), .A2(n12358), .ZN(n12366) );
  NAND2_X1 U15418 ( .A1(n12359), .A2(n12358), .ZN(n12360) );
  INV_X1 U15419 ( .A(n20358), .ZN(n12363) );
  INV_X1 U15420 ( .A(n12361), .ZN(n12362) );
  NAND2_X1 U15421 ( .A1(n12363), .A2(n12362), .ZN(n20297) );
  NAND2_X1 U15422 ( .A1(n14376), .A2(n13692), .ZN(n12365) );
  INV_X2 U15423 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20929) );
  NOR2_X2 U15424 ( .A1(n12239), .A2(n20929), .ZN(n12640) );
  AND2_X1 U15425 ( .A1(n13086), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12424) );
  INV_X1 U15426 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n12368) );
  NOR2_X1 U15427 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12716) );
  XNOR2_X1 U15428 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15153) );
  AOI21_X1 U15429 ( .B1(n13741), .B2(n15153), .A(n14428), .ZN(n12367) );
  OAI21_X1 U15430 ( .B1(n13010), .B2(n12368), .A(n12367), .ZN(n12369) );
  AOI21_X1 U15431 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n12424), .A(
        n12369), .ZN(n12370) );
  NAND2_X1 U15432 ( .A1(n14428), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12387) );
  INV_X1 U15433 ( .A(n13772), .ZN(n12386) );
  INV_X1 U15434 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n12372) );
  INV_X1 U15435 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13767) );
  OAI22_X1 U15436 ( .A1(n13010), .A2(n12372), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13767), .ZN(n12373) );
  AOI21_X1 U15437 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n12424), .A(
        n12373), .ZN(n12374) );
  NAND2_X1 U15438 ( .A1(n12375), .A2(n12374), .ZN(n13688) );
  NAND2_X1 U15439 ( .A1(n13562), .A2(n13604), .ZN(n12377) );
  NAND2_X1 U15440 ( .A1(n12377), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13556) );
  INV_X1 U15441 ( .A(n12424), .ZN(n12445) );
  NAND2_X1 U15442 ( .A1(n14429), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12380) );
  NAND2_X1 U15443 ( .A1(n20929), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12379) );
  OAI211_X1 U15444 ( .C1(n12445), .C2(n12381), .A(n12380), .B(n12379), .ZN(
        n12382) );
  AOI21_X1 U15445 ( .B1(n12378), .B2(n12640), .A(n12382), .ZN(n12383) );
  OR2_X1 U15446 ( .A1(n13556), .A2(n12383), .ZN(n13557) );
  INV_X1 U15447 ( .A(n12383), .ZN(n13558) );
  INV_X1 U15448 ( .A(n12716), .ZN(n12982) );
  OR2_X1 U15449 ( .A1(n13558), .A2(n12982), .ZN(n12384) );
  NAND2_X1 U15450 ( .A1(n13557), .A2(n12384), .ZN(n13687) );
  NAND2_X1 U15451 ( .A1(n13688), .A2(n13687), .ZN(n13686) );
  OR2_X1 U15452 ( .A1(n12280), .A2(n12088), .ZN(n12395) );
  INV_X1 U15453 ( .A(n13566), .ZN(n12393) );
  NAND2_X1 U15454 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10313), .ZN(
        n20514) );
  NAND2_X1 U15455 ( .A1(n20658), .A2(n20514), .ZN(n12392) );
  NOR3_X1 U15456 ( .A1(n20658), .A2(n13020), .A3(n20585), .ZN(n20791) );
  NAND2_X1 U15457 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20791), .ZN(
        n20831) );
  AND2_X1 U15458 ( .A1(n12392), .A2(n20831), .ZN(n20529) );
  AOI22_X1 U15459 ( .A1(n12393), .A2(n20529), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16150), .ZN(n12394) );
  XNOR2_X2 U15460 ( .A(n12391), .B(n20400), .ZN(n20527) );
  INV_X1 U15461 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12400) );
  NAND2_X1 U15462 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12399) );
  NAND2_X1 U15463 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12398) );
  OAI211_X1 U15464 ( .C1(n13879), .C2(n12400), .A(n12399), .B(n12398), .ZN(
        n12401) );
  INV_X1 U15465 ( .A(n12401), .ZN(n12405) );
  AOI22_X1 U15466 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15467 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12403) );
  NAND2_X1 U15468 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12402) );
  NAND4_X1 U15469 ( .A1(n12405), .A2(n12404), .A3(n12403), .A4(n12402), .ZN(
        n12411) );
  AOI22_X1 U15470 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U15471 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15472 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12407) );
  INV_X2 U15473 ( .A(n12102), .ZN(n12968) );
  AOI22_X1 U15474 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12406) );
  NAND4_X1 U15475 ( .A1(n12409), .A2(n12408), .A3(n12407), .A4(n12406), .ZN(
        n12410) );
  AOI22_X1 U15476 ( .A1(n13034), .A2(n14349), .B1(n13059), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12412) );
  INV_X1 U15477 ( .A(n12414), .ZN(n12415) );
  INV_X1 U15478 ( .A(n13920), .ZN(n13919) );
  NAND2_X1 U15479 ( .A1(n12415), .A2(n13919), .ZN(n12416) );
  INV_X1 U15480 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n12422) );
  INV_X1 U15481 ( .A(n12418), .ZN(n12420) );
  INV_X1 U15482 ( .A(n12466), .ZN(n12419) );
  OAI21_X1 U15483 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12420), .A(
        n12419), .ZN(n13979) );
  AOI22_X1 U15484 ( .A1(n13741), .A2(n13979), .B1(n14428), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12421) );
  OAI21_X1 U15485 ( .B1(n13010), .B2(n12422), .A(n12421), .ZN(n12423) );
  AOI21_X1 U15486 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12424), .A(
        n12423), .ZN(n12425) );
  INV_X1 U15487 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12428) );
  NAND2_X1 U15488 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12427) );
  NAND2_X1 U15489 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12426) );
  OAI211_X1 U15490 ( .C1(n13879), .C2(n12428), .A(n12427), .B(n12426), .ZN(
        n12429) );
  INV_X1 U15491 ( .A(n12429), .ZN(n12433) );
  AOI22_X1 U15492 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12915), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15493 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12431) );
  NAND2_X1 U15494 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12430) );
  NAND4_X1 U15495 ( .A1(n12433), .A2(n12432), .A3(n12431), .A4(n12430), .ZN(
        n12440) );
  AOI22_X1 U15496 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n9961), .B1(
        n12702), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15497 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12753), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15498 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15499 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n9944), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12435) );
  NAND4_X1 U15500 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        n12439) );
  NAND2_X1 U15501 ( .A1(n13034), .A2(n14348), .ZN(n12442) );
  NAND2_X1 U15502 ( .A1(n13059), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12441) );
  NAND2_X1 U15503 ( .A1(n12442), .A2(n12441), .ZN(n12450) );
  XNOR2_X1 U15504 ( .A(n12449), .B(n12450), .ZN(n14341) );
  NAND2_X1 U15505 ( .A1(n14341), .A2(n12640), .ZN(n12448) );
  XNOR2_X1 U15506 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B(n12466), .ZN(
        n20192) );
  INV_X1 U15507 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13496) );
  INV_X1 U15508 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21085) );
  OAI21_X1 U15509 ( .B1(n21085), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20929), .ZN(n12444) );
  NAND2_X1 U15510 ( .A1(n14429), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12443) );
  OAI211_X1 U15511 ( .C1(n12445), .C2(n13496), .A(n12444), .B(n12443), .ZN(
        n12446) );
  OAI21_X1 U15512 ( .B1(n12982), .B2(n20192), .A(n12446), .ZN(n12447) );
  INV_X1 U15513 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12938) );
  NAND2_X1 U15514 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12452) );
  NAND2_X1 U15515 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12451) );
  OAI211_X1 U15516 ( .C1(n13879), .C2(n12938), .A(n12452), .B(n12451), .ZN(
        n12453) );
  INV_X1 U15517 ( .A(n12453), .ZN(n12457) );
  AOI22_X1 U15518 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U15519 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12455) );
  NAND2_X1 U15520 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12454) );
  NAND4_X1 U15521 ( .A1(n12457), .A2(n12456), .A3(n12455), .A4(n12454), .ZN(
        n12463) );
  AOI22_X1 U15522 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12461) );
  AOI22_X1 U15523 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U15524 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U15525 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12458) );
  NAND4_X1 U15526 ( .A1(n12461), .A2(n12460), .A3(n12459), .A4(n12458), .ZN(
        n12462) );
  NAND2_X1 U15527 ( .A1(n13034), .A2(n14359), .ZN(n12465) );
  NAND2_X1 U15528 ( .A1(n13059), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12464) );
  NAND2_X1 U15529 ( .A1(n12465), .A2(n12464), .ZN(n12476) );
  XNOR2_X1 U15530 ( .A(n12475), .B(n12476), .ZN(n14347) );
  NAND2_X1 U15531 ( .A1(n14347), .A2(n12640), .ZN(n12474) );
  INV_X1 U15532 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12471) );
  INV_X1 U15533 ( .A(n12492), .ZN(n12494) );
  INV_X1 U15534 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12468) );
  NAND2_X1 U15535 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12466), .ZN(
        n12467) );
  NAND2_X1 U15536 ( .A1(n12468), .A2(n12467), .ZN(n12469) );
  NAND2_X1 U15537 ( .A1(n12494), .A2(n12469), .ZN(n20124) );
  AOI22_X1 U15538 ( .A1(n20124), .A2(n13741), .B1(n14428), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12470) );
  OAI21_X1 U15539 ( .B1(n13010), .B2(n12471), .A(n12470), .ZN(n12472) );
  INV_X1 U15540 ( .A(n12472), .ZN(n12473) );
  NAND2_X1 U15541 ( .A1(n12474), .A2(n12473), .ZN(n13988) );
  NAND2_X1 U15542 ( .A1(n13985), .A2(n13988), .ZN(n13986) );
  INV_X1 U15543 ( .A(n13986), .ZN(n12500) );
  INV_X1 U15544 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12480) );
  NAND2_X1 U15545 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12479) );
  NAND2_X1 U15546 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12478) );
  OAI211_X1 U15547 ( .C1(n13879), .C2(n12480), .A(n12479), .B(n12478), .ZN(
        n12481) );
  INV_X1 U15548 ( .A(n12481), .ZN(n12485) );
  AOI22_X1 U15549 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12484) );
  AOI22_X1 U15550 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12483) );
  NAND2_X1 U15551 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12482) );
  NAND4_X1 U15552 ( .A1(n12485), .A2(n12484), .A3(n12483), .A4(n12482), .ZN(
        n12491) );
  AOI22_X1 U15553 ( .A1(n9944), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U15554 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15555 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15556 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12486) );
  NAND4_X1 U15557 ( .A1(n12489), .A2(n12488), .A3(n12487), .A4(n12486), .ZN(
        n12490) );
  AOI22_X1 U15558 ( .A1(n13034), .A2(n14368), .B1(n13059), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12501) );
  INV_X1 U15559 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20156) );
  INV_X1 U15560 ( .A(n12505), .ZN(n12496) );
  INV_X1 U15561 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12493) );
  NAND2_X1 U15562 ( .A1(n12494), .A2(n12493), .ZN(n12495) );
  NAND2_X1 U15563 ( .A1(n12496), .A2(n12495), .ZN(n20110) );
  AOI22_X1 U15564 ( .A1(n20110), .A2(n12716), .B1(n14428), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12497) );
  OAI21_X1 U15565 ( .B1(n13010), .B2(n20156), .A(n12497), .ZN(n12498) );
  INV_X1 U15566 ( .A(n14092), .ZN(n12499) );
  NAND2_X1 U15567 ( .A1(n12500), .A2(n12499), .ZN(n14161) );
  NAND2_X1 U15568 ( .A1(n13034), .A2(n14374), .ZN(n12503) );
  NAND2_X1 U15569 ( .A1(n13059), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12502) );
  NAND2_X1 U15570 ( .A1(n12503), .A2(n12502), .ZN(n12504) );
  INV_X1 U15571 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n14184) );
  OAI21_X1 U15572 ( .B1(n12505), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n12522), .ZN(n20098) );
  AOI22_X1 U15573 ( .A1(n20098), .A2(n12716), .B1(n14428), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12506) );
  OAI21_X1 U15574 ( .B1(n13010), .B2(n14184), .A(n12506), .ZN(n12507) );
  AOI21_X1 U15575 ( .B1(n14366), .B2(n12640), .A(n12507), .ZN(n14160) );
  NAND2_X1 U15576 ( .A1(n14429), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U15577 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12512) );
  AOI22_X1 U15578 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U15579 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12510) );
  AOI22_X1 U15580 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12509) );
  AND4_X1 U15581 ( .A1(n12512), .A2(n12511), .A3(n12510), .A4(n12509), .ZN(
        n12520) );
  AOI22_X1 U15582 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U15583 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9922), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12514) );
  NAND2_X1 U15584 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12513) );
  AND3_X1 U15585 ( .A1(n12515), .A2(n12514), .A3(n12513), .ZN(n12519) );
  AOI22_X1 U15586 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12518) );
  NAND2_X1 U15587 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12517) );
  NAND4_X1 U15588 ( .A1(n12520), .A2(n12519), .A3(n12518), .A4(n12517), .ZN(
        n12521) );
  NAND2_X1 U15589 ( .A1(n12640), .A2(n12521), .ZN(n12524) );
  XNOR2_X1 U15590 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12527), .ZN(
        n14833) );
  AOI22_X1 U15591 ( .A1(n12716), .A2(n14833), .B1(n14428), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12523) );
  XOR2_X1 U15592 ( .A(n20073), .B(n12556), .Z(n20085) );
  AOI22_X1 U15593 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9961), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U15594 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12530) );
  AOI22_X1 U15595 ( .A1(n9944), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15596 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12528) );
  AND4_X1 U15597 ( .A1(n12531), .A2(n12530), .A3(n12529), .A4(n12528), .ZN(
        n12538) );
  AOI22_X1 U15598 ( .A1(n12997), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U15599 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12533) );
  NAND2_X1 U15600 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12532) );
  AND3_X1 U15601 ( .A1(n12534), .A2(n12533), .A3(n12532), .ZN(n12537) );
  AOI22_X1 U15602 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12536) );
  NAND2_X1 U15603 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12535) );
  NAND4_X1 U15604 ( .A1(n12538), .A2(n12537), .A3(n12536), .A4(n12535), .ZN(
        n12539) );
  AOI22_X1 U15605 ( .A1(n12640), .A2(n12539), .B1(n14428), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12541) );
  NAND2_X1 U15606 ( .A1(n14429), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12540) );
  OAI211_X1 U15607 ( .C1(n20085), .C2(n12982), .A(n12541), .B(n12540), .ZN(
        n14233) );
  INV_X1 U15608 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12544) );
  NAND2_X1 U15609 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12543) );
  NAND2_X1 U15610 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12542) );
  OAI211_X1 U15611 ( .C1(n13879), .C2(n12544), .A(n12543), .B(n12542), .ZN(
        n12545) );
  INV_X1 U15612 ( .A(n12545), .ZN(n12549) );
  AOI22_X1 U15613 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15614 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U15615 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12546) );
  NAND4_X1 U15616 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12555) );
  AOI22_X1 U15617 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15618 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U15619 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U15620 ( .A1(n9944), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12550) );
  NAND4_X1 U15621 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12554) );
  NOR2_X1 U15622 ( .A1(n12555), .A2(n12554), .ZN(n12559) );
  XNOR2_X1 U15623 ( .A(n12560), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15144) );
  NAND2_X1 U15624 ( .A1(n15144), .A2(n12716), .ZN(n12558) );
  AOI22_X1 U15625 ( .A1(n14429), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n14428), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12557) );
  OAI211_X1 U15626 ( .C1(n12559), .C2(n10283), .A(n12558), .B(n12557), .ZN(
        n14309) );
  INV_X1 U15627 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12564) );
  INV_X1 U15628 ( .A(n14428), .ZN(n12563) );
  OAI21_X1 U15629 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12561), .A(
        n12590), .ZN(n16283) );
  NAND2_X1 U15630 ( .A1(n16283), .A2(n12716), .ZN(n12562) );
  OAI21_X1 U15631 ( .B1(n12564), .B2(n12563), .A(n12562), .ZN(n12565) );
  AOI21_X1 U15632 ( .B1(n14429), .B2(P1_EAX_REG_11__SCAN_IN), .A(n12565), .ZN(
        n14810) );
  AOI22_X1 U15633 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15634 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15635 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U15636 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12566) );
  AND4_X1 U15637 ( .A1(n12569), .A2(n12568), .A3(n12567), .A4(n12566), .ZN(
        n12576) );
  AOI22_X1 U15638 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12572) );
  AOI22_X1 U15639 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12571) );
  NAND2_X1 U15640 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12570) );
  AND3_X1 U15641 ( .A1(n12572), .A2(n12571), .A3(n12570), .ZN(n12575) );
  AOI22_X1 U15642 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12574) );
  NAND2_X1 U15643 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12573) );
  NAND4_X1 U15644 ( .A1(n12576), .A2(n12575), .A3(n12574), .A4(n12573), .ZN(
        n12577) );
  NAND2_X1 U15645 ( .A1(n12640), .A2(n12577), .ZN(n14900) );
  INV_X1 U15646 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14981) );
  AOI22_X1 U15647 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15648 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12751), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15649 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15650 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12915), .B1(
        n12610), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12578) );
  AND4_X1 U15651 ( .A1(n12581), .A2(n12580), .A3(n12579), .A4(n12578), .ZN(
        n12588) );
  AOI22_X1 U15652 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12997), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U15653 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n9961), .B1(n9922), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12583) );
  NAND2_X1 U15654 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12582) );
  AND3_X1 U15655 ( .A1(n12584), .A2(n12583), .A3(n12582), .ZN(n12587) );
  AOI22_X1 U15656 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12993), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U15657 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12585) );
  NAND4_X1 U15658 ( .A1(n12588), .A2(n12587), .A3(n12586), .A4(n12585), .ZN(
        n12589) );
  NAND2_X1 U15659 ( .A1(n12640), .A2(n12589), .ZN(n12593) );
  XOR2_X1 U15660 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12623), .Z(
        n16240) );
  INV_X1 U15661 ( .A(n16240), .ZN(n12591) );
  AOI22_X1 U15662 ( .A1(n14428), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n12716), .B2(n12591), .ZN(n12592) );
  OAI211_X1 U15663 ( .C1(n14981), .C2(n13010), .A(n12593), .B(n12592), .ZN(
        n14895) );
  INV_X1 U15664 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14977) );
  AOI22_X1 U15665 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15666 ( .A1(n12997), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15667 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15668 ( .A1(n9944), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12594) );
  AND4_X1 U15669 ( .A1(n12597), .A2(n12596), .A3(n12595), .A4(n12594), .ZN(
        n12604) );
  AOI22_X1 U15670 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12603) );
  AOI22_X1 U15671 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U15672 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12599) );
  NAND2_X1 U15673 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12598) );
  AND3_X1 U15674 ( .A1(n12600), .A2(n12599), .A3(n12598), .ZN(n12602) );
  NAND2_X1 U15675 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12601) );
  NAND4_X1 U15676 ( .A1(n12604), .A2(n12603), .A3(n12602), .A4(n12601), .ZN(
        n12605) );
  NAND2_X1 U15677 ( .A1(n12640), .A2(n12605), .ZN(n12608) );
  INV_X1 U15678 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14824) );
  NAND2_X1 U15679 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n12623), .ZN(
        n12606) );
  XNOR2_X1 U15680 ( .A(n14824), .B(n12606), .ZN(n15123) );
  AOI22_X1 U15681 ( .A1(n15123), .A2(n12716), .B1(n14428), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12607) );
  OAI211_X1 U15682 ( .C1(n13010), .C2(n14977), .A(n12608), .B(n12607), .ZN(
        n14814) );
  NAND2_X1 U15683 ( .A1(n14895), .A2(n14814), .ZN(n12609) );
  AOI21_X4 U15684 ( .B1(n14812), .B2(n9979), .A(n12609), .ZN(n14815) );
  INV_X1 U15685 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14974) );
  AOI22_X1 U15686 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U15687 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9957), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U15688 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U15689 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12611) );
  AND4_X1 U15690 ( .A1(n12614), .A2(n12613), .A3(n12612), .A4(n12611), .ZN(
        n12621) );
  AOI22_X1 U15691 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15692 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12616) );
  NAND2_X1 U15693 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12615) );
  AND3_X1 U15694 ( .A1(n12617), .A2(n12616), .A3(n12615), .ZN(n12620) );
  AOI22_X1 U15695 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12619) );
  NAND2_X1 U15696 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12618) );
  NAND4_X1 U15697 ( .A1(n12621), .A2(n12620), .A3(n12619), .A4(n12618), .ZN(
        n12622) );
  NAND2_X1 U15698 ( .A1(n12640), .A2(n12622), .ZN(n12625) );
  XNOR2_X1 U15699 ( .A(n12626), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15110) );
  AOI22_X1 U15700 ( .A1(n15110), .A2(n13741), .B1(n14428), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12624) );
  OAI211_X1 U15701 ( .C1(n13010), .C2(n14974), .A(n12625), .B(n12624), .ZN(
        n14796) );
  INV_X1 U15702 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16230) );
  XOR2_X1 U15703 ( .A(n16230), .B(n12643), .Z(n16271) );
  AOI22_X1 U15704 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12915), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U15705 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15706 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12628) );
  AOI22_X1 U15707 ( .A1(n9944), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12627) );
  AND4_X1 U15708 ( .A1(n12630), .A2(n12629), .A3(n12628), .A4(n12627), .ZN(
        n12638) );
  AOI22_X1 U15709 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U15710 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12632) );
  NAND2_X1 U15711 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12631) );
  AND3_X1 U15712 ( .A1(n12633), .A2(n12632), .A3(n12631), .ZN(n12637) );
  AOI22_X1 U15713 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12636) );
  NAND2_X1 U15714 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12635) );
  NAND4_X1 U15715 ( .A1(n12638), .A2(n12637), .A3(n12636), .A4(n12635), .ZN(
        n12639) );
  AOI22_X1 U15716 ( .A1(n12640), .A2(n12639), .B1(n14428), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12642) );
  NAND2_X1 U15717 ( .A1(n14429), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12641) );
  OAI211_X1 U15718 ( .C1(n16271), .C2(n12982), .A(n12642), .B(n12641), .ZN(
        n14883) );
  INV_X1 U15719 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12697) );
  XNOR2_X1 U15720 ( .A(n12739), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16194) );
  INV_X1 U15721 ( .A(n12254), .ZN(n13461) );
  NAND2_X1 U15722 ( .A1(n13461), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12979) );
  NAND2_X1 U15723 ( .A1(n12979), .A2(n12982), .ZN(n12732) );
  AOI22_X1 U15724 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9945), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12649) );
  NAND2_X1 U15725 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12645) );
  NAND2_X1 U15726 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12644) );
  AND3_X1 U15727 ( .A1(n12645), .A2(n12644), .A3(n12982), .ZN(n12648) );
  AOI22_X1 U15728 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12753), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U15729 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12752), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12646) );
  NAND4_X1 U15730 ( .A1(n12649), .A2(n12648), .A3(n12647), .A4(n12646), .ZN(
        n12655) );
  AOI22_X1 U15731 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U15732 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n9957), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U15733 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U15734 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12993), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12650) );
  NAND4_X1 U15735 ( .A1(n12653), .A2(n12652), .A3(n12651), .A4(n12650), .ZN(
        n12654) );
  OR2_X1 U15736 ( .A1(n12655), .A2(n12654), .ZN(n12657) );
  INV_X1 U15737 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14947) );
  INV_X1 U15738 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16192) );
  OAI22_X1 U15739 ( .A1(n13010), .A2(n14947), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n16192), .ZN(n12656) );
  AOI21_X1 U15740 ( .B1(n12732), .B2(n12657), .A(n12656), .ZN(n12658) );
  AOI21_X1 U15741 ( .B1(n16194), .B2(n13741), .A(n12658), .ZN(n14860) );
  INV_X1 U15742 ( .A(n14860), .ZN(n12719) );
  OAI21_X1 U15743 ( .B1(n12659), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n12739), .ZN(n15084) );
  OR2_X1 U15744 ( .A1(n15084), .A2(n12982), .ZN(n12678) );
  INV_X1 U15745 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12662) );
  NAND2_X1 U15746 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12661) );
  NAND2_X1 U15747 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12660) );
  OAI211_X1 U15748 ( .C1(n13879), .C2(n12662), .A(n12661), .B(n12660), .ZN(
        n12663) );
  INV_X1 U15749 ( .A(n12663), .ZN(n12667) );
  AOI22_X1 U15750 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12666) );
  AOI22_X1 U15751 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12665) );
  NAND2_X1 U15752 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12664) );
  NAND4_X1 U15753 ( .A1(n12667), .A2(n12666), .A3(n12665), .A4(n12664), .ZN(
        n12673) );
  AOI22_X1 U15754 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U15755 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12670) );
  AOI22_X1 U15756 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U15757 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12668) );
  NAND4_X1 U15758 ( .A1(n12671), .A2(n12670), .A3(n12669), .A4(n12668), .ZN(
        n12672) );
  NOR2_X1 U15759 ( .A1(n12673), .A2(n12672), .ZN(n12676) );
  OAI21_X1 U15760 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n21085), .A(
        n20929), .ZN(n12675) );
  NAND2_X1 U15761 ( .A1(n14429), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n12674) );
  OAI211_X1 U15762 ( .C1(n12979), .C2(n12676), .A(n12675), .B(n12674), .ZN(
        n12677) );
  AND2_X1 U15763 ( .A1(n12678), .A2(n12677), .ZN(n14769) );
  INV_X1 U15764 ( .A(n14769), .ZN(n12718) );
  INV_X1 U15765 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15091) );
  XNOR2_X1 U15766 ( .A(n12679), .B(n15091), .ZN(n16207) );
  NAND2_X1 U15767 ( .A1(n16207), .A2(n12716), .ZN(n12695) );
  AOI22_X1 U15768 ( .A1(n9944), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12915), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U15769 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U15770 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U15771 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12680) );
  NAND4_X1 U15772 ( .A1(n12683), .A2(n12682), .A3(n12681), .A4(n12680), .ZN(
        n12691) );
  AOI22_X1 U15773 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9945), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12689) );
  NAND2_X1 U15774 ( .A1(n12997), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12685) );
  NAND2_X1 U15775 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12684) );
  AND3_X1 U15776 ( .A1(n12685), .A2(n12684), .A3(n12982), .ZN(n12688) );
  AOI22_X1 U15777 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U15778 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12686) );
  NAND4_X1 U15779 ( .A1(n12689), .A2(n12688), .A3(n12687), .A4(n12686), .ZN(
        n12690) );
  OAI21_X1 U15780 ( .B1(n12691), .B2(n12690), .A(n12732), .ZN(n12693) );
  AOI22_X1 U15781 ( .A1(n14429), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20929), .ZN(n12692) );
  NAND2_X1 U15782 ( .A1(n12693), .A2(n12692), .ZN(n12694) );
  NAND2_X1 U15783 ( .A1(n12695), .A2(n12694), .ZN(n14866) );
  XOR2_X1 U15784 ( .A(n12697), .B(n12696), .Z(n16259) );
  INV_X1 U15785 ( .A(n16259), .ZN(n12717) );
  INV_X1 U15786 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12700) );
  NAND2_X1 U15787 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12699) );
  NAND2_X1 U15788 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12698) );
  OAI211_X1 U15789 ( .C1(n13879), .C2(n12700), .A(n12699), .B(n12698), .ZN(
        n12701) );
  INV_X1 U15790 ( .A(n12701), .ZN(n12706) );
  AOI22_X1 U15791 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15792 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9922), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12704) );
  NAND2_X1 U15793 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12703) );
  NAND4_X1 U15794 ( .A1(n12706), .A2(n12705), .A3(n12704), .A4(n12703), .ZN(
        n12712) );
  AOI22_X1 U15795 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12710) );
  AOI22_X1 U15796 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U15797 ( .A1(n9815), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U15798 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12707) );
  NAND4_X1 U15799 ( .A1(n12710), .A2(n12709), .A3(n12708), .A4(n12707), .ZN(
        n12711) );
  NOR2_X1 U15800 ( .A1(n12712), .A2(n12711), .ZN(n12714) );
  AOI22_X1 U15801 ( .A1(n14429), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n14428), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12713) );
  OAI21_X1 U15802 ( .B1(n12979), .B2(n12714), .A(n12713), .ZN(n12715) );
  AOI21_X1 U15803 ( .B1(n12717), .B2(n12716), .A(n12715), .ZN(n14787) );
  OR2_X1 U15804 ( .A1(n14866), .A2(n14787), .ZN(n14768) );
  INV_X1 U15805 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12720) );
  XNOR2_X1 U15806 ( .A(n12721), .B(n12720), .ZN(n16217) );
  NAND2_X1 U15807 ( .A1(n16217), .A2(n13741), .ZN(n12738) );
  AOI22_X1 U15808 ( .A1(n9944), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15809 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15810 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U15811 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12722) );
  NAND4_X1 U15812 ( .A1(n12725), .A2(n12724), .A3(n12723), .A4(n12722), .ZN(
        n12734) );
  AOI22_X1 U15813 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9945), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12731) );
  NAND2_X1 U15814 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12727) );
  NAND2_X1 U15815 ( .A1(n9957), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12726) );
  AND3_X1 U15816 ( .A1(n12727), .A2(n12726), .A3(n12982), .ZN(n12730) );
  AOI22_X1 U15817 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15818 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12728) );
  NAND4_X1 U15819 ( .A1(n12731), .A2(n12730), .A3(n12729), .A4(n12728), .ZN(
        n12733) );
  OAI21_X1 U15820 ( .B1(n12734), .B2(n12733), .A(n12732), .ZN(n12736) );
  AOI22_X1 U15821 ( .A1(n14429), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20929), .ZN(n12735) );
  NAND2_X1 U15822 ( .A1(n12736), .A2(n12735), .ZN(n12737) );
  NAND2_X1 U15823 ( .A1(n12738), .A2(n12737), .ZN(n14872) );
  INV_X1 U15824 ( .A(n12740), .ZN(n12741) );
  INV_X1 U15825 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16184) );
  NAND2_X1 U15826 ( .A1(n12741), .A2(n16184), .ZN(n12742) );
  NAND2_X1 U15827 ( .A1(n12785), .A2(n12742), .ZN(n16191) );
  OR2_X1 U15828 ( .A1(n16191), .A2(n12982), .ZN(n12764) );
  INV_X1 U15829 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12745) );
  NAND2_X1 U15830 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12744) );
  NAND2_X1 U15831 ( .A1(n12999), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12743) );
  OAI211_X1 U15832 ( .C1(n13879), .C2(n12745), .A(n12744), .B(n12743), .ZN(
        n12746) );
  INV_X1 U15833 ( .A(n12746), .ZN(n12750) );
  AOI22_X1 U15834 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U15835 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12748) );
  NAND2_X1 U15836 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12747) );
  NAND4_X1 U15837 ( .A1(n12750), .A2(n12749), .A3(n12748), .A4(n12747), .ZN(
        n12759) );
  AOI22_X1 U15838 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13000), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U15839 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U15840 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15841 ( .A1(n12997), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12754) );
  NAND4_X1 U15842 ( .A1(n12757), .A2(n12756), .A3(n12755), .A4(n12754), .ZN(
        n12758) );
  NOR2_X1 U15843 ( .A1(n12759), .A2(n12758), .ZN(n12762) );
  OAI21_X1 U15844 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n21085), .A(
        n20929), .ZN(n12761) );
  NAND2_X1 U15845 ( .A1(n14429), .A2(P1_EAX_REG_21__SCAN_IN), .ZN(n12760) );
  OAI211_X1 U15846 ( .C1(n12979), .C2(n12762), .A(n12761), .B(n12760), .ZN(
        n12763) );
  XNOR2_X1 U15847 ( .A(n12785), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15063) );
  NAND2_X1 U15848 ( .A1(n15063), .A2(n13741), .ZN(n12783) );
  INV_X1 U15849 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12767) );
  NAND2_X1 U15850 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12766) );
  NAND2_X1 U15851 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12765) );
  OAI211_X1 U15852 ( .C1(n13879), .C2(n12767), .A(n12766), .B(n12765), .ZN(
        n12768) );
  INV_X1 U15853 ( .A(n12768), .ZN(n12772) );
  AOI22_X1 U15854 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U15855 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12770) );
  NAND2_X1 U15856 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12769) );
  NAND4_X1 U15857 ( .A1(n12772), .A2(n12771), .A3(n12770), .A4(n12769), .ZN(
        n12778) );
  AOI22_X1 U15858 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n9957), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12776) );
  AOI22_X1 U15859 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12775) );
  AOI22_X1 U15860 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12774) );
  AOI22_X1 U15861 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12773) );
  NAND4_X1 U15862 ( .A1(n12776), .A2(n12775), .A3(n12774), .A4(n12773), .ZN(
        n12777) );
  NOR2_X1 U15863 ( .A1(n12778), .A2(n12777), .ZN(n12781) );
  INV_X1 U15864 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15061) );
  AOI21_X1 U15865 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15061), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12779) );
  AOI21_X1 U15866 ( .B1(n14429), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12779), .ZN(
        n12780) );
  OAI21_X1 U15867 ( .B1(n12979), .B2(n12781), .A(n12780), .ZN(n12782) );
  NAND2_X1 U15868 ( .A1(n12783), .A2(n12782), .ZN(n14757) );
  INV_X1 U15869 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14746) );
  NAND2_X1 U15870 ( .A1(n12786), .A2(n14746), .ZN(n12787) );
  NAND2_X1 U15871 ( .A1(n12843), .A2(n12787), .ZN(n15053) );
  INV_X1 U15872 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12796) );
  INV_X1 U15873 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12789) );
  OAI22_X1 U15874 ( .A1(n12956), .A2(n12789), .B1(n12986), .B2(n12788), .ZN(
        n12793) );
  INV_X1 U15875 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12791) );
  INV_X1 U15876 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12790) );
  OAI22_X1 U15877 ( .A1(n9820), .A2(n12791), .B1(n12907), .B2(n12790), .ZN(
        n12792) );
  AOI211_X1 U15878 ( .C1(n9945), .C2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n12793), .B(n12792), .ZN(n12795) );
  AOI22_X1 U15879 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12794) );
  OAI211_X1 U15880 ( .C1(n13879), .C2(n12796), .A(n12795), .B(n12794), .ZN(
        n12803) );
  AOI22_X1 U15881 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U15882 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12800) );
  AOI22_X1 U15883 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U15884 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12798) );
  NAND4_X1 U15885 ( .A1(n12801), .A2(n12800), .A3(n12799), .A4(n12798), .ZN(
        n12802) );
  NOR2_X1 U15886 ( .A1(n12803), .A2(n12802), .ZN(n12823) );
  INV_X1 U15887 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12811) );
  INV_X1 U15888 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12804) );
  OAI22_X1 U15889 ( .A1(n12850), .A2(n12804), .B1(n12434), .B2(n12985), .ZN(
        n12807) );
  INV_X1 U15890 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12990) );
  INV_X1 U15891 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12805) );
  OAI22_X1 U15892 ( .A1(n12961), .A2(n12990), .B1(n9820), .B2(n12805), .ZN(
        n12806) );
  AOI211_X1 U15893 ( .C1(n9945), .C2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n12807), .B(n12806), .ZN(n12810) );
  AOI22_X1 U15894 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12993), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12809) );
  OAI211_X1 U15895 ( .C1(n13879), .C2(n12811), .A(n12810), .B(n12809), .ZN(
        n12817) );
  AOI22_X1 U15896 ( .A1(n12997), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12815) );
  AOI22_X1 U15897 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U15898 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U15899 ( .A1(n9952), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12812) );
  NAND4_X1 U15900 ( .A1(n12815), .A2(n12814), .A3(n12813), .A4(n12812), .ZN(
        n12816) );
  NOR2_X1 U15901 ( .A1(n12817), .A2(n12816), .ZN(n12822) );
  XNOR2_X1 U15902 ( .A(n12823), .B(n12822), .ZN(n12820) );
  AOI21_X1 U15903 ( .B1(n14746), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12818) );
  AOI21_X1 U15904 ( .B1(n14429), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12818), .ZN(
        n12819) );
  OAI21_X1 U15905 ( .B1(n12820), .B2(n12979), .A(n12819), .ZN(n12821) );
  OAI21_X1 U15906 ( .B1(n15053), .B2(n12982), .A(n12821), .ZN(n14744) );
  XNOR2_X1 U15907 ( .A(n12843), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15048) );
  NOR2_X1 U15908 ( .A1(n12823), .A2(n12822), .ZN(n12867) );
  INV_X1 U15909 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U15910 ( .A1(n12855), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12825) );
  NAND2_X1 U15911 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12824) );
  OAI211_X1 U15912 ( .C1(n13879), .C2(n12826), .A(n12825), .B(n12824), .ZN(
        n12827) );
  INV_X1 U15913 ( .A(n12827), .ZN(n12831) );
  AOI22_X1 U15914 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12830) );
  AOI22_X1 U15915 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12829) );
  NAND2_X1 U15916 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12828) );
  NAND4_X1 U15917 ( .A1(n12831), .A2(n12830), .A3(n12829), .A4(n12828), .ZN(
        n12837) );
  AOI22_X1 U15918 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U15919 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U15920 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U15921 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12832) );
  NAND4_X1 U15922 ( .A1(n12835), .A2(n12834), .A3(n12833), .A4(n12832), .ZN(
        n12836) );
  OR2_X1 U15923 ( .A1(n12837), .A2(n12836), .ZN(n12866) );
  INV_X1 U15924 ( .A(n12866), .ZN(n12838) );
  XNOR2_X1 U15925 ( .A(n12867), .B(n12838), .ZN(n12841) );
  INV_X1 U15926 ( .A(n12979), .ZN(n13012) );
  INV_X1 U15927 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14930) );
  NAND2_X1 U15928 ( .A1(n20929), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12839) );
  OAI211_X1 U15929 ( .C1(n13010), .C2(n14930), .A(n12982), .B(n12839), .ZN(
        n12840) );
  AOI21_X1 U15930 ( .B1(n12841), .B2(n13012), .A(n12840), .ZN(n12842) );
  AOI21_X1 U15931 ( .B1(n15048), .B2(n13741), .A(n12842), .ZN(n14728) );
  INV_X1 U15932 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15044) );
  NAND2_X1 U15933 ( .A1(n12844), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12897) );
  INV_X1 U15934 ( .A(n12844), .ZN(n12845) );
  INV_X1 U15935 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14714) );
  NAND2_X1 U15936 ( .A1(n12845), .A2(n14714), .ZN(n12846) );
  NAND2_X1 U15937 ( .A1(n12897), .A2(n12846), .ZN(n15035) );
  INV_X1 U15938 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12858) );
  INV_X1 U15939 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12849) );
  INV_X1 U15940 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12847) );
  OAI22_X1 U15941 ( .A1(n12850), .A2(n12849), .B1(n12848), .B2(n12847), .ZN(
        n12854) );
  INV_X1 U15942 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12852) );
  INV_X1 U15943 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12851) );
  OAI22_X1 U15944 ( .A1(n12959), .A2(n12852), .B1(n12907), .B2(n12851), .ZN(
        n12853) );
  AOI211_X1 U15945 ( .C1(n9945), .C2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n12854), .B(n12853), .ZN(n12857) );
  AOI22_X1 U15946 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12855), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12856) );
  OAI211_X1 U15947 ( .C1(n13879), .C2(n12858), .A(n12857), .B(n12856), .ZN(
        n12865) );
  AOI22_X1 U15948 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9961), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12863) );
  AOI22_X1 U15949 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U15950 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12861) );
  AOI22_X1 U15951 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12860) );
  NAND4_X1 U15952 ( .A1(n12863), .A2(n12862), .A3(n12861), .A4(n12860), .ZN(
        n12864) );
  NOR2_X1 U15953 ( .A1(n12865), .A2(n12864), .ZN(n12875) );
  NAND2_X1 U15954 ( .A1(n12867), .A2(n12866), .ZN(n12874) );
  XNOR2_X1 U15955 ( .A(n12875), .B(n12874), .ZN(n12871) );
  NAND2_X1 U15956 ( .A1(n20929), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12868) );
  NAND2_X1 U15957 ( .A1(n12982), .A2(n12868), .ZN(n12869) );
  AOI21_X1 U15958 ( .B1(n14429), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12869), .ZN(
        n12870) );
  OAI21_X1 U15959 ( .B1(n12871), .B2(n12979), .A(n12870), .ZN(n12872) );
  XNOR2_X1 U15960 ( .A(n12897), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15024) );
  NAND2_X1 U15961 ( .A1(n15024), .A2(n13741), .ZN(n12896) );
  NOR2_X1 U15962 ( .A1(n12875), .A2(n12874), .ZN(n12903) );
  INV_X1 U15963 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12878) );
  NAND2_X1 U15964 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12877) );
  NAND2_X1 U15965 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12876) );
  OAI211_X1 U15966 ( .C1(n13879), .C2(n12878), .A(n12877), .B(n12876), .ZN(
        n12879) );
  INV_X1 U15967 ( .A(n12879), .ZN(n12884) );
  AOI22_X1 U15968 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12883) );
  AOI22_X1 U15969 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12882) );
  NAND2_X1 U15970 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12881) );
  NAND4_X1 U15971 ( .A1(n12884), .A2(n12883), .A3(n12882), .A4(n12881), .ZN(
        n12890) );
  AOI22_X1 U15972 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U15973 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U15974 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12886) );
  AOI22_X1 U15975 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12885) );
  NAND4_X1 U15976 ( .A1(n12888), .A2(n12887), .A3(n12886), .A4(n12885), .ZN(
        n12889) );
  OR2_X1 U15977 ( .A1(n12890), .A2(n12889), .ZN(n12902) );
  XNOR2_X1 U15978 ( .A(n12903), .B(n12902), .ZN(n12894) );
  NAND2_X1 U15979 ( .A1(n20929), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12891) );
  NAND2_X1 U15980 ( .A1(n12982), .A2(n12891), .ZN(n12892) );
  AOI21_X1 U15981 ( .B1(n14429), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12892), .ZN(
        n12893) );
  OAI21_X1 U15982 ( .B1(n12894), .B2(n12979), .A(n12893), .ZN(n12895) );
  NAND2_X1 U15983 ( .A1(n12896), .A2(n12895), .ZN(n14703) );
  INV_X1 U15984 ( .A(n12897), .ZN(n12898) );
  INV_X1 U15985 ( .A(n12899), .ZN(n12900) );
  INV_X1 U15986 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12922) );
  NAND2_X1 U15987 ( .A1(n12900), .A2(n12922), .ZN(n12901) );
  NAND2_X1 U15988 ( .A1(n12949), .A2(n12901), .ZN(n15017) );
  NAND2_X1 U15989 ( .A1(n12903), .A2(n12902), .ZN(n12928) );
  INV_X1 U15990 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12914) );
  INV_X1 U15991 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12905) );
  OAI22_X1 U15992 ( .A1(n12956), .A2(n12905), .B1(n12102), .B2(n12904), .ZN(
        n12911) );
  INV_X1 U15993 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12908) );
  INV_X1 U15994 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12906) );
  OAI22_X1 U15995 ( .A1(n9820), .A2(n12908), .B1(n12907), .B2(n12906), .ZN(
        n12910) );
  AOI211_X1 U15996 ( .C1(n9945), .C2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n12911), .B(n12910), .ZN(n12913) );
  AOI22_X1 U15997 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12993), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12912) );
  OAI211_X1 U15998 ( .C1(n12914), .C2(n13879), .A(n12913), .B(n12912), .ZN(
        n12921) );
  AOI22_X1 U15999 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12915), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12919) );
  AOI22_X1 U16000 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n9815), .B1(
        n9952), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U16001 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U16002 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12916) );
  NAND4_X1 U16003 ( .A1(n12919), .A2(n12918), .A3(n12917), .A4(n12916), .ZN(
        n12920) );
  NOR2_X1 U16004 ( .A1(n12921), .A2(n12920), .ZN(n12929) );
  XNOR2_X1 U16005 ( .A(n12928), .B(n12929), .ZN(n12925) );
  AOI21_X1 U16006 ( .B1(n12922), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12923) );
  AOI21_X1 U16007 ( .B1(n14429), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12923), .ZN(
        n12924) );
  OAI21_X1 U16008 ( .B1(n12925), .B2(n12979), .A(n12924), .ZN(n12926) );
  NAND2_X1 U16009 ( .A1(n12927), .A2(n12926), .ZN(n14686) );
  XNOR2_X1 U16010 ( .A(n12949), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14999) );
  INV_X1 U16011 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14997) );
  OAI21_X1 U16012 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14997), .A(n12982), 
        .ZN(n12947) );
  NOR2_X1 U16013 ( .A1(n12929), .A2(n12928), .ZN(n12976) );
  INV_X1 U16014 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12932) );
  NAND2_X1 U16015 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12931) );
  NAND2_X1 U16016 ( .A1(n12859), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12930) );
  OAI211_X1 U16017 ( .C1(n13879), .C2(n12932), .A(n12931), .B(n12930), .ZN(
        n12933) );
  INV_X1 U16018 ( .A(n12933), .ZN(n12937) );
  AOI22_X1 U16019 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U16020 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12935) );
  NAND2_X1 U16021 ( .A1(n9945), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12934) );
  NAND4_X1 U16022 ( .A1(n12937), .A2(n12936), .A3(n12935), .A4(n12934), .ZN(
        n12944) );
  AOI22_X1 U16023 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U16024 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12941) );
  AOI22_X1 U16025 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U16026 ( .A1(n12753), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12939) );
  NAND4_X1 U16027 ( .A1(n12942), .A2(n12941), .A3(n12940), .A4(n12939), .ZN(
        n12943) );
  OR2_X1 U16028 ( .A1(n12944), .A2(n12943), .ZN(n12975) );
  XNOR2_X1 U16029 ( .A(n12976), .B(n12975), .ZN(n12945) );
  NOR2_X1 U16030 ( .A1(n12945), .A2(n12979), .ZN(n12946) );
  AOI211_X1 U16031 ( .C1(n14429), .C2(P1_EAX_REG_28__SCAN_IN), .A(n12947), .B(
        n12946), .ZN(n12948) );
  AOI21_X1 U16032 ( .B1(n14999), .B2(n13741), .A(n12948), .ZN(n14672) );
  INV_X1 U16033 ( .A(n12949), .ZN(n12950) );
  NAND2_X1 U16034 ( .A1(n12951), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13744) );
  INV_X1 U16035 ( .A(n12951), .ZN(n12953) );
  INV_X1 U16036 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12952) );
  NAND2_X1 U16037 ( .A1(n12953), .A2(n12952), .ZN(n12954) );
  NAND2_X1 U16038 ( .A1(n13744), .A2(n12954), .ZN(n14992) );
  INV_X1 U16039 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12966) );
  INV_X1 U16040 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12957) );
  INV_X1 U16041 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12955) );
  OAI22_X1 U16042 ( .A1(n12988), .A2(n12957), .B1(n12956), .B2(n12955), .ZN(
        n12963) );
  INV_X1 U16043 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12958) );
  OAI22_X1 U16044 ( .A1(n12961), .A2(n12960), .B1(n12959), .B2(n12958), .ZN(
        n12962) );
  AOI211_X1 U16045 ( .C1(n9945), .C2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12963), .B(n12962), .ZN(n12965) );
  AOI22_X1 U16046 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12964) );
  OAI211_X1 U16047 ( .C1(n13879), .C2(n12966), .A(n12965), .B(n12964), .ZN(
        n12974) );
  AOI22_X1 U16048 ( .A1(n9961), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9957), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16049 ( .A1(n12751), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12752), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U16050 ( .A1(n9922), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12967), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U16051 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12969) );
  NAND4_X1 U16052 ( .A1(n12972), .A2(n12971), .A3(n12970), .A4(n12969), .ZN(
        n12973) );
  NOR2_X1 U16053 ( .A1(n12974), .A2(n12973), .ZN(n12984) );
  NAND2_X1 U16054 ( .A1(n12976), .A2(n12975), .ZN(n12983) );
  XNOR2_X1 U16055 ( .A(n12984), .B(n12983), .ZN(n12980) );
  AOI21_X1 U16056 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20929), .A(
        n13741), .ZN(n12978) );
  NAND2_X1 U16057 ( .A1(n14429), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12977) );
  OAI211_X1 U16058 ( .C1(n12980), .C2(n12979), .A(n12978), .B(n12977), .ZN(
        n12981) );
  OAI21_X1 U16059 ( .B1(n14992), .B2(n12982), .A(n12981), .ZN(n14660) );
  XNOR2_X1 U16060 ( .A(n13744), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14650) );
  NOR2_X1 U16061 ( .A1(n12984), .A2(n12983), .ZN(n13008) );
  INV_X1 U16062 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12996) );
  INV_X1 U16063 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12987) );
  OAI22_X1 U16064 ( .A1(n12988), .A2(n12987), .B1(n12986), .B2(n12985), .ZN(
        n12992) );
  OAI22_X1 U16065 ( .A1(n12294), .A2(n12990), .B1(n12102), .B2(n12989), .ZN(
        n12991) );
  AOI211_X1 U16066 ( .C1(n9945), .C2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n12992), .B(n12991), .ZN(n12995) );
  AOI22_X1 U16067 ( .A1(n12993), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12859), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12994) );
  OAI211_X1 U16068 ( .C1(n13879), .C2(n12996), .A(n12995), .B(n12994), .ZN(
        n13006) );
  AOI22_X1 U16069 ( .A1(n12915), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9957), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U16070 ( .A1(n9962), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12997), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U16071 ( .A1(n12752), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12999), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U16072 ( .A1(n13000), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9922), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13001) );
  NAND4_X1 U16073 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        n13005) );
  NOR2_X1 U16074 ( .A1(n13006), .A2(n13005), .ZN(n13007) );
  XNOR2_X1 U16075 ( .A(n13008), .B(n13007), .ZN(n13013) );
  INV_X1 U16076 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13098) );
  OAI21_X1 U16077 ( .B1(n21085), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n20929), .ZN(n13009) );
  OAI21_X1 U16078 ( .B1(n13010), .B2(n13098), .A(n13009), .ZN(n13011) );
  AOI21_X1 U16079 ( .B1(n13013), .B2(n13012), .A(n13011), .ZN(n13014) );
  AOI21_X1 U16080 ( .B1(n14650), .B2(n13741), .A(n13014), .ZN(n14427) );
  AOI21_X1 U16081 ( .B1(n12253), .B2(n13587), .A(n12187), .ZN(n13447) );
  NAND2_X1 U16082 ( .A1(n12254), .A2(n13751), .ZN(n13017) );
  NAND3_X1 U16083 ( .A1(n13447), .A2(n13016), .A3(n13017), .ZN(n13590) );
  NOR2_X1 U16084 ( .A1(n13590), .A2(n14631), .ZN(n13541) );
  XNOR2_X1 U16085 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13032) );
  NAND2_X1 U16086 ( .A1(n20690), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13036) );
  INV_X1 U16087 ( .A(n13036), .ZN(n13031) );
  NAND2_X1 U16088 ( .A1(n13032), .A2(n13031), .ZN(n13019) );
  NAND2_X1 U16089 ( .A1(n20585), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13018) );
  NAND2_X1 U16090 ( .A1(n13019), .A2(n13018), .ZN(n13028) );
  MUX2_X1 U16091 ( .A(n13020), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13027) );
  NAND2_X1 U16092 ( .A1(n13028), .A2(n13027), .ZN(n13022) );
  NAND2_X1 U16093 ( .A1(n13020), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13021) );
  NAND2_X1 U16094 ( .A1(n13022), .A2(n13021), .ZN(n13026) );
  XNOR2_X1 U16095 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13025) );
  NOR2_X1 U16096 ( .A1(n12088), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13023) );
  AOI21_X1 U16097 ( .B1(n13026), .B2(n13025), .A(n13023), .ZN(n13057) );
  INV_X1 U16098 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16140) );
  NAND2_X1 U16099 ( .A1(n16140), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13024) );
  NOR2_X1 U16100 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16140), .ZN(
        n13056) );
  AOI21_X1 U16101 ( .B1(n13057), .B2(n13024), .A(n13056), .ZN(n13075) );
  NAND2_X1 U16102 ( .A1(n13055), .A2(n13075), .ZN(n13066) );
  NAND2_X1 U16103 ( .A1(n13075), .A2(n13034), .ZN(n13065) );
  XNOR2_X1 U16104 ( .A(n13026), .B(n13025), .ZN(n13072) );
  XNOR2_X1 U16105 ( .A(n13028), .B(n13027), .ZN(n13071) );
  INV_X1 U16106 ( .A(n13048), .ZN(n13051) );
  OR2_X1 U16107 ( .A1(n13029), .A2(n12268), .ZN(n13050) );
  INV_X1 U16108 ( .A(n13071), .ZN(n13030) );
  OAI21_X1 U16109 ( .B1(n13030), .B2(n13052), .A(n13050), .ZN(n13047) );
  XNOR2_X1 U16110 ( .A(n13032), .B(n13031), .ZN(n13070) );
  NOR2_X1 U16111 ( .A1(n12241), .A2(n20932), .ZN(n13033) );
  INV_X1 U16112 ( .A(n13044), .ZN(n13035) );
  NOR2_X1 U16113 ( .A1(n13070), .A2(n13035), .ZN(n13042) );
  OAI21_X1 U16114 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20690), .A(
        n13036), .ZN(n13038) );
  NOR2_X1 U16115 ( .A1(n13037), .A2(n13038), .ZN(n13041) );
  INV_X1 U16116 ( .A(n12221), .ZN(n13564) );
  INV_X1 U16117 ( .A(n13038), .ZN(n13039) );
  OAI211_X1 U16118 ( .C1(n13751), .C2(n13564), .A(n13050), .B(n13039), .ZN(
        n13040) );
  OAI21_X1 U16119 ( .B1(n13055), .B2(n13041), .A(n13040), .ZN(n13043) );
  NAND2_X1 U16120 ( .A1(n13042), .A2(n13043), .ZN(n13046) );
  NAND2_X1 U16121 ( .A1(n13044), .A2(n12268), .ZN(n13061) );
  OAI211_X1 U16122 ( .C1(n13044), .C2(n13043), .A(n13070), .B(n13061), .ZN(
        n13045) );
  OAI211_X1 U16123 ( .C1(n13048), .C2(n13047), .A(n13046), .B(n13045), .ZN(
        n13049) );
  OAI21_X1 U16124 ( .B1(n13051), .B2(n13050), .A(n13049), .ZN(n13054) );
  NAND2_X1 U16125 ( .A1(n13052), .A2(n13072), .ZN(n13053) );
  AOI22_X1 U16126 ( .A1(n13055), .A2(n13072), .B1(n13054), .B2(n13053), .ZN(
        n13063) );
  AND2_X1 U16127 ( .A1(n13057), .A2(n13056), .ZN(n13073) );
  INV_X1 U16128 ( .A(n13073), .ZN(n13058) );
  NOR2_X1 U16129 ( .A1(n13059), .A2(n13058), .ZN(n13062) );
  NAND2_X1 U16130 ( .A1(n13059), .A2(n13073), .ZN(n13060) );
  OAI22_X1 U16131 ( .A1(n13063), .A2(n13062), .B1(n13061), .B2(n13060), .ZN(
        n13064) );
  INV_X1 U16132 ( .A(n13067), .ZN(n13068) );
  NAND2_X1 U16133 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20936) );
  AOI22_X1 U16134 ( .A1(n13541), .A2(n16153), .B1(n13068), .B2(n16142), .ZN(
        n13077) );
  INV_X1 U16135 ( .A(n13069), .ZN(n13494) );
  NOR4_X1 U16136 ( .A1(n13073), .A2(n13072), .A3(n13071), .A4(n13070), .ZN(
        n13074) );
  OR2_X1 U16137 ( .A1(n13075), .A2(n13074), .ZN(n14624) );
  INV_X1 U16138 ( .A(n14624), .ZN(n13573) );
  NAND3_X1 U16139 ( .A1(n13494), .A2(n13573), .A3(n20936), .ZN(n13076) );
  NAND2_X1 U16140 ( .A1(n13077), .A2(n13076), .ZN(n13439) );
  OR2_X1 U16141 ( .A1(n16150), .A2(n20932), .ZN(n14634) );
  INV_X1 U16142 ( .A(n14634), .ZN(n13585) );
  INV_X1 U16143 ( .A(n13078), .ZN(n13081) );
  OR2_X1 U16144 ( .A1(n12301), .A2(n14634), .ZN(n13079) );
  NOR2_X1 U16145 ( .A1(n13079), .A2(n13015), .ZN(n13080) );
  AND3_X1 U16146 ( .A1(n13081), .A2(n13881), .A3(n13080), .ZN(n13990) );
  NAND2_X1 U16147 ( .A1(n13990), .A2(n9938), .ZN(n13082) );
  NAND2_X1 U16148 ( .A1(n13084), .A2(n13015), .ZN(n13769) );
  INV_X1 U16149 ( .A(n14987), .ZN(n13085) );
  INV_X1 U16150 ( .A(n13086), .ZN(n13575) );
  NOR4_X1 U16151 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13090) );
  NOR4_X1 U16152 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13089) );
  NOR4_X1 U16153 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13088) );
  NOR4_X1 U16154 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13087) );
  AND4_X1 U16155 ( .A1(n13090), .A2(n13089), .A3(n13088), .A4(n13087), .ZN(
        n13095) );
  NOR4_X1 U16156 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13093) );
  NOR4_X1 U16157 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13092) );
  NOR4_X1 U16158 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13091) );
  INV_X1 U16159 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20871) );
  AND4_X1 U16160 ( .A1(n13093), .A2(n13092), .A3(n13091), .A4(n20871), .ZN(
        n13094) );
  NAND2_X1 U16161 ( .A1(n13095), .A2(n13094), .ZN(n13096) );
  INV_X1 U16162 ( .A(n20236), .ZN(n20235) );
  NOR2_X1 U16163 ( .A1(n13575), .A2(n20235), .ZN(n13097) );
  NAND2_X1 U16164 ( .A1(n14983), .A2(n13097), .ZN(n14957) );
  NOR2_X1 U16165 ( .A1(n14983), .A2(n13098), .ZN(n13102) );
  NOR3_X2 U16166 ( .A1(n14965), .A2(n20236), .A3(n13575), .ZN(n14968) );
  INV_X1 U16167 ( .A(n14968), .ZN(n14951) );
  INV_X1 U16168 ( .A(DATAI_30_), .ZN(n13100) );
  INV_X1 U16169 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16640) );
  NOR2_X1 U16170 ( .A1(n20235), .A2(n16640), .ZN(n13099) );
  AOI21_X1 U16171 ( .B1(DATAI_14_), .B2(n20235), .A(n13099), .ZN(n14975) );
  NAND3_X1 U16172 ( .A1(n14983), .A2(n10059), .A3(n13015), .ZN(n14948) );
  OAI22_X1 U16173 ( .A1(n14951), .A2(n13100), .B1(n14975), .B2(n14948), .ZN(
        n13101) );
  AOI211_X1 U16174 ( .C1(n14966), .C2(BUF1_REG_30__SCAN_IN), .A(n13102), .B(
        n13101), .ZN(n13103) );
  AOI211_X1 U16175 ( .C1(n13108), .C2(n13107), .A(n13106), .B(n13105), .ZN(
        n14419) );
  NAND2_X1 U16176 ( .A1(n18886), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19023) );
  INV_X2 U16177 ( .A(n19023), .ZN(n18955) );
  NAND2_X1 U16178 ( .A1(n18955), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18951) );
  OAI211_X1 U16179 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18886), .B(n18944), .ZN(n19012) );
  OAI21_X1 U16180 ( .B1(n13109), .B2(n18375), .A(n19012), .ZN(n13110) );
  NAND2_X1 U16181 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19015) );
  OAI21_X1 U16182 ( .B1(n13111), .B2(n13110), .A(n19015), .ZN(n16716) );
  OAI22_X1 U16183 ( .A1(n13113), .A2(n13112), .B1(n13115), .B2(n16716), .ZN(
        n13114) );
  AOI22_X1 U16184 ( .A1(n18797), .A2(n13115), .B1(n16172), .B2(n13114), .ZN(
        n13116) );
  NAND2_X1 U16185 ( .A1(n18791), .A2(n18326), .ZN(n18350) );
  NOR2_X2 U16186 ( .A1(n17524), .A2(n18350), .ZN(n18250) );
  NAND2_X1 U16187 ( .A1(n13117), .A2(n18250), .ZN(n13138) );
  NAND2_X1 U16188 ( .A1(n17524), .A2(n18791), .ZN(n18226) );
  INV_X1 U16189 ( .A(n18226), .ZN(n18044) );
  NAND2_X1 U16190 ( .A1(n18326), .A2(n18044), .ZN(n18199) );
  INV_X1 U16191 ( .A(n18199), .ZN(n18266) );
  OAI21_X1 U16192 ( .B1(n18973), .B2(n18991), .A(n18329), .ZN(n18321) );
  INV_X1 U16193 ( .A(n18321), .ZN(n18255) );
  INV_X1 U16194 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18280) );
  NAND3_X1 U16195 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18283) );
  OR2_X1 U16196 ( .A1(n18284), .A2(n18283), .ZN(n18254) );
  OR3_X1 U16197 ( .A1(n18263), .A2(n18280), .A3(n18254), .ZN(n13118) );
  NOR2_X1 U16198 ( .A1(n18255), .A2(n13118), .ZN(n18181) );
  NAND2_X1 U16199 ( .A1(n13119), .A2(n18181), .ZN(n18101) );
  NOR2_X1 U16200 ( .A1(n18804), .A2(n18101), .ZN(n16608) );
  NOR3_X1 U16201 ( .A1(n18329), .A2(n18973), .A3(n13118), .ZN(n18182) );
  NAND2_X1 U16202 ( .A1(n13119), .A2(n18182), .ZN(n18100) );
  INV_X1 U16203 ( .A(n18100), .ZN(n18159) );
  OAI221_X1 U16204 ( .B1(n16608), .B2(n18159), .C1(n16608), .C2(n18812), .A(
        n17683), .ZN(n13122) );
  INV_X1 U16205 ( .A(n13120), .ZN(n16609) );
  NAND3_X1 U16206 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17770), .A3(
        n18159), .ZN(n18118) );
  NOR2_X1 U16207 ( .A1(n16609), .A2(n18118), .ZN(n18039) );
  INV_X1 U16208 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18049) );
  NAND3_X1 U16209 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18057) );
  NOR2_X1 U16210 ( .A1(n18049), .A2(n18057), .ZN(n13123) );
  NAND3_X1 U16211 ( .A1(n18039), .A2(n13123), .A3(n18817), .ZN(n13121) );
  AOI211_X1 U16212 ( .C1(n13122), .C2(n13121), .A(n18344), .B(n16094), .ZN(
        n16096) );
  INV_X1 U16213 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17686) );
  INV_X1 U16214 ( .A(n13123), .ZN(n18038) );
  NOR2_X1 U16215 ( .A1(n17686), .A2(n18038), .ZN(n17662) );
  NAND2_X1 U16216 ( .A1(n17683), .A2(n18159), .ZN(n13126) );
  INV_X1 U16217 ( .A(n17683), .ZN(n13124) );
  INV_X1 U16218 ( .A(n18804), .ZN(n18822) );
  OAI21_X1 U16219 ( .B1(n13124), .B2(n18101), .A(n18822), .ZN(n18046) );
  INV_X1 U16220 ( .A(n18046), .ZN(n13125) );
  AOI211_X1 U16221 ( .C1(n18812), .C2(n13126), .A(n13125), .B(n18344), .ZN(
        n13127) );
  OAI221_X1 U16222 ( .B1(n18809), .B2(n18039), .C1(n18809), .C2(n17662), .A(
        n13127), .ZN(n16097) );
  INV_X1 U16223 ( .A(n18297), .ZN(n13129) );
  OAI221_X1 U16224 ( .B1(n16097), .B2(n13129), .C1(n16097), .C2(n13128), .A(
        n18345), .ZN(n16162) );
  NOR2_X1 U16225 ( .A1(n18344), .A2(n18297), .ZN(n18260) );
  INV_X1 U16226 ( .A(n18260), .ZN(n18331) );
  AOI221_X1 U16227 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16162), 
        .C1(n18331), .C2(n16162), .A(n18974), .ZN(n13131) );
  AOI211_X1 U16228 ( .C1(n13132), .C2(n16096), .A(n13131), .B(n13130), .ZN(
        n13133) );
  OAI21_X1 U16229 ( .B1(n13134), .B2(n18352), .A(n13133), .ZN(n13135) );
  AOI21_X1 U16230 ( .B1(n13136), .B2(n18266), .A(n13135), .ZN(n13137) );
  NAND2_X1 U16231 ( .A1(n13138), .A2(n13137), .ZN(P3_U2831) );
  INV_X1 U16232 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21261) );
  NOR3_X1 U16233 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n21261), .ZN(n13140) );
  NOR4_X1 U16234 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13139)
         );
  NAND4_X1 U16235 ( .A1(n20236), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13140), .A4(
        n13139), .ZN(U214) );
  NOR2_X1 U16236 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13142) );
  NOR4_X1 U16237 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13141) );
  NAND4_X1 U16238 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13142), .A4(n13141), .ZN(n13162) );
  NOR2_X1 U16239 ( .A1(n14137), .A2(n13162), .ZN(n16615) );
  NAND2_X1 U16240 ( .A1(n16615), .A2(U214), .ZN(U212) );
  NAND2_X1 U16241 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17718), .ZN(
        n13145) );
  INV_X1 U16242 ( .A(n13145), .ZN(n13146) );
  NAND3_X1 U16243 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(n13146), .ZN(n17669) );
  NAND2_X1 U16244 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17667), .ZN(
        n16742) );
  INV_X1 U16245 ( .A(n16742), .ZN(n13143) );
  AOI21_X1 U16246 ( .B1(n17695), .B2(n17669), .A(n13143), .ZN(n17697) );
  INV_X1 U16247 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17721) );
  NOR2_X1 U16248 ( .A1(n17721), .A2(n13145), .ZN(n13144) );
  OAI21_X1 U16249 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n13144), .A(
        n17669), .ZN(n17708) );
  INV_X1 U16250 ( .A(n17708), .ZN(n16797) );
  AOI21_X1 U16251 ( .B1(n17721), .B2(n13145), .A(n13144), .ZN(n17728) );
  INV_X1 U16252 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18027) );
  NOR2_X1 U16253 ( .A1(n18027), .A2(n17730), .ZN(n13148) );
  INV_X1 U16254 ( .A(n13148), .ZN(n17707) );
  AOI21_X1 U16255 ( .B1(n17745), .B2(n17707), .A(n13146), .ZN(n17737) );
  INV_X1 U16256 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17764) );
  NAND2_X1 U16257 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9967), .ZN(
        n13147) );
  XOR2_X1 U16258 ( .A(n17764), .B(n13147), .Z(n17773) );
  INV_X1 U16259 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17817) );
  NOR3_X1 U16260 ( .A1(n18027), .A2(n10603), .A3(n17817), .ZN(n17793) );
  NAND3_X1 U16261 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n17793), .ZN(n17747) );
  AOI22_X1 U16262 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9967), .B1(
        n17777), .B2(n17747), .ZN(n17781) );
  INV_X1 U16263 ( .A(n17747), .ZN(n16855) );
  NOR2_X1 U16264 ( .A1(n18027), .A2(n10021), .ZN(n17828) );
  NAND2_X1 U16265 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17828), .ZN(
        n16900) );
  OAI21_X1 U16266 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16900), .A(
        n16960), .ZN(n16891) );
  INV_X1 U16267 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17762) );
  NAND3_X1 U16268 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9967), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n13149) );
  AOI21_X1 U16269 ( .B1(n17762), .B2(n13149), .A(n13148), .ZN(n17752) );
  NOR2_X1 U16270 ( .A1(n17737), .A2(n16816), .ZN(n16815) );
  NOR2_X1 U16271 ( .A1(n16815), .A2(n17047), .ZN(n16809) );
  NOR2_X1 U16272 ( .A1(n17728), .A2(n16809), .ZN(n16808) );
  NOR2_X1 U16273 ( .A1(n16808), .A2(n17047), .ZN(n16796) );
  NOR2_X1 U16274 ( .A1(n16797), .A2(n16796), .ZN(n16795) );
  NOR2_X1 U16275 ( .A1(n16795), .A2(n17047), .ZN(n13150) );
  NOR2_X1 U16276 ( .A1(n17697), .A2(n13150), .ZN(n16743) );
  NOR4_X4 U16277 ( .A1(n18972), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(
        P3_STATE2_REG_0__SCAN_IN), .A4(P3_STATEBS16_REG_SCAN_IN), .ZN(n17069)
         );
  INV_X1 U16278 ( .A(n17069), .ZN(n18866) );
  AOI211_X1 U16279 ( .C1(n17697), .C2(n13150), .A(n16743), .B(n18866), .ZN(
        n13161) );
  NOR3_X1 U16280 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17062) );
  NAND2_X1 U16281 ( .A1(n17062), .A2(n17374), .ZN(n17055) );
  NOR2_X1 U16282 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17055), .ZN(n17034) );
  INV_X1 U16283 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17026) );
  NAND2_X1 U16284 ( .A1(n17034), .A2(n17026), .ZN(n17025) );
  NOR2_X1 U16285 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17025), .ZN(n17014) );
  INV_X1 U16286 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17362) );
  NAND2_X1 U16287 ( .A1(n17014), .A2(n17362), .ZN(n17003) );
  NOR2_X1 U16288 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17003), .ZN(n16978) );
  INV_X1 U16289 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16980) );
  NAND2_X1 U16290 ( .A1(n16978), .A2(n16980), .ZN(n16963) );
  NOR2_X1 U16291 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16963), .ZN(n16962) );
  INV_X1 U16292 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17297) );
  NAND2_X1 U16293 ( .A1(n16962), .A2(n17297), .ZN(n16955) );
  NOR2_X1 U16294 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16955), .ZN(n16936) );
  INV_X1 U16295 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16935) );
  NAND2_X1 U16296 ( .A1(n16936), .A2(n16935), .ZN(n16932) );
  NOR2_X1 U16297 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16932), .ZN(n16913) );
  INV_X1 U16298 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16906) );
  NAND2_X1 U16299 ( .A1(n16913), .A2(n16906), .ZN(n16902) );
  NOR2_X1 U16300 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16902), .ZN(n16888) );
  INV_X1 U16301 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16884) );
  NAND2_X1 U16302 ( .A1(n16888), .A2(n16884), .ZN(n16883) );
  NOR2_X1 U16303 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16883), .ZN(n16866) );
  INV_X1 U16304 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16857) );
  NAND2_X1 U16305 ( .A1(n16866), .A2(n16857), .ZN(n16856) );
  NOR2_X1 U16306 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16856), .ZN(n16845) );
  INV_X1 U16307 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17192) );
  NAND2_X1 U16308 ( .A1(n16845), .A2(n17192), .ZN(n16839) );
  NOR2_X1 U16309 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16839), .ZN(n16831) );
  INV_X1 U16310 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16821) );
  NAND2_X1 U16311 ( .A1(n16831), .A2(n16821), .ZN(n16820) );
  NOR2_X1 U16312 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16820), .ZN(n16805) );
  INV_X1 U16313 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17099) );
  NAND2_X1 U16314 ( .A1(n16805), .A2(n17099), .ZN(n16801) );
  NOR2_X1 U16315 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16801), .ZN(n16787) );
  NAND2_X1 U16316 ( .A1(n19009), .A2(n16172), .ZN(n16712) );
  NAND2_X1 U16317 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18375), .ZN(n13152) );
  AOI211_X4 U16318 ( .C1(n19013), .C2(n19015), .A(n19028), .B(n13152), .ZN(
        n17056) );
  AOI211_X1 U16319 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16801), .A(n16787), .B(
        n17091), .ZN(n13160) );
  NAND2_X1 U16320 ( .A1(n18354), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18732) );
  OR2_X1 U16321 ( .A1(n18862), .A2(n18732), .ZN(n18854) );
  INV_X1 U16322 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17100) );
  INV_X1 U16323 ( .A(n19015), .ZN(n18858) );
  AOI211_X1 U16324 ( .C1(n19014), .C2(n19012), .A(n18858), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n13153) );
  AOI211_X4 U16325 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18375), .A(n13153), .B(
        n19028), .ZN(n17078) );
  OAI22_X1 U16326 ( .A1(n17695), .A2(n17080), .B1(n17100), .B2(n17090), .ZN(
        n13159) );
  INV_X1 U16327 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18936) );
  INV_X1 U16328 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18933) );
  INV_X1 U16329 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18915) );
  INV_X1 U16330 ( .A(n13153), .ZN(n18850) );
  INV_X1 U16331 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18908) );
  INV_X1 U16332 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18900) );
  INV_X1 U16333 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18896) );
  INV_X1 U16334 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18894) );
  NAND3_X1 U16335 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17033) );
  NOR3_X1 U16336 ( .A1(n18896), .A2(n18894), .A3(n17033), .ZN(n17002) );
  NAND2_X1 U16337 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17002), .ZN(n16997) );
  NOR2_X1 U16338 ( .A1(n18900), .A2(n16997), .ZN(n16987) );
  NAND2_X1 U16339 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16987), .ZN(n16967) );
  NAND2_X1 U16340 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16952) );
  NOR3_X1 U16341 ( .A1(n18908), .A2(n16967), .A3(n16952), .ZN(n16943) );
  NAND2_X1 U16342 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16943), .ZN(n13154) );
  NAND2_X1 U16343 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16931), .ZN(n16916) );
  INV_X1 U16344 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18930) );
  INV_X1 U16345 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18926) );
  INV_X1 U16346 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18921) );
  INV_X1 U16347 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18918) );
  INV_X1 U16348 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18916) );
  NOR3_X1 U16349 ( .A1(n18921), .A2(n18918), .A3(n18916), .ZN(n16854) );
  INV_X1 U16350 ( .A(n16854), .ZN(n16861) );
  NAND2_X1 U16351 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16862) );
  NOR3_X1 U16352 ( .A1(n18926), .A2(n16861), .A3(n16862), .ZN(n16826) );
  NAND2_X1 U16353 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16826), .ZN(n16830) );
  NOR2_X1 U16354 ( .A1(n18930), .A2(n16830), .ZN(n13155) );
  NAND2_X1 U16355 ( .A1(n16897), .A2(n13155), .ZN(n16814) );
  NOR2_X1 U16356 ( .A1(n18933), .A2(n16814), .ZN(n16811) );
  NAND2_X1 U16357 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16811), .ZN(n16735) );
  NOR2_X1 U16358 ( .A1(n18936), .A2(n16735), .ZN(n13157) );
  INV_X1 U16359 ( .A(n16923), .ZN(n17092) );
  INV_X1 U16360 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18934) );
  INV_X1 U16361 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18912) );
  NAND2_X1 U16362 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17094), .ZN(n16914) );
  NOR3_X1 U16363 ( .A1(n18912), .A2(n13154), .A3(n16914), .ZN(n16887) );
  NAND3_X1 U16364 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n13155), .A3(n16887), 
        .ZN(n16807) );
  NOR2_X1 U16365 ( .A1(n18934), .A2(n16807), .ZN(n16794) );
  NAND3_X1 U16366 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n16794), .ZN(n16736) );
  NAND2_X1 U16367 ( .A1(n17092), .A2(n16736), .ZN(n16792) );
  INV_X1 U16368 ( .A(n16792), .ZN(n13156) );
  MUX2_X1 U16369 ( .A(n13157), .B(n13156), .S(P3_REIP_REG_26__SCAN_IN), .Z(
        n13158) );
  OR4_X1 U16370 ( .A1(n13161), .A2(n13160), .A3(n13159), .A4(n13158), .ZN(
        P3_U2645) );
  NOR2_X1 U16371 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13162), .ZN(n16699)
         );
  AOI21_X1 U16372 ( .B1(n13174), .B2(n16459), .A(n13163), .ZN(n16451) );
  AOI21_X1 U16373 ( .B1(n16472), .B2(n13172), .A(n13164), .ZN(n16460) );
  AOI21_X1 U16374 ( .B1(n16485), .B2(n13171), .A(n13165), .ZN(n16478) );
  AOI21_X1 U16375 ( .B1(n16494), .B2(n13166), .A(n13167), .ZN(n16486) );
  AOI21_X1 U16376 ( .B1(n16507), .B2(n13169), .A(n10007), .ZN(n16495) );
  AOI21_X1 U16377 ( .B1(n14015), .B2(n13168), .A(n13170), .ZN(n14147) );
  OAI22_X1 U16378 ( .A1(n19032), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n14267) );
  INV_X1 U16379 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14269) );
  OAI22_X1 U16380 ( .A1(n19032), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14269), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14266) );
  AND2_X1 U16381 ( .A1(n14267), .A2(n14266), .ZN(n14252) );
  OAI21_X1 U16382 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13168), .ZN(n14254) );
  NAND2_X1 U16383 ( .A1(n14252), .A2(n14254), .ZN(n14145) );
  NOR2_X1 U16384 ( .A1(n14147), .A2(n14145), .ZN(n19205) );
  OAI21_X1 U16385 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13170), .A(
        n13169), .ZN(n19340) );
  NAND2_X1 U16386 ( .A1(n19205), .A2(n19340), .ZN(n14097) );
  NOR2_X1 U16387 ( .A1(n16495), .A2(n14097), .ZN(n19186) );
  OAI21_X1 U16388 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10007), .A(
        n13166), .ZN(n19187) );
  NAND2_X1 U16389 ( .A1(n19186), .A2(n19187), .ZN(n14066) );
  NOR2_X1 U16390 ( .A1(n16486), .A2(n14066), .ZN(n19173) );
  OAI21_X1 U16391 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13167), .A(
        n13171), .ZN(n19174) );
  NAND2_X1 U16392 ( .A1(n19173), .A2(n19174), .ZN(n14110) );
  NOR2_X1 U16393 ( .A1(n16478), .A2(n14110), .ZN(n19160) );
  OAI21_X1 U16394 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13165), .A(
        n13172), .ZN(n19161) );
  NAND2_X1 U16395 ( .A1(n19160), .A2(n19161), .ZN(n14078) );
  NOR2_X1 U16396 ( .A1(n16460), .A2(n14078), .ZN(n19146) );
  OR2_X1 U16397 ( .A1(n13164), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13173) );
  NAND2_X1 U16398 ( .A1(n13174), .A2(n13173), .ZN(n19147) );
  NAND2_X1 U16399 ( .A1(n19146), .A2(n19147), .ZN(n13177) );
  NOR2_X1 U16400 ( .A1(n16451), .A2(n13177), .ZN(n19132) );
  INV_X1 U16401 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13175) );
  INV_X1 U16402 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14588) );
  INV_X1 U16403 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20039) );
  NAND4_X1 U16404 ( .A1(n20039), .A2(n19032), .A3(n19629), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19895) );
  INV_X1 U16405 ( .A(n19895), .ZN(n19191) );
  NAND2_X1 U16406 ( .A1(n10206), .A2(n19191), .ZN(n19093) );
  AOI211_X1 U16407 ( .C1(n16451), .C2(n13177), .A(n19132), .B(n19093), .ZN(
        n13204) );
  NAND3_X1 U16408 ( .A1(n11491), .A2(n13828), .A3(n13178), .ZN(n13255) );
  OR2_X1 U16409 ( .A1(n13255), .A2(n13179), .ZN(n13329) );
  INV_X1 U16410 ( .A(n13250), .ZN(n13795) );
  NOR2_X1 U16411 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13795), .ZN(n13196) );
  NOR2_X1 U16412 ( .A1(n13329), .A2(n13196), .ZN(n15358) );
  INV_X1 U16413 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13180) );
  NAND2_X1 U16414 ( .A1(n20046), .A2(n19629), .ZN(n13193) );
  NAND2_X1 U16415 ( .A1(n13180), .A2(n13193), .ZN(n13181) );
  NOR2_X1 U16416 ( .A1(n13255), .A2(n13181), .ZN(n13182) );
  INV_X1 U16417 ( .A(n19168), .ZN(n19215) );
  INV_X1 U16418 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n14022) );
  NOR2_X1 U16419 ( .A1(n20012), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19398) );
  INV_X1 U16420 ( .A(n19398), .ZN(n19891) );
  NOR2_X1 U16421 ( .A1(n19898), .A2(n19891), .ZN(n16574) );
  INV_X1 U16422 ( .A(n16574), .ZN(n13183) );
  NAND2_X1 U16423 ( .A1(n19895), .A2(n13183), .ZN(n13184) );
  NOR2_X1 U16424 ( .A1(n19328), .A2(n13184), .ZN(n13185) );
  NAND2_X1 U16425 ( .A1(n19220), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19155) );
  OAI22_X1 U16426 ( .A1(n19215), .A2(n14022), .B1(n16459), .B2(n19155), .ZN(
        n13203) );
  INV_X1 U16427 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19938) );
  NAND3_X1 U16428 ( .A1(n20026), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n13193), 
        .ZN(n13186) );
  INV_X1 U16429 ( .A(n19217), .ZN(n19110) );
  AOI22_X1 U16430 ( .A1(n13187), .A2(n19110), .B1(n16451), .B2(n19228), .ZN(
        n13188) );
  OAI211_X1 U16431 ( .C1(n19938), .C2(n19220), .A(n13188), .B(n19181), .ZN(
        n13202) );
  INV_X1 U16432 ( .A(n13189), .ZN(n13192) );
  INV_X1 U16433 ( .A(n13190), .ZN(n13940) );
  AOI21_X1 U16434 ( .B1(n13192), .B2(n13940), .A(n13191), .ZN(n16523) );
  INV_X1 U16435 ( .A(n16523), .ZN(n13200) );
  INV_X1 U16436 ( .A(n13193), .ZN(n13194) );
  NAND2_X1 U16437 ( .A1(n20026), .A2(n13194), .ZN(n13195) );
  OR2_X1 U16438 ( .A1(n20043), .A2(n13195), .ZN(n19202) );
  NAND2_X1 U16439 ( .A1(n13197), .A2(n13196), .ZN(n13847) );
  NAND2_X1 U16440 ( .A1(n13632), .A2(n13198), .ZN(n13199) );
  NAND2_X1 U16441 ( .A1(n13199), .A2(n10006), .ZN(n19244) );
  OAI22_X1 U16442 ( .A1(n13200), .A2(n19202), .B1(n19214), .B2(n19244), .ZN(
        n13201) );
  OR4_X1 U16443 ( .A1(n13204), .A2(n13203), .A3(n13202), .A4(n13201), .ZN(
        P2_U2842) );
  AOI21_X1 U16444 ( .B1(n15608), .B2(n13207), .A(n13206), .ZN(n16424) );
  OAI21_X1 U16445 ( .B1(n10022), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n13207), .ZN(n15619) );
  INV_X1 U16446 ( .A(n15619), .ZN(n15382) );
  AOI21_X1 U16447 ( .B1(n13209), .B2(n10204), .A(n10022), .ZN(n15628) );
  OAI21_X1 U16448 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n13208), .A(
        n13209), .ZN(n16103) );
  AOI21_X1 U16449 ( .B1(n13216), .B2(n13211), .A(n13210), .ZN(n19071) );
  AOI21_X1 U16450 ( .B1(n15705), .B2(n13215), .A(n13212), .ZN(n19096) );
  AOI21_X1 U16451 ( .B1(n16445), .B2(n13214), .A(n13213), .ZN(n19124) );
  OAI21_X1 U16452 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13163), .A(
        n13214), .ZN(n19133) );
  NAND2_X1 U16453 ( .A1(n19132), .A2(n19133), .ZN(n19122) );
  NOR2_X1 U16454 ( .A1(n19124), .A2(n19122), .ZN(n19114) );
  OAI21_X1 U16455 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13213), .A(
        n13215), .ZN(n19115) );
  NAND2_X1 U16456 ( .A1(n19114), .A2(n19115), .ZN(n19095) );
  NOR2_X1 U16457 ( .A1(n19096), .A2(n19095), .ZN(n19094) );
  OAI21_X1 U16458 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13212), .A(
        n13216), .ZN(n19085) );
  NAND2_X1 U16459 ( .A1(n19094), .A2(n19085), .ZN(n19069) );
  NOR2_X1 U16460 ( .A1(n19071), .A2(n19069), .ZN(n19065) );
  OAI21_X1 U16461 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n13210), .A(
        n13217), .ZN(n19068) );
  NAND2_X1 U16462 ( .A1(n19065), .A2(n19068), .ZN(n15410) );
  NAND2_X1 U16463 ( .A1(n15663), .A2(n13217), .ZN(n13219) );
  INV_X1 U16464 ( .A(n13208), .ZN(n13218) );
  AND2_X1 U16465 ( .A1(n13219), .A2(n13218), .ZN(n15665) );
  NOR2_X1 U16466 ( .A1(n15628), .A2(n15398), .ZN(n15397) );
  NOR2_X1 U16467 ( .A1(n19206), .A2(n16422), .ZN(n13221) );
  OAI21_X1 U16468 ( .B1(n13206), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15354), .ZN(n15596) );
  INV_X1 U16469 ( .A(n15596), .ZN(n13220) );
  NOR2_X1 U16470 ( .A1(n13220), .A2(n13221), .ZN(n15357) );
  AOI211_X1 U16471 ( .C1(n13221), .C2(n13220), .A(n19895), .B(n15357), .ZN(
        n13236) );
  OR2_X1 U16472 ( .A1(n13223), .A2(n13224), .ZN(n13225) );
  NAND2_X1 U16473 ( .A1(n13222), .A2(n13225), .ZN(n15779) );
  NOR2_X1 U16474 ( .A1(n15779), .A2(n19202), .ZN(n13235) );
  AOI211_X1 U16475 ( .C1(P2_EBX_REG_26__SCAN_IN), .C2(n13226), .A(n19217), .B(
        n14573), .ZN(n13234) );
  INV_X1 U16476 ( .A(n13227), .ZN(n13230) );
  INV_X1 U16477 ( .A(n13228), .ZN(n13229) );
  OAI21_X1 U16478 ( .B1(n13230), .B2(n13229), .A(n15511), .ZN(n15784) );
  AOI22_X1 U16479 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19199), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19168), .ZN(n13232) );
  NAND2_X1 U16480 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19229), .ZN(
        n13231) );
  OAI211_X1 U16481 ( .C1(n15784), .C2(n19214), .A(n13232), .B(n13231), .ZN(
        n13233) );
  OR4_X1 U16482 ( .A1(n13236), .A2(n13235), .A3(n13234), .A4(n13233), .ZN(
        P2_U2829) );
  MUX2_X1 U16483 ( .A(n15889), .B(n13370), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13244) );
  OAI21_X1 U16484 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19216), .A(
        n13368), .ZN(n13409) );
  NOR2_X1 U16485 ( .A1(n16552), .A2(n13409), .ZN(n13243) );
  OAI21_X1 U16486 ( .B1(n13238), .B2(n13237), .A(n11526), .ZN(n19254) );
  OAI22_X1 U16487 ( .A1(n16544), .A2(n19254), .B1(n13414), .B2(n15976), .ZN(
        n13242) );
  AOI22_X1 U16488 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13240), .B1(
        n13239), .B2(n13367), .ZN(n13405) );
  NAND2_X1 U16489 ( .A1(n19172), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13407) );
  OAI21_X1 U16490 ( .B1(n15966), .B2(n13405), .A(n13407), .ZN(n13241) );
  OR4_X1 U16491 ( .A1(n13244), .A2(n13243), .A3(n13242), .A4(n13241), .ZN(
        P2_U3046) );
  NOR2_X1 U16492 ( .A1(n11484), .A2(n16580), .ZN(n13328) );
  NAND2_X1 U16493 ( .A1(n13328), .A2(n13828), .ZN(n19203) );
  INV_X1 U16494 ( .A(n19203), .ZN(n19227) );
  INV_X1 U16495 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13246) );
  AND2_X1 U16496 ( .A1(n19990), .A2(n14396), .ZN(n13247) );
  INV_X1 U16497 ( .A(n13247), .ZN(n13245) );
  OAI211_X1 U16498 ( .C1(n19227), .C2(n13246), .A(n13255), .B(n13245), .ZN(
        P2_U2814) );
  INV_X1 U16499 ( .A(n11703), .ZN(n20037) );
  OAI21_X1 U16500 ( .B1(n13247), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n20043), 
        .ZN(n13248) );
  OAI21_X1 U16501 ( .B1(n20037), .B2(n20043), .A(n13248), .ZN(P2_U3612) );
  INV_X1 U16502 ( .A(n13249), .ZN(n13251) );
  NOR3_X1 U16503 ( .A1(n13252), .A2(n13251), .A3(n13250), .ZN(n13834) );
  NOR2_X1 U16504 ( .A1(n13834), .A2(n16580), .ZN(n20032) );
  OAI21_X1 U16505 ( .B1(n20032), .B2(n11121), .A(n13253), .ZN(P2_U2819) );
  NAND2_X1 U16506 ( .A1(n11507), .A2(n20046), .ZN(n13254) );
  OR2_X1 U16507 ( .A1(n13255), .A2(n13254), .ZN(n13308) );
  NAND2_X1 U16508 ( .A1(n13297), .A2(n13929), .ZN(n13302) );
  INV_X1 U16509 ( .A(n13255), .ZN(n13256) );
  OAI21_X1 U16510 ( .B1(n19356), .B2(n20046), .A(n13256), .ZN(n13264) );
  NAND2_X1 U16511 ( .A1(n13264), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13257) );
  OAI211_X1 U16512 ( .C1(n12077), .C2(n13329), .A(n13302), .B(n13257), .ZN(
        P2_U2966) );
  AOI22_X1 U16513 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n13264), .B1(n13305), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13258) );
  AOI22_X1 U16514 ( .A1(n14135), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14137), .ZN(n19362) );
  INV_X1 U16515 ( .A(n19362), .ZN(n14202) );
  NAND2_X1 U16516 ( .A1(n13297), .A2(n14202), .ZN(n13283) );
  NAND2_X1 U16517 ( .A1(n13258), .A2(n13283), .ZN(P2_U2954) );
  AOI22_X1 U16518 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n13264), .B1(n13305), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13259) );
  INV_X1 U16519 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16654) );
  INV_X1 U16520 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18404) );
  AOI22_X1 U16521 ( .A1(n14135), .A2(n16654), .B1(n18404), .B2(n14137), .ZN(
        n19245) );
  NAND2_X1 U16522 ( .A1(n13297), .A2(n19245), .ZN(n13267) );
  NAND2_X1 U16523 ( .A1(n13259), .A2(n13267), .ZN(P2_U2959) );
  AOI22_X1 U16524 ( .A1(P2_UWORD_REG_8__SCAN_IN), .A2(n13264), .B1(n13305), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n13261) );
  AOI22_X1 U16525 ( .A1(n14135), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n14137), .ZN(n15533) );
  INV_X1 U16526 ( .A(n15533), .ZN(n13260) );
  NAND2_X1 U16527 ( .A1(n13297), .A2(n13260), .ZN(n13281) );
  NAND2_X1 U16528 ( .A1(n13261), .A2(n13281), .ZN(P2_U2960) );
  AOI22_X1 U16529 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n13264), .B1(n13305), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13262) );
  AOI22_X1 U16530 ( .A1(n14135), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14137), .ZN(n19374) );
  INV_X1 U16531 ( .A(n19374), .ZN(n14285) );
  NAND2_X1 U16532 ( .A1(n13297), .A2(n14285), .ZN(n13270) );
  NAND2_X1 U16533 ( .A1(n13262), .A2(n13270), .ZN(P2_U2956) );
  AOI22_X1 U16534 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n13264), .B1(n13305), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13263) );
  AOI22_X1 U16535 ( .A1(n14135), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14137), .ZN(n19357) );
  INV_X1 U16536 ( .A(n19357), .ZN(n15565) );
  NAND2_X1 U16537 ( .A1(n13297), .A2(n15565), .ZN(n13291) );
  NAND2_X1 U16538 ( .A1(n13263), .A2(n13291), .ZN(P2_U2953) );
  CLKBUF_X2 U16539 ( .A(n13264), .Z(n13306) );
  AOI22_X1 U16540 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13265) );
  AOI22_X1 U16541 ( .A1(n14135), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14137), .ZN(n19385) );
  INV_X1 U16542 ( .A(n19385), .ZN(n15543) );
  NAND2_X1 U16543 ( .A1(n13297), .A2(n15543), .ZN(n13274) );
  NAND2_X1 U16544 ( .A1(n13265), .A2(n13274), .ZN(P2_U2958) );
  AOI22_X1 U16545 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13266) );
  AOI22_X1 U16546 ( .A1(n14135), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14137), .ZN(n19381) );
  INV_X1 U16547 ( .A(n19381), .ZN(n15549) );
  NAND2_X1 U16548 ( .A1(n13297), .A2(n15549), .ZN(n13279) );
  NAND2_X1 U16549 ( .A1(n13266), .A2(n13279), .ZN(P2_U2957) );
  AOI22_X1 U16550 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13268) );
  NAND2_X1 U16551 ( .A1(n13268), .A2(n13267), .ZN(P2_U2974) );
  AOI22_X1 U16552 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n13269) );
  AOI22_X1 U16553 ( .A1(n14135), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14137), .ZN(n19292) );
  INV_X1 U16554 ( .A(n19292), .ZN(n14049) );
  NAND2_X1 U16555 ( .A1(n13297), .A2(n14049), .ZN(n13287) );
  NAND2_X1 U16556 ( .A1(n13269), .A2(n13287), .ZN(P2_U2952) );
  AOI22_X1 U16557 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13271) );
  NAND2_X1 U16558 ( .A1(n13271), .A2(n13270), .ZN(P2_U2971) );
  AOI22_X1 U16559 ( .A1(P2_LWORD_REG_10__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n13272) );
  MUX2_X1 U16560 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n14137), .Z(n15521) );
  NAND2_X1 U16561 ( .A1(n13297), .A2(n15521), .ZN(n13285) );
  NAND2_X1 U16562 ( .A1(n13272), .A2(n13285), .ZN(P2_U2977) );
  AOI22_X1 U16563 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13273) );
  AOI22_X1 U16564 ( .A1(n14135), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14137), .ZN(n19368) );
  INV_X1 U16565 ( .A(n19368), .ZN(n15557) );
  NAND2_X1 U16566 ( .A1(n13297), .A2(n15557), .ZN(n13277) );
  NAND2_X1 U16567 ( .A1(n13273), .A2(n13277), .ZN(P2_U2955) );
  AOI22_X1 U16568 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13275) );
  NAND2_X1 U16569 ( .A1(n13275), .A2(n13274), .ZN(P2_U2973) );
  AOI22_X1 U16570 ( .A1(P2_LWORD_REG_12__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n13276) );
  MUX2_X1 U16571 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n14137), .Z(n15506) );
  NAND2_X1 U16572 ( .A1(n13297), .A2(n15506), .ZN(n13289) );
  NAND2_X1 U16573 ( .A1(n13276), .A2(n13289), .ZN(P2_U2979) );
  AOI22_X1 U16574 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13278) );
  NAND2_X1 U16575 ( .A1(n13278), .A2(n13277), .ZN(P2_U2970) );
  AOI22_X1 U16576 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13280) );
  NAND2_X1 U16577 ( .A1(n13280), .A2(n13279), .ZN(P2_U2972) );
  AOI22_X1 U16578 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13282) );
  NAND2_X1 U16579 ( .A1(n13282), .A2(n13281), .ZN(P2_U2975) );
  AOI22_X1 U16580 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13284) );
  NAND2_X1 U16581 ( .A1(n13284), .A2(n13283), .ZN(P2_U2969) );
  AOI22_X1 U16582 ( .A1(P2_UWORD_REG_10__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n13286) );
  NAND2_X1 U16583 ( .A1(n13286), .A2(n13285), .ZN(P2_U2962) );
  AOI22_X1 U16584 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13288) );
  NAND2_X1 U16585 ( .A1(n13288), .A2(n13287), .ZN(P2_U2967) );
  AOI22_X1 U16586 ( .A1(P2_UWORD_REG_12__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n13290) );
  NAND2_X1 U16587 ( .A1(n13290), .A2(n13289), .ZN(P2_U2964) );
  AOI22_X1 U16588 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13292) );
  NAND2_X1 U16589 ( .A1(n13292), .A2(n13291), .ZN(P2_U2968) );
  INV_X1 U16590 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19299) );
  MUX2_X1 U16591 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n14137), .Z(n19241) );
  NAND2_X1 U16592 ( .A1(n13297), .A2(n19241), .ZN(n13300) );
  NAND2_X1 U16593 ( .A1(n13306), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13293) );
  OAI211_X1 U16594 ( .C1(n19299), .C2(n13329), .A(n13300), .B(n13293), .ZN(
        P2_U2980) );
  INV_X1 U16595 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n13517) );
  MUX2_X1 U16596 ( .A(BUF1_REG_9__SCAN_IN), .B(BUF2_REG_9__SCAN_IN), .S(n14137), .Z(n15528) );
  NAND2_X1 U16597 ( .A1(n13297), .A2(n15528), .ZN(n13296) );
  NAND2_X1 U16598 ( .A1(n13306), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13294) );
  OAI211_X1 U16599 ( .C1(n13517), .C2(n13329), .A(n13296), .B(n13294), .ZN(
        P2_U2961) );
  INV_X1 U16600 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19307) );
  NAND2_X1 U16601 ( .A1(n13306), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13295) );
  OAI211_X1 U16602 ( .C1(n19307), .C2(n13329), .A(n13296), .B(n13295), .ZN(
        P2_U2976) );
  INV_X1 U16603 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19303) );
  MUX2_X1 U16604 ( .A(BUF1_REG_11__SCAN_IN), .B(BUF2_REG_11__SCAN_IN), .S(
        n14137), .Z(n15515) );
  NAND2_X1 U16605 ( .A1(n13297), .A2(n15515), .ZN(n13304) );
  NAND2_X1 U16606 ( .A1(n13306), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13298) );
  OAI211_X1 U16607 ( .C1(n19303), .C2(n13329), .A(n13304), .B(n13298), .ZN(
        P2_U2978) );
  INV_X1 U16608 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13510) );
  NAND2_X1 U16609 ( .A1(n13306), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13299) );
  OAI211_X1 U16610 ( .C1(n13510), .C2(n13329), .A(n13300), .B(n13299), .ZN(
        P2_U2965) );
  INV_X1 U16611 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19297) );
  NAND2_X1 U16612 ( .A1(n13306), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13301) );
  OAI211_X1 U16613 ( .C1(n19297), .C2(n13329), .A(n13302), .B(n13301), .ZN(
        P2_U2981) );
  INV_X1 U16614 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13514) );
  NAND2_X1 U16615 ( .A1(n13306), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13303) );
  OAI211_X1 U16616 ( .C1(n13514), .C2(n13329), .A(n13304), .B(n13303), .ZN(
        P2_U2963) );
  AOI22_X1 U16617 ( .A1(n14135), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14137), .ZN(n19240) );
  AOI22_X1 U16618 ( .A1(P2_LWORD_REG_15__SCAN_IN), .A2(n13306), .B1(n13305), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n13307) );
  OAI21_X1 U16619 ( .B1(n19240), .B2(n13308), .A(n13307), .ZN(P2_U2982) );
  NAND2_X1 U16620 ( .A1(n9934), .A2(n13573), .ZN(n13316) );
  INV_X1 U16621 ( .A(n13324), .ZN(n13314) );
  INV_X1 U16622 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n13313) );
  INV_X1 U16623 ( .A(n13310), .ZN(n13311) );
  NAND3_X1 U16624 ( .A1(n13311), .A2(n13585), .A3(n16153), .ZN(n13475) );
  NOR2_X2 U16625 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20790) );
  AND2_X1 U16626 ( .A1(n20790), .A2(n20849), .ZN(n14322) );
  INV_X1 U16627 ( .A(n14322), .ZN(n13312) );
  OAI211_X1 U16628 ( .C1(n13314), .C2(n13313), .A(n13475), .B(n13312), .ZN(
        P1_U2801) );
  NOR2_X1 U16629 ( .A1(n16153), .A2(n9938), .ZN(n13315) );
  AOI21_X1 U16630 ( .B1(n13316), .B2(n13310), .A(n13315), .ZN(n14633) );
  AND2_X1 U16631 ( .A1(n14633), .A2(n13585), .ZN(n13318) );
  INV_X1 U16632 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21076) );
  NAND2_X1 U16633 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14322), .ZN(n13317) );
  OAI21_X1 U16634 ( .B1(n13318), .B2(n21076), .A(n13317), .ZN(P1_U2803) );
  OR2_X1 U16635 ( .A1(n13320), .A2(n13319), .ZN(n13321) );
  NAND2_X1 U16636 ( .A1(n13322), .A2(n13321), .ZN(n19195) );
  INV_X1 U16637 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19314) );
  INV_X1 U16638 ( .A(n16430), .ZN(n15534) );
  OAI222_X1 U16639 ( .A1(n19195), .A2(n19252), .B1(n19250), .B2(n19314), .C1(
        n19291), .C2(n19385), .ZN(P2_U2913) );
  NOR2_X1 U16640 ( .A1(n14322), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13327)
         );
  NAND2_X1 U16641 ( .A1(n20934), .A2(n13325), .ZN(n13326) );
  OAI21_X1 U16642 ( .B1(n20934), .B2(n13327), .A(n13326), .ZN(P1_U3487) );
  INV_X1 U16643 ( .A(n13328), .ZN(n13330) );
  OAI21_X1 U16644 ( .B1(n13794), .B2(n13330), .A(n13329), .ZN(n13331) );
  INV_X1 U16645 ( .A(n19906), .ZN(n20034) );
  AND2_X1 U16646 ( .A1(n13331), .A2(n20034), .ZN(n19293) );
  NAND2_X1 U16647 ( .A1(n19293), .A2(n13332), .ZN(n13527) );
  NOR2_X1 U16648 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13851), .ZN(n13515) );
  AOI22_X1 U16649 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n19312), .B1(n13515), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13333) );
  OAI21_X1 U16650 ( .B1(n12077), .B2(n13527), .A(n13333), .ZN(P2_U2921) );
  INV_X1 U16651 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15504) );
  AOI22_X1 U16652 ( .A1(n13515), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19312), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13334) );
  OAI21_X1 U16653 ( .B1(n15504), .B2(n13527), .A(n13334), .ZN(P2_U2923) );
  INV_X1 U16654 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15532) );
  AOI22_X1 U16655 ( .A1(n13515), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19312), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13335) );
  OAI21_X1 U16656 ( .B1(n15532), .B2(n13527), .A(n13335), .ZN(P2_U2927) );
  INV_X1 U16657 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n15519) );
  AOI22_X1 U16658 ( .A1(n13515), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19312), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13336) );
  OAI21_X1 U16659 ( .B1(n15519), .B2(n13527), .A(n13336), .ZN(P2_U2925) );
  OAI21_X1 U16660 ( .B1(n13338), .B2(n13351), .A(n13337), .ZN(n13355) );
  INV_X1 U16661 ( .A(n13339), .ZN(n13340) );
  XNOR2_X1 U16662 ( .A(n13341), .B(n13340), .ZN(n13393) );
  NAND2_X1 U16663 ( .A1(n13393), .A2(n16566), .ZN(n13350) );
  OAI21_X1 U16664 ( .B1(n13344), .B2(n13343), .A(n13342), .ZN(n20000) );
  AOI22_X1 U16665 ( .A1(n20000), .A2(n16558), .B1(P2_REIP_REG_2__SCAN_IN), 
        .B2(n19328), .ZN(n13349) );
  OR2_X1 U16666 ( .A1(n13346), .A2(n13345), .ZN(n13389) );
  NAND3_X1 U16667 ( .A1(n16563), .A2(n13388), .A3(n13389), .ZN(n13348) );
  NAND4_X1 U16668 ( .A1(n13350), .A2(n13349), .A3(n13348), .A4(n13347), .ZN(
        n13354) );
  NOR2_X1 U16669 ( .A1(n13352), .A2(n13351), .ZN(n13353) );
  AOI211_X1 U16670 ( .C1(n13366), .C2(n13355), .A(n13354), .B(n13353), .ZN(
        n13356) );
  OAI21_X1 U16671 ( .B1(n13472), .B2(n15976), .A(n13356), .ZN(P2_U3044) );
  NAND2_X1 U16672 ( .A1(n13359), .A2(n13358), .ZN(n13360) );
  INV_X1 U16673 ( .A(n13833), .ZN(n13361) );
  INV_X1 U16674 ( .A(n13785), .ZN(n13830) );
  NAND2_X1 U16675 ( .A1(n13361), .A2(n13830), .ZN(n13798) );
  NAND2_X1 U16676 ( .A1(n13798), .A2(n11717), .ZN(n13363) );
  NAND2_X1 U16677 ( .A1(n13363), .A2(n13362), .ZN(n14224) );
  NAND2_X1 U16678 ( .A1(n14214), .A2(n13364), .ZN(n15493) );
  MUX2_X1 U16679 ( .A(n14273), .B(n13818), .S(n14214), .Z(n13365) );
  OAI21_X1 U16680 ( .B1(n20007), .B2(n15493), .A(n13365), .ZN(P2_U2886) );
  AOI211_X1 U16681 ( .C1(n14394), .C2(n13367), .A(n13366), .B(n15944), .ZN(
        n13381) );
  XNOR2_X1 U16682 ( .A(n13368), .B(n14394), .ZN(n13369) );
  XNOR2_X1 U16683 ( .A(n14271), .B(n13369), .ZN(n13395) );
  NAND2_X1 U16684 ( .A1(n13370), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13371) );
  NAND2_X1 U16685 ( .A1(n19172), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13396) );
  OAI211_X1 U16686 ( .C1(n13395), .C2(n16552), .A(n13371), .B(n13396), .ZN(
        n13380) );
  OAI21_X1 U16687 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13373), .A(
        n13372), .ZN(n13398) );
  NAND2_X1 U16688 ( .A1(n13375), .A2(n13374), .ZN(n13376) );
  NAND2_X1 U16689 ( .A1(n13377), .A2(n13376), .ZN(n20003) );
  INV_X1 U16690 ( .A(n20003), .ZN(n13378) );
  OAI22_X1 U16691 ( .A1(n13398), .A2(n15966), .B1(n16544), .B2(n13378), .ZN(
        n13379) );
  NOR3_X1 U16692 ( .A1(n13381), .A2(n13380), .A3(n13379), .ZN(n13382) );
  OAI21_X1 U16693 ( .B1(n13818), .B2(n15976), .A(n13382), .ZN(P2_U3045) );
  INV_X1 U16694 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13384) );
  AND2_X1 U16695 ( .A1(n20012), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13383) );
  OAI211_X1 U16696 ( .C1(n19356), .C2(n13384), .A(n19384), .B(n13383), .ZN(
        n13385) );
  INV_X1 U16697 ( .A(n13385), .ZN(n13386) );
  INV_X2 U16698 ( .A(n14214), .ZN(n15490) );
  MUX2_X1 U16699 ( .A(n13414), .B(n11136), .S(n15490), .Z(n13387) );
  OAI21_X1 U16700 ( .B1(n19342), .B2(n15493), .A(n13387), .ZN(P2_U2887) );
  NAND3_X1 U16701 ( .A1(n13389), .A2(n16502), .A3(n13388), .ZN(n13391) );
  AOI22_X1 U16702 ( .A1(n19329), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n19172), .B2(P2_REIP_REG_2__SCAN_IN), .ZN(n13390) );
  OAI211_X1 U16703 ( .C1(n14254), .C2(n19341), .A(n13391), .B(n13390), .ZN(
        n13392) );
  AOI21_X1 U16704 ( .B1(n13393), .B2(n16503), .A(n13392), .ZN(n13394) );
  OAI21_X1 U16705 ( .B1(n13472), .B2(n14136), .A(n13394), .ZN(P2_U3012) );
  INV_X1 U16706 ( .A(n13395), .ZN(n13400) );
  MUX2_X1 U16707 ( .A(n19341), .B(n16506), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13397) );
  OAI211_X1 U16708 ( .C1(n13398), .C2(n19332), .A(n13397), .B(n13396), .ZN(
        n13399) );
  AOI21_X1 U16709 ( .B1(n16502), .B2(n13400), .A(n13399), .ZN(n13401) );
  OAI21_X1 U16710 ( .B1(n13818), .B2(n14136), .A(n13401), .ZN(P2_U3013) );
  OAI21_X1 U16711 ( .B1(n13404), .B2(n13402), .A(n13403), .ZN(n19180) );
  INV_X1 U16712 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19309) );
  OAI222_X1 U16713 ( .A1(n19180), .A2(n19252), .B1(n15533), .B2(n19291), .C1(
        n19309), .C2(n19250), .ZN(P2_U2911) );
  INV_X1 U16714 ( .A(n13405), .ZN(n13406) );
  NAND2_X1 U16715 ( .A1(n16503), .A2(n13406), .ZN(n13408) );
  OAI211_X1 U16716 ( .C1(n13409), .C2(n19333), .A(n13408), .B(n13407), .ZN(
        n13410) );
  INV_X1 U16717 ( .A(n13410), .ZN(n13413) );
  OAI21_X1 U16718 ( .B1(n19329), .B2(n13411), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13412) );
  OAI211_X1 U16719 ( .C1(n13414), .C2(n14136), .A(n13413), .B(n13412), .ZN(
        P2_U3014) );
  AND2_X1 U16720 ( .A1(n9934), .A2(n12268), .ZN(n15345) );
  OR2_X1 U16721 ( .A1(n13415), .A2(n14378), .ZN(n13594) );
  INV_X1 U16722 ( .A(n13594), .ZN(n16143) );
  OR2_X1 U16723 ( .A1(n15345), .A2(n16143), .ZN(n13421) );
  INV_X1 U16724 ( .A(n13416), .ZN(n13418) );
  INV_X1 U16725 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n13417) );
  NAND2_X1 U16726 ( .A1(n13418), .A2(n13417), .ZN(n16165) );
  NOR2_X1 U16727 ( .A1(n16165), .A2(n14634), .ZN(n13419) );
  AND2_X1 U16728 ( .A1(n16153), .A2(n13419), .ZN(n13420) );
  NAND2_X1 U16729 ( .A1(n20144), .A2(n20243), .ZN(n13650) );
  NOR2_X1 U16730 ( .A1(n20929), .A2(n20849), .ZN(n16368) );
  NAND2_X1 U16731 ( .A1(n20932), .A2(n16368), .ZN(n20142) );
  AOI22_X1 U16732 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20164), .B1(n16167), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13422) );
  OAI21_X1 U16733 ( .B1(n14930), .B2(n13650), .A(n13422), .ZN(P1_U2912) );
  INV_X1 U16734 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n21032) );
  AOI22_X1 U16735 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20164), .B1(n16167), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13423) );
  OAI21_X1 U16736 ( .B1(n21032), .B2(n13650), .A(n13423), .ZN(P1_U2908) );
  INV_X1 U16737 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13425) );
  AOI22_X1 U16738 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20164), .B1(n16167), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13424) );
  OAI21_X1 U16739 ( .B1(n13425), .B2(n13650), .A(n13424), .ZN(P1_U2914) );
  INV_X1 U16740 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21044) );
  AOI22_X1 U16741 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20164), .B1(n16167), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13426) );
  OAI21_X1 U16742 ( .B1(n21044), .B2(n13650), .A(n13426), .ZN(P1_U2915) );
  INV_X1 U16743 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13428) );
  AOI22_X1 U16744 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20164), .B1(n16167), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13427) );
  OAI21_X1 U16745 ( .B1(n13428), .B2(n13650), .A(n13427), .ZN(P1_U2909) );
  INV_X1 U16746 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21264) );
  AOI22_X1 U16747 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20164), .B1(n16167), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13429) );
  OAI21_X1 U16748 ( .B1(n21264), .B2(n13650), .A(n13429), .ZN(P1_U2911) );
  AOI22_X1 U16749 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20164), .B1(n16167), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13430) );
  OAI21_X1 U16750 ( .B1(n14947), .B2(n13650), .A(n13430), .ZN(P1_U2916) );
  INV_X1 U16751 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14936) );
  AOI22_X1 U16752 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20164), .B1(n16167), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13431) );
  OAI21_X1 U16753 ( .B1(n14936), .B2(n13650), .A(n13431), .ZN(P1_U2913) );
  INV_X1 U16754 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13433) );
  AOI22_X1 U16755 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20164), .B1(n16167), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13432) );
  OAI21_X1 U16756 ( .B1(n13433), .B2(n13650), .A(n13432), .ZN(P1_U2917) );
  INV_X1 U16757 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n21046) );
  AOI22_X1 U16758 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20164), .B1(n16167), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13434) );
  OAI21_X1 U16759 ( .B1(n21046), .B2(n13650), .A(n13434), .ZN(P1_U2907) );
  AOI21_X1 U16760 ( .B1(n13436), .B2(n13403), .A(n13435), .ZN(n15960) );
  INV_X1 U16761 ( .A(n15960), .ZN(n13438) );
  INV_X1 U16762 ( .A(n15528), .ZN(n13437) );
  OAI222_X1 U16763 ( .A1(n13438), .A2(n19252), .B1(n19250), .B2(n19307), .C1(
        n19291), .C2(n13437), .ZN(P2_U2910) );
  INV_X1 U16764 ( .A(n13439), .ZN(n13453) );
  INV_X1 U16765 ( .A(n13590), .ZN(n13440) );
  OR2_X1 U16766 ( .A1(n9934), .A2(n13440), .ZN(n13443) );
  OAI21_X1 U16767 ( .B1(n12253), .B2(n13751), .A(n14378), .ZN(n13441) );
  NAND2_X1 U16768 ( .A1(n13442), .A2(n13441), .ZN(n13606) );
  AND2_X1 U16769 ( .A1(n13443), .A2(n13606), .ZN(n13583) );
  AND2_X1 U16770 ( .A1(n13751), .A2(n12268), .ZN(n13749) );
  NAND2_X1 U16771 ( .A1(n13749), .A2(n13578), .ZN(n13444) );
  AND2_X1 U16772 ( .A1(n13583), .A2(n13444), .ZN(n13452) );
  OR2_X1 U16773 ( .A1(n12221), .A2(n20243), .ZN(n13445) );
  NAND3_X1 U16774 ( .A1(n13447), .A2(n13446), .A3(n13445), .ZN(n13449) );
  AOI21_X1 U16775 ( .B1(n13449), .B2(n12268), .A(n13448), .ZN(n13609) );
  NAND2_X1 U16776 ( .A1(n13609), .A2(n12241), .ZN(n13458) );
  NAND2_X1 U16777 ( .A1(n12253), .A2(n12268), .ZN(n13581) );
  INV_X1 U16778 ( .A(n13415), .ZN(n13450) );
  INV_X1 U16779 ( .A(n16165), .ZN(n16141) );
  OAI211_X1 U16780 ( .C1(n15345), .C2(n13450), .A(n16141), .B(n16142), .ZN(
        n13451) );
  NAND4_X1 U16781 ( .A1(n13453), .A2(n13452), .A3(n13992), .A4(n13451), .ZN(
        n16115) );
  INV_X1 U16782 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20057) );
  NAND2_X1 U16783 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16368), .ZN(n16372) );
  NOR2_X1 U16784 ( .A1(n20057), .A2(n16372), .ZN(n13454) );
  AOI21_X1 U16785 ( .B1(n16115), .B2(n13585), .A(n13454), .ZN(n13463) );
  INV_X1 U16786 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20664) );
  NAND2_X1 U16787 ( .A1(n20932), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13455) );
  OAI22_X1 U16788 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20914), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20849), .ZN(n13456) );
  INV_X1 U16789 ( .A(n13456), .ZN(n13467) );
  INV_X1 U16790 ( .A(n13606), .ZN(n13457) );
  NOR2_X1 U16791 ( .A1(n13458), .A2(n13457), .ZN(n13460) );
  AND3_X1 U16792 ( .A1(n13460), .A2(n13459), .A3(n13069), .ZN(n15342) );
  INV_X1 U16793 ( .A(n15342), .ZN(n13892) );
  MUX2_X1 U16794 ( .A(n13461), .B(n15345), .S(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13462) );
  AOI21_X1 U16795 ( .B1(n12378), .B2(n13892), .A(n13462), .ZN(n16118) );
  INV_X1 U16796 ( .A(n16118), .ZN(n13464) );
  INV_X1 U16797 ( .A(n13553), .ZN(n20916) );
  NOR2_X1 U16798 ( .A1(n13463), .A2(n20916), .ZN(n13495) );
  NAND2_X1 U16799 ( .A1(n13464), .A2(n13495), .ZN(n13466) );
  NAND2_X1 U16800 ( .A1(n20918), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13465) );
  OAI211_X1 U16801 ( .C1(n20918), .C2(n13467), .A(n13466), .B(n13465), .ZN(
        P1_U3474) );
  MUX2_X1 U16802 ( .A(n10787), .B(n13472), .S(n14214), .Z(n13473) );
  OAI21_X1 U16803 ( .B1(n19998), .B2(n15493), .A(n13473), .ZN(P2_U2885) );
  INV_X1 U16804 ( .A(n20936), .ZN(n20859) );
  AND2_X1 U16805 ( .A1(n14378), .A2(n20859), .ZN(n13474) );
  OR2_X2 U16806 ( .A1(n13475), .A2(n13474), .ZN(n20178) );
  OR2_X1 U16807 ( .A1(n20178), .A2(n12268), .ZN(n13652) );
  NAND2_X1 U16808 ( .A1(n20178), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13478) );
  INV_X1 U16809 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16650) );
  NOR2_X1 U16810 ( .A1(n20235), .A2(n16650), .ZN(n13476) );
  AOI21_X1 U16811 ( .B1(DATAI_9_), .B2(n20235), .A(n13476), .ZN(n14925) );
  INV_X1 U16812 ( .A(n14925), .ZN(n13477) );
  NAND2_X1 U16813 ( .A1(n13682), .A2(n13477), .ZN(n20168) );
  OAI211_X1 U16814 ( .C1(n13652), .C2(n21264), .A(n13478), .B(n20168), .ZN(
        P1_U2946) );
  INV_X1 U16815 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21234) );
  NAND2_X1 U16816 ( .A1(n20178), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13479) );
  MUX2_X1 U16817 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20236), .Z(
        n14921) );
  NAND2_X1 U16818 ( .A1(n13682), .A2(n14921), .ZN(n20170) );
  OAI211_X1 U16819 ( .C1(n13652), .C2(n21234), .A(n13479), .B(n20170), .ZN(
        P1_U2947) );
  NAND2_X1 U16820 ( .A1(n20178), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13482) );
  INV_X1 U16821 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16642) );
  NOR2_X1 U16822 ( .A1(n20235), .A2(n16642), .ZN(n13480) );
  AOI21_X1 U16823 ( .B1(DATAI_13_), .B2(n20235), .A(n13480), .ZN(n14978) );
  INV_X1 U16824 ( .A(n14978), .ZN(n13481) );
  NAND2_X1 U16825 ( .A1(n13682), .A2(n13481), .ZN(n20176) );
  OAI211_X1 U16826 ( .C1(n13652), .C2(n21046), .A(n13482), .B(n20176), .ZN(
        P1_U2950) );
  NAND2_X1 U16827 ( .A1(n20178), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13484) );
  INV_X1 U16828 ( .A(n14975), .ZN(n13483) );
  NAND2_X1 U16829 ( .A1(n13682), .A2(n13483), .ZN(n20180) );
  OAI211_X1 U16830 ( .C1(n13652), .C2(n13098), .A(n13484), .B(n20180), .ZN(
        P1_U2951) );
  NAND2_X1 U16831 ( .A1(n20178), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13485) );
  MUX2_X1 U16832 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n20236), .Z(
        n14980) );
  NAND2_X1 U16833 ( .A1(n13682), .A2(n14980), .ZN(n20174) );
  OAI211_X1 U16834 ( .C1(n13652), .C2(n21032), .A(n13485), .B(n20174), .ZN(
        P1_U2949) );
  INV_X1 U16835 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14971) );
  INV_X1 U16836 ( .A(n13682), .ZN(n13488) );
  INV_X1 U16837 ( .A(DATAI_15_), .ZN(n13486) );
  NOR2_X1 U16838 ( .A1(n20236), .A2(n13486), .ZN(n13487) );
  AOI21_X1 U16839 ( .B1(n20236), .B2(BUF1_REG_15__SCAN_IN), .A(n13487), .ZN(
        n14972) );
  INV_X1 U16840 ( .A(n20178), .ZN(n13653) );
  INV_X1 U16841 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20143) );
  OAI222_X1 U16842 ( .A1(n13652), .A2(n14971), .B1(n13488), .B2(n14972), .C1(
        n13653), .C2(n20143), .ZN(P1_U2967) );
  NAND2_X1 U16843 ( .A1(n20178), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13490) );
  INV_X1 U16844 ( .A(DATAI_8_), .ZN(n21201) );
  INV_X1 U16845 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16652) );
  MUX2_X1 U16846 ( .A(n21201), .B(n16652), .S(n20236), .Z(n14931) );
  INV_X1 U16847 ( .A(n14931), .ZN(n13489) );
  NAND2_X1 U16848 ( .A1(n13682), .A2(n13489), .ZN(n13491) );
  OAI211_X1 U16849 ( .C1(n13652), .C2(n14930), .A(n13490), .B(n13491), .ZN(
        P1_U2945) );
  INV_X1 U16850 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20153) );
  NAND2_X1 U16851 ( .A1(n20178), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13492) );
  OAI211_X1 U16852 ( .C1(n13652), .C2(n20153), .A(n13492), .B(n13491), .ZN(
        P1_U2960) );
  INV_X1 U16853 ( .A(n20400), .ZN(n20654) );
  OR2_X1 U16854 ( .A1(n12391), .A2(n20654), .ZN(n13493) );
  XNOR2_X1 U16855 ( .A(n13493), .B(n13496), .ZN(n20130) );
  NAND2_X1 U16856 ( .A1(n13495), .A2(n13494), .ZN(n13497) );
  INV_X1 U16857 ( .A(n20918), .ZN(n15350) );
  OAI22_X1 U16858 ( .A1(n20130), .A2(n13497), .B1(n13496), .B2(n15350), .ZN(
        P1_U3468) );
  INV_X1 U16859 ( .A(n13498), .ZN(n13503) );
  INV_X1 U16860 ( .A(n13499), .ZN(n13501) );
  INV_X1 U16861 ( .A(n13435), .ZN(n13500) );
  NAND2_X1 U16862 ( .A1(n13501), .A2(n13500), .ZN(n13502) );
  NAND2_X1 U16863 ( .A1(n13503), .A2(n13502), .ZN(n19167) );
  INV_X1 U16864 ( .A(n15521), .ZN(n13504) );
  INV_X1 U16865 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19305) );
  OAI222_X1 U16866 ( .A1(n19167), .A2(n19252), .B1(n13504), .B2(n19291), .C1(
        n19305), .C2(n19250), .ZN(P2_U2909) );
  INV_X1 U16867 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13506) );
  AOI22_X1 U16868 ( .A1(n13515), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13505) );
  OAI21_X1 U16869 ( .B1(n13506), .B2(n13527), .A(n13505), .ZN(P2_U2929) );
  INV_X1 U16870 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n13508) );
  AOI22_X1 U16871 ( .A1(n13515), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13507) );
  OAI21_X1 U16872 ( .B1(n13508), .B2(n13527), .A(n13507), .ZN(P2_U2930) );
  AOI22_X1 U16873 ( .A1(n13515), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13509) );
  OAI21_X1 U16874 ( .B1(n13510), .B2(n13527), .A(n13509), .ZN(P2_U2922) );
  INV_X1 U16875 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13512) );
  AOI22_X1 U16876 ( .A1(n13515), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13511) );
  OAI21_X1 U16877 ( .B1(n13512), .B2(n13527), .A(n13511), .ZN(P2_U2928) );
  AOI22_X1 U16878 ( .A1(n13515), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13513) );
  OAI21_X1 U16879 ( .B1(n13514), .B2(n13527), .A(n13513), .ZN(P2_U2924) );
  AOI22_X1 U16880 ( .A1(n13515), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13516) );
  OAI21_X1 U16881 ( .B1(n13517), .B2(n13527), .A(n13516), .ZN(P2_U2926) );
  INV_X1 U16882 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13519) );
  AOI22_X1 U16883 ( .A1(n20047), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13518) );
  OAI21_X1 U16884 ( .B1(n13519), .B2(n13527), .A(n13518), .ZN(P2_U2933) );
  INV_X1 U16885 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13521) );
  AOI22_X1 U16886 ( .A1(n20047), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13520) );
  OAI21_X1 U16887 ( .B1(n13521), .B2(n13527), .A(n13520), .ZN(P2_U2935) );
  INV_X1 U16888 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13523) );
  AOI22_X1 U16889 ( .A1(n20047), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13522) );
  OAI21_X1 U16890 ( .B1(n13523), .B2(n13527), .A(n13522), .ZN(P2_U2934) );
  INV_X1 U16891 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13525) );
  AOI22_X1 U16892 ( .A1(n20047), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13524) );
  OAI21_X1 U16893 ( .B1(n13525), .B2(n13527), .A(n13524), .ZN(P2_U2931) );
  INV_X1 U16894 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13528) );
  AOI22_X1 U16895 ( .A1(n20047), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13526) );
  OAI21_X1 U16896 ( .B1(n13528), .B2(n13527), .A(n13526), .ZN(P2_U2932) );
  NOR2_X1 U16897 ( .A1(n13532), .A2(n15490), .ZN(n13533) );
  AOI21_X1 U16898 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n15490), .A(n13533), .ZN(
        n13534) );
  OAI21_X1 U16899 ( .B1(n19988), .B2(n15493), .A(n13534), .ZN(P2_U2884) );
  OR2_X1 U16900 ( .A1(n20655), .A2(n15342), .ZN(n13549) );
  INV_X1 U16901 ( .A(n13536), .ZN(n13539) );
  INV_X1 U16902 ( .A(n13537), .ZN(n13538) );
  NAND2_X1 U16903 ( .A1(n13538), .A2(n10052), .ZN(n13882) );
  NAND2_X1 U16904 ( .A1(n13539), .A2(n13882), .ZN(n13543) );
  INV_X1 U16905 ( .A(n13543), .ZN(n13551) );
  NAND2_X1 U16906 ( .A1(n13881), .A2(n13551), .ZN(n13546) );
  XNOR2_X1 U16907 ( .A(n10058), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13540) );
  NAND2_X1 U16908 ( .A1(n15345), .A2(n13540), .ZN(n13545) );
  INV_X1 U16909 ( .A(n13541), .ZN(n13542) );
  NAND2_X1 U16910 ( .A1(n14623), .A2(n13542), .ZN(n13884) );
  NAND2_X1 U16911 ( .A1(n13884), .A2(n13543), .ZN(n13544) );
  OAI211_X1 U16912 ( .C1(n13892), .C2(n13546), .A(n13545), .B(n13544), .ZN(
        n13547) );
  INV_X1 U16913 ( .A(n13547), .ZN(n13548) );
  NAND2_X1 U16914 ( .A1(n13549), .A2(n13548), .ZN(n13896) );
  INV_X1 U16915 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14525) );
  NOR2_X1 U16916 ( .A1(n20849), .A2(n14525), .ZN(n15347) );
  INV_X1 U16917 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14538) );
  INV_X1 U16918 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20214) );
  OAI22_X1 U16919 ( .A1(n14538), .A2(n20214), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15348) );
  INV_X1 U16920 ( .A(n15348), .ZN(n13552) );
  AOI222_X1 U16921 ( .A1(n13896), .A2(n13553), .B1(n15347), .B2(n13552), .C1(
        n13551), .C2(n13550), .ZN(n13554) );
  MUX2_X1 U16922 ( .A(n13554), .B(n10052), .S(n20918), .Z(n13555) );
  INV_X1 U16923 ( .A(n13555), .ZN(P1_U3472) );
  AND3_X1 U16924 ( .A1(n20932), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16364) );
  AND2_X2 U16925 ( .A1(n16364), .A2(n20790), .ZN(n20188) );
  INV_X1 U16926 ( .A(n20188), .ZN(n15135) );
  INV_X1 U16927 ( .A(n13556), .ZN(n13559) );
  OAI21_X1 U16928 ( .B1(n13559), .B2(n13558), .A(n13557), .ZN(n14020) );
  INV_X1 U16929 ( .A(n14375), .ZN(n13872) );
  NAND2_X1 U16930 ( .A1(n13751), .A2(n20268), .ZN(n13857) );
  OAI21_X1 U16931 ( .B1(n14378), .B2(n13693), .A(n13857), .ZN(n13560) );
  INV_X1 U16932 ( .A(n13560), .ZN(n13561) );
  OAI21_X1 U16933 ( .B1(n13563), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13864), .ZN(n13614) );
  NOR2_X1 U16934 ( .A1(n13590), .A2(n13564), .ZN(n13565) );
  AND2_X1 U16935 ( .A1(n13565), .A2(n16153), .ZN(n16131) );
  OR2_X1 U16936 ( .A1(n13566), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20222) );
  NAND2_X1 U16937 ( .A1(n10057), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13600) );
  INV_X1 U16938 ( .A(n20790), .ZN(n20779) );
  NAND2_X1 U16939 ( .A1(n20779), .A2(n13566), .ZN(n20935) );
  AND2_X1 U16940 ( .A1(n20935), .A2(n20932), .ZN(n13567) );
  NAND2_X1 U16941 ( .A1(n20932), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16144) );
  NAND2_X1 U16942 ( .A1(n21085), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13568) );
  NAND2_X1 U16943 ( .A1(n16144), .A2(n13568), .ZN(n13684) );
  OAI21_X1 U16944 ( .B1(n20182), .B2(n13684), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13569) );
  OAI211_X1 U16945 ( .C1(n13614), .C2(n20056), .A(n13600), .B(n13569), .ZN(
        n13570) );
  INV_X1 U16946 ( .A(n13570), .ZN(n13571) );
  OAI21_X1 U16947 ( .B1(n15135), .B2(n14020), .A(n13571), .ZN(P1_U2999) );
  AOI21_X1 U16948 ( .B1(n12268), .B2(n16165), .A(n20859), .ZN(n13572) );
  NAND2_X1 U16949 ( .A1(n13573), .A2(n13572), .ZN(n13580) );
  INV_X1 U16950 ( .A(n13753), .ZN(n13574) );
  NOR2_X1 U16951 ( .A1(n13415), .A2(n13574), .ZN(n13577) );
  NAND2_X1 U16952 ( .A1(n13575), .A2(n20243), .ZN(n13576) );
  AOI22_X1 U16953 ( .A1(n16142), .A2(n13577), .B1(n16153), .B2(n13576), .ZN(
        n13579) );
  MUX2_X1 U16954 ( .A(n13580), .B(n13579), .S(n13578), .Z(n13584) );
  OR2_X1 U16955 ( .A1(n16153), .A2(n13581), .ZN(n13582) );
  NAND3_X1 U16956 ( .A1(n13584), .A2(n13583), .A3(n13582), .ZN(n13586) );
  NOR2_X1 U16957 ( .A1(n13595), .A2(n13587), .ZN(n13591) );
  NOR2_X1 U16958 ( .A1(n12221), .A2(n9938), .ZN(n13589) );
  NOR2_X1 U16959 ( .A1(n13590), .A2(n13589), .ZN(n14626) );
  OR3_X1 U16960 ( .A1(n13592), .A2(n13591), .A3(n14626), .ZN(n13593) );
  NAND2_X1 U16961 ( .A1(n13612), .A2(n15345), .ZN(n15334) );
  NAND2_X1 U16962 ( .A1(n15330), .A2(n15334), .ZN(n13602) );
  OAI21_X1 U16963 ( .B1(n13595), .B2(n12301), .A(n13594), .ZN(n13596) );
  INV_X1 U16964 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13775) );
  NAND2_X1 U16965 ( .A1(n14517), .A2(n13775), .ZN(n13599) );
  NAND2_X1 U16966 ( .A1(n14236), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13598) );
  OAI21_X1 U16967 ( .B1(n13597), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13949), .ZN(n14021) );
  OAI21_X1 U16968 ( .B1(n20225), .B2(n14021), .A(n13600), .ZN(n13601) );
  AOI21_X1 U16969 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13602), .A(
        n13601), .ZN(n13613) );
  INV_X1 U16970 ( .A(n13603), .ZN(n13605) );
  AOI22_X1 U16971 ( .A1(n13605), .A2(n13751), .B1(n13604), .B2(n13881), .ZN(
        n13608) );
  NAND4_X1 U16972 ( .A1(n13609), .A2(n13608), .A3(n13607), .A4(n13606), .ZN(
        n13610) );
  NAND2_X1 U16973 ( .A1(n13612), .A2(n13610), .ZN(n14523) );
  INV_X1 U16974 ( .A(n14623), .ZN(n13611) );
  OAI21_X1 U16975 ( .B1(n14539), .B2(n20221), .A(n14525), .ZN(n15329) );
  OAI211_X1 U16976 ( .C1(n13614), .C2(n16326), .A(n13613), .B(n15329), .ZN(
        P1_U3031) );
  INV_X1 U16977 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13615) );
  NOR2_X1 U16978 ( .A1(n13616), .A2(n13615), .ZN(n13620) );
  NAND2_X1 U16979 ( .A1(n13617), .A2(n13620), .ZN(n13706) );
  INV_X1 U16980 ( .A(n13620), .ZN(n13621) );
  NAND3_X1 U16981 ( .A1(n13618), .A2(n13619), .A3(n13621), .ZN(n13622) );
  NAND2_X1 U16982 ( .A1(n13706), .A2(n13622), .ZN(n19262) );
  NAND2_X1 U16983 ( .A1(n13624), .A2(n13623), .ZN(n13626) );
  INV_X1 U16984 ( .A(n13625), .ZN(n13637) );
  AND2_X1 U16985 ( .A1(n13626), .A2(n13637), .ZN(n19336) );
  INV_X1 U16986 ( .A(n19336), .ZN(n19201) );
  MUX2_X1 U16987 ( .A(n19201), .B(n19196), .S(n15490), .Z(n13627) );
  OAI21_X1 U16988 ( .B1(n19262), .B2(n15493), .A(n13627), .ZN(P2_U2883) );
  NOR2_X1 U16989 ( .A1(n13498), .A2(n13628), .ZN(n13629) );
  NOR2_X1 U16990 ( .A1(n13634), .A2(n13629), .ZN(n16530) );
  INV_X1 U16991 ( .A(n16530), .ZN(n13631) );
  INV_X1 U16992 ( .A(n15515), .ZN(n13630) );
  OAI222_X1 U16993 ( .A1(n13631), .A2(n19252), .B1(n13630), .B2(n19291), .C1(
        n19303), .C2(n19250), .ZN(P2_U2908) );
  OAI21_X1 U16994 ( .B1(n13634), .B2(n13633), .A(n13632), .ZN(n19154) );
  INV_X1 U16995 ( .A(n15506), .ZN(n13635) );
  INV_X1 U16996 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19301) );
  OAI222_X1 U16997 ( .A1(n19154), .A2(n19252), .B1(n13635), .B2(n19291), .C1(
        n19301), .C2(n19250), .ZN(P2_U2907) );
  INV_X1 U16998 ( .A(n13706), .ZN(n13708) );
  XNOR2_X1 U16999 ( .A(n13708), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13642) );
  INV_X1 U17000 ( .A(n13636), .ZN(n13638) );
  NAND2_X1 U17001 ( .A1(n13638), .A2(n13637), .ZN(n13639) );
  AND2_X1 U17002 ( .A1(n13639), .A2(n13700), .ZN(n16564) );
  NOR2_X1 U17003 ( .A1(n14214), .A2(n11306), .ZN(n13640) );
  AOI21_X1 U17004 ( .B1(n16564), .B2(n14214), .A(n13640), .ZN(n13641) );
  OAI21_X1 U17005 ( .B1(n13642), .B2(n15493), .A(n13641), .ZN(P2_U2882) );
  AOI22_X1 U17006 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20164), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20163), .ZN(n13643) );
  OAI21_X1 U17007 ( .B1(n13098), .B2(n13650), .A(n13643), .ZN(P1_U2906) );
  INV_X1 U17008 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13645) );
  AOI22_X1 U17009 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13644) );
  OAI21_X1 U17010 ( .B1(n13645), .B2(n13650), .A(n13644), .ZN(P1_U2918) );
  INV_X1 U17011 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13647) );
  AOI22_X1 U17012 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13646) );
  OAI21_X1 U17013 ( .B1(n13647), .B2(n13650), .A(n13646), .ZN(P1_U2920) );
  AOI22_X1 U17014 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13648) );
  OAI21_X1 U17015 ( .B1(n21234), .B2(n13650), .A(n13648), .ZN(P1_U2910) );
  INV_X1 U17016 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13651) );
  AOI22_X1 U17017 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13649) );
  OAI21_X1 U17018 ( .B1(n13651), .B2(n13650), .A(n13649), .ZN(P1_U2919) );
  AOI22_X1 U17019 ( .A1(n20179), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20178), .ZN(n13654) );
  MUX2_X1 U17020 ( .A(DATAI_3_), .B(BUF1_REG_3__SCAN_IN), .S(n20236), .Z(
        n20269) );
  NAND2_X1 U17021 ( .A1(n13682), .A2(n20269), .ZN(n13678) );
  NAND2_X1 U17022 ( .A1(n13654), .A2(n13678), .ZN(P1_U2955) );
  AOI22_X1 U17023 ( .A1(n20179), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20178), .ZN(n13655) );
  MUX2_X1 U17024 ( .A(DATAI_2_), .B(BUF1_REG_2__SCAN_IN), .S(n20236), .Z(
        n20264) );
  NAND2_X1 U17025 ( .A1(n13682), .A2(n20264), .ZN(n13657) );
  NAND2_X1 U17026 ( .A1(n13655), .A2(n13657), .ZN(P1_U2954) );
  AOI22_X1 U17027 ( .A1(n20179), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20178), .ZN(n13656) );
  MUX2_X1 U17028 ( .A(DATAI_4_), .B(BUF1_REG_4__SCAN_IN), .S(n20236), .Z(
        n20273) );
  NAND2_X1 U17029 ( .A1(n13682), .A2(n20273), .ZN(n13662) );
  NAND2_X1 U17030 ( .A1(n13656), .A2(n13662), .ZN(P1_U2941) );
  AOI22_X1 U17031 ( .A1(n20179), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20178), .ZN(n13658) );
  NAND2_X1 U17032 ( .A1(n13658), .A2(n13657), .ZN(P1_U2939) );
  AOI22_X1 U17033 ( .A1(n20179), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20178), .ZN(n13661) );
  INV_X1 U17034 ( .A(DATAI_7_), .ZN(n13660) );
  NAND2_X1 U17035 ( .A1(n20236), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13659) );
  OAI21_X1 U17036 ( .B1(n20236), .B2(n13660), .A(n13659), .ZN(n20291) );
  NAND2_X1 U17037 ( .A1(n13682), .A2(n20291), .ZN(n13676) );
  NAND2_X1 U17038 ( .A1(n13661), .A2(n13676), .ZN(P1_U2944) );
  AOI22_X1 U17039 ( .A1(n20179), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20178), .ZN(n13663) );
  NAND2_X1 U17040 ( .A1(n13663), .A2(n13662), .ZN(P1_U2956) );
  AOI22_X1 U17041 ( .A1(n20179), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20178), .ZN(n13664) );
  MUX2_X1 U17042 ( .A(DATAI_1_), .B(BUF1_REG_1__SCAN_IN), .S(n20236), .Z(
        n20259) );
  NAND2_X1 U17043 ( .A1(n13682), .A2(n20259), .ZN(n13666) );
  NAND2_X1 U17044 ( .A1(n13664), .A2(n13666), .ZN(P1_U2938) );
  AOI22_X1 U17045 ( .A1(n20179), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20178), .ZN(n13665) );
  MUX2_X1 U17046 ( .A(DATAI_0_), .B(BUF1_REG_0__SCAN_IN), .S(n20236), .Z(
        n20250) );
  NAND2_X1 U17047 ( .A1(n13682), .A2(n20250), .ZN(n13670) );
  NAND2_X1 U17048 ( .A1(n13665), .A2(n13670), .ZN(P1_U2952) );
  AOI22_X1 U17049 ( .A1(n20179), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20178), .ZN(n13667) );
  NAND2_X1 U17050 ( .A1(n13667), .A2(n13666), .ZN(P1_U2953) );
  AOI22_X1 U17051 ( .A1(n20179), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20178), .ZN(n13668) );
  MUX2_X1 U17052 ( .A(DATAI_5_), .B(BUF1_REG_5__SCAN_IN), .S(n20236), .Z(
        n20277) );
  NAND2_X1 U17053 ( .A1(n13682), .A2(n20277), .ZN(n13672) );
  NAND2_X1 U17054 ( .A1(n13668), .A2(n13672), .ZN(P1_U2942) );
  AOI22_X1 U17055 ( .A1(n20179), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20178), .ZN(n13669) );
  MUX2_X1 U17056 ( .A(DATAI_6_), .B(BUF1_REG_6__SCAN_IN), .S(n20236), .Z(
        n20281) );
  NAND2_X1 U17057 ( .A1(n13682), .A2(n20281), .ZN(n13674) );
  NAND2_X1 U17058 ( .A1(n13669), .A2(n13674), .ZN(P1_U2943) );
  AOI22_X1 U17059 ( .A1(n20179), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20178), .ZN(n13671) );
  NAND2_X1 U17060 ( .A1(n13671), .A2(n13670), .ZN(P1_U2937) );
  AOI22_X1 U17061 ( .A1(n20179), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20178), .ZN(n13673) );
  NAND2_X1 U17062 ( .A1(n13673), .A2(n13672), .ZN(P1_U2957) );
  AOI22_X1 U17063 ( .A1(n20179), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20178), .ZN(n13675) );
  NAND2_X1 U17064 ( .A1(n13675), .A2(n13674), .ZN(P1_U2958) );
  AOI22_X1 U17065 ( .A1(n20179), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20178), .ZN(n13677) );
  NAND2_X1 U17066 ( .A1(n13677), .A2(n13676), .ZN(P1_U2959) );
  AOI22_X1 U17067 ( .A1(n20179), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20178), .ZN(n13679) );
  NAND2_X1 U17068 ( .A1(n13679), .A2(n13678), .ZN(P1_U2940) );
  AOI22_X1 U17069 ( .A1(n20179), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20178), .ZN(n13683) );
  INV_X1 U17070 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16646) );
  NOR2_X1 U17071 ( .A1(n20235), .A2(n16646), .ZN(n13680) );
  AOI21_X1 U17072 ( .B1(DATAI_11_), .B2(n20235), .A(n13680), .ZN(n14985) );
  INV_X1 U17073 ( .A(n14985), .ZN(n13681) );
  NAND2_X1 U17074 ( .A1(n13682), .A2(n13681), .ZN(n20172) );
  NAND2_X1 U17075 ( .A1(n13683), .A2(n20172), .ZN(P1_U2948) );
  INV_X1 U17076 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13685) );
  OR2_X1 U17077 ( .A1(n20222), .A2(n13685), .ZN(n15328) );
  OAI21_X1 U17078 ( .B1(n15131), .B2(n13767), .A(n15328), .ZN(n13691) );
  OR2_X1 U17079 ( .A1(n13688), .A2(n13687), .ZN(n13689) );
  NAND2_X1 U17080 ( .A1(n13686), .A2(n13689), .ZN(n14006) );
  NOR2_X1 U17081 ( .A1(n14006), .A2(n15135), .ZN(n13690) );
  AOI211_X1 U17082 ( .C1(n16270), .C2(n13767), .A(n13691), .B(n13690), .ZN(
        n13699) );
  NAND2_X1 U17083 ( .A1(n13692), .A2(n13693), .ZN(n13870) );
  OAI21_X1 U17084 ( .B1(n13693), .B2(n13692), .A(n13870), .ZN(n13694) );
  OAI211_X1 U17085 ( .C1(n13694), .C2(n14378), .A(n13016), .B(n12241), .ZN(
        n13695) );
  INV_X1 U17086 ( .A(n13695), .ZN(n13696) );
  OR2_X1 U17087 ( .A1(n13697), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15327) );
  NAND2_X1 U17088 ( .A1(n13697), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13866) );
  NAND3_X1 U17089 ( .A1(n15327), .A2(n9937), .A3(n20189), .ZN(n13698) );
  NAND2_X1 U17090 ( .A1(n13699), .A2(n13698), .ZN(P1_U2998) );
  NAND2_X1 U17091 ( .A1(n13701), .A2(n13700), .ZN(n13704) );
  INV_X1 U17092 ( .A(n13702), .ZN(n13703) );
  NAND2_X1 U17093 ( .A1(n13704), .A2(n13703), .ZN(n19189) );
  NOR2_X1 U17094 ( .A1(n13706), .A2(n13705), .ZN(n13709) );
  NAND2_X1 U17095 ( .A1(n13708), .A2(n13707), .ZN(n13726) );
  OAI211_X1 U17096 ( .C1(n13709), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15481), .B(n13726), .ZN(n13711) );
  NAND2_X1 U17097 ( .A1(n15490), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13710) );
  OAI211_X1 U17098 ( .C1(n19189), .C2(n14224), .A(n13711), .B(n13710), .ZN(
        P2_U2881) );
  AOI21_X1 U17099 ( .B1(n13713), .B2(n13727), .A(n13712), .ZN(n19176) );
  INV_X1 U17100 ( .A(n19176), .ZN(n13720) );
  INV_X1 U17101 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13715) );
  OAI21_X1 U17102 ( .B1(n13726), .B2(n13715), .A(n13714), .ZN(n13717) );
  NAND3_X1 U17103 ( .A1(n13717), .A2(n15481), .A3(n13716), .ZN(n13719) );
  NAND2_X1 U17104 ( .A1(n15490), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13718) );
  OAI211_X1 U17105 ( .C1(n13720), .C2(n14224), .A(n13719), .B(n13718), .ZN(
        P2_U2879) );
  XNOR2_X1 U17106 ( .A(n13716), .B(n13721), .ZN(n13725) );
  NOR2_X1 U17107 ( .A1(n13722), .A2(n13712), .ZN(n13723) );
  NOR2_X1 U17108 ( .A1(n10018), .A2(n13723), .ZN(n16481) );
  INV_X1 U17109 ( .A(n16481), .ZN(n14115) );
  MUX2_X1 U17110 ( .A(n11324), .B(n14115), .S(n14214), .Z(n13724) );
  OAI21_X1 U17111 ( .B1(n13725), .B2(n15493), .A(n13724), .ZN(P2_U2878) );
  XOR2_X1 U17112 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13726), .Z(n13730)
         );
  OAI21_X1 U17113 ( .B1(n13728), .B2(n13702), .A(n13727), .ZN(n16488) );
  MUX2_X1 U17114 ( .A(n16488), .B(n11315), .S(n15490), .Z(n13729) );
  OAI21_X1 U17115 ( .B1(n13730), .B2(n15493), .A(n13729), .ZN(P2_U2880) );
  OAI211_X1 U17116 ( .C1(n10028), .C2(n13733), .A(n13732), .B(n15481), .ZN(
        n13738) );
  NOR2_X1 U17117 ( .A1(n10018), .A2(n13735), .ZN(n13736) );
  NOR2_X1 U17118 ( .A1(n13734), .A2(n13736), .ZN(n19163) );
  NAND2_X1 U17119 ( .A1(n19163), .A2(n14214), .ZN(n13737) );
  OAI211_X1 U17120 ( .C1(n14214), .C2(n13739), .A(n13738), .B(n13737), .ZN(
        P2_U2877) );
  AND2_X1 U17121 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20932), .ZN(n13740) );
  NOR2_X1 U17122 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13906) );
  INV_X1 U17123 ( .A(n13906), .ZN(n20931) );
  NOR2_X1 U17124 ( .A1(n20664), .A2(n20931), .ZN(n16154) );
  AOI22_X1 U17125 ( .A1(n13741), .A2(n13740), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n16154), .ZN(n13742) );
  NAND2_X1 U17126 ( .A1(n20222), .A2(n13742), .ZN(n13743) );
  INV_X1 U17127 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14557) );
  INV_X1 U17128 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14643) );
  XNOR2_X1 U17129 ( .A(n13745), .B(n14643), .ZN(n14615) );
  NAND2_X1 U17130 ( .A1(n14831), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13746) );
  OAI21_X1 U17131 ( .B1(n14631), .B2(n13752), .A(n14809), .ZN(n20135) );
  INV_X1 U17132 ( .A(n20135), .ZN(n13984) );
  INV_X1 U17133 ( .A(n13746), .ZN(n13747) );
  INV_X1 U17134 ( .A(n13752), .ZN(n13750) );
  NAND2_X1 U17135 ( .A1(n13750), .A2(n13749), .ZN(n20129) );
  NOR2_X1 U17136 ( .A1(n13752), .A2(n13751), .ZN(n13761) );
  AND2_X1 U17137 ( .A1(n20936), .A2(n21085), .ZN(n13758) );
  AND2_X1 U17138 ( .A1(n13753), .A2(n13758), .ZN(n13757) );
  NAND2_X1 U17139 ( .A1(n12268), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13759) );
  INV_X1 U17140 ( .A(n13759), .ZN(n13754) );
  NOR2_X1 U17141 ( .A1(n13757), .A2(n13754), .ZN(n13755) );
  NAND2_X1 U17142 ( .A1(n13761), .A2(n13755), .ZN(n20104) );
  OAI22_X1 U17143 ( .A1(n20115), .A2(n13767), .B1(n13685), .B2(n14831), .ZN(
        n13756) );
  AOI21_X1 U17144 ( .B1(n20127), .B2(P1_EBX_REG_1__SCAN_IN), .A(n13756), .ZN(
        n13765) );
  NOR2_X1 U17145 ( .A1(n13759), .A2(n13758), .ZN(n13760) );
  INV_X1 U17146 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n21099) );
  NAND2_X1 U17147 ( .A1(n9811), .A2(n20214), .ZN(n13762) );
  OAI211_X1 U17148 ( .C1(n14630), .C2(P1_EBX_REG_1__SCAN_IN), .A(n13762), .B(
        n14517), .ZN(n13763) );
  AOI22_X1 U17149 ( .A1(n13685), .A2(n14839), .B1(n20126), .B2(n13948), .ZN(
        n13764) );
  OAI211_X1 U17150 ( .C1(n20528), .C2(n20129), .A(n13765), .B(n13764), .ZN(
        n13766) );
  AOI21_X1 U17151 ( .B1(n20084), .B2(n13767), .A(n13766), .ZN(n13768) );
  OAI21_X1 U17152 ( .B1(n13984), .B2(n14006), .A(n13768), .ZN(P1_U2839) );
  INV_X1 U17153 ( .A(n20250), .ZN(n13770) );
  INV_X1 U17154 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20167) );
  OAI222_X1 U17155 ( .A1(n14020), .A2(n14987), .B1(n14986), .B2(n13770), .C1(
        n14983), .C2(n20167), .ZN(P1_U2904) );
  INV_X1 U17156 ( .A(n20259), .ZN(n13771) );
  OAI222_X1 U17157 ( .A1(n14006), .A2(n14987), .B1(n14986), .B2(n13771), .C1(
        n14983), .C2(n12372), .ZN(P1_U2903) );
  NAND2_X1 U17158 ( .A1(n13772), .A2(n13686), .ZN(n13773) );
  INV_X1 U17159 ( .A(n20264), .ZN(n13774) );
  OAI222_X1 U17160 ( .A1(n15148), .A2(n14987), .B1(n14986), .B2(n13774), .C1(
        n14983), .C2(n12368), .ZN(P1_U2902) );
  INV_X1 U17161 ( .A(n14831), .ZN(n14688) );
  OR2_X1 U17162 ( .A1(n14839), .A2(n14688), .ZN(n14719) );
  OAI22_X1 U17163 ( .A1(n20080), .A2(n14021), .B1(n13775), .B2(n20104), .ZN(
        n13777) );
  INV_X1 U17164 ( .A(n12378), .ZN(n13909) );
  NOR2_X1 U17165 ( .A1(n13909), .A2(n20129), .ZN(n13776) );
  AOI211_X1 U17166 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n14719), .A(n13777), .B(
        n13776), .ZN(n13779) );
  OAI21_X1 U17167 ( .B1(n20084), .B2(n20133), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13778) );
  OAI211_X1 U17168 ( .C1(n13984), .C2(n14020), .A(n13779), .B(n13778), .ZN(
        P1_U2840) );
  INV_X1 U17169 ( .A(n13817), .ZN(n13821) );
  INV_X1 U17170 ( .A(n11118), .ZN(n13780) );
  NAND2_X1 U17171 ( .A1(n10759), .A2(n13780), .ZN(n13803) );
  NAND2_X1 U17172 ( .A1(n13781), .A2(n11717), .ZN(n13782) );
  NAND2_X1 U17173 ( .A1(n13782), .A2(n13787), .ZN(n13804) );
  NOR2_X1 U17174 ( .A1(n13783), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13786) );
  NOR2_X1 U17175 ( .A1(n13804), .A2(n13786), .ZN(n13790) );
  INV_X1 U17176 ( .A(n13784), .ZN(n13832) );
  NAND2_X1 U17177 ( .A1(n13832), .A2(n13785), .ZN(n13806) );
  INV_X1 U17178 ( .A(n13804), .ZN(n13789) );
  INV_X1 U17179 ( .A(n13786), .ZN(n13805) );
  NAND2_X1 U17180 ( .A1(n13787), .A2(n13805), .ZN(n13788) );
  OAI22_X1 U17181 ( .A1(n13790), .A2(n13806), .B1(n13789), .B2(n13788), .ZN(
        n13791) );
  OAI21_X1 U17182 ( .B1(n10157), .B2(n13803), .A(n13791), .ZN(n13793) );
  AOI21_X1 U17183 ( .B1(n14262), .B2(n13821), .A(n13793), .ZN(n15983) );
  INV_X1 U17184 ( .A(n13794), .ZN(n13797) );
  NOR2_X1 U17185 ( .A1(n11484), .A2(n13795), .ZN(n13796) );
  NAND2_X1 U17186 ( .A1(n13797), .A2(n13796), .ZN(n13801) );
  AND4_X1 U17187 ( .A1(n13801), .A2(n13800), .A3(n13799), .A4(n13798), .ZN(
        n14243) );
  INV_X1 U17188 ( .A(n14243), .ZN(n13826) );
  MUX2_X1 U17189 ( .A(n13802), .B(n15983), .S(n13826), .Z(n13841) );
  AND3_X1 U17190 ( .A1(n13804), .A2(n13805), .A3(n13803), .ZN(n13808) );
  AOI22_X1 U17191 ( .A1(n13806), .A2(n13805), .B1(n9927), .B2(n10759), .ZN(
        n13807) );
  MUX2_X1 U17192 ( .A(n13808), .B(n13807), .S(n13827), .Z(n13811) );
  INV_X1 U17193 ( .A(n13809), .ZN(n13810) );
  NAND2_X1 U17194 ( .A1(n13811), .A2(n13810), .ZN(n13812) );
  AOI21_X1 U17195 ( .B1(n10813), .B2(n13821), .A(n13812), .ZN(n15987) );
  OAI22_X1 U17196 ( .A1(n13841), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15987), .ZN(n13813) );
  INV_X1 U17197 ( .A(n13813), .ZN(n13825) );
  NOR2_X1 U17198 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19457) );
  INV_X1 U17199 ( .A(n19457), .ZN(n19455) );
  NAND2_X1 U17200 ( .A1(n13815), .A2(n13814), .ZN(n13819) );
  OAI21_X1 U17201 ( .B1(n13818), .B2(n13817), .A(n13816), .ZN(n14398) );
  INV_X1 U17202 ( .A(n14398), .ZN(n13822) );
  MUX2_X1 U17203 ( .A(n13819), .B(n10759), .S(n9932), .Z(n13820) );
  AOI21_X1 U17204 ( .B1(n19224), .B2(n13821), .A(n13820), .ZN(n14246) );
  OAI211_X1 U17205 ( .C1(n13822), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n14246), .ZN(n13823) );
  OAI21_X1 U17206 ( .B1(n14398), .B2(n20011), .A(n13823), .ZN(n13824) );
  AOI211_X1 U17207 ( .C1(n13825), .C2(n19455), .A(n14243), .B(n13824), .ZN(
        n13845) );
  MUX2_X1 U17208 ( .A(n13827), .B(n15987), .S(n13826), .Z(n13842) );
  OAI22_X1 U17209 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13842), .B1(
        n19455), .B2(n13841), .ZN(n13844) );
  INV_X1 U17210 ( .A(n13828), .ZN(n13829) );
  AOI22_X1 U17211 ( .A1(n13833), .A2(n13830), .B1(n11695), .B2(n13829), .ZN(
        n13831) );
  OAI21_X1 U17212 ( .B1(n13833), .B2(n13832), .A(n13831), .ZN(n20024) );
  OAI21_X1 U17213 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n13834), .ZN(n13837) );
  INV_X1 U17214 ( .A(n11484), .ZN(n13835) );
  NAND3_X1 U17215 ( .A1(n13835), .A2(n19356), .A3(n16089), .ZN(n13836) );
  OAI211_X1 U17216 ( .C1(n20035), .C2(n13838), .A(n13837), .B(n13836), .ZN(
        n13839) );
  AOI211_X1 U17217 ( .C1(n14243), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n20024), .B(n13839), .ZN(n13840) );
  OAI21_X1 U17218 ( .B1(n13842), .B2(n13841), .A(n13840), .ZN(n13843) );
  AOI221_X1 U17219 ( .B1(n13845), .B2(n16171), .C1(n13844), .C2(n16171), .A(
        n13843), .ZN(n16581) );
  AOI21_X1 U17220 ( .B1(n14396), .B2(n16581), .A(n19032), .ZN(n13850) );
  NOR2_X1 U17221 ( .A1(n13846), .A2(n20039), .ZN(n20044) );
  OAI21_X1 U17222 ( .B1(n13848), .B2(n13847), .A(n20044), .ZN(n13849) );
  NOR2_X1 U17223 ( .A1(n13850), .A2(n13849), .ZN(n19894) );
  OAI21_X1 U17224 ( .B1(n19894), .B2(n19032), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13853) );
  NOR2_X1 U17225 ( .A1(n19032), .A2(n13851), .ZN(n16170) );
  INV_X1 U17226 ( .A(n16170), .ZN(n13852) );
  NAND2_X1 U17227 ( .A1(n13853), .A2(n13852), .ZN(P2_U3593) );
  INV_X1 U17228 ( .A(n20269), .ZN(n13856) );
  OAI222_X1 U17229 ( .A1(n14173), .A2(n14987), .B1(n14986), .B2(n13856), .C1(
        n14983), .C2(n12422), .ZN(P1_U2901) );
  NAND2_X1 U17230 ( .A1(n13914), .A2(n14375), .ZN(n13861) );
  XNOR2_X1 U17231 ( .A(n13870), .B(n13869), .ZN(n13859) );
  INV_X1 U17232 ( .A(n13857), .ZN(n13858) );
  AOI21_X1 U17233 ( .B1(n13859), .B2(n20930), .A(n13858), .ZN(n13860) );
  INV_X1 U17234 ( .A(n13862), .ZN(n13863) );
  OR2_X1 U17235 ( .A1(n13864), .A2(n13863), .ZN(n13865) );
  NAND2_X1 U17236 ( .A1(n13866), .A2(n13865), .ZN(n13867) );
  INV_X1 U17237 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20232) );
  NAND2_X1 U17238 ( .A1(n13867), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13868) );
  INV_X1 U17239 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14520) );
  NAND2_X1 U17240 ( .A1(n13870), .A2(n13869), .ZN(n14351) );
  XNOR2_X1 U17241 ( .A(n14351), .B(n14349), .ZN(n13871) );
  OAI22_X1 U17242 ( .A1(n20238), .A2(n13872), .B1(n14378), .B2(n13871), .ZN(
        n13874) );
  OAI21_X1 U17243 ( .B1(n13873), .B2(n13874), .A(n14340), .ZN(n13875) );
  INV_X1 U17244 ( .A(n13875), .ZN(n20206) );
  NAND2_X1 U17245 ( .A1(n20206), .A2(n20189), .ZN(n13878) );
  NOR2_X1 U17246 ( .A1(n20222), .A2(n20870), .ZN(n20203) );
  NOR2_X1 U17247 ( .A1(n20193), .A2(n13979), .ZN(n13876) );
  AOI211_X1 U17248 ( .C1(n20182), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20203), .B(n13876), .ZN(n13877) );
  OAI211_X1 U17249 ( .C1(n15135), .C2(n14173), .A(n13878), .B(n13877), .ZN(
        P1_U2996) );
  NAND2_X1 U17250 ( .A1(n20527), .A2(n13892), .ZN(n13895) );
  OAI21_X1 U17251 ( .B1(n13536), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13879), .ZN(n20915) );
  INV_X1 U17252 ( .A(n20915), .ZN(n13880) );
  NAND2_X1 U17253 ( .A1(n13881), .A2(n13880), .ZN(n13891) );
  XNOR2_X1 U17254 ( .A(n13882), .B(n12088), .ZN(n13883) );
  NAND2_X1 U17255 ( .A1(n13884), .A2(n13883), .ZN(n13890) );
  MUX2_X1 U17256 ( .A(n13885), .B(n12088), .S(n10058), .Z(n13887) );
  NOR2_X1 U17257 ( .A1(n13887), .A2(n13886), .ZN(n13888) );
  NAND2_X1 U17258 ( .A1(n15345), .A2(n13888), .ZN(n13889) );
  OAI211_X1 U17259 ( .C1(n13892), .C2(n13891), .A(n13890), .B(n13889), .ZN(
        n13893) );
  INV_X1 U17260 ( .A(n13893), .ZN(n13894) );
  NAND2_X1 U17261 ( .A1(n13895), .A2(n13894), .ZN(n20913) );
  MUX2_X1 U17262 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20913), .S(
        n16115), .Z(n16126) );
  NAND2_X1 U17263 ( .A1(n16126), .A2(n20849), .ZN(n13899) );
  NOR2_X1 U17264 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20849), .ZN(n13903) );
  NAND2_X1 U17265 ( .A1(n13903), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13898) );
  MUX2_X1 U17266 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13896), .S(
        n16115), .Z(n16123) );
  AOI22_X1 U17267 ( .A1(n20849), .A2(n16123), .B1(n13903), .B2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13897) );
  AOI21_X1 U17268 ( .B1(n13899), .B2(n13898), .A(n13897), .ZN(n16138) );
  INV_X1 U17269 ( .A(n9951), .ZN(n13901) );
  NAND2_X1 U17270 ( .A1(n16138), .A2(n13901), .ZN(n13908) );
  NOR2_X1 U17271 ( .A1(n20130), .A2(n13069), .ZN(n13902) );
  MUX2_X1 U17272 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n13902), .S(
        n16115), .Z(n13905) );
  AND2_X1 U17273 ( .A1(n13903), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13904) );
  AOI21_X1 U17274 ( .B1(n13905), .B2(n20849), .A(n13904), .ZN(n16136) );
  AND3_X1 U17275 ( .A1(n13908), .A2(n20057), .A3(n16136), .ZN(n13907) );
  OAI21_X1 U17276 ( .B1(n13907), .B2(n16372), .A(n20406), .ZN(n20234) );
  NAND3_X1 U17277 ( .A1(n13908), .A2(n16136), .A3(n16368), .ZN(n16148) );
  INV_X1 U17278 ( .A(n16148), .ZN(n13911) );
  NAND2_X1 U17279 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20664), .ZN(n13923) );
  INV_X1 U17280 ( .A(n13923), .ZN(n15340) );
  OAI22_X1 U17281 ( .A1(n13562), .A2(n20779), .B1(n13909), .B2(n15340), .ZN(
        n13910) );
  OAI21_X1 U17282 ( .B1(n13911), .B2(n13910), .A(n20234), .ZN(n13912) );
  OAI21_X1 U17283 ( .B1(n20234), .B2(n20690), .A(n13912), .ZN(P1_U3478) );
  NOR2_X1 U17284 ( .A1(n20655), .A2(n15340), .ZN(n13917) );
  NAND2_X1 U17285 ( .A1(n13913), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13921) );
  NOR2_X1 U17286 ( .A1(n13921), .A2(n20779), .ZN(n13915) );
  MUX2_X1 U17287 ( .A(n13915), .B(n20787), .S(n13914), .Z(n13916) );
  OAI21_X1 U17288 ( .B1(n13917), .B2(n13916), .A(n20234), .ZN(n13918) );
  OAI21_X1 U17289 ( .B1(n13020), .B2(n20234), .A(n13918), .ZN(P1_U3476) );
  INV_X1 U17290 ( .A(n20234), .ZN(n13928) );
  NAND2_X1 U17291 ( .A1(n13914), .A2(n13919), .ZN(n20497) );
  INV_X1 U17292 ( .A(n20497), .ZN(n20429) );
  OAI22_X1 U17293 ( .A1(n20429), .A2(n13921), .B1(n20719), .B2(n13913), .ZN(
        n13922) );
  NAND2_X1 U17294 ( .A1(n13922), .A2(n20629), .ZN(n13925) );
  AOI21_X1 U17295 ( .B1(n20238), .B2(n21085), .A(n20779), .ZN(n13924) );
  AOI22_X1 U17296 ( .A1(n13925), .A2(n13924), .B1(n13923), .B2(n20527), .ZN(
        n13927) );
  NAND2_X1 U17297 ( .A1(n13928), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13926) );
  OAI21_X1 U17298 ( .B1(n13928), .B2(n13927), .A(n13926), .ZN(P1_U3475) );
  INV_X1 U17299 ( .A(n13929), .ZN(n13932) );
  XNOR2_X1 U17300 ( .A(n13930), .B(n10006), .ZN(n19138) );
  INV_X1 U17301 ( .A(n19138), .ZN(n13931) );
  OAI222_X1 U17302 ( .A1(n19250), .A2(n19297), .B1(n13932), .B2(n19291), .C1(
        n13931), .C2(n19252), .ZN(P2_U2905) );
  XNOR2_X1 U17303 ( .A(n13732), .B(n13933), .ZN(n13939) );
  INV_X1 U17304 ( .A(n13934), .ZN(n13935) );
  NOR2_X1 U17305 ( .A1(n13734), .A2(n13936), .ZN(n13937) );
  NOR2_X1 U17306 ( .A1(n13935), .A2(n13937), .ZN(n16533) );
  INV_X1 U17307 ( .A(n16533), .ZN(n14083) );
  MUX2_X1 U17308 ( .A(n10190), .B(n14083), .S(n14214), .Z(n13938) );
  OAI21_X1 U17309 ( .B1(n13939), .B2(n15493), .A(n13938), .ZN(P2_U2876) );
  OAI21_X1 U17310 ( .B1(n13935), .B2(n13941), .A(n13940), .ZN(n19149) );
  INV_X1 U17311 ( .A(n13942), .ZN(n13945) );
  OAI211_X1 U17312 ( .C1(n13945), .C2(n13944), .A(n15481), .B(n14057), .ZN(
        n13947) );
  NAND2_X1 U17313 ( .A1(n15490), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13946) );
  OAI211_X1 U17314 ( .C1(n19149), .C2(n15490), .A(n13947), .B(n13946), .ZN(
        P2_U2875) );
  INV_X1 U17315 ( .A(n20129), .ZN(n13982) );
  INV_X1 U17316 ( .A(n20655), .ZN(n20247) );
  INV_X1 U17317 ( .A(n13993), .ZN(n14467) );
  NAND2_X1 U17318 ( .A1(n13948), .A2(n14467), .ZN(n13953) );
  INV_X1 U17319 ( .A(n13949), .ZN(n13950) );
  OR2_X1 U17320 ( .A1(n13951), .A2(n13950), .ZN(n13952) );
  INV_X1 U17321 ( .A(n14236), .ZN(n14465) );
  INV_X1 U17322 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13954) );
  MUX2_X1 U17323 ( .A(n14465), .B(n14500), .S(n13954), .Z(n13956) );
  NAND2_X1 U17324 ( .A1(n14465), .A2(n14630), .ZN(n14489) );
  OAI21_X1 U17325 ( .B1(n14467), .B2(n20232), .A(n14489), .ZN(n13955) );
  NOR2_X1 U17326 ( .A1(n13956), .A2(n13955), .ZN(n13958) );
  NAND2_X1 U17327 ( .A1(n13959), .A2(n13958), .ZN(n13960) );
  NAND2_X1 U17328 ( .A1(n13973), .A2(n13960), .ZN(n20224) );
  INV_X1 U17329 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20223) );
  AOI21_X1 U17330 ( .B1(n14839), .B2(n13685), .A(n14688), .ZN(n13964) );
  NAND2_X1 U17331 ( .A1(n20133), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13963) );
  NOR2_X1 U17332 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n20075), .ZN(n13961) );
  NAND2_X1 U17333 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(n13961), .ZN(n13962) );
  OAI211_X1 U17334 ( .C1(n20223), .C2(n13964), .A(n13963), .B(n13962), .ZN(
        n13965) );
  AOI21_X1 U17335 ( .B1(n20127), .B2(P1_EBX_REG_2__SCAN_IN), .A(n13965), .ZN(
        n13966) );
  OAI21_X1 U17336 ( .B1(n20080), .B2(n20224), .A(n13966), .ZN(n13968) );
  NOR2_X1 U17337 ( .A1(n20140), .A2(n15153), .ZN(n13967) );
  AOI211_X1 U17338 ( .C1(n13982), .C2(n20247), .A(n13968), .B(n13967), .ZN(
        n13969) );
  OAI21_X1 U17339 ( .B1(n13984), .B2(n15148), .A(n13969), .ZN(P1_U2838) );
  NAND3_X1 U17340 ( .A1(n14839), .A2(P1_REIP_REG_2__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n20134) );
  MUX2_X1 U17341 ( .A(n14510), .B(n14517), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13971) );
  INV_X1 U17342 ( .A(n13597), .ZN(n14511) );
  NAND2_X1 U17343 ( .A1(n14511), .A2(n14520), .ZN(n13970) );
  NAND2_X1 U17344 ( .A1(n13971), .A2(n13970), .ZN(n13972) );
  AND2_X1 U17345 ( .A1(n13973), .A2(n13972), .ZN(n13974) );
  NOR2_X1 U17346 ( .A1(n14090), .A2(n13974), .ZN(n20204) );
  INV_X1 U17347 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14174) );
  OAI221_X1 U17348 ( .B1(n20075), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n20075), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n14831), .ZN(n13975) );
  AOI22_X1 U17349 ( .A1(n20133), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13975), .ZN(n13976) );
  OAI21_X1 U17350 ( .B1(n20104), .B2(n14174), .A(n13976), .ZN(n13977) );
  AOI21_X1 U17351 ( .B1(n20126), .B2(n20204), .A(n13977), .ZN(n13978) );
  OAI21_X1 U17352 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n20134), .A(n13978), .ZN(
        n13981) );
  NOR2_X1 U17353 ( .A1(n20140), .A2(n13979), .ZN(n13980) );
  AOI211_X1 U17354 ( .C1(n13982), .C2(n20527), .A(n13981), .B(n13980), .ZN(
        n13983) );
  OAI21_X1 U17355 ( .B1(n13984), .B2(n14173), .A(n13983), .ZN(P1_U2837) );
  OAI21_X1 U17356 ( .B1(n13985), .B2(n13988), .A(n13987), .ZN(n16299) );
  INV_X1 U17357 ( .A(n20277), .ZN(n13989) );
  OAI222_X1 U17358 ( .A1(n16299), .A2(n14987), .B1(n14986), .B2(n13989), .C1(
        n14983), .C2(n12471), .ZN(P1_U2899) );
  NAND2_X1 U17359 ( .A1(n13990), .A2(n14467), .ZN(n13991) );
  OAI21_X4 U17360 ( .B1(n13992), .B2(n14634), .A(n13991), .ZN(n14897) );
  NAND2_X2 U17361 ( .A1(n13015), .A2(n14897), .ZN(n14908) );
  MUX2_X1 U17362 ( .A(n14514), .B(n14236), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13996) );
  NAND2_X1 U17363 ( .A1(n14630), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13994) );
  AND2_X1 U17364 ( .A1(n14489), .A2(n13994), .ZN(n13995) );
  NAND2_X1 U17365 ( .A1(n13996), .A2(n13995), .ZN(n14089) );
  INV_X1 U17366 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13997) );
  NAND2_X1 U17367 ( .A1(n14504), .A2(n13997), .ZN(n14000) );
  NAND2_X1 U17368 ( .A1(n14480), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13998) );
  OAI211_X1 U17369 ( .C1(n14630), .C2(P1_EBX_REG_5__SCAN_IN), .A(n14236), .B(
        n13998), .ZN(n13999) );
  AOI21_X1 U17370 ( .B1(n14090), .B2(n14089), .A(n14001), .ZN(n14003) );
  NOR2_X1 U17371 ( .A1(n14003), .A2(n14170), .ZN(n20117) );
  AOI22_X1 U17372 ( .A1(n20117), .A2(n14906), .B1(n14905), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n14004) );
  OAI21_X1 U17373 ( .B1(n16299), .B2(n14908), .A(n14004), .ZN(P1_U2867) );
  XNOR2_X1 U17374 ( .A(n13948), .B(n14467), .ZN(n15333) );
  AOI22_X1 U17375 ( .A1(n14906), .A2(n15333), .B1(n14905), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n14005) );
  OAI21_X1 U17376 ( .B1(n14006), .B2(n14908), .A(n14005), .ZN(P1_U2871) );
  INV_X1 U17377 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20159) );
  INV_X1 U17378 ( .A(n20273), .ZN(n14949) );
  INV_X1 U17379 ( .A(n14007), .ZN(n14008) );
  INV_X1 U17380 ( .A(n20187), .ZN(n14091) );
  OAI222_X1 U17381 ( .A1(n14983), .A2(n20159), .B1(n14986), .B2(n14949), .C1(
        n14987), .C2(n14091), .ZN(P1_U2900) );
  XOR2_X1 U17382 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n14009), .Z(
        n14010) );
  XNOR2_X1 U17383 ( .A(n14011), .B(n14010), .ZN(n14037) );
  XOR2_X1 U17384 ( .A(n14013), .B(n14012), .Z(n14035) );
  INV_X1 U17385 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n14014) );
  OAI22_X1 U17386 ( .A1(n16506), .A2(n14015), .B1(n14014), .B2(n19181), .ZN(
        n14016) );
  AOI21_X1 U17387 ( .B1(n16496), .B2(n14147), .A(n14016), .ZN(n14017) );
  OAI21_X1 U17388 ( .B1(n13532), .B2(n14136), .A(n14017), .ZN(n14018) );
  AOI21_X1 U17389 ( .B1(n14035), .B2(n16503), .A(n14018), .ZN(n14019) );
  OAI21_X1 U17390 ( .B1(n14037), .B2(n19333), .A(n14019), .ZN(P2_U3011) );
  OAI222_X1 U17391 ( .A1(n14021), .A2(n14898), .B1(n14897), .B2(n13775), .C1(
        n14020), .C2(n14908), .ZN(P1_U2872) );
  XNOR2_X1 U17392 ( .A(n14057), .B(n14056), .ZN(n14025) );
  NOR2_X1 U17393 ( .A1(n14214), .A2(n14022), .ZN(n14023) );
  AOI21_X1 U17394 ( .B1(n16523), .B2(n14214), .A(n14023), .ZN(n14024) );
  OAI21_X1 U17395 ( .B1(n14025), .B2(n15493), .A(n14024), .ZN(P2_U2874) );
  XNOR2_X1 U17396 ( .A(n14027), .B(n14026), .ZN(n19266) );
  NOR2_X1 U17397 ( .A1(n14014), .A2(n19181), .ZN(n14028) );
  AOI221_X1 U17398 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14031), .C1(
        n14030), .C2(n14029), .A(n14028), .ZN(n14033) );
  NAND2_X1 U17399 ( .A1(n10813), .A2(n16565), .ZN(n14032) );
  OAI211_X1 U17400 ( .C1(n19266), .C2(n16544), .A(n14033), .B(n14032), .ZN(
        n14034) );
  AOI21_X1 U17401 ( .B1(n16566), .B2(n14035), .A(n14034), .ZN(n14036) );
  OAI21_X1 U17402 ( .B1(n16552), .B2(n14037), .A(n14036), .ZN(P2_U3043) );
  INV_X1 U17403 ( .A(n14039), .ZN(n14040) );
  AOI21_X1 U17404 ( .B1(n14041), .B2(n14038), .A(n14040), .ZN(n14211) );
  INV_X1 U17405 ( .A(n14042), .ZN(n14048) );
  INV_X1 U17406 ( .A(n14043), .ZN(n14046) );
  INV_X1 U17407 ( .A(n14044), .ZN(n14045) );
  NAND2_X1 U17408 ( .A1(n14046), .A2(n14045), .ZN(n14047) );
  NAND2_X1 U17409 ( .A1(n14048), .A2(n14047), .ZN(n19121) );
  AOI22_X1 U17410 ( .A1(n19233), .A2(BUF2_REG_16__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n14051) );
  AOI22_X1 U17411 ( .A1(n16430), .A2(n14049), .B1(n19284), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n14050) );
  OAI211_X1 U17412 ( .C1(n15552), .C2(n19121), .A(n14051), .B(n14050), .ZN(
        n14052) );
  AOI21_X1 U17413 ( .B1(n14211), .B2(n19286), .A(n14052), .ZN(n14053) );
  INV_X1 U17414 ( .A(n14053), .ZN(P2_U2903) );
  AND2_X1 U17415 ( .A1(n13943), .A2(n14054), .ZN(n14177) );
  INV_X1 U17416 ( .A(n14177), .ZN(n14059) );
  OAI21_X1 U17417 ( .B1(n14057), .B2(n14056), .A(n14055), .ZN(n14058) );
  NAND3_X1 U17418 ( .A1(n14059), .A2(n15481), .A3(n14058), .ZN(n14064) );
  NOR2_X1 U17419 ( .A1(n13191), .A2(n14061), .ZN(n14062) );
  NOR2_X1 U17420 ( .A1(n14060), .A2(n14062), .ZN(n19139) );
  NAND2_X1 U17421 ( .A1(n19139), .A2(n14214), .ZN(n14063) );
  OAI211_X1 U17422 ( .C1(n14214), .C2(n14065), .A(n14064), .B(n14063), .ZN(
        P2_U2873) );
  NAND2_X1 U17423 ( .A1(n10206), .A2(n14066), .ZN(n14067) );
  XNOR2_X1 U17424 ( .A(n16486), .B(n14067), .ZN(n14076) );
  AOI22_X1 U17425 ( .A1(n14068), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19229), .ZN(n14069) );
  OAI21_X1 U17426 ( .B1(n19215), .B2(n11315), .A(n14069), .ZN(n14070) );
  AOI211_X1 U17427 ( .C1(n19199), .C2(P2_REIP_REG_7__SCAN_IN), .A(n19328), .B(
        n14070), .ZN(n14074) );
  AOI21_X1 U17428 ( .B1(n14072), .B2(n14071), .A(n13402), .ZN(n19246) );
  INV_X1 U17429 ( .A(n19214), .ZN(n19200) );
  NAND2_X1 U17430 ( .A1(n19246), .A2(n19200), .ZN(n14073) );
  OAI211_X1 U17431 ( .C1(n16488), .C2(n19202), .A(n14074), .B(n14073), .ZN(
        n14075) );
  AOI21_X1 U17432 ( .B1(n14076), .B2(n19191), .A(n14075), .ZN(n14077) );
  INV_X1 U17433 ( .A(n14077), .ZN(P2_U2848) );
  NAND2_X1 U17434 ( .A1(n10206), .A2(n14078), .ZN(n14079) );
  XNOR2_X1 U17435 ( .A(n16460), .B(n14079), .ZN(n14080) );
  NAND2_X1 U17436 ( .A1(n14080), .A2(n19191), .ZN(n14087) );
  INV_X1 U17437 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17438 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19229), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n19168), .ZN(n14081) );
  OAI211_X1 U17439 ( .C1(n19220), .C2(n14082), .A(n14081), .B(n19181), .ZN(
        n14085) );
  NOR2_X1 U17440 ( .A1(n14083), .A2(n19202), .ZN(n14084) );
  AOI211_X1 U17441 ( .C1(n19200), .C2(n16530), .A(n14085), .B(n14084), .ZN(
        n14086) );
  OAI211_X1 U17442 ( .C1(n19217), .C2(n14088), .A(n14087), .B(n14086), .ZN(
        P2_U2844) );
  XNOR2_X1 U17443 ( .A(n14090), .B(n14089), .ZN(n20125) );
  INV_X1 U17444 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21267) );
  OAI222_X1 U17445 ( .A1(n14908), .A2(n14091), .B1(n14898), .B2(n20125), .C1(
        n14897), .C2(n21267), .ZN(P1_U2868) );
  XOR2_X1 U17446 ( .A(n13987), .B(n14092), .Z(n20107) );
  INV_X1 U17447 ( .A(n20107), .ZN(n14143) );
  MUX2_X1 U17448 ( .A(n14514), .B(n14236), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n14095) );
  NAND2_X1 U17449 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14630), .ZN(
        n14093) );
  AND2_X1 U17450 ( .A1(n14489), .A2(n14093), .ZN(n14094) );
  NAND2_X1 U17451 ( .A1(n14095), .A2(n14094), .ZN(n14169) );
  XOR2_X1 U17452 ( .A(n14170), .B(n14169), .Z(n20100) );
  INV_X1 U17453 ( .A(n20100), .ZN(n14096) );
  INV_X1 U17454 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21296) );
  OAI222_X1 U17455 ( .A1(n14908), .A2(n14143), .B1(n14898), .B2(n14096), .C1(
        n14897), .C2(n21296), .ZN(P1_U2866) );
  NAND2_X1 U17456 ( .A1(n10206), .A2(n14097), .ZN(n14098) );
  XNOR2_X1 U17457 ( .A(n16495), .B(n14098), .ZN(n14099) );
  NAND2_X1 U17458 ( .A1(n14099), .A2(n19191), .ZN(n14108) );
  OAI21_X1 U17459 ( .B1(n14102), .B2(n14101), .A(n14100), .ZN(n19251) );
  INV_X1 U17460 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19924) );
  OAI21_X1 U17461 ( .B1(n19924), .B2(n19220), .A(n19181), .ZN(n14104) );
  NOR2_X1 U17462 ( .A1(n19155), .A2(n16507), .ZN(n14103) );
  AOI211_X1 U17463 ( .C1(n19168), .C2(P2_EBX_REG_5__SCAN_IN), .A(n14104), .B(
        n14103), .ZN(n14105) );
  OAI21_X1 U17464 ( .B1(n19214), .B2(n19251), .A(n14105), .ZN(n14106) );
  AOI21_X1 U17465 ( .B1(n16564), .B2(n19223), .A(n14106), .ZN(n14107) );
  OAI211_X1 U17466 ( .C1(n19217), .C2(n14109), .A(n14108), .B(n14107), .ZN(
        P2_U2850) );
  NAND2_X1 U17467 ( .A1(n10206), .A2(n14110), .ZN(n14111) );
  XNOR2_X1 U17468 ( .A(n16478), .B(n14111), .ZN(n14112) );
  NAND2_X1 U17469 ( .A1(n14112), .A2(n19191), .ZN(n14119) );
  INV_X1 U17470 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U17471 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n19229), .B1(
        P2_EBX_REG_9__SCAN_IN), .B2(n19168), .ZN(n14113) );
  OAI211_X1 U17472 ( .C1(n19220), .C2(n14114), .A(n14113), .B(n19181), .ZN(
        n14117) );
  NOR2_X1 U17473 ( .A1(n14115), .A2(n19202), .ZN(n14116) );
  AOI211_X1 U17474 ( .C1(n15960), .C2(n19200), .A(n14117), .B(n14116), .ZN(
        n14118) );
  OAI211_X1 U17475 ( .C1(n19217), .C2(n14120), .A(n14119), .B(n14118), .ZN(
        P2_U2846) );
  NOR2_X1 U17476 ( .A1(n14122), .A2(n14121), .ZN(n14129) );
  AOI21_X1 U17477 ( .B1(n19750), .B2(n19779), .A(n19629), .ZN(n14123) );
  AOI21_X1 U17478 ( .B1(n14129), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n14123), .ZN(n14127) );
  NAND3_X1 U17479 ( .A1(n20011), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19751) );
  NOR2_X1 U17480 ( .A1(n19751), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19745) );
  INV_X1 U17481 ( .A(n19745), .ZN(n14139) );
  OAI211_X1 U17482 ( .C1(n14124), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n14139), 
        .B(n19599), .ZN(n14125) );
  NAND2_X1 U17483 ( .A1(n14125), .A2(n19833), .ZN(n14126) );
  INV_X1 U17484 ( .A(n19747), .ZN(n19733) );
  INV_X1 U17485 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14142) );
  INV_X1 U17486 ( .A(n14128), .ZN(n14131) );
  INV_X1 U17487 ( .A(n14129), .ZN(n19489) );
  OAI21_X1 U17488 ( .B1(n10956), .B2(n19745), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14130) );
  OAI21_X1 U17489 ( .B1(n14131), .B2(n19489), .A(n14130), .ZN(n19746) );
  INV_X1 U17490 ( .A(n19390), .ZN(n14133) );
  NAND2_X1 U17491 ( .A1(n14134), .A2(n14133), .ZN(n19343) );
  AOI22_X1 U17492 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19388), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19389), .ZN(n19763) );
  AOI22_X1 U17493 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19389), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19388), .ZN(n19843) );
  INV_X1 U17494 ( .A(n19843), .ZN(n19760) );
  AOI22_X1 U17495 ( .A1(n19742), .A2(n19840), .B1(n19784), .B2(n19760), .ZN(
        n14138) );
  OAI21_X1 U17496 ( .B1(n19343), .B2(n14139), .A(n14138), .ZN(n14140) );
  AOI21_X1 U17497 ( .B1(n19746), .B2(n14132), .A(n14140), .ZN(n14141) );
  OAI21_X1 U17498 ( .B1(n19733), .B2(n14142), .A(n14141), .ZN(P2_U3144) );
  INV_X1 U17499 ( .A(n20281), .ZN(n14144) );
  OAI222_X1 U17500 ( .A1(n14983), .A2(n20156), .B1(n14986), .B2(n14144), .C1(
        n14987), .C2(n14143), .ZN(P1_U2898) );
  NAND2_X1 U17501 ( .A1(n10206), .A2(n14145), .ZN(n14146) );
  XNOR2_X1 U17502 ( .A(n14147), .B(n14146), .ZN(n14157) );
  NOR2_X1 U17503 ( .A1(n19988), .A2(n19203), .ZN(n14156) );
  OAI22_X1 U17504 ( .A1(n19215), .A2(n14148), .B1(n14014), .B2(n19220), .ZN(
        n14149) );
  INV_X1 U17505 ( .A(n14149), .ZN(n14154) );
  INV_X1 U17506 ( .A(n14150), .ZN(n14152) );
  OAI22_X1 U17507 ( .A1(n19214), .A2(n19266), .B1(n19155), .B2(n14015), .ZN(
        n14151) );
  AOI21_X1 U17508 ( .B1(n14152), .B2(n19110), .A(n14151), .ZN(n14153) );
  OAI211_X1 U17509 ( .C1(n13532), .C2(n19202), .A(n14154), .B(n14153), .ZN(
        n14155) );
  AOI211_X1 U17510 ( .C1(n14157), .C2(n19191), .A(n14156), .B(n14155), .ZN(
        n14158) );
  INV_X1 U17511 ( .A(n14158), .ZN(P2_U2852) );
  INV_X1 U17512 ( .A(n14159), .ZN(n14208) );
  NAND2_X1 U17513 ( .A1(n14161), .A2(n14160), .ZN(n14162) );
  AND2_X1 U17514 ( .A1(n14208), .A2(n14162), .ZN(n20095) );
  INV_X1 U17515 ( .A(n20095), .ZN(n14186) );
  INV_X1 U17516 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14163) );
  NAND2_X1 U17517 ( .A1(n14504), .A2(n14163), .ZN(n14166) );
  NAND2_X1 U17518 ( .A1(n14517), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14164) );
  OAI211_X1 U17519 ( .C1(n14630), .C2(P1_EBX_REG_7__SCAN_IN), .A(n14236), .B(
        n14164), .ZN(n14165) );
  AND2_X1 U17520 ( .A1(n14166), .A2(n14165), .ZN(n14168) );
  AOI21_X1 U17521 ( .B1(n14170), .B2(n14169), .A(n14168), .ZN(n14171) );
  NOR2_X1 U17522 ( .A1(n10226), .A2(n14171), .ZN(n20094) );
  AOI22_X1 U17523 ( .A1(n20094), .A2(n14906), .B1(n14905), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n14172) );
  OAI21_X1 U17524 ( .B1(n14186), .B2(n14908), .A(n14172), .ZN(P1_U2865) );
  INV_X1 U17525 ( .A(n20204), .ZN(n14175) );
  OAI222_X1 U17526 ( .A1(n14175), .A2(n14898), .B1(n14897), .B2(n14174), .C1(
        n14908), .C2(n14173), .ZN(P1_U2869) );
  OAI222_X1 U17527 ( .A1(n20224), .A2(n14898), .B1(n14897), .B2(n13954), .C1(
        n14908), .C2(n15148), .ZN(P1_U2870) );
  XNOR2_X1 U17528 ( .A(n14177), .B(n14176), .ZN(n14183) );
  INV_X1 U17529 ( .A(n14060), .ZN(n14180) );
  INV_X1 U17530 ( .A(n14178), .ZN(n14179) );
  AOI21_X1 U17531 ( .B1(n14180), .B2(n14179), .A(n14212), .ZN(n19128) );
  NOR2_X1 U17532 ( .A1(n14214), .A2(n11343), .ZN(n14181) );
  AOI21_X1 U17533 ( .B1(n19128), .B2(n14214), .A(n14181), .ZN(n14182) );
  OAI21_X1 U17534 ( .B1(n14183), .B2(n15493), .A(n14182), .ZN(P2_U2872) );
  INV_X1 U17535 ( .A(n20291), .ZN(n14185) );
  OAI222_X1 U17536 ( .A1(n14186), .A2(n14987), .B1(n14986), .B2(n14185), .C1(
        n14184), .C2(n14983), .ZN(P1_U2897) );
  XNOR2_X1 U17537 ( .A(n9910), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14188) );
  XNOR2_X1 U17538 ( .A(n14188), .B(n14187), .ZN(n19331) );
  XOR2_X1 U17539 ( .A(n14189), .B(n14190), .Z(n19330) );
  NAND2_X1 U17540 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19172), .ZN(n14191) );
  OAI221_X1 U17541 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16554), .C1(
        n16556), .C2(n16571), .A(n14191), .ZN(n14197) );
  INV_X1 U17542 ( .A(n14192), .ZN(n14193) );
  XNOR2_X1 U17543 ( .A(n14194), .B(n14193), .ZN(n19260) );
  INV_X1 U17544 ( .A(n19260), .ZN(n14195) );
  OAI22_X1 U17545 ( .A1(n19201), .A2(n15976), .B1(n14195), .B2(n16544), .ZN(
        n14196) );
  AOI211_X1 U17546 ( .C1(n19330), .C2(n16563), .A(n14197), .B(n14196), .ZN(
        n14198) );
  OAI21_X1 U17547 ( .B1(n15966), .B2(n19331), .A(n14198), .ZN(P2_U3042) );
  INV_X1 U17548 ( .A(n14199), .ZN(n14221) );
  NOR2_X1 U17549 ( .A1(n14039), .A2(n14221), .ZN(n14220) );
  NAND2_X1 U17550 ( .A1(n14220), .A2(n14200), .ZN(n14334) );
  OAI21_X1 U17551 ( .B1(n14220), .B2(n14200), .A(n14334), .ZN(n14392) );
  OAI21_X1 U17552 ( .B1(n15568), .B2(n14201), .A(n15558), .ZN(n19092) );
  AOI22_X1 U17553 ( .A1(n19233), .A2(BUF2_REG_18__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n14204) );
  AOI22_X1 U17554 ( .A1(n16430), .A2(n14202), .B1(n19284), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n14203) );
  OAI211_X1 U17555 ( .C1(n15552), .C2(n19092), .A(n14204), .B(n14203), .ZN(
        n14205) );
  INV_X1 U17556 ( .A(n14205), .ZN(n14206) );
  OAI21_X1 U17557 ( .B1(n14392), .B2(n19257), .A(n14206), .ZN(P2_U2901) );
  AND2_X1 U17558 ( .A1(n14208), .A2(n14207), .ZN(n14210) );
  OR2_X1 U17559 ( .A1(n14210), .A2(n14209), .ZN(n14383) );
  OAI222_X1 U17560 ( .A1(n14383), .A2(n14987), .B1(n14983), .B2(n20153), .C1(
        n14931), .C2(n14986), .ZN(P1_U2896) );
  NAND2_X1 U17561 ( .A1(n14211), .A2(n15481), .ZN(n14216) );
  OAI21_X1 U17562 ( .B1(n14213), .B2(n14212), .A(n14217), .ZN(n15905) );
  INV_X1 U17563 ( .A(n15905), .ZN(n19117) );
  NAND2_X1 U17564 ( .A1(n14214), .A2(n19117), .ZN(n14215) );
  OAI211_X1 U17565 ( .C1(n14214), .C2(n11349), .A(n14216), .B(n14215), .ZN(
        P2_U2871) );
  AND2_X1 U17566 ( .A1(n14218), .A2(n14217), .ZN(n14219) );
  OR2_X1 U17567 ( .A1(n14219), .A2(n14389), .ZN(n15890) );
  AOI21_X1 U17568 ( .B1(n14221), .B2(n14039), .A(n14220), .ZN(n15564) );
  NAND2_X1 U17569 ( .A1(n15564), .A2(n15481), .ZN(n14223) );
  NAND2_X1 U17570 ( .A1(n15490), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14222) );
  OAI211_X1 U17571 ( .C1(n15890), .C2(n14224), .A(n14223), .B(n14222), .ZN(
        P2_U2870) );
  INV_X1 U17572 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14835) );
  MUX2_X1 U17573 ( .A(n14465), .B(n14500), .S(n14835), .Z(n14227) );
  NAND2_X1 U17574 ( .A1(n14630), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14225) );
  NAND2_X1 U17575 ( .A1(n14489), .A2(n14225), .ZN(n14226) );
  NOR2_X1 U17576 ( .A1(n14227), .A2(n14226), .ZN(n14228) );
  NAND2_X1 U17577 ( .A1(n14229), .A2(n14228), .ZN(n14230) );
  AND2_X1 U17578 ( .A1(n14239), .A2(n14230), .ZN(n16341) );
  INV_X1 U17579 ( .A(n16341), .ZN(n14231) );
  OAI222_X1 U17580 ( .A1(n14231), .A2(n14898), .B1(n14897), .B2(n14835), .C1(
        n14908), .C2(n14383), .ZN(P1_U2864) );
  NOR2_X1 U17581 ( .A1(n14209), .A2(n14233), .ZN(n14234) );
  OR2_X1 U17582 ( .A1(n14232), .A2(n14234), .ZN(n14408) );
  NAND2_X1 U17583 ( .A1(n14517), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14235) );
  OAI211_X1 U17584 ( .C1(n14630), .C2(P1_EBX_REG_9__SCAN_IN), .A(n14236), .B(
        n14235), .ZN(n14237) );
  OAI21_X1 U17585 ( .B1(n14510), .B2(P1_EBX_REG_9__SCAN_IN), .A(n14237), .ZN(
        n14238) );
  AND2_X1 U17586 ( .A1(n14239), .A2(n14238), .ZN(n14240) );
  OR2_X1 U17587 ( .A1(n14316), .A2(n14240), .ZN(n20079) );
  INV_X1 U17588 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n21252) );
  OAI22_X1 U17589 ( .A1(n20079), .A2(n14898), .B1(n21252), .B2(n14897), .ZN(
        n14241) );
  INV_X1 U17590 ( .A(n14241), .ZN(n14242) );
  OAI21_X1 U17591 ( .B1(n14408), .B2(n14908), .A(n14242), .ZN(P1_U2863) );
  OAI22_X1 U17592 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20012), .B1(n14243), 
        .B2(n16580), .ZN(n14244) );
  AOI21_X1 U17593 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16170), .A(n14244), .ZN(
        n15989) );
  INV_X1 U17594 ( .A(n15989), .ZN(n16093) );
  NOR2_X1 U17595 ( .A1(n11782), .A2(n15988), .ZN(n14248) );
  INV_X1 U17596 ( .A(n19033), .ZN(n19985) );
  INV_X1 U17597 ( .A(n14267), .ZN(n19226) );
  AOI22_X1 U17598 ( .A1(n19206), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19226), .B2(n10206), .ZN(n14397) );
  INV_X1 U17599 ( .A(n14397), .ZN(n14245) );
  OAI22_X1 U17600 ( .A1(n14246), .A2(n19985), .B1(n14396), .B2(n14245), .ZN(
        n14247) );
  OAI21_X1 U17601 ( .B1(n14248), .B2(n14247), .A(n16093), .ZN(n14249) );
  OAI21_X1 U17602 ( .B1(n16093), .B2(n14250), .A(n14249), .ZN(P2_U3601) );
  INV_X1 U17603 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14251) );
  OAI222_X1 U17604 ( .A1(n14408), .A2(n14987), .B1(n14986), .B2(n14925), .C1(
        n14251), .C2(n14983), .ZN(P1_U2895) );
  INV_X1 U17605 ( .A(n14254), .ZN(n14255) );
  INV_X1 U17606 ( .A(n14265), .ZN(n14253) );
  AOI221_X1 U17607 ( .B1(n14255), .B2(n14265), .C1(n14254), .C2(n14253), .A(
        n19895), .ZN(n14256) );
  INV_X1 U17608 ( .A(n14256), .ZN(n14264) );
  AOI22_X1 U17609 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19229), .B1(
        n19200), .B2(n20000), .ZN(n14257) );
  OAI21_X1 U17610 ( .B1(n19215), .B2(n10787), .A(n14257), .ZN(n14258) );
  AOI21_X1 U17611 ( .B1(P2_REIP_REG_2__SCAN_IN), .B2(n19199), .A(n14258), .ZN(
        n14259) );
  OAI21_X1 U17612 ( .B1(n14260), .B2(n19217), .A(n14259), .ZN(n14261) );
  AOI21_X1 U17613 ( .B1(n14262), .B2(n19223), .A(n14261), .ZN(n14263) );
  OAI211_X1 U17614 ( .C1(n19998), .C2(n19203), .A(n14264), .B(n14263), .ZN(
        P2_U2853) );
  OAI21_X1 U17615 ( .B1(n14267), .B2(n14266), .A(n14265), .ZN(n14393) );
  NOR2_X1 U17616 ( .A1(n19155), .A2(n14269), .ZN(n14268) );
  AOI21_X1 U17617 ( .B1(n14269), .B2(n19228), .A(n14268), .ZN(n14270) );
  OAI21_X1 U17618 ( .B1(n14271), .B2(n19217), .A(n14270), .ZN(n14275) );
  AOI22_X1 U17619 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19199), .B1(n19200), 
        .B2(n20003), .ZN(n14272) );
  OAI21_X1 U17620 ( .B1(n19215), .B2(n14273), .A(n14272), .ZN(n14274) );
  AOI211_X1 U17621 ( .C1(n19223), .C2(n11777), .A(n14275), .B(n14274), .ZN(
        n14277) );
  NAND2_X1 U17622 ( .A1(n19986), .A2(n19227), .ZN(n14276) );
  OAI211_X1 U17623 ( .C1(n14393), .C2(n19895), .A(n14277), .B(n14276), .ZN(
        P2_U2854) );
  INV_X1 U17624 ( .A(n14278), .ZN(n14335) );
  NOR2_X1 U17625 ( .A1(n14334), .A2(n14335), .ZN(n14333) );
  INV_X1 U17626 ( .A(n14279), .ZN(n14280) );
  OAI21_X1 U17627 ( .B1(n14333), .B2(n14281), .A(n14280), .ZN(n15494) );
  OAI21_X1 U17628 ( .B1(n14284), .B2(n14282), .A(n15416), .ZN(n19059) );
  AOI22_X1 U17629 ( .A1(n19233), .A2(BUF2_REG_20__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n14287) );
  AOI22_X1 U17630 ( .A1(n16430), .A2(n14285), .B1(n19284), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n14286) );
  OAI211_X1 U17631 ( .C1(n15552), .C2(n19059), .A(n14287), .B(n14286), .ZN(
        n14288) );
  INV_X1 U17632 ( .A(n14288), .ZN(n14289) );
  OAI21_X1 U17633 ( .B1(n15494), .B2(n19257), .A(n14289), .ZN(P2_U2899) );
  OAI21_X1 U17634 ( .B1(n14290), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14291), .ZN(n14307) );
  XOR2_X1 U17635 ( .A(n14292), .B(n14293), .Z(n14305) );
  AND2_X1 U17636 ( .A1(n14294), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14301) );
  NAND2_X1 U17637 ( .A1(n14296), .A2(n14295), .ZN(n14299) );
  INV_X1 U17638 ( .A(n19195), .ZN(n14297) );
  AOI22_X1 U17639 ( .A1(n16558), .A2(n14297), .B1(n19172), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n14298) );
  OAI211_X1 U17640 ( .C1(n19189), .C2(n15976), .A(n14299), .B(n14298), .ZN(
        n14300) );
  AOI211_X1 U17641 ( .C1(n14305), .C2(n16563), .A(n14301), .B(n14300), .ZN(
        n14302) );
  OAI21_X1 U17642 ( .B1(n15966), .B2(n14307), .A(n14302), .ZN(P2_U3040) );
  INV_X1 U17643 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19926) );
  OAI22_X1 U17644 ( .A1(n19926), .A2(n19181), .B1(n19341), .B2(n19187), .ZN(
        n14304) );
  OAI22_X1 U17645 ( .A1(n14136), .A2(n19189), .B1(n16506), .B2(n10215), .ZN(
        n14303) );
  AOI211_X1 U17646 ( .C1(n14305), .C2(n16502), .A(n14304), .B(n14303), .ZN(
        n14306) );
  OAI21_X1 U17647 ( .B1(n19332), .B2(n14307), .A(n14306), .ZN(P2_U3008) );
  OAI21_X1 U17648 ( .B1(n14232), .B2(n14309), .A(n14308), .ZN(n15142) );
  INV_X1 U17649 ( .A(n14986), .ZN(n14310) );
  AOI22_X1 U17650 ( .A1(n14310), .A2(n14921), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14965), .ZN(n14311) );
  OAI21_X1 U17651 ( .B1(n15142), .B2(n14987), .A(n14311), .ZN(P1_U2894) );
  INV_X1 U17652 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21276) );
  INV_X1 U17653 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20870) );
  INV_X1 U17654 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21228) );
  NOR4_X1 U17655 ( .A1(n20870), .A2(n21228), .A3(n13685), .A4(n20223), .ZN(
        n14838) );
  INV_X1 U17656 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21246) );
  NAND3_X1 U17657 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n14840) );
  NOR2_X1 U17658 ( .A1(n21246), .A2(n14840), .ZN(n14832) );
  NAND2_X1 U17659 ( .A1(n14838), .A2(n14832), .ZN(n20074) );
  NOR2_X1 U17660 ( .A1(n21276), .A2(n20074), .ZN(n14318) );
  NAND2_X1 U17661 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n14318), .ZN(n14776) );
  NOR2_X1 U17662 ( .A1(n14688), .A2(n14776), .ZN(n14821) );
  NOR2_X1 U17663 ( .A1(n20112), .A2(n14821), .ZN(n16247) );
  INV_X1 U17664 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n21204) );
  NAND2_X1 U17665 ( .A1(n14500), .A2(n21204), .ZN(n14314) );
  INV_X1 U17666 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16275) );
  NAND2_X1 U17667 ( .A1(n14236), .A2(n16275), .ZN(n14312) );
  OAI211_X1 U17668 ( .C1(n14630), .C2(P1_EBX_REG_10__SCAN_IN), .A(n14312), .B(
        n14517), .ZN(n14313) );
  NAND2_X1 U17669 ( .A1(n14314), .A2(n14313), .ZN(n14315) );
  OR2_X1 U17670 ( .A1(n14316), .A2(n14315), .ZN(n14317) );
  NAND2_X1 U17671 ( .A1(n14903), .A2(n14317), .ZN(n15315) );
  INV_X1 U17672 ( .A(n14318), .ZN(n14319) );
  NOR3_X1 U17673 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n20075), .A3(n14319), 
        .ZN(n14320) );
  AOI21_X1 U17674 ( .B1(n20127), .B2(P1_EBX_REG_10__SCAN_IN), .A(n14320), .ZN(
        n14321) );
  OAI21_X1 U17675 ( .B1(n20080), .B2(n15315), .A(n14321), .ZN(n14323) );
  NAND2_X1 U17676 ( .A1(n14322), .A2(n14831), .ZN(n20113) );
  INV_X1 U17677 ( .A(n20113), .ZN(n20132) );
  AOI211_X1 U17678 ( .C1(n20133), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n14323), .B(n20132), .ZN(n14324) );
  OAI21_X1 U17679 ( .B1(n20140), .B2(n15144), .A(n14324), .ZN(n14325) );
  AOI21_X1 U17680 ( .B1(n16247), .B2(P1_REIP_REG_10__SCAN_IN), .A(n14325), 
        .ZN(n14326) );
  OAI21_X1 U17681 ( .B1(n15142), .B2(n14809), .A(n14326), .ZN(P1_U2830) );
  OAI22_X1 U17682 ( .A1(n15315), .A2(n14898), .B1(n21204), .B2(n14897), .ZN(
        n14327) );
  INV_X1 U17683 ( .A(n14327), .ZN(n14328) );
  OAI21_X1 U17684 ( .B1(n15142), .B2(n14908), .A(n14328), .ZN(P1_U2862) );
  INV_X1 U17685 ( .A(n14329), .ZN(n15488) );
  NAND2_X1 U17686 ( .A1(n14330), .A2(n14331), .ZN(n14332) );
  NAND2_X1 U17687 ( .A1(n15488), .A2(n14332), .ZN(n19075) );
  AOI21_X1 U17688 ( .B1(n14335), .B2(n14334), .A(n14333), .ZN(n15556) );
  NAND2_X1 U17689 ( .A1(n15556), .A2(n15481), .ZN(n14337) );
  NAND2_X1 U17690 ( .A1(n15490), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14336) );
  OAI211_X1 U17691 ( .C1(n19075), .C2(n15490), .A(n14337), .B(n14336), .ZN(
        P2_U2868) );
  NAND2_X1 U17692 ( .A1(n14338), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14339) );
  INV_X1 U17693 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14521) );
  NAND2_X1 U17694 ( .A1(n14341), .A2(n14375), .ZN(n14345) );
  NAND2_X1 U17695 ( .A1(n14351), .A2(n14349), .ZN(n14342) );
  XNOR2_X1 U17696 ( .A(n14342), .B(n14348), .ZN(n14343) );
  NAND2_X1 U17697 ( .A1(n14343), .A2(n20930), .ZN(n14344) );
  NAND2_X1 U17698 ( .A1(n14345), .A2(n14344), .ZN(n20185) );
  NAND2_X1 U17699 ( .A1(n14347), .A2(n14375), .ZN(n14354) );
  AND2_X1 U17700 ( .A1(n14349), .A2(n14348), .ZN(n14350) );
  NAND2_X1 U17701 ( .A1(n14351), .A2(n14350), .ZN(n14358) );
  XNOR2_X1 U17702 ( .A(n14358), .B(n14359), .ZN(n14352) );
  NAND2_X1 U17703 ( .A1(n14352), .A2(n20930), .ZN(n14353) );
  NAND2_X1 U17704 ( .A1(n14354), .A2(n14353), .ZN(n14355) );
  INV_X1 U17705 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16362) );
  XNOR2_X1 U17706 ( .A(n14355), .B(n16362), .ZN(n16296) );
  NAND3_X1 U17707 ( .A1(n14356), .A2(n14357), .A3(n14375), .ZN(n14363) );
  INV_X1 U17708 ( .A(n14358), .ZN(n14360) );
  NAND2_X1 U17709 ( .A1(n14360), .A2(n14359), .ZN(n14367) );
  XNOR2_X1 U17710 ( .A(n14367), .B(n14368), .ZN(n14361) );
  NAND2_X1 U17711 ( .A1(n14361), .A2(n20930), .ZN(n14362) );
  NAND2_X1 U17712 ( .A1(n14363), .A2(n14362), .ZN(n16291) );
  OR2_X1 U17713 ( .A1(n16291), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14364) );
  NAND2_X1 U17714 ( .A1(n16291), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14365) );
  NAND2_X1 U17715 ( .A1(n14366), .A2(n14375), .ZN(n14372) );
  INV_X1 U17716 ( .A(n14367), .ZN(n14369) );
  NAND2_X1 U17717 ( .A1(n14369), .A2(n14368), .ZN(n14380) );
  XNOR2_X1 U17718 ( .A(n14380), .B(n14374), .ZN(n14370) );
  NAND2_X1 U17719 ( .A1(n14370), .A2(n20930), .ZN(n14371) );
  NAND2_X1 U17720 ( .A1(n14372), .A2(n14371), .ZN(n14373) );
  NAND2_X1 U17721 ( .A1(n14373), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16285) );
  AND3_X1 U17722 ( .A1(n14376), .A2(n14375), .A3(n14374), .ZN(n14377) );
  NAND2_X4 U17723 ( .A1(n14356), .A2(n14377), .ZN(n15140) );
  OR3_X1 U17724 ( .A1(n14380), .A2(n14379), .A3(n14378), .ZN(n14381) );
  NAND2_X1 U17725 ( .A1(n15140), .A2(n14381), .ZN(n14403) );
  XNOR2_X1 U17726 ( .A(n14403), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14382) );
  XNOR2_X1 U17727 ( .A(n14402), .B(n14382), .ZN(n16340) );
  INV_X1 U17728 ( .A(n16340), .ZN(n14387) );
  INV_X1 U17729 ( .A(n14383), .ZN(n14830) );
  AOI22_X1 U17730 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n10057), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14384) );
  OAI21_X1 U17731 ( .B1(n14833), .B2(n20193), .A(n14384), .ZN(n14385) );
  AOI21_X1 U17732 ( .B1(n14830), .B2(n20188), .A(n14385), .ZN(n14386) );
  OAI21_X1 U17733 ( .B1(n14387), .B2(n20056), .A(n14386), .ZN(P1_U2991) );
  OR2_X1 U17734 ( .A1(n14389), .A2(n14388), .ZN(n14390) );
  NAND2_X1 U17735 ( .A1(n14330), .A2(n14390), .ZN(n19087) );
  INV_X1 U17736 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n19081) );
  MUX2_X1 U17737 ( .A(n19087), .B(n19081), .S(n15490), .Z(n14391) );
  OAI21_X1 U17738 ( .B1(n14392), .B2(n15493), .A(n14391), .ZN(P2_U2869) );
  INV_X1 U17739 ( .A(n15988), .ZN(n16576) );
  OAI21_X1 U17740 ( .B1(n10206), .B2(n14394), .A(n14393), .ZN(n14395) );
  INV_X1 U17741 ( .A(n14395), .ZN(n15985) );
  NOR2_X1 U17742 ( .A1(n14397), .A2(n14396), .ZN(n15982) );
  AOI222_X1 U17743 ( .A1(n19986), .A2(n16576), .B1(n14398), .B2(n19033), .C1(
        n15985), .C2(n15982), .ZN(n14400) );
  NAND2_X1 U17744 ( .A1(n15989), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14399) );
  OAI21_X1 U17745 ( .B1(n15989), .B2(n14400), .A(n14399), .ZN(P2_U3600) );
  OR2_X1 U17746 ( .A1(n14403), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14401) );
  NAND2_X1 U17747 ( .A1(n14403), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14404) );
  INV_X1 U17748 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14406) );
  NOR2_X1 U17749 ( .A1(n15140), .A2(n14406), .ZN(n14434) );
  NAND2_X1 U17750 ( .A1(n15140), .A2(n14406), .ZN(n14436) );
  NOR2_X1 U17751 ( .A1(n14434), .A2(n10049), .ZN(n14407) );
  XNOR2_X1 U17752 ( .A(n14433), .B(n14407), .ZN(n16327) );
  INV_X1 U17753 ( .A(n14408), .ZN(n20082) );
  INV_X1 U17754 ( .A(n20085), .ZN(n14410) );
  AOI22_X1 U17755 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n10057), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14409) );
  OAI21_X1 U17756 ( .B1(n14410), .B2(n20193), .A(n14409), .ZN(n14411) );
  AOI21_X1 U17757 ( .B1(n20082), .B2(n20188), .A(n14411), .ZN(n14412) );
  OAI21_X1 U17758 ( .B1(n16327), .B2(n20056), .A(n14412), .ZN(P1_U2990) );
  INV_X1 U17759 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14422) );
  OAI21_X1 U17760 ( .B1(n18825), .B2(n18969), .A(n14422), .ZN(n14413) );
  NAND2_X1 U17761 ( .A1(n18827), .A2(n14413), .ZN(n18841) );
  NOR2_X1 U17762 ( .A1(n18967), .A2(n18841), .ZN(n14421) );
  NAND2_X1 U17763 ( .A1(n18797), .A2(n14414), .ZN(n15995) );
  AOI21_X1 U17764 ( .B1(n18848), .B2(n19014), .A(n14415), .ZN(n14416) );
  NOR2_X1 U17765 ( .A1(n14416), .A2(n19012), .ZN(n17553) );
  INV_X1 U17766 ( .A(n16176), .ZN(n14417) );
  OAI211_X1 U17767 ( .C1(n17553), .C2(n14417), .A(n16172), .B(n19015), .ZN(
        n14418) );
  NAND3_X1 U17768 ( .A1(n14419), .A2(n15995), .A3(n14418), .ZN(n18832) );
  INV_X1 U17769 ( .A(n18832), .ZN(n18846) );
  NAND2_X1 U17770 ( .A1(n18859), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18364) );
  INV_X1 U17771 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18356) );
  NAND3_X1 U17772 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18961)
         );
  OR2_X1 U17773 ( .A1(n18356), .A2(n18961), .ZN(n14420) );
  OAI211_X1 U17774 ( .C1(n18856), .C2(n18846), .A(n18364), .B(n14420), .ZN(
        n18992) );
  MUX2_X1 U17775 ( .A(n14421), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18995), .Z(P3_U3284) );
  OAI211_X1 U17776 ( .C1(n18825), .C2(n18969), .A(n17166), .B(n14422), .ZN(
        n18355) );
  NOR2_X1 U17777 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18355), .ZN(n14423) );
  OAI21_X1 U17778 ( .B1(n14423), .B2(n18961), .A(n18707), .ZN(n18362) );
  INV_X1 U17779 ( .A(n18362), .ZN(n14424) );
  NOR2_X1 U17780 ( .A1(n19008), .A2(n17993), .ZN(n16086) );
  AOI21_X1 U17781 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n16086), .ZN(n16087) );
  NOR2_X1 U17782 ( .A1(n14424), .A2(n16087), .ZN(n14426) );
  INV_X1 U17783 ( .A(n18611), .ZN(n18358) );
  NOR2_X1 U17784 ( .A1(n18963), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18411) );
  OR2_X1 U17785 ( .A1(n18411), .A2(n14424), .ZN(n16085) );
  OR2_X1 U17786 ( .A1(n18358), .A2(n16085), .ZN(n14425) );
  MUX2_X1 U17787 ( .A(n14426), .B(n14425), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  INV_X1 U17788 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16616) );
  AOI22_X1 U17789 ( .A1(n14429), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n14428), .ZN(n14430) );
  NAND3_X1 U17790 ( .A1(n14637), .A2(n12187), .A3(n14983), .ZN(n14432) );
  AOI22_X1 U17791 ( .A1(n14968), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14965), .ZN(n14431) );
  OAI211_X1 U17792 ( .C1(n14957), .C2(n16616), .A(n14432), .B(n14431), .ZN(
        P1_U2873) );
  INV_X1 U17793 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15296) );
  OR2_X1 U17794 ( .A1(n15140), .A2(n15296), .ZN(n15104) );
  NAND2_X1 U17795 ( .A1(n15140), .A2(n15296), .ZN(n14437) );
  INV_X1 U17796 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14466) );
  NAND2_X1 U17797 ( .A1(n15140), .A2(n14466), .ZN(n15119) );
  NAND2_X1 U17798 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14438) );
  NAND2_X1 U17799 ( .A1(n15140), .A2(n14438), .ZN(n15116) );
  NAND2_X1 U17800 ( .A1(n15119), .A2(n15116), .ZN(n14439) );
  INV_X1 U17801 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15283) );
  NAND2_X1 U17802 ( .A1(n15140), .A2(n15283), .ZN(n14440) );
  OR2_X1 U17803 ( .A1(n15140), .A2(n15283), .ZN(n14441) );
  INV_X1 U17804 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15272) );
  OR2_X1 U17805 ( .A1(n15140), .A2(n15272), .ZN(n16267) );
  XNOR2_X1 U17806 ( .A(n15140), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15096) );
  NAND2_X1 U17807 ( .A1(n15140), .A2(n15272), .ZN(n16266) );
  NAND2_X1 U17808 ( .A1(n15096), .A2(n16266), .ZN(n14442) );
  OAI21_X1 U17809 ( .B1(n16276), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16252), .ZN(n14448) );
  NOR2_X1 U17810 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14444) );
  OR2_X1 U17811 ( .A1(n15140), .A2(n14466), .ZN(n15118) );
  NOR2_X1 U17812 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14443) );
  OR2_X1 U17813 ( .A1(n15140), .A2(n14443), .ZN(n15114) );
  OAI21_X1 U17814 ( .B1(n14444), .B2(n15140), .A(n15103), .ZN(n14446) );
  INV_X1 U17815 ( .A(n15089), .ZN(n14450) );
  NOR2_X1 U17816 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14449) );
  INV_X1 U17817 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14452) );
  INV_X1 U17818 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14451) );
  NAND3_X1 U17819 ( .A1(n9999), .A2(n14452), .A3(n14451), .ZN(n14453) );
  XNOR2_X1 U17820 ( .A(n15140), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15088) );
  INV_X1 U17821 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15247) );
  NAND2_X1 U17822 ( .A1(n15066), .A2(n10317), .ZN(n14454) );
  INV_X1 U17823 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15212) );
  INV_X1 U17824 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15033) );
  NAND2_X1 U17825 ( .A1(n15212), .A2(n15033), .ZN(n15002) );
  OAI21_X1 U17826 ( .B1(n15031), .B2(n15002), .A(n16276), .ZN(n15022) );
  NAND3_X1 U17827 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15190) );
  INV_X1 U17828 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14546) );
  NAND2_X1 U17829 ( .A1(n15012), .A2(n15030), .ZN(n14455) );
  INV_X1 U17830 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15183) );
  INV_X1 U17831 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15006) );
  NAND2_X1 U17832 ( .A1(n15183), .A2(n15006), .ZN(n15173) );
  NOR2_X1 U17833 ( .A1(n15140), .A2(n15173), .ZN(n14456) );
  NAND2_X1 U17834 ( .A1(n14553), .A2(n14554), .ZN(n14459) );
  AND2_X1 U17835 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14547) );
  AND2_X1 U17836 ( .A1(n15140), .A2(n14547), .ZN(n14457) );
  INV_X1 U17837 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15163) );
  NAND2_X1 U17838 ( .A1(n14552), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14458) );
  AOI22_X1 U17839 ( .A1(n13597), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14630), .ZN(n14561) );
  NAND2_X1 U17840 ( .A1(n14517), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14461) );
  OAI211_X1 U17841 ( .C1(n14630), .C2(P1_EBX_REG_11__SCAN_IN), .A(n14236), .B(
        n14461), .ZN(n14463) );
  OAI21_X1 U17842 ( .B1(n14510), .B2(P1_EBX_REG_11__SCAN_IN), .A(n14463), .ZN(
        n14904) );
  INV_X1 U17843 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14464) );
  MUX2_X1 U17844 ( .A(n14465), .B(n14500), .S(n14464), .Z(n14469) );
  OAI21_X1 U17845 ( .B1(n14467), .B2(n14466), .A(n14489), .ZN(n14468) );
  NOR2_X1 U17846 ( .A1(n14469), .A2(n14468), .ZN(n14891) );
  MUX2_X1 U17847 ( .A(n14510), .B(n14517), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14471) );
  NAND2_X1 U17848 ( .A1(n14511), .A2(n15296), .ZN(n14470) );
  NAND2_X1 U17849 ( .A1(n14471), .A2(n14470), .ZN(n14817) );
  INV_X1 U17850 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n21255) );
  NAND2_X1 U17851 ( .A1(n14500), .A2(n21255), .ZN(n14474) );
  NAND2_X1 U17852 ( .A1(n14236), .A2(n15283), .ZN(n14472) );
  OAI211_X1 U17853 ( .C1(n14630), .C2(P1_EBX_REG_14__SCAN_IN), .A(n14472), .B(
        n14480), .ZN(n14473) );
  NAND2_X1 U17854 ( .A1(n14474), .A2(n14473), .ZN(n14802) );
  MUX2_X1 U17855 ( .A(n14510), .B(n14517), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n14476) );
  NAND2_X1 U17856 ( .A1(n14511), .A2(n15272), .ZN(n14475) );
  AND2_X1 U17857 ( .A1(n14476), .A2(n14475), .ZN(n14880) );
  INV_X1 U17858 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21202) );
  NAND2_X1 U17859 ( .A1(n14500), .A2(n21202), .ZN(n14479) );
  INV_X1 U17860 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16255) );
  NAND2_X1 U17861 ( .A1(n14236), .A2(n16255), .ZN(n14477) );
  OAI211_X1 U17862 ( .C1(n14630), .C2(P1_EBX_REG_16__SCAN_IN), .A(n14477), .B(
        n14517), .ZN(n14478) );
  AND2_X1 U17863 ( .A1(n14479), .A2(n14478), .ZN(n14875) );
  MUX2_X1 U17864 ( .A(n14510), .B(n14480), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14482) );
  INV_X1 U17865 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16302) );
  NAND2_X1 U17866 ( .A1(n14511), .A2(n16302), .ZN(n14481) );
  NAND2_X1 U17867 ( .A1(n14482), .A2(n14481), .ZN(n14788) );
  INV_X1 U17868 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21289) );
  NAND2_X1 U17869 ( .A1(n14500), .A2(n21289), .ZN(n14485) );
  INV_X1 U17870 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15259) );
  NAND2_X1 U17871 ( .A1(n9811), .A2(n15259), .ZN(n14483) );
  OAI211_X1 U17872 ( .C1(n14630), .C2(P1_EBX_REG_18__SCAN_IN), .A(n14483), .B(
        n14517), .ZN(n14484) );
  AND2_X1 U17873 ( .A1(n14485), .A2(n14484), .ZN(n14772) );
  NAND2_X1 U17874 ( .A1(n14517), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14486) );
  OAI211_X1 U17875 ( .C1(n14630), .C2(P1_EBX_REG_19__SCAN_IN), .A(n9811), .B(
        n14486), .ZN(n14487) );
  OAI21_X1 U17876 ( .B1(n14510), .B2(P1_EBX_REG_19__SCAN_IN), .A(n14487), .ZN(
        n14775) );
  MUX2_X1 U17877 ( .A(n14514), .B(n9811), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n14491) );
  NAND2_X1 U17878 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n14630), .ZN(
        n14488) );
  AND2_X1 U17879 ( .A1(n14489), .A2(n14488), .ZN(n14490) );
  NAND2_X1 U17880 ( .A1(n14491), .A2(n14490), .ZN(n14861) );
  MUX2_X1 U17881 ( .A(n14510), .B(n14517), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n14492) );
  OAI21_X1 U17882 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13597), .A(
        n14492), .ZN(n14854) );
  MUX2_X1 U17883 ( .A(n14514), .B(n9811), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14494) );
  NAND2_X1 U17884 ( .A1(n14630), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14493) );
  NAND2_X1 U17885 ( .A1(n14494), .A2(n14493), .ZN(n14738) );
  INV_X1 U17886 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21216) );
  NAND2_X1 U17887 ( .A1(n14504), .A2(n21216), .ZN(n14497) );
  NAND2_X1 U17888 ( .A1(n14517), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14495) );
  OAI211_X1 U17889 ( .C1(n14630), .C2(P1_EBX_REG_23__SCAN_IN), .A(n14236), .B(
        n14495), .ZN(n14496) );
  AND2_X1 U17890 ( .A1(n14497), .A2(n14496), .ZN(n14739) );
  NAND2_X1 U17891 ( .A1(n14738), .A2(n14739), .ZN(n14498) );
  INV_X1 U17892 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14499) );
  NAND2_X1 U17893 ( .A1(n14500), .A2(n14499), .ZN(n14503) );
  NAND2_X1 U17894 ( .A1(n14236), .A2(n15212), .ZN(n14501) );
  OAI211_X1 U17895 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n14630), .A(n14501), .B(
        n14517), .ZN(n14502) );
  AND2_X1 U17896 ( .A1(n14503), .A2(n14502), .ZN(n14733) );
  INV_X1 U17897 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21023) );
  NAND2_X1 U17898 ( .A1(n14504), .A2(n21023), .ZN(n14507) );
  NAND2_X1 U17899 ( .A1(n14517), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14505) );
  OAI211_X1 U17900 ( .C1(n14630), .C2(P1_EBX_REG_25__SCAN_IN), .A(n9811), .B(
        n14505), .ZN(n14506) );
  AND2_X1 U17901 ( .A1(n14507), .A2(n14506), .ZN(n14713) );
  MUX2_X1 U17902 ( .A(n14514), .B(n9811), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14509) );
  NAND2_X1 U17903 ( .A1(n14630), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14508) );
  NAND2_X1 U17904 ( .A1(n14509), .A2(n14508), .ZN(n14698) );
  MUX2_X1 U17905 ( .A(n14510), .B(n14517), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14513) );
  NAND2_X1 U17906 ( .A1(n14511), .A2(n15183), .ZN(n14512) );
  AND2_X1 U17907 ( .A1(n14513), .A2(n14512), .ZN(n14683) );
  MUX2_X1 U17908 ( .A(n14514), .B(n14236), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n14516) );
  NAND2_X1 U17909 ( .A1(n14630), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14515) );
  AND2_X1 U17910 ( .A1(n14516), .A2(n14515), .ZN(n14677) );
  OAI22_X1 U17911 ( .A1(n13597), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n14630), .ZN(n14560) );
  MUX2_X1 U17912 ( .A(P1_EBX_REG_29__SCAN_IN), .B(n14560), .S(n14517), .Z(
        n14662) );
  NOR2_X2 U17913 ( .A1(n14679), .A2(n14662), .ZN(n14661) );
  MUX2_X1 U17914 ( .A(n14517), .B(n14561), .S(n14661), .Z(n14519) );
  AOI22_X1 U17915 ( .A1(n13597), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14630), .ZN(n14518) );
  NOR2_X1 U17916 ( .A1(n14636), .A2(n20225), .ZN(n14550) );
  INV_X1 U17917 ( .A(n16338), .ZN(n15269) );
  NOR2_X1 U17918 ( .A1(n14521), .A2(n14520), .ZN(n20201) );
  NAND2_X1 U17919 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20201), .ZN(
        n14524) );
  NOR2_X1 U17920 ( .A1(n20232), .A2(n20214), .ZN(n15277) );
  INV_X1 U17921 ( .A(n15277), .ZN(n16333) );
  NOR2_X1 U17922 ( .A1(n14524), .A2(n16333), .ZN(n15316) );
  NAND3_X1 U17923 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15318) );
  NAND2_X1 U17924 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15320) );
  NOR2_X1 U17925 ( .A1(n15318), .A2(n15320), .ZN(n15303) );
  AND3_X1 U17926 ( .A1(n15316), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n15303), .ZN(n15307) );
  NAND2_X1 U17927 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15307), .ZN(
        n14541) );
  NOR2_X1 U17928 ( .A1(n15296), .A2(n14541), .ZN(n14522) );
  NOR2_X1 U17929 ( .A1(n16334), .A2(n14522), .ZN(n15257) );
  OR2_X1 U17930 ( .A1(n15257), .A2(n20212), .ZN(n15281) );
  NOR4_X1 U17931 ( .A1(n15272), .A2(n15283), .A3(n16302), .A4(n16255), .ZN(
        n15258) );
  INV_X1 U17932 ( .A(n15258), .ZN(n14542) );
  NOR2_X1 U17933 ( .A1(n15259), .A2(n14542), .ZN(n14528) );
  INV_X1 U17934 ( .A(n14524), .ZN(n15279) );
  OAI21_X1 U17935 ( .B1(n14525), .B2(n20214), .A(n20232), .ZN(n20218) );
  NAND2_X1 U17936 ( .A1(n15279), .A2(n20218), .ZN(n16336) );
  INV_X1 U17937 ( .A(n16336), .ZN(n15317) );
  AND3_X1 U17938 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15317), .A3(
        n15303), .ZN(n15254) );
  AND2_X1 U17939 ( .A1(n15254), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14540) );
  NAND3_X1 U17940 ( .A1(n14540), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n14528), .ZN(n14526) );
  NAND2_X1 U17941 ( .A1(n20221), .A2(n14526), .ZN(n14527) );
  OAI21_X1 U17942 ( .B1(n16334), .B2(n14528), .A(n14527), .ZN(n14529) );
  NOR2_X1 U17943 ( .A1(n15281), .A2(n14529), .ZN(n15248) );
  OAI21_X1 U17944 ( .B1(n14451), .B2(n15247), .A(n16338), .ZN(n14530) );
  NAND2_X1 U17945 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14544) );
  INV_X1 U17946 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15221) );
  AND2_X1 U17947 ( .A1(n20221), .A2(n15221), .ZN(n14531) );
  INV_X1 U17948 ( .A(n15190), .ZN(n14534) );
  NAND2_X1 U17949 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15187) );
  NAND2_X1 U17950 ( .A1(n14539), .A2(n15187), .ZN(n14533) );
  NAND2_X1 U17951 ( .A1(n20221), .A2(n15212), .ZN(n14532) );
  OAI211_X1 U17952 ( .C1(n14534), .C2(n15334), .A(n14533), .B(n14532), .ZN(
        n14535) );
  NAND2_X1 U17953 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14536) );
  NAND2_X1 U17954 ( .A1(n16338), .A2(n14536), .ZN(n14537) );
  OAI21_X1 U17955 ( .B1(n14547), .B2(n15269), .A(n15180), .ZN(n15159) );
  AOI211_X1 U17956 ( .C1(n15163), .C2(n16338), .A(n14554), .B(n15159), .ZN(
        n14564) );
  AOI211_X1 U17957 ( .C1(n15269), .C2(n15197), .A(n14538), .B(n14564), .ZN(
        n14549) );
  INV_X1 U17958 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21083) );
  NOR2_X1 U17959 ( .A1(n20222), .A2(n21083), .ZN(n14613) );
  NOR2_X1 U17960 ( .A1(n15334), .A2(n14541), .ZN(n15292) );
  NAND2_X1 U17961 ( .A1(n14539), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15205) );
  INV_X1 U17962 ( .A(n14540), .ZN(n15282) );
  OAI22_X1 U17963 ( .A1(n14541), .A2(n15205), .B1(n20196), .B2(n15282), .ZN(
        n15293) );
  AND2_X1 U17964 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14543) );
  NAND2_X1 U17965 ( .A1(n15260), .A2(n14543), .ZN(n15239) );
  INV_X1 U17966 ( .A(n14544), .ZN(n14545) );
  NAND2_X1 U17967 ( .A1(n15236), .A2(n14545), .ZN(n15211) );
  INV_X1 U17968 ( .A(n14547), .ZN(n15174) );
  NOR2_X1 U17969 ( .A1(n15172), .A2(n15174), .ZN(n15164) );
  NAND2_X1 U17970 ( .A1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15164), .ZN(
        n14565) );
  NOR3_X1 U17971 ( .A1(n14554), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14565), .ZN(n14548) );
  NOR4_X1 U17972 ( .A1(n14550), .A2(n14549), .A3(n14613), .A4(n14548), .ZN(
        n14551) );
  OAI21_X1 U17973 ( .B1(n14618), .B2(n16326), .A(n14551), .ZN(P1_U3000) );
  NOR2_X1 U17974 ( .A1(n14553), .A2(n14552), .ZN(n14555) );
  XNOR2_X1 U17975 ( .A(n14555), .B(n14554), .ZN(n14569) );
  NAND2_X1 U17976 ( .A1(n14650), .A2(n16270), .ZN(n14556) );
  NAND2_X1 U17977 ( .A1(n10057), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14563) );
  OAI211_X1 U17978 ( .C1(n14557), .C2(n15131), .A(n14556), .B(n14563), .ZN(
        n14558) );
  AOI21_X1 U17979 ( .B1(n14649), .B2(n20188), .A(n14558), .ZN(n14559) );
  OAI21_X1 U17980 ( .B1(n14569), .B2(n20056), .A(n14559), .ZN(P1_U2969) );
  OAI22_X1 U17981 ( .A1(n14661), .A2(n14517), .B1(n14560), .B2(n14679), .ZN(
        n14562) );
  XNOR2_X1 U17982 ( .A(n14562), .B(n14561), .ZN(n14845) );
  INV_X1 U17983 ( .A(n14563), .ZN(n14567) );
  AOI21_X1 U17984 ( .B1(n14565), .B2(n14554), .A(n14564), .ZN(n14566) );
  AOI211_X1 U17985 ( .C1(n14845), .C2(n20205), .A(n14567), .B(n14566), .ZN(
        n14568) );
  OAI21_X1 U17986 ( .B1(n14569), .B2(n16326), .A(n14568), .ZN(P1_U3001) );
  INV_X1 U17987 ( .A(n14573), .ZN(n14577) );
  NOR2_X1 U17988 ( .A1(n14574), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14576) );
  MUX2_X1 U17989 ( .A(n14577), .B(n14576), .S(n14575), .Z(n15363) );
  NAND2_X1 U17990 ( .A1(n15363), .A2(n14578), .ZN(n14579) );
  XNOR2_X1 U17991 ( .A(n14579), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14580) );
  XNOR2_X1 U17992 ( .A(n14581), .B(n14580), .ZN(n14612) );
  NAND2_X1 U17993 ( .A1(n15578), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14582) );
  NAND2_X1 U17994 ( .A1(n14605), .A2(n16566), .ZN(n14604) );
  OAI21_X1 U17995 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15944), .A(
        n14583), .ZN(n14602) );
  AOI22_X1 U17996 ( .A1(n11383), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14587) );
  NAND2_X1 U17997 ( .A1(n14585), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14586) );
  OAI211_X1 U17998 ( .C1(n9960), .C2(n14588), .A(n14587), .B(n14586), .ZN(
        n14589) );
  INV_X1 U17999 ( .A(n14589), .ZN(n14590) );
  AOI222_X1 U18000 ( .A1(n9948), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n14593), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11538), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14594) );
  INV_X1 U18001 ( .A(n14594), .ZN(n14595) );
  NOR4_X1 U18002 ( .A1(n15770), .A2(n15744), .A3(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A4(n14597), .ZN(n14598) );
  INV_X1 U18003 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n15361) );
  NOR2_X1 U18004 ( .A1(n19181), .A2(n15361), .ZN(n14606) );
  OAI21_X1 U18005 ( .B1(n15366), .B2(n15976), .A(n14600), .ZN(n14601) );
  OAI211_X1 U18006 ( .C1(n14612), .C2(n16552), .A(n14604), .B(n14603), .ZN(
        P2_U3015) );
  NAND2_X1 U18007 ( .A1(n14605), .A2(n16503), .ZN(n14611) );
  AOI21_X1 U18008 ( .B1(n19329), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14606), .ZN(n14607) );
  OAI21_X1 U18009 ( .B1(n19341), .B2(n14608), .A(n14607), .ZN(n14609) );
  AOI21_X1 U18010 ( .B1(n15425), .B2(n19337), .A(n14609), .ZN(n14610) );
  OAI211_X1 U18011 ( .C1(n14612), .C2(n19333), .A(n14611), .B(n14610), .ZN(
        P2_U2983) );
  AOI21_X1 U18012 ( .B1(n20182), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14613), .ZN(n14614) );
  OAI21_X1 U18013 ( .B1(n14615), .B2(n20193), .A(n14614), .ZN(n14616) );
  OAI21_X1 U18014 ( .B1(n14618), .B2(n20056), .A(n14617), .ZN(P1_U2968) );
  NOR2_X1 U18015 ( .A1(n15379), .A2(n15490), .ZN(n14619) );
  AOI21_X1 U18016 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15490), .A(n14619), .ZN(
        n14620) );
  MUX2_X1 U18017 ( .A(n14623), .B(n14622), .S(n14625), .Z(n14628) );
  AOI22_X1 U18018 ( .A1(n14626), .A2(n14625), .B1(n9934), .B2(n14624), .ZN(
        n14627) );
  NAND2_X1 U18019 ( .A1(n14628), .A2(n14627), .ZN(n14629) );
  NAND2_X1 U18020 ( .A1(n14629), .A2(n13015), .ZN(n16134) );
  INV_X1 U18021 ( .A(n16134), .ZN(n14635) );
  NAND3_X1 U18022 ( .A1(n14631), .A2(n14630), .A3(n16165), .ZN(n14632) );
  NAND2_X1 U18023 ( .A1(n14632), .A2(n20936), .ZN(n20928) );
  AND2_X1 U18024 ( .A1(n14633), .A2(n20928), .ZN(n16133) );
  NOR2_X1 U18025 ( .A1(n16133), .A2(n14634), .ZN(n20058) );
  MUX2_X1 U18026 ( .A(P1_MORE_REG_SCAN_IN), .B(n14635), .S(n20058), .Z(
        P1_U3484) );
  NAND2_X1 U18027 ( .A1(n14637), .A2(n20106), .ZN(n14648) );
  AND2_X1 U18028 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14641) );
  INV_X1 U18029 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20893) );
  INV_X1 U18030 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n16196) );
  AND4_X1 U18031 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .A4(P1_REIP_REG_12__SCAN_IN), .ZN(n14799) );
  NAND4_X1 U18032 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14799), .A3(
        P1_REIP_REG_15__SCAN_IN), .A4(P1_REIP_REG_16__SCAN_IN), .ZN(n16204) );
  INV_X1 U18033 ( .A(n16204), .ZN(n14780) );
  NAND3_X1 U18034 ( .A1(n14780), .A2(P1_REIP_REG_18__SCAN_IN), .A3(
        P1_REIP_REG_19__SCAN_IN), .ZN(n16197) );
  NOR3_X1 U18035 ( .A1(n16196), .A2(n14776), .A3(n16197), .ZN(n16181) );
  NAND2_X1 U18036 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n16181), .ZN(n14758) );
  NOR2_X1 U18037 ( .A1(n20893), .A2(n14758), .ZN(n14745) );
  NAND2_X1 U18038 ( .A1(n14745), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14717) );
  NAND3_X1 U18039 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .A3(P1_REIP_REG_26__SCAN_IN), .ZN(n14638) );
  OR2_X1 U18040 ( .A1(n14717), .A2(n14638), .ZN(n14687) );
  NAND2_X1 U18041 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14639) );
  NOR2_X1 U18042 ( .A1(n14687), .A2(n14639), .ZN(n14640) );
  NOR2_X1 U18043 ( .A1(n20075), .A2(n14640), .ZN(n14673) );
  NOR2_X1 U18044 ( .A1(n14673), .A2(n14688), .ZN(n14676) );
  OAI21_X1 U18045 ( .B1(n14641), .B2(n20075), .A(n14676), .ZN(n14651) );
  NAND2_X1 U18046 ( .A1(n14839), .A2(n14640), .ZN(n14664) );
  INV_X1 U18047 ( .A(n14641), .ZN(n14642) );
  NOR3_X1 U18048 ( .A1(n14664), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14642), 
        .ZN(n14646) );
  INV_X1 U18049 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14644) );
  OAI22_X1 U18050 ( .A1(n20104), .A2(n14644), .B1(n14643), .B2(n20115), .ZN(
        n14645) );
  AOI211_X1 U18051 ( .C1(n14651), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14646), 
        .B(n14645), .ZN(n14647) );
  OAI211_X1 U18052 ( .C1(n14636), .C2(n20080), .A(n14648), .B(n14647), .ZN(
        P1_U2809) );
  INV_X1 U18053 ( .A(n14650), .ZN(n14655) );
  AOI22_X1 U18054 ( .A1(n20127), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20133), .ZN(n14654) );
  INV_X1 U18055 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21249) );
  NOR2_X1 U18056 ( .A1(n14664), .A2(n21249), .ZN(n14652) );
  OAI21_X1 U18057 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14652), .A(n14651), 
        .ZN(n14653) );
  OAI211_X1 U18058 ( .C1(n20140), .C2(n14655), .A(n14654), .B(n14653), .ZN(
        n14656) );
  AOI21_X1 U18059 ( .B1(n14845), .B2(n20126), .A(n14656), .ZN(n14657) );
  OAI21_X1 U18060 ( .B1(n14847), .B2(n14809), .A(n14657), .ZN(P1_U2810) );
  AOI21_X1 U18061 ( .B1(n14660), .B2(n14658), .A(n14659), .ZN(n14994) );
  INV_X1 U18062 ( .A(n14994), .ZN(n14913) );
  AOI21_X1 U18063 ( .B1(n14662), .B2(n14679), .A(n14661), .ZN(n14848) );
  INV_X1 U18064 ( .A(n14676), .ZN(n14666) );
  AOI22_X1 U18065 ( .A1(n20127), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20133), .ZN(n14663) );
  OAI21_X1 U18066 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n14664), .A(n14663), 
        .ZN(n14665) );
  AOI21_X1 U18067 ( .B1(n14666), .B2(P1_REIP_REG_29__SCAN_IN), .A(n14665), 
        .ZN(n14667) );
  OAI21_X1 U18068 ( .B1(n20140), .B2(n14992), .A(n14667), .ZN(n14668) );
  AOI21_X1 U18069 ( .B1(n14848), .B2(n20126), .A(n14668), .ZN(n14669) );
  OAI21_X1 U18070 ( .B1(n14913), .B2(n14809), .A(n14669), .ZN(P1_U2811) );
  OAI21_X1 U18071 ( .B1(n14671), .B2(n14672), .A(n14658), .ZN(n15009) );
  INV_X1 U18072 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14996) );
  AOI22_X1 U18073 ( .A1(n20127), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20133), .ZN(n14675) );
  INV_X1 U18074 ( .A(n14687), .ZN(n14689) );
  NAND3_X1 U18075 ( .A1(n14673), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14689), 
        .ZN(n14674) );
  OAI211_X1 U18076 ( .C1(n14676), .C2(n14996), .A(n14675), .B(n14674), .ZN(
        n14681) );
  NAND2_X1 U18077 ( .A1(n9963), .A2(n14677), .ZN(n14678) );
  NAND2_X1 U18078 ( .A1(n14679), .A2(n14678), .ZN(n15168) );
  NOR2_X1 U18079 ( .A1(n15168), .A2(n20080), .ZN(n14680) );
  AOI211_X1 U18080 ( .C1(n20084), .C2(n14999), .A(n14681), .B(n14680), .ZN(
        n14682) );
  OAI21_X1 U18081 ( .B1(n15009), .B2(n14809), .A(n14682), .ZN(P1_U2812) );
  OR2_X1 U18082 ( .A1(n14700), .A2(n14683), .ZN(n14684) );
  NAND2_X1 U18083 ( .A1(n9963), .A2(n14684), .ZN(n15178) );
  AOI21_X1 U18084 ( .B1(n14686), .B2(n14685), .A(n14671), .ZN(n15019) );
  NAND2_X1 U18085 ( .A1(n15019), .A2(n20106), .ZN(n14696) );
  INV_X1 U18086 ( .A(n15017), .ZN(n14694) );
  OAI21_X1 U18087 ( .B1(n14688), .B2(n14687), .A(n14719), .ZN(n14705) );
  INV_X1 U18088 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14692) );
  AOI22_X1 U18089 ( .A1(n20127), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20133), .ZN(n14691) );
  NAND3_X1 U18090 ( .A1(n14839), .A2(n14689), .A3(n14692), .ZN(n14690) );
  OAI211_X1 U18091 ( .C1(n14705), .C2(n14692), .A(n14691), .B(n14690), .ZN(
        n14693) );
  AOI21_X1 U18092 ( .B1(n20084), .B2(n14694), .A(n14693), .ZN(n14695) );
  OAI211_X1 U18093 ( .C1(n20080), .C2(n15178), .A(n14696), .B(n14695), .ZN(
        P1_U2813) );
  NOR2_X1 U18094 ( .A1(n14697), .A2(n14698), .ZN(n14699) );
  OR2_X1 U18095 ( .A1(n14700), .A2(n14699), .ZN(n15189) );
  INV_X1 U18096 ( .A(n14685), .ZN(n14702) );
  AOI21_X1 U18097 ( .B1(n14703), .B2(n14701), .A(n14702), .ZN(n15028) );
  NAND2_X1 U18098 ( .A1(n15028), .A2(n20106), .ZN(n14709) );
  INV_X1 U18099 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21232) );
  NOR3_X1 U18100 ( .A1(n20075), .A2(n21232), .A3(n14717), .ZN(n14716) );
  AOI21_X1 U18101 ( .B1(n14716), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_26__SCAN_IN), .ZN(n14706) );
  AOI22_X1 U18102 ( .A1(n20127), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20133), .ZN(n14704) );
  OAI21_X1 U18103 ( .B1(n14706), .B2(n14705), .A(n14704), .ZN(n14707) );
  AOI21_X1 U18104 ( .B1(n20084), .B2(n15024), .A(n14707), .ZN(n14708) );
  OAI211_X1 U18105 ( .C1(n20080), .C2(n15189), .A(n14709), .B(n14708), .ZN(
        P1_U2814) );
  OAI21_X1 U18106 ( .B1(n14710), .B2(n14711), .A(n14701), .ZN(n15039) );
  INV_X1 U18107 ( .A(n14697), .ZN(n14712) );
  OAI21_X1 U18108 ( .B1(n14713), .B2(n14735), .A(n14712), .ZN(n15198) );
  INV_X1 U18109 ( .A(n15198), .ZN(n14724) );
  INV_X1 U18110 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21128) );
  OAI22_X1 U18111 ( .A1(n20104), .A2(n21023), .B1(n14714), .B2(n20115), .ZN(
        n14715) );
  AOI21_X1 U18112 ( .B1(n14716), .B2(n21128), .A(n14715), .ZN(n14722) );
  INV_X1 U18113 ( .A(n14717), .ZN(n14729) );
  NAND2_X1 U18114 ( .A1(n14831), .A2(n14729), .ZN(n14718) );
  NAND2_X1 U18115 ( .A1(n14719), .A2(n14718), .ZN(n14750) );
  OAI21_X1 U18116 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n20075), .A(n14750), 
        .ZN(n14720) );
  NAND2_X1 U18117 ( .A1(n14720), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14721) );
  OAI211_X1 U18118 ( .C1(n20140), .C2(n15035), .A(n14722), .B(n14721), .ZN(
        n14723) );
  AOI21_X1 U18119 ( .B1(n14724), .B2(n20126), .A(n14723), .ZN(n14725) );
  OAI21_X1 U18120 ( .B1(n15039), .B2(n14809), .A(n14725), .ZN(P1_U2815) );
  INV_X1 U18121 ( .A(n14710), .ZN(n14727) );
  OAI21_X1 U18122 ( .B1(n14728), .B2(n14726), .A(n14727), .ZN(n15045) );
  AOI22_X1 U18123 ( .A1(n20127), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20133), .ZN(n14731) );
  NAND3_X1 U18124 ( .A1(n14839), .A2(n14729), .A3(n21232), .ZN(n14730) );
  OAI211_X1 U18125 ( .C1(n14750), .C2(n21232), .A(n14731), .B(n14730), .ZN(
        n14732) );
  AOI21_X1 U18126 ( .B1(n20084), .B2(n15048), .A(n14732), .ZN(n14737) );
  AND2_X1 U18127 ( .A1(n14741), .A2(n14733), .ZN(n14734) );
  NOR2_X1 U18128 ( .A1(n14735), .A2(n14734), .ZN(n15210) );
  NAND2_X1 U18129 ( .A1(n15210), .A2(n20126), .ZN(n14736) );
  OAI211_X1 U18130 ( .C1(n15045), .C2(n14809), .A(n14737), .B(n14736), .ZN(
        P1_U2816) );
  INV_X1 U18131 ( .A(n14738), .ZN(n14759) );
  INV_X1 U18132 ( .A(n14739), .ZN(n14740) );
  OAI21_X1 U18133 ( .B1(n14856), .B2(n14759), .A(n14740), .ZN(n14742) );
  NAND2_X1 U18134 ( .A1(n14742), .A2(n14741), .ZN(n15219) );
  AOI21_X1 U18135 ( .B1(n14744), .B2(n14743), .A(n14726), .ZN(n15055) );
  NAND2_X1 U18136 ( .A1(n15055), .A2(n20106), .ZN(n14754) );
  INV_X1 U18137 ( .A(n15053), .ZN(n14752) );
  AOI21_X1 U18138 ( .B1(n14839), .B2(n14745), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14749) );
  OAI22_X1 U18139 ( .A1(n20104), .A2(n21216), .B1(n14746), .B2(n20115), .ZN(
        n14747) );
  INV_X1 U18140 ( .A(n14747), .ZN(n14748) );
  OAI21_X1 U18141 ( .B1(n14750), .B2(n14749), .A(n14748), .ZN(n14751) );
  AOI21_X1 U18142 ( .B1(n20084), .B2(n14752), .A(n14751), .ZN(n14753) );
  OAI211_X1 U18143 ( .C1(n20080), .C2(n15219), .A(n14754), .B(n14753), .ZN(
        P1_U2817) );
  AOI21_X1 U18144 ( .B1(n14757), .B2(n14756), .A(n12784), .ZN(n15060) );
  NOR3_X1 U18145 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n20075), .A3(n14758), 
        .ZN(n14765) );
  XNOR2_X1 U18146 ( .A(n14856), .B(n14759), .ZN(n15227) );
  OAI21_X1 U18147 ( .B1(n20075), .B2(n16181), .A(n14831), .ZN(n16198) );
  NOR2_X1 U18148 ( .A1(n20075), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16182) );
  OAI21_X1 U18149 ( .B1(n16198), .B2(n16182), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14763) );
  AOI22_X1 U18150 ( .A1(n20084), .A2(n15063), .B1(n20127), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n14760) );
  OAI21_X1 U18151 ( .B1(n15061), .B2(n20115), .A(n14760), .ZN(n14761) );
  INV_X1 U18152 ( .A(n14761), .ZN(n14762) );
  OAI211_X1 U18153 ( .C1(n15227), .C2(n20080), .A(n14763), .B(n14762), .ZN(
        n14764) );
  AOI211_X1 U18154 ( .C1(n15060), .C2(n20106), .A(n14765), .B(n14764), .ZN(
        n14766) );
  INV_X1 U18155 ( .A(n14766), .ZN(P1_U2818) );
  NOR2_X1 U18156 ( .A1(n14874), .A2(n14767), .ZN(n14859) );
  NOR2_X1 U18157 ( .A1(n14874), .A2(n14768), .ZN(n14770) );
  NOR2_X1 U18158 ( .A1(n14770), .A2(n14769), .ZN(n14771) );
  INV_X1 U18159 ( .A(n14772), .ZN(n14867) );
  NAND2_X1 U18160 ( .A1(n14868), .A2(n14867), .ZN(n14774) );
  AOI21_X1 U18161 ( .B1(n14775), .B2(n14774), .A(n14773), .ZN(n15250) );
  INV_X1 U18162 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n16205) );
  INV_X1 U18163 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21219) );
  NOR2_X1 U18164 ( .A1(n16205), .A2(n21219), .ZN(n14779) );
  INV_X1 U18165 ( .A(n14776), .ZN(n14777) );
  OAI211_X1 U18166 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(P1_REIP_REG_19__SCAN_IN), .A(n14780), .B(n16242), .ZN(n14778) );
  OAI22_X1 U18167 ( .A1(n14779), .A2(n14778), .B1(n15084), .B2(n20140), .ZN(
        n14784) );
  INV_X1 U18168 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14782) );
  AOI21_X1 U18169 ( .B1(n14780), .B2(n14821), .A(n20112), .ZN(n16208) );
  AOI22_X1 U18170 ( .A1(n16208), .A2(P1_REIP_REG_19__SCAN_IN), .B1(n20127), 
        .B2(P1_EBX_REG_19__SCAN_IN), .ZN(n14781) );
  OAI211_X1 U18171 ( .C1(n20115), .C2(n14782), .A(n14781), .B(n20113), .ZN(
        n14783) );
  AOI211_X1 U18172 ( .C1(n20126), .C2(n15250), .A(n14784), .B(n14783), .ZN(
        n14785) );
  OAI21_X1 U18173 ( .B1(n15082), .B2(n14809), .A(n14785), .ZN(P1_U2821) );
  INV_X1 U18174 ( .A(n14865), .ZN(n14786) );
  AOI21_X1 U18175 ( .B1(n14787), .B2(n14874), .A(n14786), .ZN(n16260) );
  INV_X1 U18176 ( .A(n16260), .ZN(n14964) );
  INV_X1 U18177 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n21283) );
  AOI21_X1 U18178 ( .B1(n14788), .B2(n14877), .A(n14868), .ZN(n16305) );
  NAND2_X1 U18179 ( .A1(n16305), .A2(n20126), .ZN(n14790) );
  AOI21_X1 U18180 ( .B1(n20133), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n20132), .ZN(n14789) );
  OAI211_X1 U18181 ( .C1(n21283), .C2(n20104), .A(n14790), .B(n14789), .ZN(
        n14791) );
  AOI21_X1 U18182 ( .B1(n20084), .B2(n16259), .A(n14791), .ZN(n14795) );
  NAND2_X1 U18183 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14792) );
  INV_X1 U18184 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20882) );
  NAND2_X1 U18185 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n14820) );
  NOR3_X1 U18186 ( .A1(n20882), .A2(n14820), .A3(n16246), .ZN(n14800) );
  NAND2_X1 U18187 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n14800), .ZN(n16224) );
  INV_X1 U18188 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21073) );
  OAI21_X1 U18189 ( .B1(n14792), .B2(n16224), .A(n21073), .ZN(n14793) );
  NAND2_X1 U18190 ( .A1(n14793), .A2(n16208), .ZN(n14794) );
  OAI211_X1 U18191 ( .C1(n14964), .C2(n14809), .A(n14795), .B(n14794), .ZN(
        P1_U2823) );
  INV_X1 U18192 ( .A(n14796), .ZN(n14798) );
  INV_X1 U18193 ( .A(n14815), .ZN(n14797) );
  AOI21_X1 U18194 ( .B1(n14798), .B2(n14797), .A(n14884), .ZN(n15112) );
  INV_X1 U18195 ( .A(n15112), .ZN(n14976) );
  AOI21_X1 U18196 ( .B1(n14799), .B2(n14821), .A(n20112), .ZN(n16228) );
  OAI21_X1 U18197 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n14800), .A(n16228), 
        .ZN(n14808) );
  INV_X1 U18198 ( .A(n15110), .ZN(n14806) );
  NOR2_X1 U18199 ( .A1(n14819), .A2(n14802), .ZN(n14803) );
  OR2_X1 U18200 ( .A1(n14801), .A2(n14803), .ZN(n15286) );
  AOI22_X1 U18201 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20133), .B1(
        n20127), .B2(P1_EBX_REG_14__SCAN_IN), .ZN(n14804) );
  OAI211_X1 U18202 ( .C1(n15286), .C2(n20080), .A(n14804), .B(n20113), .ZN(
        n14805) );
  AOI21_X1 U18203 ( .B1(n20084), .B2(n14806), .A(n14805), .ZN(n14807) );
  OAI211_X1 U18204 ( .C1(n14976), .C2(n14809), .A(n14808), .B(n14807), .ZN(
        P1_U2826) );
  NAND2_X1 U18205 ( .A1(n14308), .A2(n14810), .ZN(n14811) );
  NAND2_X1 U18206 ( .A1(n14812), .A2(n14811), .ZN(n14899) );
  OR2_X1 U18207 ( .A1(n14899), .A2(n14900), .ZN(n14813) );
  NAND2_X1 U18208 ( .A1(n14813), .A2(n14812), .ZN(n14896) );
  NAND2_X1 U18209 ( .A1(n14896), .A2(n14895), .ZN(n14894) );
  INV_X1 U18210 ( .A(n14814), .ZN(n14816) );
  AOI21_X1 U18211 ( .B1(n14894), .B2(n14816), .A(n14815), .ZN(n15125) );
  NOR3_X1 U18212 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14820), .A3(n16246), 
        .ZN(n14828) );
  AND2_X1 U18213 ( .A1(n14893), .A2(n14817), .ZN(n14818) );
  NOR2_X1 U18214 ( .A1(n14819), .A2(n14818), .ZN(n15299) );
  INV_X1 U18215 ( .A(n14820), .ZN(n14822) );
  AOI21_X1 U18216 ( .B1(n14822), .B2(n14821), .A(n20112), .ZN(n16241) );
  AOI22_X1 U18217 ( .A1(n20127), .A2(P1_EBX_REG_13__SCAN_IN), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n16241), .ZN(n14823) );
  OAI211_X1 U18218 ( .C1(n20115), .C2(n14824), .A(n14823), .B(n20113), .ZN(
        n14825) );
  AOI21_X1 U18219 ( .B1(n15299), .B2(n20126), .A(n14825), .ZN(n14826) );
  OAI21_X1 U18220 ( .B1(n20140), .B2(n15123), .A(n14826), .ZN(n14827) );
  AOI211_X1 U18221 ( .C1(n15125), .C2(n20106), .A(n14828), .B(n14827), .ZN(
        n14829) );
  INV_X1 U18222 ( .A(n14829), .ZN(P1_U2827) );
  NAND2_X1 U18223 ( .A1(n14830), .A2(n20106), .ZN(n14844) );
  AND2_X1 U18224 ( .A1(n14831), .A2(n14838), .ZN(n20111) );
  AOI21_X1 U18225 ( .B1(n14832), .B2(n20111), .A(n20112), .ZN(n20083) );
  AOI22_X1 U18226 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20133), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20083), .ZN(n14843) );
  INV_X1 U18227 ( .A(n14833), .ZN(n14837) );
  NAND2_X1 U18228 ( .A1(n16341), .A2(n20126), .ZN(n14834) );
  OAI211_X1 U18229 ( .C1(n20104), .C2(n14835), .A(n14834), .B(n20113), .ZN(
        n14836) );
  AOI21_X1 U18230 ( .B1(n20084), .B2(n14837), .A(n14836), .ZN(n14842) );
  NAND2_X1 U18231 ( .A1(n14839), .A2(n14838), .ZN(n20120) );
  OR3_X1 U18232 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14840), .A3(n20120), .ZN(
        n14841) );
  NAND4_X1 U18233 ( .A1(n14844), .A2(n14843), .A3(n14842), .A4(n14841), .ZN(
        P1_U2832) );
  OAI22_X1 U18234 ( .A1(n14636), .A2(n14898), .B1(n14644), .B2(n14897), .ZN(
        P1_U2841) );
  AOI22_X1 U18235 ( .A1(n14845), .A2(n14906), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n14905), .ZN(n14846) );
  OAI21_X1 U18236 ( .B1(n14847), .B2(n14908), .A(n14846), .ZN(P1_U2842) );
  INV_X1 U18237 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n21260) );
  INV_X1 U18238 ( .A(n14848), .ZN(n15161) );
  OAI222_X1 U18239 ( .A1(n21260), .A2(n14897), .B1(n14898), .B2(n15161), .C1(
        n14913), .C2(n14908), .ZN(P1_U2843) );
  INV_X1 U18240 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n21294) );
  OAI222_X1 U18241 ( .A1(n21294), .A2(n14897), .B1(n14898), .B2(n15168), .C1(
        n15009), .C2(n14908), .ZN(P1_U2844) );
  INV_X1 U18242 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14849) );
  INV_X1 U18243 ( .A(n15019), .ZN(n14920) );
  OAI222_X1 U18244 ( .A1(n14849), .A2(n14897), .B1(n14898), .B2(n15178), .C1(
        n14920), .C2(n14908), .ZN(P1_U2845) );
  INV_X1 U18245 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21038) );
  INV_X1 U18246 ( .A(n15028), .ZN(n14924) );
  OAI222_X1 U18247 ( .A1(n21038), .A2(n14897), .B1(n14898), .B2(n15189), .C1(
        n14924), .C2(n14908), .ZN(P1_U2846) );
  OAI222_X1 U18248 ( .A1(n21023), .A2(n14897), .B1(n14898), .B2(n15198), .C1(
        n15039), .C2(n14908), .ZN(P1_U2847) );
  AOI22_X1 U18249 ( .A1(n15210), .A2(n14906), .B1(n14905), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n14850) );
  OAI21_X1 U18250 ( .B1(n15045), .B2(n14908), .A(n14850), .ZN(P1_U2848) );
  INV_X1 U18251 ( .A(n15055), .ZN(n14940) );
  OAI222_X1 U18252 ( .A1(n21216), .A2(n14897), .B1(n14898), .B2(n15219), .C1(
        n14940), .C2(n14908), .ZN(P1_U2849) );
  INV_X1 U18253 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14851) );
  INV_X1 U18254 ( .A(n15060), .ZN(n14943) );
  OAI222_X1 U18255 ( .A1(n14851), .A2(n14897), .B1(n14898), .B2(n15227), .C1(
        n14908), .C2(n14943), .ZN(P1_U2850) );
  OAI21_X1 U18256 ( .B1(n14852), .B2(n14853), .A(n14756), .ZN(n15070) );
  INV_X1 U18257 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14857) );
  NAND2_X1 U18258 ( .A1(n14863), .A2(n14854), .ZN(n14855) );
  NAND2_X1 U18259 ( .A1(n14856), .A2(n14855), .ZN(n16186) );
  OAI222_X1 U18260 ( .A1(n14908), .A2(n15070), .B1(n14897), .B2(n14857), .C1(
        n16186), .C2(n14898), .ZN(P1_U2851) );
  INV_X1 U18261 ( .A(n14852), .ZN(n14858) );
  OAI21_X1 U18262 ( .B1(n14860), .B2(n14859), .A(n14858), .ZN(n16195) );
  INV_X1 U18263 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n21215) );
  OR2_X1 U18264 ( .A1(n14773), .A2(n14861), .ZN(n14862) );
  NAND2_X1 U18265 ( .A1(n14863), .A2(n14862), .ZN(n16203) );
  OAI222_X1 U18266 ( .A1(n14908), .A2(n16195), .B1(n14897), .B2(n21215), .C1(
        n16203), .C2(n14898), .ZN(P1_U2852) );
  AOI22_X1 U18267 ( .A1(n15250), .A2(n14906), .B1(n14905), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n14864) );
  OAI21_X1 U18268 ( .B1(n15082), .B2(n14908), .A(n14864), .ZN(P1_U2853) );
  XOR2_X1 U18269 ( .A(n14866), .B(n14865), .Z(n16211) );
  INV_X1 U18270 ( .A(n16211), .ZN(n14961) );
  XNOR2_X1 U18271 ( .A(n14868), .B(n14867), .ZN(n16209) );
  OAI22_X1 U18272 ( .A1(n16209), .A2(n14898), .B1(n21289), .B2(n14897), .ZN(
        n14869) );
  INV_X1 U18273 ( .A(n14869), .ZN(n14870) );
  OAI21_X1 U18274 ( .B1(n14961), .B2(n14908), .A(n14870), .ZN(P1_U2854) );
  AOI22_X1 U18275 ( .A1(n16305), .A2(n14906), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14905), .ZN(n14871) );
  OAI21_X1 U18276 ( .B1(n14964), .B2(n14908), .A(n14871), .ZN(P1_U2855) );
  NAND2_X1 U18277 ( .A1(n14886), .A2(n14872), .ZN(n14873) );
  NAND2_X1 U18278 ( .A1(n14874), .A2(n14873), .ZN(n16216) );
  NAND2_X1 U18279 ( .A1(n14882), .A2(n14875), .ZN(n14876) );
  NAND2_X1 U18280 ( .A1(n14877), .A2(n14876), .ZN(n16227) );
  OAI22_X1 U18281 ( .A1(n16227), .A2(n14898), .B1(n21202), .B2(n14897), .ZN(
        n14878) );
  INV_X1 U18282 ( .A(n14878), .ZN(n14879) );
  OAI21_X1 U18283 ( .B1(n16216), .B2(n14908), .A(n14879), .ZN(P1_U2856) );
  OR2_X1 U18284 ( .A1(n14801), .A2(n14880), .ZN(n14881) );
  NAND2_X1 U18285 ( .A1(n14882), .A2(n14881), .ZN(n16311) );
  INV_X1 U18286 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14887) );
  OR2_X1 U18287 ( .A1(n14884), .A2(n14883), .ZN(n14885) );
  AND2_X1 U18288 ( .A1(n14886), .A2(n14885), .ZN(n16272) );
  INV_X1 U18289 ( .A(n16272), .ZN(n14973) );
  OAI222_X1 U18290 ( .A1(n16311), .A2(n14898), .B1(n14897), .B2(n14887), .C1(
        n14908), .C2(n14973), .ZN(P1_U2857) );
  OAI22_X1 U18291 ( .A1(n15286), .A2(n14898), .B1(n21255), .B2(n14897), .ZN(
        n14888) );
  INV_X1 U18292 ( .A(n14888), .ZN(n14889) );
  OAI21_X1 U18293 ( .B1(n14976), .B2(n14908), .A(n14889), .ZN(P1_U2858) );
  INV_X1 U18294 ( .A(n15125), .ZN(n14979) );
  AOI22_X1 U18295 ( .A1(n15299), .A2(n14906), .B1(n14905), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14890) );
  OAI21_X1 U18296 ( .B1(n14979), .B2(n14908), .A(n14890), .ZN(P1_U2859) );
  NAND2_X1 U18297 ( .A1(n14901), .A2(n14891), .ZN(n14892) );
  NAND2_X1 U18298 ( .A1(n14893), .A2(n14892), .ZN(n16236) );
  OAI222_X1 U18299 ( .A1(n16236), .A2(n14898), .B1(n14897), .B2(n14464), .C1(
        n14908), .C2(n16238), .ZN(P1_U2860) );
  XOR2_X1 U18300 ( .A(n14900), .B(n14899), .Z(n16280) );
  INV_X1 U18301 ( .A(n16280), .ZN(n14988) );
  INV_X1 U18302 ( .A(n14901), .ZN(n14902) );
  AOI21_X1 U18303 ( .B1(n14904), .B2(n14903), .A(n14902), .ZN(n16318) );
  AOI22_X1 U18304 ( .A1(n16318), .A2(n14906), .B1(n14905), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n14907) );
  OAI21_X1 U18305 ( .B1(n14988), .B2(n14908), .A(n14907), .ZN(P1_U2861) );
  INV_X1 U18306 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16620) );
  NOR2_X1 U18307 ( .A1(n14957), .A2(n16620), .ZN(n14911) );
  INV_X1 U18308 ( .A(DATAI_29_), .ZN(n14909) );
  OAI22_X1 U18309 ( .A1(n14951), .A2(n14909), .B1(n14978), .B2(n14948), .ZN(
        n14910) );
  AOI211_X1 U18310 ( .C1(n14965), .C2(P1_EAX_REG_29__SCAN_IN), .A(n14911), .B(
        n14910), .ZN(n14912) );
  OAI21_X1 U18311 ( .B1(n14913), .B2(n14987), .A(n14912), .ZN(P1_U2875) );
  AOI22_X1 U18312 ( .A1(n14966), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14965), .ZN(n14915) );
  AOI22_X1 U18313 ( .A1(n14968), .A2(DATAI_28_), .B1(n14967), .B2(n14980), 
        .ZN(n14914) );
  OAI211_X1 U18314 ( .C1(n15009), .C2(n14987), .A(n14915), .B(n14914), .ZN(
        P1_U2876) );
  INV_X1 U18315 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19366) );
  NOR2_X1 U18316 ( .A1(n14957), .A2(n19366), .ZN(n14918) );
  INV_X1 U18317 ( .A(DATAI_27_), .ZN(n14916) );
  OAI22_X1 U18318 ( .A1(n14951), .A2(n14916), .B1(n14985), .B2(n14948), .ZN(
        n14917) );
  AOI211_X1 U18319 ( .C1(n14965), .C2(P1_EAX_REG_27__SCAN_IN), .A(n14918), .B(
        n14917), .ZN(n14919) );
  OAI21_X1 U18320 ( .B1(n14920), .B2(n14987), .A(n14919), .ZN(P1_U2877) );
  AOI22_X1 U18321 ( .A1(n14966), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14965), .ZN(n14923) );
  AOI22_X1 U18322 ( .A1(n14968), .A2(DATAI_26_), .B1(n14967), .B2(n14921), 
        .ZN(n14922) );
  OAI211_X1 U18323 ( .C1(n14924), .C2(n14987), .A(n14923), .B(n14922), .ZN(
        P1_U2878) );
  INV_X1 U18324 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16626) );
  NOR2_X1 U18325 ( .A1(n14957), .A2(n16626), .ZN(n14928) );
  INV_X1 U18326 ( .A(DATAI_25_), .ZN(n14926) );
  OAI22_X1 U18327 ( .A1(n14951), .A2(n14926), .B1(n14925), .B2(n14948), .ZN(
        n14927) );
  AOI211_X1 U18328 ( .C1(n14965), .C2(P1_EAX_REG_25__SCAN_IN), .A(n14928), .B(
        n14927), .ZN(n14929) );
  OAI21_X1 U18329 ( .B1(n15039), .B2(n14987), .A(n14929), .ZN(P1_U2879) );
  NOR2_X1 U18330 ( .A1(n14983), .A2(n14930), .ZN(n14934) );
  INV_X1 U18331 ( .A(DATAI_24_), .ZN(n14932) );
  OAI22_X1 U18332 ( .A1(n14951), .A2(n14932), .B1(n14948), .B2(n14931), .ZN(
        n14933) );
  AOI211_X1 U18333 ( .C1(BUF1_REG_24__SCAN_IN), .C2(n14966), .A(n14934), .B(
        n14933), .ZN(n14935) );
  OAI21_X1 U18334 ( .B1(n15045), .B2(n14987), .A(n14935), .ZN(P1_U2880) );
  INV_X1 U18335 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20286) );
  OAI22_X1 U18336 ( .A1(n14957), .A2(n20286), .B1(n14936), .B2(n14983), .ZN(
        n14937) );
  INV_X1 U18337 ( .A(n14937), .ZN(n14939) );
  AOI22_X1 U18338 ( .A1(n14968), .A2(DATAI_23_), .B1(n14967), .B2(n20291), 
        .ZN(n14938) );
  OAI211_X1 U18339 ( .C1(n14940), .C2(n14987), .A(n14939), .B(n14938), .ZN(
        P1_U2881) );
  AOI22_X1 U18340 ( .A1(n14966), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14965), .ZN(n14942) );
  AOI22_X1 U18341 ( .A1(n14968), .A2(DATAI_22_), .B1(n14967), .B2(n20281), 
        .ZN(n14941) );
  OAI211_X1 U18342 ( .C1(n14943), .C2(n14987), .A(n14942), .B(n14941), .ZN(
        P1_U2882) );
  INV_X1 U18343 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n19380) );
  OAI22_X1 U18344 ( .A1(n14957), .A2(n19380), .B1(n21044), .B2(n14983), .ZN(
        n14944) );
  INV_X1 U18345 ( .A(n14944), .ZN(n14946) );
  AOI22_X1 U18346 ( .A1(n14968), .A2(DATAI_21_), .B1(n14967), .B2(n20277), 
        .ZN(n14945) );
  OAI211_X1 U18347 ( .C1(n15070), .C2(n14987), .A(n14946), .B(n14945), .ZN(
        P1_U2883) );
  NOR2_X1 U18348 ( .A1(n14983), .A2(n14947), .ZN(n14953) );
  INV_X1 U18349 ( .A(DATAI_20_), .ZN(n14950) );
  OAI22_X1 U18350 ( .A1(n14951), .A2(n14950), .B1(n14949), .B2(n14948), .ZN(
        n14952) );
  AOI211_X1 U18351 ( .C1(BUF1_REG_20__SCAN_IN), .C2(n14966), .A(n14953), .B(
        n14952), .ZN(n14954) );
  OAI21_X1 U18352 ( .B1(n16195), .B2(n14987), .A(n14954), .ZN(P1_U2884) );
  AOI22_X1 U18353 ( .A1(n14966), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14965), .ZN(n14956) );
  AOI22_X1 U18354 ( .A1(n14968), .A2(DATAI_19_), .B1(n14967), .B2(n20269), 
        .ZN(n14955) );
  OAI211_X1 U18355 ( .C1(n15082), .C2(n14987), .A(n14956), .B(n14955), .ZN(
        P1_U2885) );
  INV_X1 U18356 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20262) );
  OAI22_X1 U18357 ( .A1(n14957), .A2(n20262), .B1(n13645), .B2(n14983), .ZN(
        n14958) );
  INV_X1 U18358 ( .A(n14958), .ZN(n14960) );
  AOI22_X1 U18359 ( .A1(n14968), .A2(DATAI_18_), .B1(n14967), .B2(n20264), 
        .ZN(n14959) );
  OAI211_X1 U18360 ( .C1(n14961), .C2(n14987), .A(n14960), .B(n14959), .ZN(
        P1_U2886) );
  AOI22_X1 U18361 ( .A1(n14966), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14965), .ZN(n14963) );
  AOI22_X1 U18362 ( .A1(n14968), .A2(DATAI_17_), .B1(n14967), .B2(n20259), 
        .ZN(n14962) );
  OAI211_X1 U18363 ( .C1(n14964), .C2(n14987), .A(n14963), .B(n14962), .ZN(
        P1_U2887) );
  AOI22_X1 U18364 ( .A1(n14966), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14965), .ZN(n14970) );
  AOI22_X1 U18365 ( .A1(n14968), .A2(DATAI_16_), .B1(n14967), .B2(n20250), 
        .ZN(n14969) );
  OAI211_X1 U18366 ( .C1(n16216), .C2(n14987), .A(n14970), .B(n14969), .ZN(
        P1_U2888) );
  OAI222_X1 U18367 ( .A1(n14973), .A2(n14987), .B1(n14986), .B2(n14972), .C1(
        n14983), .C2(n14971), .ZN(P1_U2889) );
  OAI222_X1 U18368 ( .A1(n14976), .A2(n14987), .B1(n14986), .B2(n14975), .C1(
        n14974), .C2(n14983), .ZN(P1_U2890) );
  OAI222_X1 U18369 ( .A1(n14979), .A2(n14987), .B1(n14986), .B2(n14978), .C1(
        n14977), .C2(n14983), .ZN(P1_U2891) );
  INV_X1 U18370 ( .A(n14980), .ZN(n14982) );
  OAI222_X1 U18371 ( .A1(n16238), .A2(n14987), .B1(n14986), .B2(n14982), .C1(
        n14981), .C2(n14983), .ZN(P1_U2892) );
  INV_X1 U18372 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14984) );
  OAI222_X1 U18373 ( .A1(n14988), .A2(n14987), .B1(n14986), .B2(n14985), .C1(
        n14984), .C2(n14983), .ZN(P1_U2893) );
  XNOR2_X1 U18374 ( .A(n14990), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15166) );
  NOR2_X1 U18375 ( .A1(n20222), .A2(n21249), .ZN(n15158) );
  AOI21_X1 U18376 ( .B1(n20182), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15158), .ZN(n14991) );
  OAI21_X1 U18377 ( .B1(n14992), .B2(n20193), .A(n14991), .ZN(n14993) );
  AOI21_X1 U18378 ( .B1(n14994), .B2(n20188), .A(n14993), .ZN(n14995) );
  OAI21_X1 U18379 ( .B1(n15166), .B2(n20056), .A(n14995), .ZN(P1_U2970) );
  NOR2_X1 U18380 ( .A1(n20222), .A2(n14996), .ZN(n15170) );
  NOR2_X1 U18381 ( .A1(n15131), .A2(n14997), .ZN(n14998) );
  AOI211_X1 U18382 ( .C1(n14999), .C2(n16270), .A(n15170), .B(n14998), .ZN(
        n15008) );
  NAND2_X1 U18383 ( .A1(n15140), .A2(n15190), .ZN(n15000) );
  NAND2_X1 U18384 ( .A1(n15051), .A2(n15000), .ZN(n15004) );
  NAND2_X1 U18385 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15001) );
  NOR2_X1 U18386 ( .A1(n15004), .A2(n15001), .ZN(n15005) );
  NOR4_X1 U18387 ( .A1(n15002), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15003) );
  OAI211_X1 U18388 ( .C1(n15009), .C2(n15135), .A(n15008), .B(n15007), .ZN(
        P1_U2971) );
  INV_X1 U18389 ( .A(n9936), .ZN(n15011) );
  NAND2_X1 U18390 ( .A1(n15012), .A2(n15011), .ZN(n15013) );
  MUX2_X1 U18391 ( .A(n15014), .B(n15013), .S(n15140), .Z(n15015) );
  XNOR2_X1 U18392 ( .A(n15015), .B(n15183), .ZN(n15186) );
  NAND2_X1 U18393 ( .A1(n10057), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15179) );
  NAND2_X1 U18394 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15016) );
  OAI211_X1 U18395 ( .C1(n15017), .C2(n20193), .A(n15179), .B(n15016), .ZN(
        n15018) );
  AOI21_X1 U18396 ( .B1(n15019), .B2(n20188), .A(n15018), .ZN(n15020) );
  OAI21_X1 U18397 ( .B1(n20056), .B2(n15186), .A(n15020), .ZN(P1_U2972) );
  INV_X1 U18398 ( .A(n15051), .ZN(n15040) );
  OAI21_X1 U18399 ( .B1(n15040), .B2(n15190), .A(n15140), .ZN(n15021) );
  NAND2_X1 U18400 ( .A1(n15022), .A2(n15021), .ZN(n15023) );
  XOR2_X1 U18401 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15023), .Z(
        n15195) );
  INV_X1 U18402 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15026) );
  NAND2_X1 U18403 ( .A1(n15024), .A2(n16270), .ZN(n15025) );
  NAND2_X1 U18404 ( .A1(n10057), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15188) );
  OAI211_X1 U18405 ( .C1(n15131), .C2(n15026), .A(n15025), .B(n15188), .ZN(
        n15027) );
  AOI21_X1 U18406 ( .B1(n15028), .B2(n20188), .A(n15027), .ZN(n15029) );
  OAI21_X1 U18407 ( .B1(n20056), .B2(n15195), .A(n15029), .ZN(P1_U2973) );
  NAND2_X1 U18408 ( .A1(n15030), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15042) );
  MUX2_X1 U18409 ( .A(n15212), .B(n15031), .S(n16276), .Z(n15032) );
  AOI21_X1 U18410 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15042), .A(
        n15032), .ZN(n15034) );
  XNOR2_X1 U18411 ( .A(n15034), .B(n15033), .ZN(n15196) );
  NAND2_X1 U18412 ( .A1(n15196), .A2(n20189), .ZN(n15038) );
  NOR2_X1 U18413 ( .A1(n20222), .A2(n21128), .ZN(n15200) );
  NOR2_X1 U18414 ( .A1(n15035), .A2(n20193), .ZN(n15036) );
  AOI211_X1 U18415 ( .C1(n20182), .C2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15200), .B(n15036), .ZN(n15037) );
  OAI211_X1 U18416 ( .C1(n15135), .C2(n15039), .A(n15038), .B(n15037), .ZN(
        P1_U2974) );
  NAND2_X1 U18417 ( .A1(n15040), .A2(n15042), .ZN(n15041) );
  MUX2_X1 U18418 ( .A(n15042), .B(n15041), .S(n16276), .Z(n15043) );
  XNOR2_X1 U18419 ( .A(n15043), .B(n15212), .ZN(n15215) );
  NAND2_X1 U18420 ( .A1(n10057), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15207) );
  OAI21_X1 U18421 ( .B1(n15131), .B2(n15044), .A(n15207), .ZN(n15047) );
  NOR2_X1 U18422 ( .A1(n15045), .A2(n15135), .ZN(n15046) );
  AOI211_X1 U18423 ( .C1(n16270), .C2(n15048), .A(n15047), .B(n15046), .ZN(
        n15049) );
  OAI21_X1 U18424 ( .B1(n20056), .B2(n15215), .A(n15049), .ZN(P1_U2975) );
  XNOR2_X1 U18425 ( .A(n15140), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15050) );
  XNOR2_X1 U18426 ( .A(n9935), .B(n15050), .ZN(n15224) );
  NAND2_X1 U18427 ( .A1(n10057), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15218) );
  NAND2_X1 U18428 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15052) );
  OAI211_X1 U18429 ( .C1(n15053), .C2(n20193), .A(n15218), .B(n15052), .ZN(
        n15054) );
  AOI21_X1 U18430 ( .B1(n15055), .B2(n20188), .A(n15054), .ZN(n15056) );
  OAI21_X1 U18431 ( .B1(n15224), .B2(n20056), .A(n15056), .ZN(P1_U2976) );
  NAND2_X1 U18432 ( .A1(n15058), .A2(n15057), .ZN(n15059) );
  XOR2_X1 U18433 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15059), .Z(
        n15231) );
  NAND2_X1 U18434 ( .A1(n15060), .A2(n20188), .ZN(n15065) );
  NOR2_X1 U18435 ( .A1(n20222), .A2(n20893), .ZN(n15225) );
  NOR2_X1 U18436 ( .A1(n15131), .A2(n15061), .ZN(n15062) );
  AOI211_X1 U18437 ( .C1(n15063), .C2(n16270), .A(n15225), .B(n15062), .ZN(
        n15064) );
  OAI211_X1 U18438 ( .C1(n15231), .C2(n20056), .A(n15065), .B(n15064), .ZN(
        P1_U2977) );
  INV_X1 U18439 ( .A(n15066), .ZN(n15067) );
  NOR2_X1 U18440 ( .A1(n15067), .A2(n16276), .ZN(n15068) );
  AOI21_X1 U18441 ( .B1(n9999), .B2(n16276), .A(n15068), .ZN(n15075) );
  NOR2_X1 U18442 ( .A1(n15075), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15074) );
  AOI22_X1 U18443 ( .A1(n15074), .A2(n16276), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n15068), .ZN(n15069) );
  XOR2_X1 U18444 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n15069), .Z(
        n15238) );
  INV_X1 U18445 ( .A(n15070), .ZN(n16188) );
  NAND2_X1 U18446 ( .A1(n10057), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15234) );
  NAND2_X1 U18447 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15071) );
  OAI211_X1 U18448 ( .C1(n16191), .C2(n20193), .A(n15234), .B(n15071), .ZN(
        n15072) );
  AOI21_X1 U18449 ( .B1(n16188), .B2(n20188), .A(n15072), .ZN(n15073) );
  OAI21_X1 U18450 ( .B1(n15238), .B2(n20056), .A(n15073), .ZN(P1_U2978) );
  AOI21_X1 U18451 ( .B1(n15075), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15074), .ZN(n15245) );
  NAND2_X1 U18452 ( .A1(n10057), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15240) );
  OAI21_X1 U18453 ( .B1(n15131), .B2(n16192), .A(n15240), .ZN(n15077) );
  NOR2_X1 U18454 ( .A1(n16195), .A2(n15135), .ZN(n15076) );
  AOI211_X1 U18455 ( .C1(n16270), .C2(n16194), .A(n15077), .B(n15076), .ZN(
        n15078) );
  OAI21_X1 U18456 ( .B1(n15245), .B2(n20056), .A(n15078), .ZN(P1_U2979) );
  NAND2_X1 U18457 ( .A1(n15079), .A2(n15259), .ZN(n15080) );
  MUX2_X1 U18458 ( .A(n15079), .B(n15080), .S(n16276), .Z(n15081) );
  XOR2_X1 U18459 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n15081), .Z(
        n15253) );
  INV_X1 U18460 ( .A(n15082), .ZN(n15086) );
  NAND2_X1 U18461 ( .A1(n10057), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15246) );
  NAND2_X1 U18462 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15083) );
  OAI211_X1 U18463 ( .C1(n15084), .C2(n20193), .A(n15246), .B(n15083), .ZN(
        n15085) );
  AOI21_X1 U18464 ( .B1(n15086), .B2(n20188), .A(n15085), .ZN(n15087) );
  OAI21_X1 U18465 ( .B1(n15253), .B2(n20056), .A(n15087), .ZN(P1_U2980) );
  OAI21_X1 U18466 ( .B1(n15089), .B2(n15088), .A(n15079), .ZN(n15265) );
  NAND2_X1 U18467 ( .A1(n16207), .A2(n16270), .ZN(n15090) );
  NAND2_X1 U18468 ( .A1(n10057), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15261) );
  OAI211_X1 U18469 ( .C1(n15131), .C2(n15091), .A(n15090), .B(n15261), .ZN(
        n15092) );
  AOI21_X1 U18470 ( .B1(n16211), .B2(n20188), .A(n15092), .ZN(n15093) );
  OAI21_X1 U18471 ( .B1(n20056), .B2(n15265), .A(n15093), .ZN(P1_U2981) );
  OAI21_X1 U18472 ( .B1(n15094), .B2(n15095), .A(n15103), .ZN(n16265) );
  OAI21_X1 U18473 ( .B1(n16265), .B2(n16253), .A(n16266), .ZN(n15097) );
  XNOR2_X1 U18474 ( .A(n15097), .B(n15096), .ZN(n15266) );
  NAND2_X1 U18475 ( .A1(n15266), .A2(n20189), .ZN(n15102) );
  INV_X1 U18476 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15098) );
  NOR2_X1 U18477 ( .A1(n20222), .A2(n15098), .ZN(n15270) );
  INV_X1 U18478 ( .A(n16217), .ZN(n15099) );
  NOR2_X1 U18479 ( .A1(n15099), .A2(n20193), .ZN(n15100) );
  AOI211_X1 U18480 ( .C1(n20182), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15270), .B(n15100), .ZN(n15101) );
  OAI211_X1 U18481 ( .C1(n15135), .C2(n16216), .A(n15102), .B(n15101), .ZN(
        P1_U2983) );
  NAND2_X1 U18482 ( .A1(n15094), .A2(n15103), .ZN(n16254) );
  INV_X1 U18483 ( .A(n15104), .ZN(n15105) );
  AOI21_X1 U18484 ( .B1(n16254), .B2(n15106), .A(n15105), .ZN(n15108) );
  XNOR2_X1 U18485 ( .A(n15140), .B(n15283), .ZN(n15107) );
  XNOR2_X1 U18486 ( .A(n15108), .B(n15107), .ZN(n15291) );
  NAND2_X1 U18487 ( .A1(n10057), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15285) );
  NAND2_X1 U18488 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15109) );
  OAI211_X1 U18489 ( .C1(n20193), .C2(n15110), .A(n15285), .B(n15109), .ZN(
        n15111) );
  AOI21_X1 U18490 ( .B1(n15112), .B2(n20188), .A(n15111), .ZN(n15113) );
  OAI21_X1 U18491 ( .B1(n15291), .B2(n20056), .A(n15113), .ZN(P1_U2985) );
  INV_X1 U18492 ( .A(n15094), .ZN(n15117) );
  INV_X1 U18493 ( .A(n15114), .ZN(n15115) );
  AOI21_X1 U18494 ( .B1(n15117), .B2(n15116), .A(n15115), .ZN(n15129) );
  AND2_X1 U18495 ( .A1(n15118), .A2(n15119), .ZN(n15128) );
  NAND2_X1 U18496 ( .A1(n15129), .A2(n15128), .ZN(n15127) );
  NAND2_X1 U18497 ( .A1(n15127), .A2(n15119), .ZN(n15121) );
  XNOR2_X1 U18498 ( .A(n15121), .B(n15120), .ZN(n15301) );
  NAND2_X1 U18499 ( .A1(n10057), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15295) );
  NAND2_X1 U18500 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15122) );
  OAI211_X1 U18501 ( .C1(n20193), .C2(n15123), .A(n15295), .B(n15122), .ZN(
        n15124) );
  AOI21_X1 U18502 ( .B1(n15125), .B2(n20188), .A(n15124), .ZN(n15126) );
  OAI21_X1 U18503 ( .B1(n15301), .B2(n20056), .A(n15126), .ZN(P1_U2986) );
  OAI21_X1 U18504 ( .B1(n15129), .B2(n15128), .A(n15127), .ZN(n15302) );
  NAND2_X1 U18505 ( .A1(n15302), .A2(n20189), .ZN(n15134) );
  INV_X1 U18506 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15130) );
  NAND2_X1 U18507 ( .A1(n10057), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15308) );
  OAI21_X1 U18508 ( .B1(n15131), .B2(n15130), .A(n15308), .ZN(n15132) );
  AOI21_X1 U18509 ( .B1(n16270), .B2(n16240), .A(n15132), .ZN(n15133) );
  OAI211_X1 U18510 ( .C1(n15135), .C2(n16238), .A(n15134), .B(n15133), .ZN(
        P1_U2987) );
  INV_X1 U18511 ( .A(n15136), .ZN(n15137) );
  NOR2_X1 U18512 ( .A1(n15137), .A2(n16275), .ZN(n15139) );
  XNOR2_X1 U18513 ( .A(n15094), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15138) );
  MUX2_X1 U18514 ( .A(n15139), .B(n15138), .S(n15140), .Z(n15141) );
  NOR3_X1 U18515 ( .A1(n15136), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15140), .ZN(n16277) );
  NOR2_X1 U18516 ( .A1(n15141), .A2(n16277), .ZN(n15326) );
  INV_X1 U18517 ( .A(n15142), .ZN(n15146) );
  AND2_X1 U18518 ( .A1(n10057), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15323) );
  AOI21_X1 U18519 ( .B1(n20182), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15323), .ZN(n15143) );
  OAI21_X1 U18520 ( .B1(n15144), .B2(n20193), .A(n15143), .ZN(n15145) );
  AOI21_X1 U18521 ( .B1(n15146), .B2(n20188), .A(n15145), .ZN(n15147) );
  OAI21_X1 U18522 ( .B1(n15326), .B2(n20056), .A(n15147), .ZN(P1_U2989) );
  INV_X1 U18523 ( .A(n15148), .ZN(n15149) );
  NAND2_X1 U18524 ( .A1(n15149), .A2(n20188), .ZN(n15157) );
  AOI22_X1 U18525 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n10057), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n15156) );
  OR2_X1 U18526 ( .A1(n15151), .A2(n15150), .ZN(n20216) );
  NAND3_X1 U18527 ( .A1(n20216), .A2(n15152), .A3(n20189), .ZN(n15155) );
  OR2_X1 U18528 ( .A1(n20193), .A2(n15153), .ZN(n15154) );
  NAND4_X1 U18529 ( .A1(n15157), .A2(n15156), .A3(n15155), .A4(n15154), .ZN(
        P1_U2997) );
  AOI21_X1 U18530 ( .B1(n15159), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15158), .ZN(n15160) );
  OAI21_X1 U18531 ( .B1(n15161), .B2(n20225), .A(n15160), .ZN(n15162) );
  AOI21_X1 U18532 ( .B1(n15164), .B2(n15163), .A(n15162), .ZN(n15165) );
  OAI21_X1 U18533 ( .B1(n15166), .B2(n16326), .A(n15165), .ZN(P1_U3002) );
  INV_X1 U18534 ( .A(n15167), .ZN(n15177) );
  INV_X1 U18535 ( .A(n15180), .ZN(n15171) );
  NOR2_X1 U18536 ( .A1(n15168), .A2(n20225), .ZN(n15169) );
  AOI211_X1 U18537 ( .C1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15171), .A(
        n15170), .B(n15169), .ZN(n15176) );
  INV_X1 U18538 ( .A(n15172), .ZN(n15184) );
  NAND3_X1 U18539 ( .A1(n15184), .A2(n15174), .A3(n15173), .ZN(n15175) );
  OAI211_X1 U18540 ( .C1(n15177), .C2(n16326), .A(n15176), .B(n15175), .ZN(
        P1_U3003) );
  NOR2_X1 U18541 ( .A1(n15178), .A2(n20225), .ZN(n15182) );
  OAI21_X1 U18542 ( .B1(n15180), .B2(n15183), .A(n15179), .ZN(n15181) );
  AOI211_X1 U18543 ( .C1(n15184), .C2(n15183), .A(n15182), .B(n15181), .ZN(
        n15185) );
  OAI21_X1 U18544 ( .B1(n15186), .B2(n16326), .A(n15185), .ZN(P1_U3004) );
  OR3_X1 U18545 ( .A1(n15211), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15187), .ZN(n15202) );
  NAND2_X1 U18546 ( .A1(n15202), .A2(n15197), .ZN(n15193) );
  OAI21_X1 U18547 ( .B1(n15189), .B2(n20225), .A(n15188), .ZN(n15192) );
  NOR3_X1 U18548 ( .A1(n15211), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15190), .ZN(n15191) );
  AOI211_X1 U18549 ( .C1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n15193), .A(
        n15192), .B(n15191), .ZN(n15194) );
  OAI21_X1 U18550 ( .B1(n15195), .B2(n16326), .A(n15194), .ZN(P1_U3005) );
  INV_X1 U18551 ( .A(n15196), .ZN(n15204) );
  INV_X1 U18552 ( .A(n15197), .ZN(n15201) );
  NOR2_X1 U18553 ( .A1(n15198), .A2(n20225), .ZN(n15199) );
  AOI211_X1 U18554 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15201), .A(
        n15200), .B(n15199), .ZN(n15203) );
  OAI211_X1 U18555 ( .C1(n15204), .C2(n16326), .A(n15203), .B(n15202), .ZN(
        P1_U3006) );
  NAND2_X1 U18556 ( .A1(n15205), .A2(n15334), .ZN(n20211) );
  AOI21_X1 U18557 ( .B1(n15221), .B2(n20211), .A(n15206), .ZN(n15208) );
  OAI21_X1 U18558 ( .B1(n15208), .B2(n15212), .A(n15207), .ZN(n15209) );
  AOI21_X1 U18559 ( .B1(n15210), .B2(n20205), .A(n15209), .ZN(n15214) );
  INV_X1 U18560 ( .A(n15211), .ZN(n15222) );
  NAND3_X1 U18561 ( .A1(n15222), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15212), .ZN(n15213) );
  OAI211_X1 U18562 ( .C1(n15215), .C2(n16326), .A(n15214), .B(n15213), .ZN(
        P1_U3007) );
  NAND2_X1 U18563 ( .A1(n15216), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15217) );
  OAI211_X1 U18564 ( .C1(n15219), .C2(n20225), .A(n15218), .B(n15217), .ZN(
        n15220) );
  AOI21_X1 U18565 ( .B1(n15222), .B2(n15221), .A(n15220), .ZN(n15223) );
  OAI21_X1 U18566 ( .B1(n15224), .B2(n16326), .A(n15223), .ZN(P1_U3008) );
  XNOR2_X1 U18567 ( .A(n14452), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15229) );
  AOI21_X1 U18568 ( .B1(n15232), .B2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15225), .ZN(n15226) );
  OAI21_X1 U18569 ( .B1(n15227), .B2(n20225), .A(n15226), .ZN(n15228) );
  AOI21_X1 U18570 ( .B1(n15236), .B2(n15229), .A(n15228), .ZN(n15230) );
  OAI21_X1 U18571 ( .B1(n15231), .B2(n16326), .A(n15230), .ZN(P1_U3009) );
  NAND2_X1 U18572 ( .A1(n15232), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15233) );
  OAI211_X1 U18573 ( .C1(n16186), .C2(n20225), .A(n15234), .B(n15233), .ZN(
        n15235) );
  AOI21_X1 U18574 ( .B1(n15236), .B2(n14452), .A(n15235), .ZN(n15237) );
  OAI21_X1 U18575 ( .B1(n15238), .B2(n16326), .A(n15237), .ZN(P1_U3010) );
  INV_X1 U18576 ( .A(n15239), .ZN(n15243) );
  OAI21_X1 U18577 ( .B1(n16203), .B2(n20225), .A(n15240), .ZN(n15242) );
  NAND3_X1 U18578 ( .A1(n15260), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15247), .ZN(n15251) );
  AOI21_X1 U18579 ( .B1(n15251), .B2(n15248), .A(n14451), .ZN(n15241) );
  AOI211_X1 U18580 ( .C1(n15243), .C2(n14451), .A(n15242), .B(n15241), .ZN(
        n15244) );
  OAI21_X1 U18581 ( .B1(n15245), .B2(n16326), .A(n15244), .ZN(P1_U3011) );
  OAI21_X1 U18582 ( .B1(n15248), .B2(n15247), .A(n15246), .ZN(n15249) );
  AOI21_X1 U18583 ( .B1(n15250), .B2(n20205), .A(n15249), .ZN(n15252) );
  OAI211_X1 U18584 ( .C1(n15253), .C2(n16326), .A(n15252), .B(n15251), .ZN(
        P1_U3012) );
  NAND2_X1 U18585 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15280) );
  INV_X1 U18586 ( .A(n15254), .ZN(n15255) );
  AND2_X1 U18587 ( .A1(n20221), .A2(n15255), .ZN(n15256) );
  OR2_X1 U18588 ( .A1(n15256), .A2(n20212), .ZN(n15306) );
  AOI211_X1 U18589 ( .C1(n20221), .C2(n15280), .A(n15257), .B(n15306), .ZN(
        n15268) );
  OAI21_X1 U18590 ( .B1(n15269), .B2(n15258), .A(n15268), .ZN(n16307) );
  NAND2_X1 U18591 ( .A1(n15260), .A2(n15259), .ZN(n15262) );
  OAI211_X1 U18592 ( .C1(n16209), .C2(n20225), .A(n15262), .B(n15261), .ZN(
        n15263) );
  AOI21_X1 U18593 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n16307), .A(
        n15263), .ZN(n15264) );
  OAI21_X1 U18594 ( .B1(n15265), .B2(n16326), .A(n15264), .ZN(P1_U3013) );
  INV_X1 U18595 ( .A(n15266), .ZN(n15276) );
  NOR2_X1 U18596 ( .A1(n15283), .A2(n16303), .ZN(n16314) );
  NAND2_X1 U18597 ( .A1(n16314), .A2(n15272), .ZN(n15267) );
  OAI211_X1 U18598 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n15269), .A(
        n15268), .B(n15267), .ZN(n16313) );
  INV_X1 U18599 ( .A(n15270), .ZN(n15271) );
  OAI21_X1 U18600 ( .B1(n16227), .B2(n20225), .A(n15271), .ZN(n15274) );
  NOR4_X1 U18601 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15283), .A3(
        n15272), .A4(n16303), .ZN(n15273) );
  AOI211_X1 U18602 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16313), .A(
        n15274), .B(n15273), .ZN(n15275) );
  OAI21_X1 U18603 ( .B1(n15276), .B2(n16326), .A(n15275), .ZN(P1_U3015) );
  INV_X1 U18604 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16339) );
  NAND2_X1 U18605 ( .A1(n20211), .A2(n15277), .ZN(n16337) );
  NAND2_X1 U18606 ( .A1(n20221), .A2(n20218), .ZN(n15278) );
  NAND2_X1 U18607 ( .A1(n16337), .A2(n15278), .ZN(n20202) );
  NAND2_X1 U18608 ( .A1(n15279), .A2(n20202), .ZN(n16356) );
  NOR2_X1 U18609 ( .A1(n16339), .A2(n16356), .ZN(n16346) );
  NAND3_X1 U18610 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n16346), .ZN(n16325) );
  NOR2_X1 U18611 ( .A1(n16325), .A2(n15320), .ZN(n16319) );
  NAND2_X1 U18612 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16319), .ZN(
        n15310) );
  NOR3_X1 U18613 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15280), .A3(
        n15310), .ZN(n15289) );
  AOI21_X1 U18614 ( .B1(n20221), .B2(n15282), .A(n15281), .ZN(n15297) );
  NAND2_X1 U18615 ( .A1(n15296), .A2(n15293), .ZN(n15284) );
  AOI21_X1 U18616 ( .B1(n15297), .B2(n15284), .A(n15283), .ZN(n15288) );
  OAI21_X1 U18617 ( .B1(n15286), .B2(n20225), .A(n15285), .ZN(n15287) );
  NOR3_X1 U18618 ( .A1(n15289), .A2(n15288), .A3(n15287), .ZN(n15290) );
  OAI21_X1 U18619 ( .B1(n15291), .B2(n16326), .A(n15290), .ZN(P1_U3017) );
  OAI21_X1 U18620 ( .B1(n15293), .B2(n15292), .A(n15296), .ZN(n15294) );
  OAI211_X1 U18621 ( .C1(n15297), .C2(n15296), .A(n15295), .B(n15294), .ZN(
        n15298) );
  AOI21_X1 U18622 ( .B1(n15299), .B2(n20205), .A(n15298), .ZN(n15300) );
  OAI21_X1 U18623 ( .B1(n15301), .B2(n16326), .A(n15300), .ZN(P1_U3018) );
  NAND2_X1 U18624 ( .A1(n15302), .A2(n20215), .ZN(n15314) );
  AND2_X1 U18625 ( .A1(n15316), .A2(n15303), .ZN(n15304) );
  NOR2_X1 U18626 ( .A1(n16334), .A2(n15304), .ZN(n15305) );
  NOR2_X1 U18627 ( .A1(n15306), .A2(n15305), .ZN(n16324) );
  INV_X1 U18628 ( .A(n16324), .ZN(n15312) );
  INV_X1 U18629 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16323) );
  NAND3_X1 U18630 ( .A1(n20211), .A2(n15307), .A3(n16323), .ZN(n15309) );
  OAI211_X1 U18631 ( .C1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15310), .A(
        n15309), .B(n15308), .ZN(n15311) );
  AOI21_X1 U18632 ( .B1(n15312), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15311), .ZN(n15313) );
  OAI211_X1 U18633 ( .C1(n20225), .C2(n16236), .A(n15314), .B(n15313), .ZN(
        P1_U3019) );
  INV_X1 U18634 ( .A(n15315), .ZN(n15324) );
  AOI21_X1 U18635 ( .B1(n15317), .B2(n16334), .A(n15316), .ZN(n15319) );
  AOI221_X1 U18636 ( .B1(n15319), .B2(n16338), .C1(n15318), .C2(n16338), .A(
        n20212), .ZN(n16332) );
  OAI21_X1 U18637 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15320), .ZN(n15321) );
  OAI22_X1 U18638 ( .A1(n16332), .A2(n16275), .B1(n16325), .B2(n15321), .ZN(
        n15322) );
  AOI211_X1 U18639 ( .C1(n20205), .C2(n15324), .A(n15323), .B(n15322), .ZN(
        n15325) );
  OAI21_X1 U18640 ( .B1(n15326), .B2(n16326), .A(n15325), .ZN(P1_U3021) );
  NAND3_X1 U18641 ( .A1(n15327), .A2(n9937), .A3(n20215), .ZN(n15338) );
  INV_X1 U18642 ( .A(n15328), .ZN(n15332) );
  AOI21_X1 U18643 ( .B1(n15330), .B2(n15329), .A(n20214), .ZN(n15331) );
  AOI211_X1 U18644 ( .C1(n20205), .C2(n15333), .A(n15332), .B(n15331), .ZN(
        n15337) );
  INV_X1 U18645 ( .A(n15334), .ZN(n15335) );
  OAI211_X1 U18646 ( .C1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n15335), .A(
        n16338), .B(n20214), .ZN(n15336) );
  NAND3_X1 U18647 ( .A1(n15338), .A2(n15337), .A3(n15336), .ZN(P1_U3030) );
  OAI21_X1 U18648 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n13913), .A(n20787), 
        .ZN(n15339) );
  OAI21_X1 U18649 ( .B1(n15340), .B2(n20528), .A(n15339), .ZN(n15341) );
  MUX2_X1 U18650 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15341), .S(
        n20234), .Z(P1_U3477) );
  NOR3_X1 U18651 ( .A1(n12254), .A2(n9951), .A3(n13537), .ZN(n15344) );
  NOR2_X1 U18652 ( .A1(n20528), .A2(n15342), .ZN(n15343) );
  AOI211_X1 U18653 ( .C1(n15345), .C2(n10058), .A(n15344), .B(n15343), .ZN(
        n16116) );
  NOR3_X1 U18654 ( .A1(n9951), .A2(n13537), .A3(n20914), .ZN(n15346) );
  AOI21_X1 U18655 ( .B1(n15348), .B2(n15347), .A(n15346), .ZN(n15349) );
  OAI21_X1 U18656 ( .B1(n16116), .B2(n20916), .A(n15349), .ZN(n15351) );
  MUX2_X1 U18657 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15351), .S(
        n15350), .Z(P1_U3473) );
  AOI21_X1 U18658 ( .B1(n16381), .B2(n15353), .A(n15352), .ZN(n16376) );
  NAND2_X1 U18659 ( .A1(n15354), .A2(n16410), .ZN(n15355) );
  AND2_X1 U18660 ( .A1(n15356), .A2(n15355), .ZN(n16403) );
  NOR2_X1 U18661 ( .A1(n19206), .A2(n16393), .ZN(n16375) );
  NOR2_X1 U18662 ( .A1(n16376), .A2(n16375), .ZN(n16374) );
  NOR2_X1 U18663 ( .A1(n19206), .A2(n16374), .ZN(n15369) );
  INV_X1 U18664 ( .A(n19093), .ZN(n19225) );
  NAND2_X1 U18665 ( .A1(n15367), .A2(n19225), .ZN(n15365) );
  NAND2_X1 U18666 ( .A1(n19234), .A2(n19200), .ZN(n15360) );
  AOI22_X1 U18667 ( .A1(n15358), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19229), .ZN(n15359) );
  OAI211_X1 U18668 ( .C1(n15361), .C2(n19220), .A(n15360), .B(n15359), .ZN(
        n15362) );
  AOI21_X1 U18669 ( .B1(n15363), .B2(n19110), .A(n15362), .ZN(n15364) );
  OAI211_X1 U18670 ( .C1(n15366), .C2(n19202), .A(n15365), .B(n15364), .ZN(
        P2_U2824) );
  INV_X1 U18671 ( .A(n15367), .ZN(n15371) );
  NAND2_X1 U18672 ( .A1(n15371), .A2(n15370), .ZN(n15378) );
  NAND2_X1 U18673 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19229), .ZN(
        n15373) );
  AOI22_X1 U18674 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19168), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19199), .ZN(n15372) );
  OAI211_X1 U18675 ( .C1(n15374), .C2(n19214), .A(n15373), .B(n15372), .ZN(
        n15375) );
  AOI21_X1 U18676 ( .B1(n15376), .B2(n19110), .A(n15375), .ZN(n15377) );
  OAI211_X1 U18677 ( .C1(n15379), .C2(n19202), .A(n15378), .B(n15377), .ZN(
        P2_U2825) );
  AOI211_X1 U18678 ( .C1(n15382), .C2(n15381), .A(n15380), .B(n19895), .ZN(
        n15385) );
  AOI22_X1 U18679 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19229), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19199), .ZN(n15383) );
  INV_X1 U18680 ( .A(n15383), .ZN(n15384) );
  AOI211_X1 U18681 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n19168), .A(n15385), .B(
        n15384), .ZN(n15394) );
  NAND2_X1 U18682 ( .A1(n15403), .A2(n15386), .ZN(n15387) );
  NAND2_X1 U18683 ( .A1(n15459), .A2(n15387), .ZN(n15811) );
  NOR2_X1 U18684 ( .A1(n15389), .A2(n15390), .ZN(n15391) );
  OR2_X1 U18685 ( .A1(n15526), .A2(n15391), .ZN(n15804) );
  OAI22_X1 U18686 ( .A1(n15811), .A2(n19202), .B1(n15804), .B2(n19214), .ZN(
        n15392) );
  INV_X1 U18687 ( .A(n15392), .ZN(n15393) );
  OAI211_X1 U18688 ( .C1(n15395), .C2(n19217), .A(n15394), .B(n15393), .ZN(
        P2_U2831) );
  INV_X1 U18689 ( .A(n15396), .ZN(n15408) );
  AOI211_X1 U18690 ( .C1(n15628), .C2(n15398), .A(n15397), .B(n19895), .ZN(
        n15400) );
  OAI22_X1 U18691 ( .A1(n19958), .A2(n19220), .B1(n10204), .B2(n19155), .ZN(
        n15399) );
  AOI211_X1 U18692 ( .C1(P2_EBX_REG_23__SCAN_IN), .C2(n19168), .A(n15400), .B(
        n15399), .ZN(n15407) );
  NAND2_X1 U18693 ( .A1(n15477), .A2(n15401), .ZN(n15402) );
  NAND2_X1 U18694 ( .A1(n15403), .A2(n15402), .ZN(n15625) );
  INV_X1 U18695 ( .A(n15625), .ZN(n15823) );
  AOI21_X1 U18696 ( .B1(n15405), .B2(n15540), .A(n15389), .ZN(n16431) );
  AOI22_X1 U18697 ( .A1(n15823), .A2(n19223), .B1(n16431), .B2(n19200), .ZN(
        n15406) );
  OAI211_X1 U18698 ( .C1(n15408), .C2(n19217), .A(n15407), .B(n15406), .ZN(
        P2_U2832) );
  NAND2_X1 U18699 ( .A1(n19225), .A2(n15410), .ZN(n19063) );
  OAI22_X1 U18700 ( .A1(n15665), .A2(n19063), .B1(n15663), .B2(n19155), .ZN(
        n15424) );
  INV_X1 U18701 ( .A(n15665), .ZN(n15409) );
  AOI211_X1 U18702 ( .C1(n10206), .C2(n15410), .A(n15409), .B(n19895), .ZN(
        n15423) );
  INV_X1 U18703 ( .A(n15411), .ZN(n15421) );
  NOR2_X1 U18704 ( .A1(n15413), .A2(n15414), .ZN(n15415) );
  OR2_X1 U18705 ( .A1(n15412), .A2(n15415), .ZN(n15667) );
  INV_X1 U18706 ( .A(n15667), .ZN(n15842) );
  INV_X1 U18707 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15485) );
  INV_X1 U18708 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19954) );
  OAI22_X1 U18709 ( .A1(n19215), .A2(n15485), .B1(n19954), .B2(n19220), .ZN(
        n15419) );
  XNOR2_X1 U18710 ( .A(n15417), .B(n15416), .ZN(n15845) );
  NOR2_X1 U18711 ( .A1(n19214), .A2(n15845), .ZN(n15418) );
  AOI211_X1 U18712 ( .C1(n15842), .C2(n19223), .A(n15419), .B(n15418), .ZN(
        n15420) );
  OAI21_X1 U18713 ( .B1(n15421), .B2(n19217), .A(n15420), .ZN(n15422) );
  OR3_X1 U18714 ( .A1(n15424), .A2(n15423), .A3(n15422), .ZN(P2_U2834) );
  MUX2_X1 U18715 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n15425), .S(n14214), .Z(
        P2_U2856) );
  NOR2_X1 U18716 ( .A1(n15427), .A2(n15426), .ZN(n15428) );
  NAND3_X1 U18717 ( .A1(n15495), .A2(n15432), .A3(n15481), .ZN(n15434) );
  NAND2_X1 U18718 ( .A1(n15490), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15433) );
  OAI211_X1 U18719 ( .C1(n16377), .C2(n15490), .A(n15434), .B(n15433), .ZN(
        P2_U2858) );
  NAND2_X1 U18720 ( .A1(n15436), .A2(n15435), .ZN(n15438) );
  XNOR2_X1 U18721 ( .A(n15438), .B(n15437), .ZN(n15509) );
  NAND2_X1 U18722 ( .A1(n15490), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15440) );
  NAND2_X1 U18723 ( .A1(n16398), .A2(n14214), .ZN(n15439) );
  OAI211_X1 U18724 ( .C1(n15509), .C2(n15493), .A(n15440), .B(n15439), .ZN(
        P2_U2859) );
  OAI21_X1 U18725 ( .B1(n15441), .B2(n15443), .A(n15442), .ZN(n15518) );
  NAND2_X1 U18726 ( .A1(n15490), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15448) );
  NAND2_X1 U18727 ( .A1(n13222), .A2(n15444), .ZN(n15445) );
  NAND2_X1 U18728 ( .A1(n16412), .A2(n14214), .ZN(n15447) );
  OAI211_X1 U18729 ( .C1(n15518), .C2(n15493), .A(n15448), .B(n15447), .ZN(
        P2_U2860) );
  AOI21_X1 U18730 ( .B1(n15449), .B2(n15451), .A(n15450), .ZN(n15452) );
  INV_X1 U18731 ( .A(n15452), .ZN(n15524) );
  NOR2_X1 U18732 ( .A1(n15779), .A2(n15490), .ZN(n15453) );
  AOI21_X1 U18733 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n15490), .A(n15453), .ZN(
        n15454) );
  OAI21_X1 U18734 ( .B1(n15524), .B2(n15493), .A(n15454), .ZN(P2_U2861) );
  OAI21_X1 U18735 ( .B1(n15457), .B2(n15456), .A(n15455), .ZN(n15531) );
  AND2_X1 U18736 ( .A1(n15459), .A2(n15458), .ZN(n15460) );
  NOR2_X1 U18737 ( .A1(n13223), .A2(n15460), .ZN(n16421) );
  INV_X1 U18738 ( .A(n16421), .ZN(n15792) );
  NOR2_X1 U18739 ( .A1(n15792), .A2(n15490), .ZN(n15461) );
  AOI21_X1 U18740 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n15490), .A(n15461), .ZN(
        n15462) );
  OAI21_X1 U18741 ( .B1(n15531), .B2(n15493), .A(n15462), .ZN(P2_U2862) );
  AOI21_X1 U18742 ( .B1(n15463), .B2(n15465), .A(n15464), .ZN(n15466) );
  XOR2_X1 U18743 ( .A(n15467), .B(n15466), .Z(n15539) );
  NOR2_X1 U18744 ( .A1(n15811), .A2(n15490), .ZN(n15468) );
  AOI21_X1 U18745 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15490), .A(n15468), .ZN(
        n15469) );
  OAI21_X1 U18746 ( .B1(n15539), .B2(n15493), .A(n15469), .ZN(P2_U2863) );
  AOI21_X1 U18747 ( .B1(n15470), .B2(n15472), .A(n15471), .ZN(n16432) );
  NAND2_X1 U18748 ( .A1(n16432), .A2(n15481), .ZN(n15474) );
  NAND2_X1 U18749 ( .A1(n15490), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15473) );
  OAI211_X1 U18750 ( .C1(n15625), .C2(n15490), .A(n15474), .B(n15473), .ZN(
        P2_U2864) );
  OR2_X1 U18751 ( .A1(n15412), .A2(n15475), .ZN(n15476) );
  NAND2_X1 U18752 ( .A1(n15477), .A2(n15476), .ZN(n16109) );
  AOI21_X1 U18753 ( .B1(n15480), .B2(n15478), .A(n15479), .ZN(n15547) );
  NAND2_X1 U18754 ( .A1(n15547), .A2(n15481), .ZN(n15483) );
  NAND2_X1 U18755 ( .A1(n15490), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15482) );
  OAI211_X1 U18756 ( .C1(n16109), .C2(n15490), .A(n15483), .B(n15482), .ZN(
        P2_U2865) );
  OAI21_X1 U18757 ( .B1(n14279), .B2(n15484), .A(n15478), .ZN(n15555) );
  MUX2_X1 U18758 ( .A(n15667), .B(n15485), .S(n15490), .Z(n15486) );
  OAI21_X1 U18759 ( .B1(n15555), .B2(n15493), .A(n15486), .ZN(P2_U2866) );
  AND2_X1 U18760 ( .A1(n15488), .A2(n15487), .ZN(n15489) );
  OR2_X1 U18761 ( .A1(n15489), .A2(n15413), .ZN(n19056) );
  MUX2_X1 U18762 ( .A(n19056), .B(n15491), .S(n15490), .Z(n15492) );
  OAI21_X1 U18763 ( .B1(n15494), .B2(n15493), .A(n15492), .ZN(P2_U2867) );
  NAND3_X1 U18764 ( .A1(n15495), .A2(n15432), .A3(n19286), .ZN(n15501) );
  AOI21_X1 U18765 ( .B1(n15497), .B2(n9992), .A(n15496), .ZN(n16388) );
  AOI22_X1 U18766 ( .A1(n16388), .A2(n19285), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n19284), .ZN(n15500) );
  AOI22_X1 U18767 ( .A1(n19233), .A2(BUF2_REG_29__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15499) );
  NAND2_X1 U18768 ( .A1(n16430), .A2(n19241), .ZN(n15498) );
  NAND4_X1 U18769 ( .A1(n15501), .A2(n15500), .A3(n15499), .A4(n15498), .ZN(
        P2_U2890) );
  OR2_X1 U18770 ( .A1(n15513), .A2(n15502), .ZN(n15503) );
  NAND2_X1 U18771 ( .A1(n9992), .A2(n15503), .ZN(n16400) );
  OAI22_X1 U18772 ( .A1(n15552), .A2(n16400), .B1(n19250), .B2(n15504), .ZN(
        n15505) );
  AOI21_X1 U18773 ( .B1(n16430), .B2(n15506), .A(n15505), .ZN(n15508) );
  AOI22_X1 U18774 ( .A1(n19233), .A2(BUF2_REG_28__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15507) );
  OAI211_X1 U18775 ( .C1(n15509), .C2(n19257), .A(n15508), .B(n15507), .ZN(
        P2_U2891) );
  AND2_X1 U18776 ( .A1(n15511), .A2(n15510), .ZN(n15512) );
  OR2_X1 U18777 ( .A1(n15513), .A2(n15512), .ZN(n15767) );
  OAI22_X1 U18778 ( .A1(n15552), .A2(n15767), .B1(n19250), .B2(n13514), .ZN(
        n15514) );
  AOI21_X1 U18779 ( .B1(n16430), .B2(n15515), .A(n15514), .ZN(n15517) );
  AOI22_X1 U18780 ( .A1(n19233), .A2(BUF2_REG_27__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15516) );
  OAI211_X1 U18781 ( .C1(n15518), .C2(n19257), .A(n15517), .B(n15516), .ZN(
        P2_U2892) );
  OAI22_X1 U18782 ( .A1(n15552), .A2(n15784), .B1(n19250), .B2(n15519), .ZN(
        n15520) );
  AOI21_X1 U18783 ( .B1(n16430), .B2(n15521), .A(n15520), .ZN(n15523) );
  AOI22_X1 U18784 ( .A1(n19233), .A2(BUF2_REG_26__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15522) );
  OAI211_X1 U18785 ( .C1(n15524), .C2(n19257), .A(n15523), .B(n15522), .ZN(
        P2_U2893) );
  OAI21_X1 U18786 ( .B1(n15526), .B2(n15525), .A(n13227), .ZN(n16419) );
  OAI22_X1 U18787 ( .A1(n15552), .A2(n16419), .B1(n19250), .B2(n13517), .ZN(
        n15527) );
  AOI21_X1 U18788 ( .B1(n16430), .B2(n15528), .A(n15527), .ZN(n15530) );
  AOI22_X1 U18789 ( .A1(n19233), .A2(BUF2_REG_25__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15529) );
  OAI211_X1 U18790 ( .C1(n15531), .C2(n19257), .A(n15530), .B(n15529), .ZN(
        P2_U2894) );
  INV_X1 U18791 ( .A(n15804), .ZN(n15536) );
  OAI22_X1 U18792 ( .A1(n15534), .A2(n15533), .B1(n19250), .B2(n15532), .ZN(
        n15535) );
  AOI21_X1 U18793 ( .B1(n19285), .B2(n15536), .A(n15535), .ZN(n15538) );
  AOI22_X1 U18794 ( .A1(n19233), .A2(BUF2_REG_24__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15537) );
  OAI211_X1 U18795 ( .C1(n15539), .C2(n19257), .A(n15538), .B(n15537), .ZN(
        P2_U2895) );
  OAI21_X1 U18796 ( .B1(n15542), .B2(n15541), .A(n15540), .ZN(n16114) );
  AOI22_X1 U18797 ( .A1(n19233), .A2(BUF2_REG_22__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15545) );
  AOI22_X1 U18798 ( .A1(n16430), .A2(n15543), .B1(n19284), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15544) );
  OAI211_X1 U18799 ( .C1(n15552), .C2(n16114), .A(n15545), .B(n15544), .ZN(
        n15546) );
  AOI21_X1 U18800 ( .B1(n15547), .B2(n19286), .A(n15546), .ZN(n15548) );
  INV_X1 U18801 ( .A(n15548), .ZN(P2_U2897) );
  AOI22_X1 U18802 ( .A1(n19233), .A2(BUF2_REG_21__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n15551) );
  AOI22_X1 U18803 ( .A1(n16430), .A2(n15549), .B1(n19284), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15550) );
  OAI211_X1 U18804 ( .C1(n15552), .C2(n15845), .A(n15551), .B(n15550), .ZN(
        n15553) );
  INV_X1 U18805 ( .A(n15553), .ZN(n15554) );
  OAI21_X1 U18806 ( .B1(n15555), .B2(n19257), .A(n15554), .ZN(P2_U2898) );
  NAND2_X1 U18807 ( .A1(n15556), .A2(n19286), .ZN(n15563) );
  AOI22_X1 U18808 ( .A1(n16430), .A2(n15557), .B1(n19284), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15562) );
  AOI22_X1 U18809 ( .A1(n19233), .A2(BUF2_REG_19__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n15561) );
  AOI21_X1 U18810 ( .B1(n15559), .B2(n15558), .A(n14282), .ZN(n19076) );
  NAND2_X1 U18811 ( .A1(n19285), .A2(n19076), .ZN(n15560) );
  NAND4_X1 U18812 ( .A1(n15563), .A2(n15562), .A3(n15561), .A4(n15560), .ZN(
        P2_U2900) );
  NAND2_X1 U18813 ( .A1(n15564), .A2(n19286), .ZN(n15572) );
  AOI22_X1 U18814 ( .A1(n16430), .A2(n15565), .B1(n19284), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n15571) );
  AOI22_X1 U18815 ( .A1(n19233), .A2(BUF2_REG_17__SCAN_IN), .B1(n19235), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n15570) );
  NOR2_X1 U18816 ( .A1(n14042), .A2(n15566), .ZN(n15567) );
  NOR2_X1 U18817 ( .A1(n15568), .A2(n15567), .ZN(n19103) );
  NAND2_X1 U18818 ( .A1(n19285), .A2(n19103), .ZN(n15569) );
  NAND4_X1 U18819 ( .A1(n15572), .A2(n15571), .A3(n15570), .A4(n15569), .ZN(
        P2_U2902) );
  NAND2_X1 U18820 ( .A1(n15574), .A2(n15573), .ZN(n15576) );
  XOR2_X1 U18821 ( .A(n15576), .B(n15575), .Z(n15754) );
  NAND2_X1 U18822 ( .A1(n19328), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15747) );
  OAI21_X1 U18823 ( .B1(n16506), .B2(n16381), .A(n15747), .ZN(n15580) );
  NOR2_X1 U18824 ( .A1(n16377), .A2(n14136), .ZN(n15579) );
  AOI211_X1 U18825 ( .C1(n16496), .C2(n16376), .A(n15580), .B(n15579), .ZN(
        n15581) );
  INV_X1 U18826 ( .A(n15582), .ZN(n15584) );
  INV_X1 U18827 ( .A(n15577), .ZN(n15583) );
  NAND2_X1 U18828 ( .A1(n16496), .A2(n16403), .ZN(n15585) );
  NAND2_X1 U18829 ( .A1(n19328), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15768) );
  OAI211_X1 U18830 ( .C1(n16506), .C2(n16410), .A(n15585), .B(n15768), .ZN(
        n15586) );
  AOI21_X1 U18831 ( .B1(n16412), .B2(n19337), .A(n15586), .ZN(n15590) );
  OR2_X1 U18832 ( .A1(n15587), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15775) );
  NAND3_X1 U18833 ( .A1(n15775), .A2(n15588), .A3(n16502), .ZN(n15589) );
  OAI211_X1 U18834 ( .C1(n15778), .C2(n19332), .A(n15590), .B(n15589), .ZN(
        P2_U2987) );
  OAI21_X1 U18835 ( .B1(n15591), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15582), .ZN(n15790) );
  INV_X1 U18836 ( .A(n15593), .ZN(n15604) );
  NOR2_X1 U18837 ( .A1(n15592), .A2(n15604), .ZN(n15595) );
  XNOR2_X1 U18838 ( .A(n15595), .B(n15594), .ZN(n15787) );
  INV_X1 U18839 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19964) );
  NOR2_X1 U18840 ( .A1(n19181), .A2(n19964), .ZN(n15780) );
  NOR2_X1 U18841 ( .A1(n19341), .A2(n15596), .ZN(n15597) );
  AOI211_X1 U18842 ( .C1(n19329), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15780), .B(n15597), .ZN(n15598) );
  OAI21_X1 U18843 ( .B1(n15779), .B2(n14136), .A(n15598), .ZN(n15599) );
  AOI21_X1 U18844 ( .B1(n15787), .B2(n16502), .A(n15599), .ZN(n15600) );
  OAI21_X1 U18845 ( .B1(n15790), .B2(n19332), .A(n15600), .ZN(P2_U2988) );
  INV_X1 U18846 ( .A(n15592), .ZN(n15605) );
  OAI21_X1 U18847 ( .B1(n15602), .B2(n15604), .A(n15601), .ZN(n15603) );
  OAI21_X1 U18848 ( .B1(n15605), .B2(n15604), .A(n15603), .ZN(n15802) );
  AOI21_X1 U18849 ( .B1(n15793), .B2(n15606), .A(n15591), .ZN(n15791) );
  NAND2_X1 U18850 ( .A1(n15791), .A2(n16503), .ZN(n15611) );
  NAND2_X1 U18851 ( .A1(n16496), .A2(n16424), .ZN(n15607) );
  NAND2_X1 U18852 ( .A1(n19328), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15796) );
  OAI211_X1 U18853 ( .C1(n16506), .C2(n15608), .A(n15607), .B(n15796), .ZN(
        n15609) );
  AOI21_X1 U18854 ( .B1(n16421), .B2(n19337), .A(n15609), .ZN(n15610) );
  OAI211_X1 U18855 ( .C1(n19333), .C2(n15802), .A(n15611), .B(n15610), .ZN(
        P2_U2989) );
  OAI21_X1 U18856 ( .B1(n11095), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15606), .ZN(n15815) );
  INV_X1 U18857 ( .A(n15615), .ZN(n15617) );
  NAND2_X1 U18858 ( .A1(n15617), .A2(n15616), .ZN(n15618) );
  XNOR2_X1 U18859 ( .A(n15614), .B(n15618), .ZN(n15813) );
  NOR2_X1 U18860 ( .A1(n19181), .A2(n19960), .ZN(n15806) );
  NOR2_X1 U18861 ( .A1(n19341), .A2(n15619), .ZN(n15620) );
  AOI211_X1 U18862 ( .C1(n19329), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15806), .B(n15620), .ZN(n15621) );
  OAI21_X1 U18863 ( .B1(n15811), .B2(n14136), .A(n15621), .ZN(n15622) );
  AOI21_X1 U18864 ( .B1(n15813), .B2(n16502), .A(n15622), .ZN(n15623) );
  OAI21_X1 U18865 ( .B1(n15815), .B2(n19332), .A(n15623), .ZN(P2_U2990) );
  OAI21_X1 U18866 ( .B1(n15624), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15613), .ZN(n15827) );
  NAND2_X1 U18867 ( .A1(n19172), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15816) );
  OAI21_X1 U18868 ( .B1(n16506), .B2(n10204), .A(n15816), .ZN(n15627) );
  NOR2_X1 U18869 ( .A1(n15625), .A2(n14136), .ZN(n15626) );
  AOI211_X1 U18870 ( .C1(n16496), .C2(n15628), .A(n15627), .B(n15626), .ZN(
        n15633) );
  OR2_X1 U18871 ( .A1(n15630), .A2(n15629), .ZN(n15824) );
  NAND3_X1 U18872 ( .A1(n15824), .A2(n16502), .A3(n15631), .ZN(n15632) );
  OAI211_X1 U18873 ( .C1(n15827), .C2(n19332), .A(n15633), .B(n15632), .ZN(
        P2_U2991) );
  INV_X1 U18874 ( .A(n15624), .ZN(n15634) );
  OAI21_X1 U18875 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n9983), .A(
        n15634), .ZN(n15837) );
  NAND2_X1 U18876 ( .A1(n15637), .A2(n15636), .ZN(n15638) );
  XNOR2_X1 U18877 ( .A(n15635), .B(n15638), .ZN(n15835) );
  INV_X1 U18878 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19956) );
  OAI22_X1 U18879 ( .A1(n19956), .A2(n19181), .B1(n19341), .B2(n16103), .ZN(
        n15640) );
  OAI22_X1 U18880 ( .A1(n16109), .A2(n14136), .B1(n10203), .B2(n16506), .ZN(
        n15639) );
  AOI211_X1 U18881 ( .C1(n15835), .C2(n16502), .A(n15640), .B(n15639), .ZN(
        n15641) );
  OAI21_X1 U18882 ( .B1(n15837), .B2(n19332), .A(n15641), .ZN(P2_U2992) );
  OAI211_X1 U18883 ( .C1(n15719), .C2(n10275), .A(n15642), .B(n16453), .ZN(
        n15643) );
  INV_X1 U18884 ( .A(n15911), .ZN(n15644) );
  INV_X1 U18885 ( .A(n15645), .ZN(n15646) );
  NAND2_X1 U18886 ( .A1(n16439), .A2(n15646), .ZN(n15647) );
  NAND2_X1 U18887 ( .A1(n15647), .A2(n16437), .ZN(n15711) );
  INV_X1 U18888 ( .A(n15710), .ZN(n15648) );
  INV_X1 U18889 ( .A(n15649), .ZN(n15650) );
  NAND2_X1 U18890 ( .A1(n15652), .A2(n15651), .ZN(n15701) );
  OR2_X1 U18891 ( .A1(n15653), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15681) );
  NAND2_X1 U18892 ( .A1(n15681), .A2(n15692), .ZN(n15654) );
  AOI21_X1 U18893 ( .B1(n15683), .B2(n15680), .A(n15654), .ZN(n15674) );
  NAND2_X1 U18894 ( .A1(n15656), .A2(n15655), .ZN(n15657) );
  AND2_X1 U18895 ( .A1(n15658), .A2(n15657), .ZN(n15673) );
  NAND2_X1 U18896 ( .A1(n15674), .A2(n15673), .ZN(n15850) );
  NAND2_X1 U18897 ( .A1(n15850), .A2(n15658), .ZN(n15661) );
  XNOR2_X1 U18898 ( .A(n15659), .B(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15660) );
  XNOR2_X1 U18899 ( .A(n15661), .B(n15660), .ZN(n15849) );
  AOI21_X1 U18900 ( .B1(n15662), .B2(n9964), .A(n9983), .ZN(n15847) );
  NAND2_X1 U18901 ( .A1(n19172), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15839) );
  OAI21_X1 U18902 ( .B1(n16506), .B2(n15663), .A(n15839), .ZN(n15664) );
  AOI21_X1 U18903 ( .B1(n16496), .B2(n15665), .A(n15664), .ZN(n15666) );
  OAI21_X1 U18904 ( .B1(n15667), .B2(n14136), .A(n15666), .ZN(n15668) );
  AOI21_X1 U18905 ( .B1(n15847), .B2(n16503), .A(n15668), .ZN(n15669) );
  OAI21_X1 U18906 ( .B1(n15849), .B2(n19333), .A(n15669), .ZN(P2_U2993) );
  INV_X1 U18907 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15672) );
  NOR2_X1 U18908 ( .A1(n15671), .A2(n15672), .ZN(n15866) );
  OAI21_X1 U18909 ( .B1(n15866), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n9964), .ZN(n15860) );
  OR2_X1 U18910 ( .A1(n15674), .A2(n15673), .ZN(n15851) );
  NAND3_X1 U18911 ( .A1(n15851), .A2(n15850), .A3(n16502), .ZN(n15679) );
  INV_X1 U18912 ( .A(n19056), .ZN(n15677) );
  NOR2_X1 U18913 ( .A1(n19181), .A2(n19952), .ZN(n15852) );
  AOI21_X1 U18914 ( .B1(n19329), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15852), .ZN(n15675) );
  OAI21_X1 U18915 ( .B1(n19341), .B2(n19068), .A(n15675), .ZN(n15676) );
  AOI21_X1 U18916 ( .B1(n15677), .B2(n19337), .A(n15676), .ZN(n15678) );
  OAI211_X1 U18917 ( .C1(n15860), .C2(n19332), .A(n15679), .B(n15678), .ZN(
        P2_U2994) );
  NAND2_X1 U18918 ( .A1(n15681), .A2(n15680), .ZN(n15685) );
  INV_X1 U18919 ( .A(n15692), .ZN(n15682) );
  NOR2_X1 U18920 ( .A1(n15683), .A2(n15682), .ZN(n15684) );
  XOR2_X1 U18921 ( .A(n15685), .B(n15684), .Z(n15871) );
  AOI22_X1 U18922 ( .A1(n19329), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n19328), .ZN(n15686) );
  OAI21_X1 U18923 ( .B1(n19075), .B2(n14136), .A(n15686), .ZN(n15688) );
  NOR2_X1 U18924 ( .A1(n9824), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15867) );
  NOR3_X1 U18925 ( .A1(n15867), .A2(n15866), .A3(n19332), .ZN(n15687) );
  AOI211_X1 U18926 ( .C1(n16496), .C2(n19071), .A(n15688), .B(n15687), .ZN(
        n15689) );
  OAI21_X1 U18927 ( .B1(n19333), .B2(n15871), .A(n15689), .ZN(P2_U2995) );
  NOR2_X1 U18928 ( .A1(n15691), .A2(n15873), .ZN(n15702) );
  OAI21_X1 U18929 ( .B1(n15702), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15671), .ZN(n15883) );
  NAND2_X1 U18930 ( .A1(n15693), .A2(n15692), .ZN(n15695) );
  XOR2_X1 U18931 ( .A(n15695), .B(n15694), .Z(n15881) );
  INV_X1 U18932 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19948) );
  OAI22_X1 U18933 ( .A1(n19948), .A2(n19181), .B1(n19341), .B2(n19085), .ZN(
        n15698) );
  INV_X1 U18934 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15696) );
  OAI22_X1 U18935 ( .A1(n19087), .A2(n14136), .B1(n15696), .B2(n16506), .ZN(
        n15697) );
  AOI211_X1 U18936 ( .C1(n15881), .C2(n16502), .A(n15698), .B(n15697), .ZN(
        n15699) );
  OAI21_X1 U18937 ( .B1(n19332), .B2(n15883), .A(n15699), .ZN(P2_U2996) );
  XOR2_X1 U18938 ( .A(n15701), .B(n15700), .Z(n15891) );
  NOR2_X1 U18939 ( .A1(n15691), .A2(n16513), .ZN(n15894) );
  NAND2_X1 U18940 ( .A1(n15894), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15884) );
  INV_X1 U18941 ( .A(n15884), .ZN(n15704) );
  INV_X1 U18942 ( .A(n15702), .ZN(n15703) );
  OAI211_X1 U18943 ( .C1(n15704), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16503), .B(n15703), .ZN(n15709) );
  INV_X1 U18944 ( .A(n15890), .ZN(n19104) );
  INV_X1 U18945 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19946) );
  NOR2_X1 U18946 ( .A1(n19946), .A2(n19181), .ZN(n15707) );
  INV_X1 U18947 ( .A(n19096), .ZN(n19108) );
  OAI22_X1 U18948 ( .A1(n15705), .A2(n16506), .B1(n19341), .B2(n19108), .ZN(
        n15706) );
  AOI211_X1 U18949 ( .C1(n19104), .C2(n19337), .A(n15707), .B(n15706), .ZN(
        n15708) );
  OAI211_X1 U18950 ( .C1(n15891), .C2(n19333), .A(n15709), .B(n15708), .ZN(
        P2_U2997) );
  XNOR2_X1 U18951 ( .A(n15711), .B(n15710), .ZN(n15901) );
  INV_X1 U18952 ( .A(n15901), .ZN(n15716) );
  OAI211_X1 U18953 ( .C1(n15894), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15884), .B(n16503), .ZN(n15715) );
  INV_X1 U18954 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19944) );
  NOR2_X1 U18955 ( .A1(n19944), .A2(n19181), .ZN(n15713) );
  OAI22_X1 U18956 ( .A1(n10220), .A2(n16506), .B1(n19341), .B2(n19115), .ZN(
        n15712) );
  AOI211_X1 U18957 ( .C1(n19117), .C2(n19337), .A(n15713), .B(n15712), .ZN(
        n15714) );
  OAI211_X1 U18958 ( .C1(n15716), .C2(n19333), .A(n15715), .B(n15714), .ZN(
        P2_U2998) );
  INV_X1 U18959 ( .A(n15717), .ZN(n15936) );
  INV_X1 U18960 ( .A(n15917), .ZN(n15915) );
  XNOR2_X1 U18961 ( .A(n16468), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15935) );
  NAND2_X1 U18962 ( .A1(n15719), .A2(n15718), .ZN(n15723) );
  NAND2_X1 U18963 ( .A1(n15721), .A2(n15720), .ZN(n15722) );
  XNOR2_X1 U18964 ( .A(n15723), .B(n15722), .ZN(n15933) );
  INV_X1 U18965 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19936) );
  NOR2_X1 U18966 ( .A1(n19181), .A2(n19936), .ZN(n15928) );
  NOR2_X1 U18967 ( .A1(n19341), .A2(n19147), .ZN(n15724) );
  AOI211_X1 U18968 ( .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n19329), .A(
        n15928), .B(n15724), .ZN(n15725) );
  OAI21_X1 U18969 ( .B1(n19149), .B2(n14136), .A(n15725), .ZN(n15726) );
  AOI21_X1 U18970 ( .B1(n15933), .B2(n16502), .A(n15726), .ZN(n15727) );
  OAI21_X1 U18971 ( .B1(n15935), .B2(n19332), .A(n15727), .ZN(P2_U3002) );
  INV_X1 U18972 ( .A(n15731), .ZN(n16549) );
  NAND2_X1 U18973 ( .A1(n15732), .A2(n15967), .ZN(n15733) );
  NAND2_X1 U18974 ( .A1(n15733), .A2(n15968), .ZN(n15737) );
  AND2_X1 U18975 ( .A1(n15735), .A2(n15734), .ZN(n15736) );
  XNOR2_X1 U18976 ( .A(n15737), .B(n15736), .ZN(n16553) );
  AOI22_X1 U18977 ( .A1(n19176), .A2(n19337), .B1(n19329), .B2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15740) );
  INV_X1 U18978 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19930) );
  OAI22_X1 U18979 ( .A1(n19930), .A2(n19181), .B1(n19341), .B2(n19174), .ZN(
        n15738) );
  INV_X1 U18980 ( .A(n15738), .ZN(n15739) );
  OAI211_X1 U18981 ( .C1(n16553), .C2(n19333), .A(n15740), .B(n15739), .ZN(
        n15741) );
  AOI21_X1 U18982 ( .B1(n16549), .B2(n16503), .A(n15741), .ZN(n15742) );
  INV_X1 U18983 ( .A(n15742), .ZN(P2_U3006) );
  NAND2_X1 U18984 ( .A1(n15743), .A2(n16566), .ZN(n15753) );
  INV_X1 U18985 ( .A(n15772), .ZN(n15751) );
  NOR2_X1 U18986 ( .A1(n16377), .A2(n15976), .ZN(n15750) );
  INV_X1 U18987 ( .A(n16388), .ZN(n15748) );
  INV_X1 U18988 ( .A(n15770), .ZN(n15756) );
  OAI211_X1 U18989 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15745), .A(
        n15756), .B(n15744), .ZN(n15746) );
  OAI211_X1 U18990 ( .C1(n15748), .C2(n16544), .A(n15747), .B(n15746), .ZN(
        n15749) );
  AOI211_X1 U18991 ( .C1(n15751), .C2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15750), .B(n15749), .ZN(n15752) );
  OAI211_X1 U18992 ( .C1(n15754), .C2(n16552), .A(n15753), .B(n15752), .ZN(
        P2_U3017) );
  XOR2_X1 U18993 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n15755) );
  NAND2_X1 U18994 ( .A1(n15756), .A2(n15755), .ZN(n15757) );
  OAI211_X1 U18995 ( .C1(n16544), .C2(n16400), .A(n15758), .B(n15757), .ZN(
        n15761) );
  NOR2_X1 U18996 ( .A1(n15772), .A2(n15759), .ZN(n15760) );
  AOI211_X1 U18997 ( .C1(n16398), .C2(n16565), .A(n15761), .B(n15760), .ZN(
        n15765) );
  INV_X1 U18998 ( .A(n15762), .ZN(n15763) );
  NAND2_X1 U18999 ( .A1(n15763), .A2(n16563), .ZN(n15764) );
  OAI211_X1 U19000 ( .C1(n15766), .C2(n15966), .A(n15765), .B(n15764), .ZN(
        P2_U3018) );
  INV_X1 U19001 ( .A(n15767), .ZN(n16416) );
  NAND2_X1 U19002 ( .A1(n16558), .A2(n16416), .ZN(n15769) );
  OAI211_X1 U19003 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15770), .A(
        n15769), .B(n15768), .ZN(n15774) );
  NOR2_X1 U19004 ( .A1(n15772), .A2(n15771), .ZN(n15773) );
  AOI211_X1 U19005 ( .C1(n16412), .C2(n16565), .A(n15774), .B(n15773), .ZN(
        n15777) );
  NAND3_X1 U19006 ( .A1(n15775), .A2(n15588), .A3(n16563), .ZN(n15776) );
  OAI211_X1 U19007 ( .C1(n15778), .C2(n15966), .A(n15777), .B(n15776), .ZN(
        P2_U3019) );
  NOR2_X1 U19008 ( .A1(n15779), .A2(n15976), .ZN(n15786) );
  INV_X1 U19009 ( .A(n15780), .ZN(n15783) );
  OAI211_X1 U19010 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15794), .B(n15781), .ZN(
        n15782) );
  OAI211_X1 U19011 ( .C1(n16544), .C2(n15784), .A(n15783), .B(n15782), .ZN(
        n15785) );
  AOI211_X1 U19012 ( .C1(n15799), .C2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15786), .B(n15785), .ZN(n15789) );
  NAND2_X1 U19013 ( .A1(n15787), .A2(n16563), .ZN(n15788) );
  OAI211_X1 U19014 ( .C1(n15790), .C2(n15966), .A(n15789), .B(n15788), .ZN(
        P2_U3020) );
  NAND2_X1 U19015 ( .A1(n15791), .A2(n16566), .ZN(n15801) );
  NOR2_X1 U19016 ( .A1(n15792), .A2(n15976), .ZN(n15798) );
  NAND2_X1 U19017 ( .A1(n15794), .A2(n15793), .ZN(n15795) );
  OAI211_X1 U19018 ( .C1(n16544), .C2(n16419), .A(n15796), .B(n15795), .ZN(
        n15797) );
  AOI211_X1 U19019 ( .C1(n15799), .C2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15798), .B(n15797), .ZN(n15800) );
  OAI211_X1 U19020 ( .C1(n15802), .C2(n16552), .A(n15801), .B(n15800), .ZN(
        P2_U3021) );
  NAND2_X1 U19021 ( .A1(n15803), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15810) );
  NOR2_X1 U19022 ( .A1(n16544), .A2(n15804), .ZN(n15805) );
  AOI211_X1 U19023 ( .C1(n15808), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        n15809) );
  OAI211_X1 U19024 ( .C1(n15811), .C2(n15976), .A(n15810), .B(n15809), .ZN(
        n15812) );
  AOI21_X1 U19025 ( .B1(n15813), .B2(n16563), .A(n15812), .ZN(n15814) );
  OAI21_X1 U19026 ( .B1(n15815), .B2(n15966), .A(n15814), .ZN(P2_U3022) );
  OAI21_X1 U19027 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n15831), .ZN(n15818) );
  NAND2_X1 U19028 ( .A1(n16558), .A2(n16431), .ZN(n15817) );
  OAI211_X1 U19029 ( .C1(n15819), .C2(n15818), .A(n15817), .B(n15816), .ZN(
        n15822) );
  NOR2_X1 U19030 ( .A1(n15828), .A2(n15820), .ZN(n15821) );
  AOI211_X1 U19031 ( .C1(n15823), .C2(n16565), .A(n15822), .B(n15821), .ZN(
        n15826) );
  NAND3_X1 U19032 ( .A1(n15824), .A2(n16563), .A3(n15631), .ZN(n15825) );
  OAI211_X1 U19033 ( .C1(n15827), .C2(n15966), .A(n15826), .B(n15825), .ZN(
        P2_U3023) );
  NOR2_X1 U19034 ( .A1(n15828), .A2(n11094), .ZN(n15834) );
  NOR2_X1 U19035 ( .A1(n19956), .A2(n19181), .ZN(n15830) );
  NOR2_X1 U19036 ( .A1(n16544), .A2(n16114), .ZN(n15829) );
  AOI211_X1 U19037 ( .C1(n15831), .C2(n11094), .A(n15830), .B(n15829), .ZN(
        n15832) );
  OAI21_X1 U19038 ( .B1(n15976), .B2(n16109), .A(n15832), .ZN(n15833) );
  AOI211_X1 U19039 ( .C1(n15835), .C2(n16563), .A(n15834), .B(n15833), .ZN(
        n15836) );
  OAI21_X1 U19040 ( .B1(n15837), .B2(n15966), .A(n15836), .ZN(P2_U3024) );
  NAND2_X1 U19041 ( .A1(n15838), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15844) );
  OAI21_X1 U19042 ( .B1(n15840), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15839), .ZN(n15841) );
  AOI21_X1 U19043 ( .B1(n15842), .B2(n16565), .A(n15841), .ZN(n15843) );
  OAI211_X1 U19044 ( .C1(n16544), .C2(n15845), .A(n15844), .B(n15843), .ZN(
        n15846) );
  AOI21_X1 U19045 ( .B1(n15847), .B2(n16566), .A(n15846), .ZN(n15848) );
  OAI21_X1 U19046 ( .B1(n15849), .B2(n16552), .A(n15848), .ZN(P2_U3025) );
  NAND3_X1 U19047 ( .A1(n15851), .A2(n15850), .A3(n16563), .ZN(n15859) );
  NOR2_X1 U19048 ( .A1(n19056), .A2(n15976), .ZN(n15857) );
  INV_X1 U19049 ( .A(n15852), .ZN(n15855) );
  OAI211_X1 U19050 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15861), .B(n15853), .ZN(
        n15854) );
  OAI211_X1 U19051 ( .C1(n16544), .C2(n19059), .A(n15855), .B(n15854), .ZN(
        n15856) );
  AOI211_X1 U19052 ( .C1(n15872), .C2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15857), .B(n15856), .ZN(n15858) );
  OAI211_X1 U19053 ( .C1(n15860), .C2(n15966), .A(n15859), .B(n15858), .ZN(
        P2_U3026) );
  INV_X1 U19054 ( .A(n15861), .ZN(n15863) );
  NAND2_X1 U19055 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n19172), .ZN(n15862) );
  OAI21_X1 U19056 ( .B1(n15863), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15862), .ZN(n15864) );
  AOI21_X1 U19057 ( .B1(n16558), .B2(n19076), .A(n15864), .ZN(n15865) );
  OAI21_X1 U19058 ( .B1(n19075), .B2(n15976), .A(n15865), .ZN(n15869) );
  NOR3_X1 U19059 ( .A1(n15867), .A2(n15866), .A3(n15966), .ZN(n15868) );
  AOI211_X1 U19060 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15872), .A(
        n15869), .B(n15868), .ZN(n15870) );
  OAI21_X1 U19061 ( .B1(n16552), .B2(n15871), .A(n15870), .ZN(P2_U3027) );
  NAND2_X1 U19062 ( .A1(n15872), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15879) );
  NOR2_X1 U19063 ( .A1(n15873), .A2(n16512), .ZN(n15877) );
  NOR2_X1 U19064 ( .A1(n19948), .A2(n19181), .ZN(n15875) );
  NOR2_X1 U19065 ( .A1(n16544), .A2(n19092), .ZN(n15874) );
  AOI211_X1 U19066 ( .C1(n15877), .C2(n15876), .A(n15875), .B(n15874), .ZN(
        n15878) );
  OAI211_X1 U19067 ( .C1(n19087), .C2(n15976), .A(n15879), .B(n15878), .ZN(
        n15880) );
  AOI21_X1 U19068 ( .B1(n15881), .B2(n16563), .A(n15880), .ZN(n15882) );
  OAI21_X1 U19069 ( .B1(n15966), .B2(n15883), .A(n15882), .ZN(P2_U3028) );
  OAI21_X1 U19070 ( .B1(n16566), .B2(n15885), .A(n15884), .ZN(n15887) );
  AOI21_X1 U19071 ( .B1(n15913), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15944), .ZN(n15886) );
  NOR2_X1 U19072 ( .A1(n15916), .A2(n15886), .ZN(n16514) );
  OAI211_X1 U19073 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15888), .A(
        n15887), .B(n16514), .ZN(n15900) );
  AOI21_X1 U19074 ( .B1(n15909), .B2(n15889), .A(n15900), .ZN(n15899) );
  OAI22_X1 U19075 ( .A1(n15976), .A2(n15890), .B1(n19946), .B2(n19181), .ZN(
        n15893) );
  NOR2_X1 U19076 ( .A1(n15891), .A2(n16552), .ZN(n15892) );
  AOI211_X1 U19077 ( .C1(n16558), .C2(n19103), .A(n15893), .B(n15892), .ZN(
        n15897) );
  INV_X1 U19078 ( .A(n15894), .ZN(n15895) );
  OAI22_X1 U19079 ( .A1(n15895), .A2(n15966), .B1(n16513), .B2(n16512), .ZN(
        n15907) );
  NAND3_X1 U19080 ( .A1(n15907), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15898), .ZN(n15896) );
  OAI211_X1 U19081 ( .C1(n15899), .C2(n15898), .A(n15897), .B(n15896), .ZN(
        P2_U3029) );
  INV_X1 U19082 ( .A(n15900), .ZN(n15910) );
  NAND2_X1 U19083 ( .A1(n15901), .A2(n16563), .ZN(n15904) );
  INV_X1 U19084 ( .A(n19121), .ZN(n15902) );
  AOI22_X1 U19085 ( .A1(n16558), .A2(n15902), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n19328), .ZN(n15903) );
  OAI211_X1 U19086 ( .C1(n15976), .C2(n15905), .A(n15904), .B(n15903), .ZN(
        n15906) );
  AOI21_X1 U19087 ( .B1(n15907), .B2(n15909), .A(n15906), .ZN(n15908) );
  OAI21_X1 U19088 ( .B1(n15910), .B2(n15909), .A(n15908), .ZN(P2_U3030) );
  OAI21_X1 U19089 ( .B1(n9981), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15691), .ZN(n16447) );
  NAND2_X1 U19090 ( .A1(n15911), .A2(n16438), .ZN(n15912) );
  AOI22_X1 U19091 ( .A1(n19139), .A2(n16565), .B1(n16558), .B2(n19138), .ZN(
        n15923) );
  NAND2_X1 U19092 ( .A1(n15913), .A2(n15914), .ZN(n15920) );
  INV_X1 U19093 ( .A(n15914), .ZN(n15958) );
  NOR2_X1 U19094 ( .A1(n15915), .A2(n15958), .ZN(n16521) );
  NAND2_X1 U19095 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15918) );
  INV_X1 U19096 ( .A(n15916), .ZN(n15963) );
  OAI21_X1 U19097 ( .B1(n15917), .B2(n15944), .A(n15963), .ZN(n15926) );
  AOI21_X1 U19098 ( .B1(n16521), .B2(n15918), .A(n15926), .ZN(n16529) );
  NAND2_X1 U19099 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19172), .ZN(n15919) );
  OAI221_X1 U19100 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15920), 
        .C1(n11243), .C2(n16529), .A(n15919), .ZN(n15921) );
  INV_X1 U19101 ( .A(n15921), .ZN(n15922) );
  OAI211_X1 U19102 ( .C1(n16446), .C2(n16552), .A(n15923), .B(n15922), .ZN(
        n15924) );
  INV_X1 U19103 ( .A(n15924), .ZN(n15925) );
  OAI21_X1 U19104 ( .B1(n16447), .B2(n15966), .A(n15925), .ZN(P2_U3032) );
  NAND2_X1 U19105 ( .A1(n15926), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15931) );
  NOR2_X1 U19106 ( .A1(n16544), .A2(n19154), .ZN(n15927) );
  AOI211_X1 U19107 ( .C1(n16521), .C2(n15929), .A(n15928), .B(n15927), .ZN(
        n15930) );
  OAI211_X1 U19108 ( .C1(n19149), .C2(n15976), .A(n15931), .B(n15930), .ZN(
        n15932) );
  AOI21_X1 U19109 ( .B1(n15933), .B2(n16563), .A(n15932), .ZN(n15934) );
  OAI21_X1 U19110 ( .B1(n15935), .B2(n15966), .A(n15934), .ZN(P2_U3034) );
  OAI21_X1 U19111 ( .B1(n15936), .B2(n15962), .A(n15946), .ZN(n15937) );
  NAND3_X1 U19112 ( .A1(n15717), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16469) );
  NAND2_X1 U19113 ( .A1(n15937), .A2(n16469), .ZN(n16474) );
  NAND2_X1 U19114 ( .A1(n9914), .A2(n15938), .ZN(n15955) );
  INV_X1 U19115 ( .A(n15939), .ZN(n15953) );
  NOR2_X1 U19116 ( .A1(n15955), .A2(n15953), .ZN(n16465) );
  INV_X1 U19117 ( .A(n15940), .ZN(n15952) );
  OR2_X1 U19118 ( .A1(n16465), .A2(n15952), .ZN(n15943) );
  AND2_X1 U19119 ( .A1(n16464), .A2(n15941), .ZN(n15942) );
  XNOR2_X1 U19120 ( .A(n15943), .B(n15942), .ZN(n16473) );
  NOR2_X1 U19121 ( .A1(n15962), .A2(n15958), .ZN(n16536) );
  OAI21_X1 U19122 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15944), .A(
        n15963), .ZN(n16531) );
  INV_X1 U19123 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19933) );
  NOR2_X1 U19124 ( .A1(n19933), .A2(n19181), .ZN(n15945) );
  AOI221_X1 U19125 ( .B1(n16536), .B2(n15946), .C1(n16531), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15945), .ZN(n15949) );
  INV_X1 U19126 ( .A(n19167), .ZN(n15947) );
  AOI22_X1 U19127 ( .A1(n19163), .A2(n16565), .B1(n16558), .B2(n15947), .ZN(
        n15948) );
  OAI211_X1 U19128 ( .C1(n16473), .C2(n16552), .A(n15949), .B(n15948), .ZN(
        n15950) );
  INV_X1 U19129 ( .A(n15950), .ZN(n15951) );
  OAI21_X1 U19130 ( .B1(n16474), .B2(n15966), .A(n15951), .ZN(P2_U3036) );
  XNOR2_X1 U19131 ( .A(n15717), .B(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16479) );
  NOR2_X1 U19132 ( .A1(n15953), .A2(n15952), .ZN(n15954) );
  XNOR2_X1 U19133 ( .A(n15955), .B(n15954), .ZN(n16480) );
  NAND2_X1 U19134 ( .A1(n16565), .A2(n16481), .ZN(n15957) );
  NAND2_X1 U19135 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19172), .ZN(n15956) );
  OAI211_X1 U19136 ( .C1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15958), .A(
        n15957), .B(n15956), .ZN(n15959) );
  AOI21_X1 U19137 ( .B1(n16558), .B2(n15960), .A(n15959), .ZN(n15961) );
  OAI21_X1 U19138 ( .B1(n15963), .B2(n15962), .A(n15961), .ZN(n15964) );
  AOI21_X1 U19139 ( .B1(n16480), .B2(n16563), .A(n15964), .ZN(n15965) );
  OAI21_X1 U19140 ( .B1(n16479), .B2(n15966), .A(n15965), .ZN(P2_U3037) );
  NAND2_X1 U19141 ( .A1(n15968), .A2(n15967), .ZN(n15969) );
  XOR2_X1 U19142 ( .A(n15969), .B(n15732), .Z(n16489) );
  NOR2_X1 U19143 ( .A1(n15971), .A2(n15972), .ZN(n16487) );
  INV_X1 U19144 ( .A(n16487), .ZN(n15975) );
  NAND3_X1 U19145 ( .A1(n15975), .A2(n16566), .A3(n15974), .ZN(n15981) );
  NOR2_X1 U19146 ( .A1(n15976), .A2(n16488), .ZN(n15979) );
  NAND2_X1 U19147 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19172), .ZN(n15977) );
  OAI221_X1 U19148 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16541), .C1(
        n16543), .C2(n16546), .A(n15977), .ZN(n15978) );
  AOI211_X1 U19149 ( .C1(n16558), .C2(n19246), .A(n15979), .B(n15978), .ZN(
        n15980) );
  OAI211_X1 U19150 ( .C1(n16489), .C2(n16552), .A(n15981), .B(n15980), .ZN(
        P2_U3039) );
  INV_X1 U19151 ( .A(n15982), .ZN(n15984) );
  OAI222_X1 U19152 ( .A1(n15985), .A2(n15984), .B1(n19985), .B2(n15983), .C1(
        n15988), .C2(n19998), .ZN(n15986) );
  MUX2_X1 U19153 ( .A(n15986), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15989), .Z(P2_U3599) );
  OAI22_X1 U19154 ( .A1(n19988), .A2(n15988), .B1(n15987), .B2(n19985), .ZN(
        n15990) );
  MUX2_X1 U19155 ( .A(n15990), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15989), .Z(P2_U3596) );
  NAND4_X1 U19156 ( .A1(n17367), .A2(n15993), .A3(n15992), .A4(n15991), .ZN(
        n15994) );
  AOI21_X2 U19157 ( .B1(n15995), .B2(n15994), .A(n18856), .ZN(n16173) );
  INV_X1 U19158 ( .A(n17382), .ZN(n17397) );
  NAND2_X1 U19159 ( .A1(n17367), .A2(n17397), .ZN(n17391) );
  INV_X1 U19160 ( .A(n17391), .ZN(n17393) );
  NAND2_X1 U19161 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17098) );
  INV_X1 U19162 ( .A(n17367), .ZN(n18402) );
  INV_X1 U19163 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n15996) );
  INV_X1 U19164 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17037) );
  NAND3_X1 U19165 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17373) );
  NOR4_X4 U19166 ( .A1(n17037), .A2(n17374), .A3(n17382), .A4(n17373), .ZN(
        n17377) );
  NAND3_X1 U19167 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17377), .ZN(n17361) );
  AND3_X1 U19168 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .ZN(n17255) );
  NAND3_X1 U19169 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17258), .A3(n17255), 
        .ZN(n17219) );
  NOR2_X2 U19170 ( .A1(n15996), .A2(n17219), .ZN(n17232) );
  NAND2_X1 U19171 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17204), .ZN(n17193) );
  NAND2_X1 U19172 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17164), .ZN(n17158) );
  NOR2_X2 U19173 ( .A1(n16821), .A2(n17158), .ZN(n17163) );
  NOR2_X1 U19174 ( .A1(n17394), .A2(n17140), .ZN(n17147) );
  INV_X1 U19175 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16774) );
  AOI22_X1 U19176 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16000) );
  AOI22_X1 U19177 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15999) );
  AOI22_X1 U19178 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15998) );
  AOI22_X1 U19179 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15997) );
  NAND4_X1 U19180 ( .A1(n16000), .A2(n15999), .A3(n15998), .A4(n15997), .ZN(
        n16006) );
  AOI22_X1 U19181 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10358), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16004) );
  AOI22_X1 U19182 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16003) );
  AOI22_X1 U19183 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16002) );
  AOI22_X1 U19184 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16001) );
  NAND4_X1 U19185 ( .A1(n16004), .A2(n16003), .A3(n16002), .A4(n16001), .ZN(
        n16005) );
  NOR2_X1 U19186 ( .A1(n16006), .A2(n16005), .ZN(n16069) );
  AOI22_X1 U19187 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16010) );
  AOI22_X1 U19188 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16009) );
  AOI22_X1 U19189 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16008) );
  AOI22_X1 U19190 ( .A1(n17113), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16007) );
  NAND4_X1 U19191 ( .A1(n16010), .A2(n16009), .A3(n16008), .A4(n16007), .ZN(
        n16016) );
  AOI22_X1 U19192 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16014) );
  AOI22_X1 U19193 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16013) );
  AOI22_X1 U19194 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16012) );
  AOI22_X1 U19195 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16011) );
  NAND4_X1 U19196 ( .A1(n16014), .A2(n16013), .A3(n16012), .A4(n16011), .ZN(
        n16015) );
  NOR2_X1 U19197 ( .A1(n16016), .A2(n16015), .ZN(n17146) );
  AOI22_X1 U19198 ( .A1(n17347), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16020) );
  AOI22_X1 U19199 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16019) );
  AOI22_X1 U19200 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16018) );
  AOI22_X1 U19201 ( .A1(n17113), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16017) );
  NAND4_X1 U19202 ( .A1(n16020), .A2(n16019), .A3(n16018), .A4(n16017), .ZN(
        n16026) );
  AOI22_X1 U19203 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10356), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16024) );
  AOI22_X1 U19204 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n16023) );
  AOI22_X1 U19205 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16022) );
  AOI22_X1 U19206 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16021) );
  NAND4_X1 U19207 ( .A1(n16024), .A2(n16023), .A3(n16022), .A4(n16021), .ZN(
        n16025) );
  NOR2_X1 U19208 ( .A1(n16026), .A2(n16025), .ZN(n17155) );
  AOI22_X1 U19209 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16036) );
  AOI22_X1 U19210 ( .A1(n17347), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16035) );
  AOI22_X1 U19211 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16027) );
  OAI21_X1 U19212 ( .B1(n17121), .B2(n17344), .A(n16027), .ZN(n16033) );
  AOI22_X1 U19213 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16031) );
  AOI22_X1 U19214 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16030) );
  AOI22_X1 U19215 ( .A1(n17113), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16029) );
  AOI22_X1 U19216 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16028) );
  NAND4_X1 U19217 ( .A1(n16031), .A2(n16030), .A3(n16029), .A4(n16028), .ZN(
        n16032) );
  AOI211_X1 U19218 ( .C1(n9832), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n16033), .B(n16032), .ZN(n16034) );
  NAND3_X1 U19219 ( .A1(n16036), .A2(n16035), .A3(n16034), .ZN(n17160) );
  AOI22_X1 U19220 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16046) );
  AOI22_X1 U19221 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16045) );
  AOI22_X1 U19222 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17325), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n9821), .ZN(n16037) );
  OAI21_X1 U19223 ( .B1(n17364), .B2(n17166), .A(n16037), .ZN(n16043) );
  AOI22_X1 U19224 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17347), .B1(
        n10356), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16041) );
  AOI22_X1 U19225 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17340), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16040) );
  AOI22_X1 U19226 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n9813), .B1(n9832), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16039) );
  AOI22_X1 U19227 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17326), .ZN(n16038) );
  NAND4_X1 U19228 ( .A1(n16041), .A2(n16040), .A3(n16039), .A4(n16038), .ZN(
        n16042) );
  AOI211_X1 U19229 ( .C1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .C2(n17167), .A(
        n16043), .B(n16042), .ZN(n16044) );
  NAND3_X1 U19230 ( .A1(n16046), .A2(n16045), .A3(n16044), .ZN(n17161) );
  NAND2_X1 U19231 ( .A1(n17160), .A2(n17161), .ZN(n17159) );
  NOR2_X1 U19232 ( .A1(n17155), .A2(n17159), .ZN(n17152) );
  AOI22_X1 U19233 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16056) );
  AOI22_X1 U19234 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10358), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16055) );
  AOI22_X1 U19235 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16047) );
  OAI21_X1 U19236 ( .B1(n17121), .B2(n17387), .A(n16047), .ZN(n16053) );
  AOI22_X1 U19237 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16051) );
  AOI22_X1 U19238 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16050) );
  AOI22_X1 U19239 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16049) );
  AOI22_X1 U19240 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16048) );
  NAND4_X1 U19241 ( .A1(n16051), .A2(n16050), .A3(n16049), .A4(n16048), .ZN(
        n16052) );
  AOI211_X1 U19242 ( .C1(n17113), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n16053), .B(n16052), .ZN(n16054) );
  NAND3_X1 U19243 ( .A1(n16056), .A2(n16055), .A3(n16054), .ZN(n17151) );
  NAND2_X1 U19244 ( .A1(n17152), .A2(n17151), .ZN(n17150) );
  NOR2_X1 U19245 ( .A1(n17146), .A2(n17150), .ZN(n17145) );
  AOI22_X1 U19246 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9813), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16068) );
  AOI22_X1 U19247 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10358), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16067) );
  INV_X1 U19248 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16058) );
  AOI22_X1 U19249 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10356), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16057) );
  OAI21_X1 U19250 ( .B1(n16059), .B2(n16058), .A(n16057), .ZN(n16065) );
  AOI22_X1 U19251 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16063) );
  AOI22_X1 U19252 ( .A1(n17299), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16062) );
  AOI22_X1 U19253 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16061) );
  AOI22_X1 U19254 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16060) );
  NAND4_X1 U19255 ( .A1(n16063), .A2(n16062), .A3(n16061), .A4(n16060), .ZN(
        n16064) );
  AOI211_X1 U19256 ( .C1(n9835), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n16065), .B(n16064), .ZN(n16066) );
  NAND3_X1 U19257 ( .A1(n16068), .A2(n16067), .A3(n16066), .ZN(n17142) );
  NAND2_X1 U19258 ( .A1(n17145), .A2(n17142), .ZN(n17141) );
  NOR2_X1 U19259 ( .A1(n16069), .A2(n17141), .ZN(n17410) );
  AOI21_X1 U19260 ( .B1(n16069), .B2(n17141), .A(n17410), .ZN(n17416) );
  AND2_X1 U19261 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17140), .ZN(n17144) );
  AOI22_X1 U19262 ( .A1(n17416), .A2(n17394), .B1(n17144), .B2(n16774), .ZN(
        n16070) );
  OAI21_X1 U19263 ( .B1(n17137), .B2(n16774), .A(n16070), .ZN(P3_U2675) );
  AOI22_X1 U19264 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16075) );
  AOI22_X1 U19265 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16074) );
  AOI22_X1 U19266 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16073) );
  AOI22_X1 U19267 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16072) );
  NAND4_X1 U19268 ( .A1(n16075), .A2(n16074), .A3(n16073), .A4(n16072), .ZN(
        n16081) );
  AOI22_X1 U19269 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16079) );
  AOI22_X1 U19270 ( .A1(n10378), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16078) );
  AOI22_X1 U19271 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16077) );
  AOI22_X1 U19272 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16076) );
  NAND4_X1 U19273 ( .A1(n16079), .A2(n16078), .A3(n16077), .A4(n16076), .ZN(
        n16080) );
  NOR2_X1 U19274 ( .A1(n16081), .A2(n16080), .ZN(n17496) );
  INV_X2 U19275 ( .A(n17394), .ZN(n17388) );
  INV_X1 U19276 ( .A(n17295), .ZN(n16082) );
  OAI33_X1 U19277 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18402), .A3(n17295), 
        .B1(n16935), .B2(n17394), .B3(n16082), .ZN(n16083) );
  INV_X1 U19278 ( .A(n16083), .ZN(n16084) );
  OAI21_X1 U19279 ( .B1(n17496), .B2(n17388), .A(n16084), .ZN(P3_U2690) );
  NAND2_X1 U19280 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18588) );
  AOI221_X1 U19281 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18588), .C1(n16086), 
        .C2(n18588), .A(n16085), .ZN(n18361) );
  NOR2_X1 U19282 ( .A1(n16087), .A2(n18636), .ZN(n16088) );
  OAI21_X1 U19283 ( .B1(n16088), .B2(n18358), .A(n18362), .ZN(n18359) );
  AOI22_X1 U19284 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18361), .B1(
        n18359), .B2(n18367), .ZN(P3_U2865) );
  INV_X1 U19285 ( .A(n16089), .ZN(n16090) );
  NOR4_X1 U19286 ( .A1(n11484), .A2(n16090), .A3(n11507), .A4(n19985), .ZN(
        n16091) );
  NAND2_X1 U19287 ( .A1(n16093), .A2(n16091), .ZN(n16092) );
  OAI21_X1 U19288 ( .B1(n16093), .B2(n11119), .A(n16092), .ZN(P2_U3595) );
  NOR2_X1 U19289 ( .A1(n18043), .A2(n16094), .ZN(n16603) );
  INV_X1 U19290 ( .A(n16605), .ZN(n16586) );
  NOR2_X1 U19291 ( .A1(n16586), .A2(n18352), .ZN(n16095) );
  AOI211_X1 U19292 ( .C1(n18266), .C2(n16603), .A(n16096), .B(n16095), .ZN(
        n16158) );
  AOI21_X1 U19293 ( .B1(n18202), .B2(n17686), .A(n16097), .ZN(n16604) );
  OAI22_X1 U19294 ( .A1(n18352), .A2(n16585), .B1(n18199), .B2(n16589), .ZN(
        n16098) );
  INV_X1 U19295 ( .A(n16098), .ZN(n16163) );
  OAI21_X1 U19296 ( .B1(n9828), .B2(n16604), .A(n16163), .ZN(n16099) );
  AOI21_X1 U19297 ( .B1(n18260), .B2(n17661), .A(n16099), .ZN(n16101) );
  OAI221_X1 U19298 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16158), 
        .C1(n9871), .C2(n16101), .A(n16100), .ZN(P3_U2833) );
  INV_X1 U19299 ( .A(n16103), .ZN(n16105) );
  INV_X1 U19300 ( .A(n16102), .ZN(n16104) );
  AOI221_X1 U19301 ( .B1(n16105), .B2(n16104), .C1(n16103), .C2(n16102), .A(
        n19895), .ZN(n16108) );
  INV_X1 U19302 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16106) );
  OAI22_X1 U19303 ( .A1(n19215), .A2(n16106), .B1(n19956), .B2(n19220), .ZN(
        n16107) );
  AOI211_X1 U19304 ( .C1(n19229), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16108), .B(n16107), .ZN(n16113) );
  OAI22_X1 U19305 ( .A1(n16110), .A2(n19217), .B1(n16109), .B2(n19202), .ZN(
        n16111) );
  INV_X1 U19306 ( .A(n16111), .ZN(n16112) );
  OAI211_X1 U19307 ( .C1(n16114), .C2(n19214), .A(n16113), .B(n16112), .ZN(
        P2_U2833) );
  INV_X1 U19308 ( .A(n16126), .ZN(n16130) );
  INV_X1 U19309 ( .A(n16115), .ZN(n16117) );
  NOR2_X1 U19310 ( .A1(n16117), .A2(n16116), .ZN(n16121) );
  INV_X1 U19311 ( .A(n16121), .ZN(n16119) );
  OAI211_X1 U19312 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n16119), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16118), .ZN(n16120) );
  OAI21_X1 U19313 ( .B1(n20585), .B2(n16121), .A(n16120), .ZN(n16125) );
  NAND2_X1 U19314 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16125), .ZN(
        n16122) );
  NAND2_X1 U19315 ( .A1(n16123), .A2(n16122), .ZN(n16124) );
  OAI21_X1 U19316 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16125), .A(
        n16124), .ZN(n16127) );
  INV_X1 U19317 ( .A(n16127), .ZN(n16129) );
  OAI21_X1 U19318 ( .B1(n16127), .B2(n16126), .A(n20658), .ZN(n16128) );
  OAI21_X1 U19319 ( .B1(n16130), .B2(n16129), .A(n16128), .ZN(n16139) );
  INV_X1 U19320 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21189) );
  NAND2_X1 U19321 ( .A1(n20057), .A2(n21189), .ZN(n16132) );
  AOI21_X1 U19322 ( .B1(n16133), .B2(n16132), .A(n16131), .ZN(n16135) );
  NAND3_X1 U19323 ( .A1(n16136), .A2(n16135), .A3(n16134), .ZN(n16137) );
  AOI211_X1 U19324 ( .C1(n16140), .C2(n16139), .A(n16138), .B(n16137), .ZN(
        n16151) );
  AOI21_X1 U19325 ( .B1(n16151), .B2(P1_STATE2_REG_0__SCAN_IN), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16147) );
  NAND4_X1 U19326 ( .A1(n16143), .A2(n16142), .A3(n16141), .A4(n21085), .ZN(
        n16146) );
  OAI21_X1 U19327 ( .B1(n16144), .B2(n20936), .A(n16150), .ZN(n16145) );
  NAND2_X1 U19328 ( .A1(n16146), .A2(n16145), .ZN(n16367) );
  NOR2_X1 U19329 ( .A1(n16147), .A2(n16367), .ZN(n16371) );
  AOI21_X1 U19330 ( .B1(n20859), .B2(n20929), .A(n16154), .ZN(n16149) );
  OAI211_X1 U19331 ( .C1(n16151), .C2(n16150), .A(n16149), .B(n16148), .ZN(
        n16152) );
  NOR2_X1 U19332 ( .A1(n16371), .A2(n16152), .ZN(n16157) );
  NAND2_X1 U19333 ( .A1(n16154), .A2(n16153), .ZN(n16155) );
  NAND2_X1 U19334 ( .A1(n20932), .A2(n16155), .ZN(n16156) );
  OAI22_X1 U19335 ( .A1(n16157), .A2(n20932), .B1(n16371), .B2(n16156), .ZN(
        P1_U3161) );
  NOR3_X1 U19336 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16158), .A3(
        n9871), .ZN(n16159) );
  INV_X1 U19337 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20867) );
  INV_X1 U19338 ( .A(HOLD), .ZN(n21248) );
  NOR2_X1 U19339 ( .A1(n20867), .A2(n21248), .ZN(n20855) );
  AOI22_X1 U19340 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n16166) );
  NAND2_X1 U19341 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20859), .ZN(n20860) );
  OAI211_X1 U19342 ( .C1(n20855), .C2(n16166), .A(n16165), .B(n20860), .ZN(
        P1_U3195) );
  AND2_X1 U19343 ( .A1(n16167), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U19344 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16169) );
  NOR2_X1 U19345 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16168) );
  NOR3_X1 U19346 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19032), .A3(n20046), 
        .ZN(n16573) );
  NOR4_X1 U19347 ( .A1(n16169), .A2(n16168), .A3(n16573), .A4(n16170), .ZN(
        P2_U3178) );
  INV_X1 U19348 ( .A(n20021), .ZN(n20018) );
  NOR2_X1 U19349 ( .A1(n16171), .A2(n20018), .ZN(P2_U3047) );
  NAND3_X1 U19350 ( .A1(n16172), .A2(n19009), .A3(n19015), .ZN(n17591) );
  NAND3_X1 U19351 ( .A1(n19014), .A2(n16174), .A3(n16173), .ZN(n16175) );
  INV_X1 U19352 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17625) );
  NAND2_X1 U19353 ( .A1(n17367), .A2(n17401), .ZN(n17445) );
  NAND2_X1 U19354 ( .A1(n17401), .A2(n16177), .ZN(n17539) );
  NAND2_X1 U19355 ( .A1(n16178), .A2(n17401), .ZN(n17536) );
  AOI22_X1 U19356 ( .A1(n17547), .A2(BUF2_REG_0__SCAN_IN), .B1(n17546), .B2(
        n16179), .ZN(n16180) );
  OAI221_X1 U19357 ( .B1(n17550), .B2(n17625), .C1(n17550), .C2(n17445), .A(
        n16180), .ZN(P3_U2735) );
  AOI22_X1 U19358 ( .A1(n16182), .A2(n16181), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n20127), .ZN(n16183) );
  OAI21_X1 U19359 ( .B1(n16184), .B2(n20115), .A(n16183), .ZN(n16185) );
  AOI21_X1 U19360 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n16198), .A(n16185), 
        .ZN(n16190) );
  INV_X1 U19361 ( .A(n16186), .ZN(n16187) );
  AOI22_X1 U19362 ( .A1(n16188), .A2(n20106), .B1(n16187), .B2(n20126), .ZN(
        n16189) );
  OAI211_X1 U19363 ( .C1(n16191), .C2(n20140), .A(n16190), .B(n16189), .ZN(
        P1_U2819) );
  OAI22_X1 U19364 ( .A1(n20104), .A2(n21215), .B1(n16192), .B2(n20115), .ZN(
        n16193) );
  AOI21_X1 U19365 ( .B1(n16194), .B2(n20084), .A(n16193), .ZN(n16202) );
  INV_X1 U19366 ( .A(n16195), .ZN(n16200) );
  OAI21_X1 U19367 ( .B1(n16197), .B2(n16246), .A(n16196), .ZN(n16199) );
  AOI22_X1 U19368 ( .A1(n16200), .A2(n20106), .B1(n16199), .B2(n16198), .ZN(
        n16201) );
  OAI211_X1 U19369 ( .C1(n20080), .C2(n16203), .A(n16202), .B(n16201), .ZN(
        P1_U2820) );
  NOR2_X1 U19370 ( .A1(n16204), .A2(n16246), .ZN(n16206) );
  AOI22_X1 U19371 ( .A1(n16207), .A2(n20084), .B1(n16206), .B2(n16205), .ZN(
        n16215) );
  AOI22_X1 U19372 ( .A1(n16208), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n20127), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n16214) );
  AOI21_X1 U19373 ( .B1(n20133), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20132), .ZN(n16213) );
  INV_X1 U19374 ( .A(n16209), .ZN(n16210) );
  AOI22_X1 U19375 ( .A1(n16211), .A2(n20106), .B1(n20126), .B2(n16210), .ZN(
        n16212) );
  NAND4_X1 U19376 ( .A1(n16215), .A2(n16214), .A3(n16213), .A4(n16212), .ZN(
        P1_U2822) );
  INV_X1 U19377 ( .A(n16216), .ZN(n16223) );
  INV_X1 U19378 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21225) );
  NOR3_X1 U19379 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n21225), .A3(n16224), 
        .ZN(n16221) );
  NAND2_X1 U19380 ( .A1(n20084), .A2(n16217), .ZN(n16219) );
  AOI21_X1 U19381 ( .B1(n20133), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20132), .ZN(n16218) );
  OAI211_X1 U19382 ( .C1(n20104), .C2(n21202), .A(n16219), .B(n16218), .ZN(
        n16220) );
  OR2_X1 U19383 ( .A1(n16221), .A2(n16220), .ZN(n16222) );
  AOI21_X1 U19384 ( .B1(n16223), .B2(n20106), .A(n16222), .ZN(n16226) );
  NOR2_X1 U19385 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n16224), .ZN(n16232) );
  OAI21_X1 U19386 ( .B1(n16228), .B2(n16232), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n16225) );
  OAI211_X1 U19387 ( .C1(n16227), .C2(n20080), .A(n16226), .B(n16225), .ZN(
        P1_U2824) );
  AOI22_X1 U19388 ( .A1(n16228), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_EBX_REG_15__SCAN_IN), .B2(n20127), .ZN(n16229) );
  OAI211_X1 U19389 ( .C1(n20115), .C2(n16230), .A(n16229), .B(n20113), .ZN(
        n16231) );
  AOI211_X1 U19390 ( .C1(n20084), .C2(n16271), .A(n16232), .B(n16231), .ZN(
        n16235) );
  NOR2_X1 U19391 ( .A1(n16311), .A2(n20080), .ZN(n16233) );
  AOI21_X1 U19392 ( .B1(n16272), .B2(n20106), .A(n16233), .ZN(n16234) );
  NAND2_X1 U19393 ( .A1(n16235), .A2(n16234), .ZN(P1_U2825) );
  OAI22_X1 U19394 ( .A1(n16236), .A2(n20080), .B1(n14464), .B2(n20104), .ZN(
        n16237) );
  AOI211_X1 U19395 ( .C1(n20133), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20132), .B(n16237), .ZN(n16245) );
  INV_X1 U19396 ( .A(n16238), .ZN(n16239) );
  AOI22_X1 U19397 ( .A1(n16240), .A2(n20084), .B1(n20106), .B2(n16239), .ZN(
        n16244) );
  OAI221_X1 U19398 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(P1_REIP_REG_11__SCAN_IN), .C1(P1_REIP_REG_12__SCAN_IN), .C2(n16242), .A(n16241), .ZN(n16243) );
  NAND3_X1 U19399 ( .A1(n16245), .A2(n16244), .A3(n16243), .ZN(P1_U2828) );
  INV_X1 U19400 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n21245) );
  OAI22_X1 U19401 ( .A1(n16246), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n21245), 
        .B2(n20104), .ZN(n16250) );
  AOI22_X1 U19402 ( .A1(n20126), .A2(n16318), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n16247), .ZN(n16248) );
  OAI211_X1 U19403 ( .C1(n20115), .C2(n12564), .A(n16248), .B(n20113), .ZN(
        n16249) );
  AOI211_X1 U19404 ( .C1(n20106), .C2(n16280), .A(n16250), .B(n16249), .ZN(
        n16251) );
  OAI21_X1 U19405 ( .B1(n16283), .B2(n20140), .A(n16251), .ZN(P1_U2829) );
  OAI21_X1 U19406 ( .B1(n16254), .B2(n16253), .A(n16252), .ZN(n16257) );
  NAND2_X1 U19407 ( .A1(n16257), .A2(n16255), .ZN(n16256) );
  MUX2_X1 U19408 ( .A(n16257), .B(n16256), .S(n16276), .Z(n16258) );
  XNOR2_X1 U19409 ( .A(n16258), .B(n16302), .ZN(n16310) );
  AOI22_X1 U19410 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n10057), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16262) );
  AOI22_X1 U19411 ( .A1(n16260), .A2(n20188), .B1(n16270), .B2(n16259), .ZN(
        n16261) );
  OAI211_X1 U19412 ( .C1(n20056), .C2(n16310), .A(n16262), .B(n16261), .ZN(
        P1_U2982) );
  INV_X1 U19413 ( .A(n16263), .ZN(n16264) );
  NOR2_X1 U19414 ( .A1(n16265), .A2(n16264), .ZN(n16269) );
  NAND2_X1 U19415 ( .A1(n16267), .A2(n16266), .ZN(n16268) );
  XNOR2_X1 U19416 ( .A(n16269), .B(n16268), .ZN(n16317) );
  AOI22_X1 U19417 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n10057), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16274) );
  AOI22_X1 U19418 ( .A1(n16272), .A2(n20188), .B1(n16271), .B2(n16270), .ZN(
        n16273) );
  OAI211_X1 U19419 ( .C1(n16317), .C2(n20056), .A(n16274), .B(n16273), .ZN(
        P1_U2984) );
  AOI22_X1 U19420 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n10057), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16282) );
  NOR3_X1 U19421 ( .A1(n15094), .A2(n16276), .A3(n16275), .ZN(n16278) );
  NOR2_X1 U19422 ( .A1(n16278), .A2(n16277), .ZN(n16279) );
  XNOR2_X1 U19423 ( .A(n16279), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16320) );
  AOI22_X1 U19424 ( .A1(n20189), .A2(n16320), .B1(n20188), .B2(n16280), .ZN(
        n16281) );
  OAI211_X1 U19425 ( .C1(n20193), .C2(n16283), .A(n16282), .B(n16281), .ZN(
        P1_U2988) );
  AOI22_X1 U19426 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n10057), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16289) );
  NAND2_X1 U19427 ( .A1(n16286), .A2(n16285), .ZN(n16287) );
  XNOR2_X1 U19428 ( .A(n16284), .B(n16287), .ZN(n16347) );
  AOI22_X1 U19429 ( .A1(n16347), .A2(n20189), .B1(n20188), .B2(n20095), .ZN(
        n16288) );
  OAI211_X1 U19430 ( .C1(n20193), .C2(n20098), .A(n16289), .B(n16288), .ZN(
        P1_U2992) );
  AOI22_X1 U19431 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n10057), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16294) );
  XNOR2_X1 U19432 ( .A(n16291), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16292) );
  XNOR2_X1 U19433 ( .A(n16290), .B(n16292), .ZN(n16353) );
  AOI22_X1 U19434 ( .A1(n16353), .A2(n20189), .B1(n20188), .B2(n20107), .ZN(
        n16293) );
  OAI211_X1 U19435 ( .C1(n20193), .C2(n20110), .A(n16294), .B(n16293), .ZN(
        P1_U2993) );
  AOI22_X1 U19436 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n10057), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16301) );
  OAI21_X1 U19437 ( .B1(n16297), .B2(n16296), .A(n16295), .ZN(n16298) );
  INV_X1 U19438 ( .A(n16298), .ZN(n16359) );
  INV_X1 U19439 ( .A(n16299), .ZN(n20122) );
  AOI22_X1 U19440 ( .A1(n16359), .A2(n20189), .B1(n20188), .B2(n20122), .ZN(
        n16300) );
  OAI211_X1 U19441 ( .C1(n20193), .C2(n20124), .A(n16301), .B(n16300), .ZN(
        P1_U2994) );
  NAND3_X1 U19442 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16304) );
  OAI21_X1 U19443 ( .B1(n16304), .B2(n16303), .A(n16302), .ZN(n16306) );
  AOI22_X1 U19444 ( .A1(n16307), .A2(n16306), .B1(n20205), .B2(n16305), .ZN(
        n16309) );
  NAND2_X1 U19445 ( .A1(n10057), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16308) );
  OAI211_X1 U19446 ( .C1(n16310), .C2(n16326), .A(n16309), .B(n16308), .ZN(
        P1_U3014) );
  INV_X1 U19447 ( .A(n16311), .ZN(n16312) );
  AOI22_X1 U19448 ( .A1(n16312), .A2(n20205), .B1(n10057), .B2(
        P1_REIP_REG_15__SCAN_IN), .ZN(n16316) );
  OAI21_X1 U19449 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16314), .A(
        n16313), .ZN(n16315) );
  OAI211_X1 U19450 ( .C1(n16317), .C2(n16326), .A(n16316), .B(n16315), .ZN(
        P1_U3016) );
  AOI22_X1 U19451 ( .A1(n16318), .A2(n20205), .B1(n10057), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16322) );
  AOI22_X1 U19452 ( .A1(n16320), .A2(n20215), .B1(n16319), .B2(n16323), .ZN(
        n16321) );
  OAI211_X1 U19453 ( .C1(n16324), .C2(n16323), .A(n16322), .B(n16321), .ZN(
        P1_U3020) );
  INV_X1 U19454 ( .A(n20079), .ZN(n16330) );
  OAI22_X1 U19455 ( .A1(n20222), .A2(n21276), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16325), .ZN(n16329) );
  NOR2_X1 U19456 ( .A1(n16327), .A2(n16326), .ZN(n16328) );
  AOI211_X1 U19457 ( .C1(n20205), .C2(n16330), .A(n16329), .B(n16328), .ZN(
        n16331) );
  OAI21_X1 U19458 ( .B1(n16332), .B2(n14406), .A(n16331), .ZN(P1_U3022) );
  NAND2_X1 U19459 ( .A1(n20201), .A2(n16362), .ZN(n16357) );
  INV_X1 U19460 ( .A(n16334), .ZN(n20213) );
  AOI21_X1 U19461 ( .B1(n20213), .B2(n16333), .A(n20212), .ZN(n20195) );
  OAI21_X1 U19462 ( .B1(n16334), .B2(n20201), .A(n20195), .ZN(n16335) );
  AOI21_X1 U19463 ( .B1(n20221), .B2(n16336), .A(n16335), .ZN(n16363) );
  OAI21_X1 U19464 ( .B1(n16337), .B2(n16357), .A(n16363), .ZN(n16352) );
  AOI21_X1 U19465 ( .B1(n16339), .B2(n16338), .A(n16352), .ZN(n16351) );
  INV_X1 U19466 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16345) );
  AOI222_X1 U19467 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n10057), .B1(n20205), 
        .B2(n16341), .C1(n20215), .C2(n16340), .ZN(n16344) );
  NAND2_X1 U19468 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16342) );
  OAI211_X1 U19469 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16346), .B(n16342), .ZN(n16343) );
  OAI211_X1 U19470 ( .C1(n16351), .C2(n16345), .A(n16344), .B(n16343), .ZN(
        P1_U3023) );
  INV_X1 U19471 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16350) );
  AOI22_X1 U19472 ( .A1(n20094), .A2(n20205), .B1(n10057), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16349) );
  AOI22_X1 U19473 ( .A1(n16347), .A2(n20215), .B1(n16346), .B2(n16350), .ZN(
        n16348) );
  OAI211_X1 U19474 ( .C1(n16351), .C2(n16350), .A(n16349), .B(n16348), .ZN(
        P1_U3024) );
  AOI22_X1 U19475 ( .A1(n20100), .A2(n20205), .B1(n10057), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16355) );
  AOI22_X1 U19476 ( .A1(n16353), .A2(n20215), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16352), .ZN(n16354) );
  OAI211_X1 U19477 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16356), .A(
        n16355), .B(n16354), .ZN(P1_U3025) );
  AOI22_X1 U19478 ( .A1(n20117), .A2(n20205), .B1(n10057), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16361) );
  INV_X1 U19479 ( .A(n16357), .ZN(n16358) );
  AOI22_X1 U19480 ( .A1(n16359), .A2(n20215), .B1(n16358), .B2(n20202), .ZN(
        n16360) );
  OAI211_X1 U19481 ( .C1(n16363), .C2(n16362), .A(n16361), .B(n16360), .ZN(
        P1_U3026) );
  INV_X1 U19482 ( .A(n16364), .ZN(n16366) );
  NAND4_X1 U19483 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20929), .A4(n20936), .ZN(n16365) );
  NAND2_X1 U19484 ( .A1(n16366), .A2(n16365), .ZN(n20850) );
  OAI21_X1 U19485 ( .B1(n16368), .B2(n20850), .A(n16367), .ZN(n16369) );
  OAI221_X1 U19486 ( .B1(n20931), .B2(n20664), .C1(n20931), .C2(n20936), .A(
        n16369), .ZN(n16370) );
  AOI221_X1 U19487 ( .B1(n16371), .B2(n20849), .C1(n20932), .C2(n20849), .A(
        n16370), .ZN(P1_U3162) );
  NOR2_X1 U19488 ( .A1(n16371), .A2(n20932), .ZN(n16373) );
  OAI21_X1 U19489 ( .B1(n16373), .B2(n20664), .A(n16372), .ZN(P1_U3466) );
  AOI211_X1 U19490 ( .C1(n16376), .C2(n16375), .A(n16374), .B(n19895), .ZN(
        n16387) );
  INV_X1 U19491 ( .A(n16377), .ZN(n16378) );
  AOI22_X1 U19492 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19199), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19168), .ZN(n16380) );
  OAI21_X1 U19493 ( .B1(n16381), .B2(n19155), .A(n16380), .ZN(n16382) );
  INV_X1 U19494 ( .A(n16382), .ZN(n16383) );
  AOI211_X1 U19495 ( .C1(n19200), .C2(n16388), .A(n16387), .B(n16386), .ZN(
        n16389) );
  INV_X1 U19496 ( .A(n16389), .ZN(P2_U2826) );
  NAND2_X1 U19497 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19229), .ZN(
        n16391) );
  AOI22_X1 U19498 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n19199), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n19168), .ZN(n16390) );
  OAI211_X1 U19499 ( .C1(n16392), .C2(n19217), .A(n16391), .B(n16390), .ZN(
        n16397) );
  AOI211_X1 U19500 ( .C1(n16395), .C2(n16394), .A(n16393), .B(n19895), .ZN(
        n16396) );
  AOI211_X1 U19501 ( .C1(n19223), .C2(n16398), .A(n16397), .B(n16396), .ZN(
        n16399) );
  OAI21_X1 U19502 ( .B1(n16400), .B2(n19214), .A(n16399), .ZN(P2_U2827) );
  AOI211_X1 U19503 ( .C1(n16403), .C2(n16402), .A(n16401), .B(n19895), .ZN(
        n16415) );
  INV_X1 U19504 ( .A(n16404), .ZN(n16406) );
  OAI211_X1 U19505 ( .C1(n16407), .C2(n16406), .A(n16405), .B(n19110), .ZN(
        n16409) );
  AOI22_X1 U19506 ( .A1(P2_REIP_REG_27__SCAN_IN), .A2(n19199), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n19168), .ZN(n16408) );
  OAI211_X1 U19507 ( .C1(n19155), .C2(n16410), .A(n16409), .B(n16408), .ZN(
        n16411) );
  AOI21_X1 U19508 ( .B1(n16412), .B2(n19223), .A(n16411), .ZN(n16413) );
  INV_X1 U19509 ( .A(n16413), .ZN(n16414) );
  AOI211_X1 U19510 ( .C1(n19200), .C2(n16416), .A(n16415), .B(n16414), .ZN(
        n16417) );
  INV_X1 U19511 ( .A(n16417), .ZN(P2_U2828) );
  AOI22_X1 U19512 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19199), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19168), .ZN(n16429) );
  AOI22_X1 U19513 ( .A1(n16418), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19229), .ZN(n16428) );
  INV_X1 U19514 ( .A(n16419), .ZN(n16420) );
  AOI22_X1 U19515 ( .A1(n16421), .A2(n19223), .B1(n16420), .B2(n19200), .ZN(
        n16427) );
  AOI21_X1 U19516 ( .B1(n16424), .B2(n16423), .A(n16422), .ZN(n16425) );
  NAND2_X1 U19517 ( .A1(n19191), .A2(n16425), .ZN(n16426) );
  NAND4_X1 U19518 ( .A1(n16429), .A2(n16428), .A3(n16427), .A4(n16426), .ZN(
        P2_U2830) );
  AOI22_X1 U19519 ( .A1(n16430), .A2(n19245), .B1(n19284), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16435) );
  AOI22_X1 U19520 ( .A1(n19235), .A2(BUF1_REG_23__SCAN_IN), .B1(n19233), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n16434) );
  AOI22_X1 U19521 ( .A1(n16432), .A2(n19286), .B1(n19285), .B2(n16431), .ZN(
        n16433) );
  NAND3_X1 U19522 ( .A1(n16435), .A2(n16434), .A3(n16433), .ZN(P2_U2896) );
  AOI22_X1 U19523 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19172), .B1(n16496), 
        .B2(n19124), .ZN(n16444) );
  NAND2_X1 U19524 ( .A1(n16437), .A2(n16436), .ZN(n16441) );
  NAND2_X1 U19525 ( .A1(n16439), .A2(n16438), .ZN(n16440) );
  XOR2_X1 U19526 ( .A(n16441), .B(n16440), .Z(n16520) );
  INV_X1 U19527 ( .A(n16520), .ZN(n16442) );
  XNOR2_X1 U19528 ( .A(n15691), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16517) );
  AOI222_X1 U19529 ( .A1(n16442), .A2(n16502), .B1(n19337), .B2(n19128), .C1(
        n16503), .C2(n16517), .ZN(n16443) );
  OAI211_X1 U19530 ( .C1(n16445), .C2(n16506), .A(n16444), .B(n16443), .ZN(
        P2_U2999) );
  AOI22_X1 U19531 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19172), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19329), .ZN(n16450) );
  OAI22_X1 U19532 ( .A1(n16447), .A2(n19332), .B1(n19333), .B2(n16446), .ZN(
        n16448) );
  AOI21_X1 U19533 ( .B1(n19337), .B2(n19139), .A(n16448), .ZN(n16449) );
  OAI211_X1 U19534 ( .C1(n19341), .C2(n19133), .A(n16450), .B(n16449), .ZN(
        P2_U3000) );
  AOI22_X1 U19535 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19172), .B1(n16496), 
        .B2(n16451), .ZN(n16458) );
  AOI21_X1 U19536 ( .B1(n16468), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16452) );
  NOR2_X1 U19537 ( .A1(n16452), .A2(n9981), .ZN(n16525) );
  NAND2_X1 U19538 ( .A1(n16454), .A2(n16453), .ZN(n16456) );
  XOR2_X1 U19539 ( .A(n16456), .B(n16455), .Z(n16524) );
  AOI222_X1 U19540 ( .A1(n16525), .A2(n16503), .B1(n16502), .B2(n16524), .C1(
        n19337), .C2(n16523), .ZN(n16457) );
  OAI211_X1 U19541 ( .C1(n16459), .C2(n16506), .A(n16458), .B(n16457), .ZN(
        P2_U3001) );
  AOI22_X1 U19542 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19172), .B1(n16496), 
        .B2(n16460), .ZN(n16471) );
  NAND2_X1 U19543 ( .A1(n16462), .A2(n16461), .ZN(n16467) );
  AOI21_X1 U19544 ( .B1(n16465), .B2(n16464), .A(n16463), .ZN(n16466) );
  XOR2_X1 U19545 ( .A(n16467), .B(n16466), .Z(n16534) );
  AOI21_X1 U19546 ( .B1(n11332), .B2(n16469), .A(n16468), .ZN(n16532) );
  OAI211_X1 U19547 ( .C1(n16472), .C2(n16506), .A(n16471), .B(n16470), .ZN(
        P2_U3003) );
  AOI22_X1 U19548 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19172), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19329), .ZN(n16477) );
  OAI22_X1 U19549 ( .A1(n16474), .A2(n19332), .B1(n16473), .B2(n19333), .ZN(
        n16475) );
  AOI21_X1 U19550 ( .B1(n19337), .B2(n19163), .A(n16475), .ZN(n16476) );
  OAI211_X1 U19551 ( .C1(n19341), .C2(n19161), .A(n16477), .B(n16476), .ZN(
        P2_U3004) );
  AOI22_X1 U19552 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19172), .B1(n16496), 
        .B2(n16478), .ZN(n16484) );
  INV_X1 U19553 ( .A(n16479), .ZN(n16482) );
  AOI222_X1 U19554 ( .A1(n16482), .A2(n16503), .B1(n19337), .B2(n16481), .C1(
        n16502), .C2(n16480), .ZN(n16483) );
  OAI211_X1 U19555 ( .C1(n16485), .C2(n16506), .A(n16484), .B(n16483), .ZN(
        P2_U3005) );
  AOI22_X1 U19556 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19172), .B1(n16496), 
        .B2(n16486), .ZN(n16493) );
  NOR2_X1 U19557 ( .A1(n16487), .A2(n19332), .ZN(n16491) );
  OAI22_X1 U19558 ( .A1(n16489), .A2(n19333), .B1(n14136), .B2(n16488), .ZN(
        n16490) );
  AOI21_X1 U19559 ( .B1(n16491), .B2(n15974), .A(n16490), .ZN(n16492) );
  OAI211_X1 U19560 ( .C1(n16494), .C2(n16506), .A(n16493), .B(n16492), .ZN(
        P2_U3007) );
  AOI22_X1 U19561 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19172), .B1(n16496), 
        .B2(n16495), .ZN(n16505) );
  NAND2_X1 U19562 ( .A1(n11040), .A2(n16497), .ZN(n16499) );
  XNOR2_X1 U19563 ( .A(n16499), .B(n16498), .ZN(n16567) );
  XOR2_X1 U19564 ( .A(n16500), .B(n16501), .Z(n16562) );
  AOI222_X1 U19565 ( .A1(n16567), .A2(n16503), .B1(n19337), .B2(n16564), .C1(
        n16502), .C2(n16562), .ZN(n16504) );
  OAI211_X1 U19566 ( .C1(n16507), .C2(n16506), .A(n16505), .B(n16504), .ZN(
        P2_U3009) );
  NOR2_X1 U19567 ( .A1(n16509), .A2(n16508), .ZN(n16510) );
  NOR2_X1 U19568 ( .A1(n16510), .A2(n14043), .ZN(n19238) );
  NAND2_X1 U19569 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19172), .ZN(n16511) );
  OAI21_X1 U19570 ( .B1(n16512), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16511), .ZN(n16516) );
  NOR2_X1 U19571 ( .A1(n16514), .A2(n16513), .ZN(n16515) );
  AOI211_X1 U19572 ( .C1(n16558), .C2(n19238), .A(n16516), .B(n16515), .ZN(
        n16519) );
  AOI22_X1 U19573 ( .A1(n16517), .A2(n16566), .B1(n16565), .B2(n19128), .ZN(
        n16518) );
  OAI211_X1 U19574 ( .C1(n16520), .C2(n16552), .A(n16519), .B(n16518), .ZN(
        P2_U3031) );
  AOI21_X1 U19575 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16521), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16528) );
  INV_X1 U19576 ( .A(n19244), .ZN(n16522) );
  AOI22_X1 U19577 ( .A1(n16558), .A2(n16522), .B1(n19328), .B2(
        P2_REIP_REG_13__SCAN_IN), .ZN(n16527) );
  AOI222_X1 U19578 ( .A1(n16525), .A2(n16566), .B1(n16563), .B2(n16524), .C1(
        n16565), .C2(n16523), .ZN(n16526) );
  OAI211_X1 U19579 ( .C1(n16529), .C2(n16528), .A(n16527), .B(n16526), .ZN(
        P2_U3033) );
  AOI22_X1 U19580 ( .A1(n16531), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16558), .B2(n16530), .ZN(n16540) );
  AOI222_X1 U19581 ( .A1(n16534), .A2(n16563), .B1(n16565), .B2(n16533), .C1(
        n16566), .C2(n16532), .ZN(n16539) );
  NAND2_X1 U19582 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19172), .ZN(n16538) );
  OAI211_X1 U19583 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16536), .B(n16535), .ZN(
        n16537) );
  NAND4_X1 U19584 ( .A1(n16540), .A2(n16539), .A3(n16538), .A4(n16537), .ZN(
        P2_U3035) );
  AOI211_X1 U19585 ( .C1(n16543), .C2(n16545), .A(n16542), .B(n16541), .ZN(
        n16548) );
  OAI22_X1 U19586 ( .A1(n16546), .A2(n16545), .B1(n16544), .B2(n19180), .ZN(
        n16547) );
  AOI211_X1 U19587 ( .C1(n19328), .C2(P2_REIP_REG_8__SCAN_IN), .A(n16548), .B(
        n16547), .ZN(n16551) );
  AOI22_X1 U19588 ( .A1(n16549), .A2(n16566), .B1(n16565), .B2(n19176), .ZN(
        n16550) );
  OAI211_X1 U19589 ( .C1(n16553), .C2(n16552), .A(n16551), .B(n16550), .ZN(
        P2_U3038) );
  AOI211_X1 U19590 ( .C1(n16556), .C2(n16570), .A(n16555), .B(n16554), .ZN(
        n16561) );
  INV_X1 U19591 ( .A(n19251), .ZN(n16557) );
  NAND2_X1 U19592 ( .A1(n16558), .A2(n16557), .ZN(n16559) );
  OAI21_X1 U19593 ( .B1(n19924), .B2(n19181), .A(n16559), .ZN(n16560) );
  NOR2_X1 U19594 ( .A1(n16561), .A2(n16560), .ZN(n16569) );
  AOI222_X1 U19595 ( .A1(n16567), .A2(n16566), .B1(n16565), .B2(n16564), .C1(
        n16563), .C2(n16562), .ZN(n16568) );
  OAI211_X1 U19596 ( .C1(n16571), .C2(n16570), .A(n16569), .B(n16568), .ZN(
        P2_U3041) );
  INV_X1 U19597 ( .A(n19894), .ZN(n19892) );
  OR2_X1 U19598 ( .A1(n16572), .A2(n20039), .ZN(n20013) );
  NAND2_X1 U19599 ( .A1(n19892), .A2(n20013), .ZN(n16575) );
  AOI211_X1 U19600 ( .C1(P2_STATE2_REG_0__SCAN_IN), .C2(n16575), .A(n16574), 
        .B(n16573), .ZN(n16579) );
  OAI21_X1 U19601 ( .B1(n16576), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n20038), 
        .ZN(n16577) );
  OAI21_X1 U19602 ( .B1(n19892), .B2(n20046), .A(n16577), .ZN(n16578) );
  OAI211_X1 U19603 ( .C1(n16581), .C2(n16580), .A(n16579), .B(n16578), .ZN(
        P2_U3176) );
  AOI21_X1 U19604 ( .B1(n10020), .B2(n18738), .A(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16582) );
  INV_X1 U19605 ( .A(n16582), .ZN(n16583) );
  AOI22_X1 U19606 ( .A1(n9828), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n16584), 
        .B2(n16583), .ZN(n16596) );
  AOI211_X1 U19607 ( .C1(n9871), .C2(n16586), .A(n16585), .B(n18036), .ZN(
        n16587) );
  AOI21_X1 U19608 ( .B1(n17926), .B2(n16588), .A(n16587), .ZN(n16595) );
  INV_X1 U19609 ( .A(n16589), .ZN(n16590) );
  OAI211_X1 U19610 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16603), .A(
        n17943), .B(n16590), .ZN(n16594) );
  AOI21_X1 U19611 ( .B1(n16763), .B2(n16740), .A(n16591), .ZN(n16762) );
  OAI21_X1 U19612 ( .B1(n16592), .B2(n17890), .A(n16762), .ZN(n16593) );
  NAND4_X1 U19613 ( .A1(n16596), .A2(n16595), .A3(n16594), .A4(n16593), .ZN(
        P3_U2801) );
  NAND2_X1 U19614 ( .A1(n16598), .A2(n16597), .ZN(n17665) );
  OAI221_X1 U19615 ( .B1(n9969), .B2(n16599), .C1(n9969), .C2(n17665), .A(
        n18250), .ZN(n16612) );
  OAI211_X1 U19616 ( .C1(n16601), .C2(n17680), .A(n18791), .B(n16600), .ZN(
        n16602) );
  OAI22_X1 U19617 ( .A1(n16603), .A2(n18226), .B1(n17664), .B2(n16602), .ZN(
        n16607) );
  OAI21_X1 U19618 ( .B1(n16605), .B2(n18225), .A(n16604), .ZN(n16606) );
  OAI211_X1 U19619 ( .C1(n16607), .C2(n16606), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18345), .ZN(n16611) );
  NAND2_X1 U19620 ( .A1(n9828), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17670) );
  AOI22_X1 U19621 ( .A1(n18790), .A2(n18224), .B1(n18227), .B2(n18044), .ZN(
        n18146) );
  OAI21_X1 U19622 ( .B1(n18809), .B2(n18991), .A(n18802), .ZN(n18318) );
  AOI21_X1 U19623 ( .B1(n18159), .B2(n18318), .A(n16608), .ZN(n18070) );
  OAI21_X1 U19624 ( .B1(n18146), .B2(n18147), .A(n18070), .ZN(n18106) );
  NAND3_X1 U19625 ( .A1(n18326), .A2(n17770), .A3(n18106), .ZN(n18138) );
  NOR2_X1 U19626 ( .A1(n16609), .A2(n18138), .ZN(n18087) );
  NAND3_X1 U19627 ( .A1(n17662), .A2(n18087), .A3(n17661), .ZN(n16610) );
  NAND4_X1 U19628 ( .A1(n16612), .A2(n16611), .A3(n17670), .A4(n16610), .ZN(
        P3_U2834) );
  NOR3_X1 U19629 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16614) );
  NOR4_X1 U19630 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16613) );
  NAND4_X1 U19631 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16614), .A3(n16613), .A4(
        U215), .ZN(U213) );
  INV_X1 U19632 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16706) );
  INV_X1 U19633 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16707) );
  OAI222_X1 U19634 ( .A1(U212), .A2(n16706), .B1(n16670), .B2(n16616), .C1(
        U214), .C2(n16707), .ZN(U216) );
  INV_X1 U19635 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16618) );
  AOI22_X1 U19636 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16655), .ZN(n16617) );
  OAI21_X1 U19637 ( .B1(n16618), .B2(n16670), .A(n16617), .ZN(U217) );
  AOI22_X1 U19638 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16655), .ZN(n16619) );
  OAI21_X1 U19639 ( .B1(n16620), .B2(n16670), .A(n16619), .ZN(U218) );
  INV_X1 U19640 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n19371) );
  AOI22_X1 U19641 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16655), .ZN(n16621) );
  OAI21_X1 U19642 ( .B1(n19371), .B2(n16670), .A(n16621), .ZN(U219) );
  AOI22_X1 U19643 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16655), .ZN(n16622) );
  OAI21_X1 U19644 ( .B1(n19366), .B2(n16670), .A(n16622), .ZN(U220) );
  INV_X1 U19645 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16624) );
  AOI22_X1 U19646 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16655), .ZN(n16623) );
  OAI21_X1 U19647 ( .B1(n16624), .B2(n16670), .A(n16623), .ZN(U221) );
  AOI22_X1 U19648 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16655), .ZN(n16625) );
  OAI21_X1 U19649 ( .B1(n16626), .B2(n16670), .A(n16625), .ZN(U222) );
  INV_X1 U19650 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16628) );
  AOI22_X1 U19651 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16655), .ZN(n16627) );
  OAI21_X1 U19652 ( .B1(n16628), .B2(n16670), .A(n16627), .ZN(U223) );
  AOI22_X1 U19653 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16655), .ZN(n16629) );
  OAI21_X1 U19654 ( .B1(n20286), .B2(n16670), .A(n16629), .ZN(U224) );
  INV_X1 U19655 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20280) );
  AOI22_X1 U19656 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16655), .ZN(n16630) );
  OAI21_X1 U19657 ( .B1(n20280), .B2(n16670), .A(n16630), .ZN(U225) );
  AOI22_X1 U19658 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16655), .ZN(n16631) );
  OAI21_X1 U19659 ( .B1(n19380), .B2(n16670), .A(n16631), .ZN(U226) );
  INV_X1 U19660 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20272) );
  AOI22_X1 U19661 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16655), .ZN(n16632) );
  OAI21_X1 U19662 ( .B1(n20272), .B2(n16670), .A(n16632), .ZN(U227) );
  INV_X1 U19663 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20267) );
  AOI22_X1 U19664 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16655), .ZN(n16633) );
  OAI21_X1 U19665 ( .B1(n20267), .B2(n16670), .A(n16633), .ZN(U228) );
  AOI22_X1 U19666 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16655), .ZN(n16634) );
  OAI21_X1 U19667 ( .B1(n20262), .B2(n16670), .A(n16634), .ZN(U229) );
  INV_X1 U19668 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20258) );
  AOI22_X1 U19669 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16655), .ZN(n16635) );
  OAI21_X1 U19670 ( .B1(n20258), .B2(n16670), .A(n16635), .ZN(U230) );
  INV_X1 U19671 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20237) );
  AOI22_X1 U19672 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16655), .ZN(n16636) );
  OAI21_X1 U19673 ( .B1(n20237), .B2(n16670), .A(n16636), .ZN(U231) );
  INV_X1 U19674 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16638) );
  AOI22_X1 U19675 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16655), .ZN(n16637) );
  OAI21_X1 U19676 ( .B1(n16638), .B2(n16670), .A(n16637), .ZN(U232) );
  AOI22_X1 U19677 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16655), .ZN(n16639) );
  OAI21_X1 U19678 ( .B1(n16640), .B2(n16670), .A(n16639), .ZN(U233) );
  AOI22_X1 U19679 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16655), .ZN(n16641) );
  OAI21_X1 U19680 ( .B1(n16642), .B2(n16670), .A(n16641), .ZN(U234) );
  INV_X1 U19681 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16644) );
  AOI22_X1 U19682 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16655), .ZN(n16643) );
  OAI21_X1 U19683 ( .B1(n16644), .B2(n16670), .A(n16643), .ZN(U235) );
  AOI22_X1 U19684 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16655), .ZN(n16645) );
  OAI21_X1 U19685 ( .B1(n16646), .B2(n16670), .A(n16645), .ZN(U236) );
  INV_X1 U19686 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16648) );
  AOI22_X1 U19687 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16655), .ZN(n16647) );
  OAI21_X1 U19688 ( .B1(n16648), .B2(n16670), .A(n16647), .ZN(U237) );
  AOI22_X1 U19689 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16655), .ZN(n16649) );
  OAI21_X1 U19690 ( .B1(n16650), .B2(n16670), .A(n16649), .ZN(U238) );
  AOI22_X1 U19691 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16655), .ZN(n16651) );
  OAI21_X1 U19692 ( .B1(n16652), .B2(n16670), .A(n16651), .ZN(U239) );
  AOI22_X1 U19693 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16655), .ZN(n16653) );
  OAI21_X1 U19694 ( .B1(n16654), .B2(n16670), .A(n16653), .ZN(U240) );
  INV_X1 U19695 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16657) );
  AOI22_X1 U19696 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16655), .ZN(n16656) );
  OAI21_X1 U19697 ( .B1(n16657), .B2(n16670), .A(n16656), .ZN(U241) );
  INV_X1 U19698 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16659) );
  AOI22_X1 U19699 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16655), .ZN(n16658) );
  OAI21_X1 U19700 ( .B1(n16659), .B2(n16670), .A(n16658), .ZN(U242) );
  INV_X1 U19701 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16661) );
  AOI22_X1 U19702 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16655), .ZN(n16660) );
  OAI21_X1 U19703 ( .B1(n16661), .B2(n16670), .A(n16660), .ZN(U243) );
  INV_X1 U19704 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16663) );
  AOI22_X1 U19705 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16655), .ZN(n16662) );
  OAI21_X1 U19706 ( .B1(n16663), .B2(n16670), .A(n16662), .ZN(U244) );
  INV_X1 U19707 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16665) );
  AOI22_X1 U19708 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16655), .ZN(n16664) );
  OAI21_X1 U19709 ( .B1(n16665), .B2(n16670), .A(n16664), .ZN(U245) );
  INV_X1 U19710 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16667) );
  AOI22_X1 U19711 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16655), .ZN(n16666) );
  OAI21_X1 U19712 ( .B1(n16667), .B2(n16670), .A(n16666), .ZN(U246) );
  INV_X1 U19713 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16671) );
  AOI22_X1 U19714 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16668), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16655), .ZN(n16669) );
  OAI21_X1 U19715 ( .B1(n16671), .B2(n16670), .A(n16669), .ZN(U247) );
  OAI22_X1 U19716 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16704), .ZN(n16672) );
  INV_X1 U19717 ( .A(n16672), .ZN(U251) );
  OAI22_X1 U19718 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16704), .ZN(n16673) );
  INV_X1 U19719 ( .A(n16673), .ZN(U252) );
  OAI22_X1 U19720 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16704), .ZN(n16674) );
  INV_X1 U19721 ( .A(n16674), .ZN(U253) );
  OAI22_X1 U19722 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16704), .ZN(n16675) );
  INV_X1 U19723 ( .A(n16675), .ZN(U254) );
  OAI22_X1 U19724 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16704), .ZN(n16676) );
  INV_X1 U19725 ( .A(n16676), .ZN(U255) );
  OAI22_X1 U19726 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16704), .ZN(n16677) );
  INV_X1 U19727 ( .A(n16677), .ZN(U256) );
  OAI22_X1 U19728 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16704), .ZN(n16678) );
  INV_X1 U19729 ( .A(n16678), .ZN(U257) );
  OAI22_X1 U19730 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16704), .ZN(n16679) );
  INV_X1 U19731 ( .A(n16679), .ZN(U258) );
  OAI22_X1 U19732 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16704), .ZN(n16680) );
  INV_X1 U19733 ( .A(n16680), .ZN(U259) );
  OAI22_X1 U19734 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16699), .ZN(n16681) );
  INV_X1 U19735 ( .A(n16681), .ZN(U260) );
  OAI22_X1 U19736 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16699), .ZN(n16682) );
  INV_X1 U19737 ( .A(n16682), .ZN(U261) );
  OAI22_X1 U19738 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16704), .ZN(n16683) );
  INV_X1 U19739 ( .A(n16683), .ZN(U262) );
  OAI22_X1 U19740 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16704), .ZN(n16684) );
  INV_X1 U19741 ( .A(n16684), .ZN(U263) );
  OAI22_X1 U19742 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16704), .ZN(n16685) );
  INV_X1 U19743 ( .A(n16685), .ZN(U264) );
  OAI22_X1 U19744 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16704), .ZN(n16686) );
  INV_X1 U19745 ( .A(n16686), .ZN(U265) );
  OAI22_X1 U19746 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16699), .ZN(n16687) );
  INV_X1 U19747 ( .A(n16687), .ZN(U266) );
  OAI22_X1 U19748 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16699), .ZN(n16688) );
  INV_X1 U19749 ( .A(n16688), .ZN(U267) );
  OAI22_X1 U19750 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16699), .ZN(n16689) );
  INV_X1 U19751 ( .A(n16689), .ZN(U268) );
  OAI22_X1 U19752 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16699), .ZN(n16690) );
  INV_X1 U19753 ( .A(n16690), .ZN(U269) );
  OAI22_X1 U19754 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16699), .ZN(n16691) );
  INV_X1 U19755 ( .A(n16691), .ZN(U270) );
  OAI22_X1 U19756 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16699), .ZN(n16692) );
  INV_X1 U19757 ( .A(n16692), .ZN(U271) );
  OAI22_X1 U19758 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16704), .ZN(n16693) );
  INV_X1 U19759 ( .A(n16693), .ZN(U272) );
  OAI22_X1 U19760 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16704), .ZN(n16694) );
  INV_X1 U19761 ( .A(n16694), .ZN(U273) );
  OAI22_X1 U19762 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16699), .ZN(n16695) );
  INV_X1 U19763 ( .A(n16695), .ZN(U274) );
  OAI22_X1 U19764 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16704), .ZN(n16696) );
  INV_X1 U19765 ( .A(n16696), .ZN(U275) );
  OAI22_X1 U19766 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16704), .ZN(n16697) );
  INV_X1 U19767 ( .A(n16697), .ZN(U276) );
  OAI22_X1 U19768 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16704), .ZN(n16698) );
  INV_X1 U19769 ( .A(n16698), .ZN(U277) );
  OAI22_X1 U19770 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16699), .ZN(n16700) );
  INV_X1 U19771 ( .A(n16700), .ZN(U278) );
  OAI22_X1 U19772 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16704), .ZN(n16701) );
  INV_X1 U19773 ( .A(n16701), .ZN(U279) );
  OAI22_X1 U19774 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16704), .ZN(n16702) );
  INV_X1 U19775 ( .A(n16702), .ZN(U280) );
  OAI22_X1 U19776 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16704), .ZN(n16703) );
  INV_X1 U19777 ( .A(n16703), .ZN(U281) );
  INV_X1 U19778 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18406) );
  AOI22_X1 U19779 ( .A1(n16704), .A2(n16706), .B1(n18406), .B2(U215), .ZN(U282) );
  INV_X1 U19780 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16705) );
  AOI222_X1 U19781 ( .A1(n16707), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16706), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16705), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16708) );
  INV_X1 U19782 ( .A(n16710), .ZN(n16709) );
  INV_X1 U19783 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18907) );
  INV_X1 U19784 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19934) );
  AOI22_X1 U19785 ( .A1(n16709), .A2(n18907), .B1(n19934), .B2(n16710), .ZN(
        U347) );
  INV_X1 U19786 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18905) );
  INV_X1 U19787 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19932) );
  AOI22_X1 U19788 ( .A1(n16709), .A2(n18905), .B1(n19932), .B2(n16710), .ZN(
        U348) );
  INV_X1 U19789 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18902) );
  INV_X1 U19790 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19931) );
  AOI22_X1 U19791 ( .A1(n16709), .A2(n18902), .B1(n19931), .B2(n16710), .ZN(
        U349) );
  INV_X1 U19792 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18901) );
  INV_X1 U19793 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19929) );
  AOI22_X1 U19794 ( .A1(n16709), .A2(n18901), .B1(n19929), .B2(n16710), .ZN(
        U350) );
  INV_X1 U19795 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18899) );
  INV_X1 U19796 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19927) );
  AOI22_X1 U19797 ( .A1(n16709), .A2(n18899), .B1(n19927), .B2(n16710), .ZN(
        U351) );
  INV_X1 U19798 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18897) );
  INV_X1 U19799 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19925) );
  AOI22_X1 U19800 ( .A1(n16709), .A2(n18897), .B1(n19925), .B2(n16710), .ZN(
        U352) );
  INV_X1 U19801 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18895) );
  INV_X1 U19802 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19923) );
  AOI22_X1 U19803 ( .A1(n16709), .A2(n18895), .B1(n19923), .B2(n16710), .ZN(
        U353) );
  INV_X1 U19804 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18893) );
  AOI22_X1 U19805 ( .A1(n16709), .A2(n18893), .B1(n19921), .B2(n16710), .ZN(
        U354) );
  INV_X1 U19806 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18946) );
  INV_X1 U19807 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19971) );
  AOI22_X1 U19808 ( .A1(n16709), .A2(n18946), .B1(n19971), .B2(n16710), .ZN(
        U356) );
  INV_X1 U19809 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18942) );
  INV_X1 U19810 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19969) );
  AOI22_X1 U19811 ( .A1(n16709), .A2(n18942), .B1(n19969), .B2(n16710), .ZN(
        U357) );
  INV_X1 U19812 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18941) );
  INV_X1 U19813 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19966) );
  AOI22_X1 U19814 ( .A1(n16709), .A2(n18941), .B1(n19966), .B2(n16710), .ZN(
        U358) );
  INV_X1 U19815 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18939) );
  INV_X1 U19816 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19965) );
  AOI22_X1 U19817 ( .A1(n16709), .A2(n18939), .B1(n19965), .B2(n16710), .ZN(
        U359) );
  INV_X1 U19818 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18937) );
  INV_X1 U19819 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19963) );
  AOI22_X1 U19820 ( .A1(n16709), .A2(n18937), .B1(n19963), .B2(n16710), .ZN(
        U360) );
  INV_X1 U19821 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18935) );
  INV_X1 U19822 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19961) );
  AOI22_X1 U19823 ( .A1(n16709), .A2(n18935), .B1(n19961), .B2(n16710), .ZN(
        U361) );
  INV_X1 U19824 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18932) );
  INV_X1 U19825 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19959) );
  AOI22_X1 U19826 ( .A1(n16709), .A2(n18932), .B1(n19959), .B2(n16710), .ZN(
        U362) );
  INV_X1 U19827 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18931) );
  INV_X1 U19828 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19957) );
  AOI22_X1 U19829 ( .A1(n16709), .A2(n18931), .B1(n19957), .B2(n16710), .ZN(
        U363) );
  INV_X1 U19830 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18929) );
  INV_X1 U19831 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19955) );
  AOI22_X1 U19832 ( .A1(n16709), .A2(n18929), .B1(n19955), .B2(n16710), .ZN(
        U364) );
  INV_X1 U19833 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18891) );
  INV_X1 U19834 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19919) );
  AOI22_X1 U19835 ( .A1(n16709), .A2(n18891), .B1(n19919), .B2(n16710), .ZN(
        U365) );
  INV_X1 U19836 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18927) );
  INV_X1 U19837 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19953) );
  AOI22_X1 U19838 ( .A1(n16709), .A2(n18927), .B1(n19953), .B2(n16710), .ZN(
        U366) );
  INV_X1 U19839 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18925) );
  INV_X1 U19840 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19951) );
  AOI22_X1 U19841 ( .A1(n16709), .A2(n18925), .B1(n19951), .B2(n16710), .ZN(
        U367) );
  INV_X1 U19842 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18923) );
  INV_X1 U19843 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19949) );
  AOI22_X1 U19844 ( .A1(n16709), .A2(n18923), .B1(n19949), .B2(n16710), .ZN(
        U368) );
  INV_X1 U19845 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18920) );
  INV_X1 U19846 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19947) );
  AOI22_X1 U19847 ( .A1(n16709), .A2(n18920), .B1(n19947), .B2(n16710), .ZN(
        U369) );
  INV_X1 U19848 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18919) );
  INV_X1 U19849 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19945) );
  AOI22_X1 U19850 ( .A1(n16709), .A2(n18919), .B1(n19945), .B2(n16710), .ZN(
        U370) );
  INV_X1 U19851 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18917) );
  INV_X1 U19852 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19943) );
  AOI22_X1 U19853 ( .A1(n16709), .A2(n18917), .B1(n19943), .B2(n16710), .ZN(
        U371) );
  INV_X1 U19854 ( .A(n16710), .ZN(n21320) );
  INV_X1 U19855 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18914) );
  INV_X1 U19856 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19941) );
  AOI22_X1 U19857 ( .A1(n21320), .A2(n18914), .B1(n19941), .B2(n16710), .ZN(
        U372) );
  INV_X1 U19858 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18913) );
  INV_X1 U19859 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19939) );
  AOI22_X1 U19860 ( .A1(n21320), .A2(n18913), .B1(n19939), .B2(n16710), .ZN(
        U373) );
  INV_X1 U19861 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18911) );
  INV_X1 U19862 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19937) );
  AOI22_X1 U19863 ( .A1(n21320), .A2(n18911), .B1(n19937), .B2(n16710), .ZN(
        U374) );
  INV_X1 U19864 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18909) );
  INV_X1 U19865 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19935) );
  AOI22_X1 U19866 ( .A1(n21320), .A2(n18909), .B1(n19935), .B2(n16710), .ZN(
        U375) );
  INV_X1 U19867 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18889) );
  INV_X1 U19868 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19918) );
  AOI22_X1 U19869 ( .A1(n21320), .A2(n18889), .B1(n19918), .B2(n16710), .ZN(
        U376) );
  INV_X1 U19870 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18873) );
  NOR2_X1 U19871 ( .A1(n18873), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18878) );
  OAI22_X1 U19872 ( .A1(n18886), .A2(n18878), .B1(n18873), .B2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18871) );
  INV_X1 U19873 ( .A(n18871), .ZN(n18960) );
  AOI21_X1 U19874 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18960), .ZN(n16711) );
  INV_X1 U19875 ( .A(n16711), .ZN(P3_U2633) );
  OAI21_X1 U19876 ( .B1(n16718), .B2(n16712), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16713) );
  OAI21_X1 U19877 ( .B1(n16714), .B2(n18862), .A(n16713), .ZN(P3_U2634) );
  INV_X1 U19878 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18888) );
  AOI21_X1 U19879 ( .B1(n18886), .B2(n18888), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16715) );
  AOI22_X1 U19880 ( .A1(n18955), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16715), 
        .B2(n19023), .ZN(P3_U2635) );
  NOR2_X1 U19881 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18874) );
  OAI21_X1 U19882 ( .B1(n18874), .B2(BS16), .A(n18960), .ZN(n18958) );
  OAI21_X1 U19883 ( .B1(n18960), .B2(n19013), .A(n18958), .ZN(P3_U2636) );
  INV_X1 U19884 ( .A(n16716), .ZN(n16717) );
  NOR3_X1 U19885 ( .A1(n16718), .A2(n16717), .A3(n18793), .ZN(n18840) );
  NOR2_X1 U19886 ( .A1(n18840), .A2(n18856), .ZN(n19006) );
  OAI21_X1 U19887 ( .B1(n19006), .B2(n18356), .A(n16719), .ZN(P3_U2637) );
  NOR4_X1 U19888 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16723) );
  NOR4_X1 U19889 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16722) );
  NOR4_X1 U19890 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16721) );
  NOR4_X1 U19891 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16720) );
  NAND4_X1 U19892 ( .A1(n16723), .A2(n16722), .A3(n16721), .A4(n16720), .ZN(
        n16729) );
  NOR4_X1 U19893 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16727) );
  AOI211_X1 U19894 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16726) );
  NOR4_X1 U19895 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16725) );
  NOR4_X1 U19896 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16724) );
  NAND4_X1 U19897 ( .A1(n16727), .A2(n16726), .A3(n16725), .A4(n16724), .ZN(
        n16728) );
  NOR2_X1 U19898 ( .A1(n16729), .A2(n16728), .ZN(n19000) );
  INV_X1 U19899 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16731) );
  NOR3_X1 U19900 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16732) );
  OAI21_X1 U19901 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16732), .A(n19000), .ZN(
        n16730) );
  OAI21_X1 U19902 ( .B1(n19000), .B2(n16731), .A(n16730), .ZN(P3_U2638) );
  INV_X1 U19903 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18996) );
  INV_X1 U19904 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18959) );
  AOI21_X1 U19905 ( .B1(n18996), .B2(n18959), .A(n16732), .ZN(n16734) );
  INV_X1 U19906 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16733) );
  INV_X1 U19907 ( .A(n19000), .ZN(n19003) );
  AOI22_X1 U19908 ( .A1(n19000), .A2(n16734), .B1(n16733), .B2(n19003), .ZN(
        P3_U2639) );
  INV_X1 U19909 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16786) );
  NAND2_X1 U19910 ( .A1(n16787), .A2(n16786), .ZN(n16785) );
  NOR2_X1 U19911 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16785), .ZN(n16773) );
  INV_X1 U19912 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17138) );
  NAND2_X1 U19913 ( .A1(n16773), .A2(n17138), .ZN(n16753) );
  NOR2_X1 U19914 ( .A1(n17091), .A2(n16753), .ZN(n16757) );
  INV_X1 U19915 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17107) );
  AOI22_X1 U19916 ( .A1(n17078), .A2(P3_EBX_REG_31__SCAN_IN), .B1(n16757), 
        .B2(n17107), .ZN(n16748) );
  INV_X1 U19917 ( .A(n16735), .ZN(n16799) );
  NAND3_X1 U19918 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n16799), .ZN(n16793) );
  NAND4_X1 U19919 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16780), .ZN(n16739) );
  NOR2_X1 U19920 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16739), .ZN(n16756) );
  INV_X1 U19921 ( .A(n16756), .ZN(n16738) );
  NAND3_X1 U19922 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16737) );
  OAI21_X1 U19923 ( .B1(n16737), .B2(n16736), .A(n17092), .ZN(n16769) );
  AOI21_X1 U19924 ( .B1(n16738), .B2(n16769), .A(n18948), .ZN(n16746) );
  NOR3_X1 U19925 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18950), .A3(n16739), 
        .ZN(n16745) );
  NOR2_X1 U19926 ( .A1(n10071), .A2(n16742), .ZN(n16741) );
  OAI21_X1 U19927 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16741), .A(
        n16740), .ZN(n17672) );
  INV_X1 U19928 ( .A(n17672), .ZN(n16772) );
  AOI21_X1 U19929 ( .B1(n10071), .B2(n16742), .A(n16741), .ZN(n17684) );
  NOR2_X1 U19930 ( .A1(n16743), .A2(n17047), .ZN(n16784) );
  NAND2_X1 U19931 ( .A1(n16960), .A2(n17069), .ZN(n17081) );
  NOR3_X1 U19932 ( .A1(n16750), .A2(n16752), .A3(n17081), .ZN(n16744) );
  OAI211_X1 U19933 ( .C1(n16749), .C2(n17080), .A(n16748), .B(n16747), .ZN(
        P3_U2640) );
  NAND2_X1 U19934 ( .A1(n17056), .A2(n16753), .ZN(n16764) );
  OAI22_X1 U19935 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16764), .B1(n16754), 
        .B2(n17080), .ZN(n16755) );
  OAI21_X1 U19936 ( .B1(n17078), .B2(n16757), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16758) );
  NAND3_X1 U19937 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16780), .ZN(n16770) );
  INV_X1 U19938 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18945) );
  INV_X1 U19939 ( .A(n16759), .ZN(n16760) );
  AOI211_X1 U19940 ( .C1(n16762), .C2(n16761), .A(n16760), .B(n18866), .ZN(
        n16767) );
  NOR2_X1 U19941 ( .A1(n16773), .A2(n17138), .ZN(n16765) );
  OAI22_X1 U19942 ( .A1(n16765), .A2(n16764), .B1(n16763), .B2(n17080), .ZN(
        n16766) );
  AOI211_X1 U19943 ( .C1(n17078), .C2(P3_EBX_REG_29__SCAN_IN), .A(n16767), .B(
        n16766), .ZN(n16768) );
  OAI221_X1 U19944 ( .B1(P3_REIP_REG_29__SCAN_IN), .B2(n16770), .C1(n18945), 
        .C2(n16769), .A(n16768), .ZN(P3_U2642) );
  INV_X1 U19945 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18943) );
  AOI211_X1 U19946 ( .C1(n16772), .C2(n10005), .A(n16771), .B(n18866), .ZN(
        n16778) );
  AOI211_X1 U19947 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16785), .A(n16773), .B(
        n17091), .ZN(n16777) );
  OAI22_X1 U19948 ( .A1(n16775), .A2(n17080), .B1(n16774), .B2(n17090), .ZN(
        n16776) );
  NOR3_X1 U19949 ( .A1(n16778), .A2(n16777), .A3(n16776), .ZN(n16782) );
  NAND2_X1 U19950 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16779) );
  OAI211_X1 U19951 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16780), .B(n16779), .ZN(n16781) );
  OAI211_X1 U19952 ( .C1(n18943), .C2(n16792), .A(n16782), .B(n16781), .ZN(
        P3_U2643) );
  INV_X1 U19953 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18940) );
  AOI211_X1 U19954 ( .C1(n17684), .C2(n16784), .A(n16783), .B(n18866), .ZN(
        n16790) );
  OAI211_X1 U19955 ( .C1(n16787), .C2(n16786), .A(n17056), .B(n16785), .ZN(
        n16788) );
  OAI21_X1 U19956 ( .B1(n17080), .B2(n10071), .A(n16788), .ZN(n16789) );
  AOI211_X1 U19957 ( .C1(n17078), .C2(P3_EBX_REG_27__SCAN_IN), .A(n16790), .B(
        n16789), .ZN(n16791) );
  OAI221_X1 U19958 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16793), .C1(n18940), 
        .C2(n16792), .A(n16791), .ZN(P3_U2644) );
  AOI22_X1 U19959 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17043), .B1(
        P3_EBX_REG_25__SCAN_IN), .B2(n17078), .ZN(n16804) );
  NOR2_X1 U19960 ( .A1(n16923), .A2(n16794), .ZN(n16800) );
  AOI211_X1 U19961 ( .C1(n16797), .C2(n16796), .A(n16795), .B(n18866), .ZN(
        n16798) );
  AOI221_X1 U19962 ( .B1(n16800), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n16799), 
        .C2(n18936), .A(n16798), .ZN(n16803) );
  OAI211_X1 U19963 ( .C1(n16805), .C2(n17099), .A(n17056), .B(n16801), .ZN(
        n16802) );
  NAND3_X1 U19964 ( .A1(n16804), .A2(n16803), .A3(n16802), .ZN(P3_U2646) );
  AOI211_X1 U19965 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16820), .A(n16805), .B(
        n17091), .ZN(n16806) );
  AOI21_X1 U19966 ( .B1(n17078), .B2(P3_EBX_REG_24__SCAN_IN), .A(n16806), .ZN(
        n16813) );
  AND2_X1 U19967 ( .A1(n17092), .A2(n16807), .ZN(n16819) );
  AOI211_X1 U19968 ( .C1(n17728), .C2(n16809), .A(n16808), .B(n18866), .ZN(
        n16810) );
  AOI221_X1 U19969 ( .B1(n16819), .B2(P3_REIP_REG_24__SCAN_IN), .C1(n16811), 
        .C2(n18934), .A(n16810), .ZN(n16812) );
  OAI211_X1 U19970 ( .C1(n17721), .C2(n17080), .A(n16813), .B(n16812), .ZN(
        P3_U2647) );
  AOI22_X1 U19971 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17043), .B1(
        P3_EBX_REG_23__SCAN_IN), .B2(n17078), .ZN(n16824) );
  INV_X1 U19972 ( .A(n16814), .ZN(n16818) );
  AOI211_X1 U19973 ( .C1(n17737), .C2(n16816), .A(n16815), .B(n18866), .ZN(
        n16817) );
  AOI221_X1 U19974 ( .B1(n16819), .B2(P3_REIP_REG_23__SCAN_IN), .C1(n16818), 
        .C2(n18933), .A(n16817), .ZN(n16823) );
  OAI211_X1 U19975 ( .C1(n16831), .C2(n16821), .A(n17056), .B(n16820), .ZN(
        n16822) );
  NAND3_X1 U19976 ( .A1(n16824), .A2(n16823), .A3(n16822), .ZN(P3_U2648) );
  AOI21_X1 U19977 ( .B1(n16826), .B2(n16887), .A(n16923), .ZN(n16825) );
  INV_X1 U19978 ( .A(n16825), .ZN(n16853) );
  INV_X1 U19979 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18928) );
  NAND3_X1 U19980 ( .A1(n16897), .A2(n16826), .A3(n18928), .ZN(n16843) );
  INV_X1 U19981 ( .A(n16827), .ZN(n16828) );
  AOI211_X1 U19982 ( .C1(n17752), .C2(n16829), .A(n16828), .B(n18866), .ZN(
        n16835) );
  INV_X1 U19983 ( .A(n16897), .ZN(n16911) );
  NOR3_X1 U19984 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16911), .A3(n16830), 
        .ZN(n16834) );
  AOI211_X1 U19985 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16839), .A(n16831), .B(
        n17091), .ZN(n16833) );
  INV_X1 U19986 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17102) );
  OAI22_X1 U19987 ( .A1(n17762), .A2(n17080), .B1(n17102), .B2(n17090), .ZN(
        n16832) );
  NOR4_X1 U19988 ( .A1(n16835), .A2(n16834), .A3(n16833), .A4(n16832), .ZN(
        n16836) );
  OAI221_X1 U19989 ( .B1(n18930), .B2(n16853), .C1(n18930), .C2(n16843), .A(
        n16836), .ZN(P3_U2649) );
  AOI211_X1 U19990 ( .C1(n17773), .C2(n16838), .A(n16837), .B(n18866), .ZN(
        n16842) );
  OAI211_X1 U19991 ( .C1(n16845), .C2(n17192), .A(n17056), .B(n16839), .ZN(
        n16840) );
  OAI21_X1 U19992 ( .B1(n17090), .B2(n17192), .A(n16840), .ZN(n16841) );
  AOI211_X1 U19993 ( .C1(n17043), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16842), .B(n16841), .ZN(n16844) );
  OAI211_X1 U19994 ( .C1(n16853), .C2(n18928), .A(n16844), .B(n16843), .ZN(
        P3_U2650) );
  AOI211_X1 U19995 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16856), .A(n16845), .B(
        n17091), .ZN(n16846) );
  AOI21_X1 U19996 ( .B1(n17078), .B2(P3_EBX_REG_20__SCAN_IN), .A(n16846), .ZN(
        n16852) );
  NOR4_X1 U19997 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16911), .A3(n16861), 
        .A4(n16862), .ZN(n16850) );
  AOI211_X1 U19998 ( .C1(n17781), .C2(n16848), .A(n16847), .B(n18866), .ZN(
        n16849) );
  AOI211_X1 U19999 ( .C1(n17043), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16850), .B(n16849), .ZN(n16851) );
  OAI211_X1 U20000 ( .C1(n18926), .C2(n16853), .A(n16852), .B(n16851), .ZN(
        P3_U2651) );
  AOI22_X1 U20001 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17043), .B1(
        P3_EBX_REG_19__SCAN_IN), .B2(n17078), .ZN(n16865) );
  AOI21_X1 U20002 ( .B1(n16854), .B2(n16887), .A(n16923), .ZN(n16882) );
  NAND2_X1 U20003 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17793), .ZN(
        n16868) );
  OAI21_X1 U20004 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16868), .A(
        n16960), .ZN(n16870) );
  INV_X1 U20005 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17790) );
  AOI21_X1 U20006 ( .B1(n17790), .B2(n16868), .A(n16855), .ZN(n17794) );
  XOR2_X1 U20007 ( .A(n16870), .B(n17794), .Z(n16859) );
  OAI211_X1 U20008 ( .C1(n16866), .C2(n16857), .A(n17056), .B(n16856), .ZN(
        n16858) );
  OAI21_X1 U20009 ( .B1(n16859), .B2(n18866), .A(n16858), .ZN(n16860) );
  AOI211_X1 U20010 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n16882), .A(n9828), .B(
        n16860), .ZN(n16864) );
  NOR2_X1 U20011 ( .A1(n16911), .A2(n16861), .ZN(n16872) );
  OAI211_X1 U20012 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16872), .B(n16862), .ZN(n16863) );
  NAND3_X1 U20013 ( .A1(n16865), .A2(n16864), .A3(n16863), .ZN(P3_U2652) );
  AOI211_X1 U20014 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16883), .A(n16866), .B(
        n17091), .ZN(n16867) );
  AOI21_X1 U20015 ( .B1(n17043), .B2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16867), .ZN(n16875) );
  OAI21_X1 U20016 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17793), .A(
        n16868), .ZN(n17804) );
  NAND2_X1 U20017 ( .A1(n17069), .A2(n17047), .ZN(n17060) );
  INV_X1 U20018 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17807) );
  INV_X1 U20019 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17082) );
  OAI221_X1 U20020 ( .B1(n17804), .B2(n17807), .C1(n17804), .C2(n17082), .A(
        n17069), .ZN(n16869) );
  AOI22_X1 U20021 ( .A1(n17804), .A2(n16870), .B1(n17060), .B2(n16869), .ZN(
        n16871) );
  AOI211_X1 U20022 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17078), .A(n9828), .B(
        n16871), .ZN(n16874) );
  INV_X1 U20023 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18922) );
  AOI22_X1 U20024 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16882), .B1(n16872), 
        .B2(n18922), .ZN(n16873) );
  NAND3_X1 U20025 ( .A1(n16875), .A2(n16874), .A3(n16873), .ZN(P3_U2653) );
  NAND2_X1 U20026 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16896) );
  NOR2_X1 U20027 ( .A1(n16911), .A2(n16896), .ZN(n16881) );
  NAND2_X1 U20028 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16889), .ZN(
        n16876) );
  AOI21_X1 U20029 ( .B1(n17817), .B2(n16876), .A(n17793), .ZN(n17820) );
  NOR2_X1 U20030 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18027), .ZN(
        n17070) );
  AOI21_X1 U20031 ( .B1(n16889), .B2(n17070), .A(n17047), .ZN(n16878) );
  AOI21_X1 U20032 ( .B1(n17820), .B2(n16878), .A(n18866), .ZN(n16877) );
  OAI21_X1 U20033 ( .B1(n17820), .B2(n16878), .A(n16877), .ZN(n16879) );
  OAI211_X1 U20034 ( .C1(n16884), .C2(n17090), .A(n18345), .B(n16879), .ZN(
        n16880) );
  AOI221_X1 U20035 ( .B1(n16882), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16881), 
        .C2(n18921), .A(n16880), .ZN(n16886) );
  OAI211_X1 U20036 ( .C1(n16888), .C2(n16884), .A(n17056), .B(n16883), .ZN(
        n16885) );
  OAI211_X1 U20037 ( .C1(n17080), .C2(n17817), .A(n16886), .B(n16885), .ZN(
        P3_U2654) );
  OR2_X1 U20038 ( .A1(n16923), .A2(n16887), .ZN(n16915) );
  AOI211_X1 U20039 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16902), .A(n16888), .B(
        n17091), .ZN(n16895) );
  INV_X1 U20040 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U20041 ( .A1(n16893), .A2(n16900), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16889), .ZN(n16890) );
  INV_X1 U20042 ( .A(n16890), .ZN(n17833) );
  INV_X1 U20043 ( .A(n16891), .ZN(n16904) );
  OAI221_X1 U20044 ( .B1(n16891), .B2(n17833), .C1(n16904), .C2(n16890), .A(
        n17069), .ZN(n16892) );
  OAI211_X1 U20045 ( .C1(n16893), .C2(n17080), .A(n18345), .B(n16892), .ZN(
        n16894) );
  AOI211_X1 U20046 ( .C1(n17078), .C2(P3_EBX_REG_16__SCAN_IN), .A(n16895), .B(
        n16894), .ZN(n16899) );
  OAI211_X1 U20047 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16897), .B(n16896), .ZN(n16898) );
  OAI211_X1 U20048 ( .C1(n16915), .C2(n18918), .A(n16899), .B(n16898), .ZN(
        P3_U2655) );
  OAI21_X1 U20049 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17828), .A(
        n16900), .ZN(n17838) );
  NAND2_X1 U20050 ( .A1(n16960), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16901) );
  NAND2_X1 U20051 ( .A1(n17069), .A2(n16901), .ZN(n17017) );
  AOI211_X1 U20052 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16960), .A(
        n17838), .B(n17017), .ZN(n16909) );
  INV_X1 U20053 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17841) );
  OAI211_X1 U20054 ( .C1(n16913), .C2(n16906), .A(n17056), .B(n16902), .ZN(
        n16903) );
  OAI21_X1 U20055 ( .B1(n17080), .B2(n17841), .A(n16903), .ZN(n16908) );
  NAND3_X1 U20056 ( .A1(n17069), .A2(n16904), .A3(n17838), .ZN(n16905) );
  OAI211_X1 U20057 ( .C1(n16906), .C2(n17090), .A(n18345), .B(n16905), .ZN(
        n16907) );
  NOR3_X1 U20058 ( .A1(n16909), .A2(n16908), .A3(n16907), .ZN(n16910) );
  OAI221_X1 U20059 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16911), .C1(n18916), 
        .C2(n16915), .A(n16910), .ZN(P3_U2656) );
  INV_X1 U20060 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16922) );
  NOR2_X1 U20061 ( .A1(n18027), .A2(n17866), .ZN(n17864) );
  NAND2_X1 U20062 ( .A1(n17867), .A2(n17864), .ZN(n16925) );
  AOI21_X1 U20063 ( .B1(n16922), .B2(n16925), .A(n17828), .ZN(n17853) );
  OAI21_X1 U20064 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16925), .A(
        n16960), .ZN(n16924) );
  XNOR2_X1 U20065 ( .A(n17853), .B(n16924), .ZN(n16912) );
  AOI21_X1 U20066 ( .B1(n16912), .B2(n17069), .A(n9828), .ZN(n16921) );
  AOI211_X1 U20067 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16932), .A(n16913), .B(
        n17091), .ZN(n16919) );
  INV_X1 U20068 ( .A(n16914), .ZN(n16917) );
  OAI22_X1 U20069 ( .A1(n16917), .A2(n16916), .B1(n18915), .B2(n16915), .ZN(
        n16918) );
  AOI211_X1 U20070 ( .C1(n17078), .C2(P3_EBX_REG_14__SCAN_IN), .A(n16919), .B(
        n16918), .ZN(n16920) );
  OAI211_X1 U20071 ( .C1(n16922), .C2(n17080), .A(n16921), .B(n16920), .ZN(
        P3_U2657) );
  AOI21_X1 U20072 ( .B1(n17094), .B2(n16943), .A(n16923), .ZN(n16954) );
  INV_X1 U20073 ( .A(n16954), .ZN(n16947) );
  OAI21_X1 U20074 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17084), .A(n16947), 
        .ZN(n16930) );
  NOR2_X1 U20075 ( .A1(n16924), .A2(n18866), .ZN(n16927) );
  INV_X1 U20076 ( .A(n17864), .ZN(n16949) );
  NOR2_X1 U20077 ( .A1(n17882), .A2(n16949), .ZN(n16938) );
  OAI21_X1 U20078 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16938), .A(
        n16925), .ZN(n17869) );
  AOI211_X1 U20079 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16960), .A(
        n17869), .B(n17017), .ZN(n16926) );
  AOI211_X1 U20080 ( .C1(n16927), .C2(n17869), .A(n9828), .B(n16926), .ZN(
        n16928) );
  OAI21_X1 U20081 ( .B1(n17868), .B2(n17080), .A(n16928), .ZN(n16929) );
  AOI221_X1 U20082 ( .B1(n16931), .B2(n18912), .C1(n16930), .C2(
        P3_REIP_REG_13__SCAN_IN), .A(n16929), .ZN(n16934) );
  OAI211_X1 U20083 ( .C1(n16936), .C2(n16935), .A(n17056), .B(n16932), .ZN(
        n16933) );
  OAI211_X1 U20084 ( .C1(n17090), .C2(n16935), .A(n16934), .B(n16933), .ZN(
        P3_U2658) );
  INV_X1 U20085 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18910) );
  AOI22_X1 U20086 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17043), .B1(
        P3_EBX_REG_12__SCAN_IN), .B2(n17078), .ZN(n16946) );
  NOR2_X1 U20087 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17084), .ZN(n16944) );
  AOI211_X1 U20088 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16955), .A(n16936), .B(
        n17091), .ZN(n16942) );
  INV_X1 U20089 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17911) );
  INV_X1 U20090 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17940) );
  NAND3_X1 U20091 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16937), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16998) );
  NOR2_X1 U20092 ( .A1(n17940), .A2(n16998), .ZN(n16988) );
  NAND2_X1 U20093 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16988), .ZN(
        n16972) );
  NOR2_X1 U20094 ( .A1(n17911), .A2(n16972), .ZN(n16959) );
  AND2_X1 U20095 ( .A1(n17082), .A2(n16959), .ZN(n16948) );
  AOI21_X1 U20096 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16948), .A(
        n17047), .ZN(n16939) );
  AOI21_X1 U20097 ( .B1(n17882), .B2(n16949), .A(n16938), .ZN(n17889) );
  XNOR2_X1 U20098 ( .A(n16939), .B(n17889), .ZN(n16940) );
  OAI21_X1 U20099 ( .B1(n18866), .B2(n16940), .A(n18345), .ZN(n16941) );
  AOI211_X1 U20100 ( .C1(n16944), .C2(n16943), .A(n16942), .B(n16941), .ZN(
        n16945) );
  OAI211_X1 U20101 ( .C1(n18910), .C2(n16947), .A(n16946), .B(n16945), .ZN(
        P3_U2659) );
  NOR2_X1 U20102 ( .A1(n16948), .A2(n17047), .ZN(n16950) );
  OAI21_X1 U20103 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16959), .A(
        n16949), .ZN(n17895) );
  XNOR2_X1 U20104 ( .A(n16950), .B(n17895), .ZN(n16951) );
  AOI22_X1 U20105 ( .A1(n17069), .A2(n16951), .B1(P3_EBX_REG_11__SCAN_IN), 
        .B2(n17078), .ZN(n16958) );
  INV_X1 U20106 ( .A(n16967), .ZN(n16985) );
  NAND2_X1 U20107 ( .A1(n17067), .A2(n16985), .ZN(n16966) );
  OAI21_X1 U20108 ( .B1(n16952), .B2(n16966), .A(n18908), .ZN(n16953) );
  AOI22_X1 U20109 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17043), .B1(
        n16954), .B2(n16953), .ZN(n16957) );
  OAI211_X1 U20110 ( .C1(n16962), .C2(n17297), .A(n17056), .B(n16955), .ZN(
        n16956) );
  NAND4_X1 U20111 ( .A1(n16958), .A2(n16957), .A3(n18345), .A4(n16956), .ZN(
        P3_U2660) );
  AOI21_X1 U20112 ( .B1(n17911), .B2(n16972), .A(n16959), .ZN(n17913) );
  OAI21_X1 U20113 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16972), .A(
        n16960), .ZN(n16971) );
  XNOR2_X1 U20114 ( .A(n17913), .B(n16971), .ZN(n16961) );
  AOI22_X1 U20115 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17043), .B1(
        n17069), .B2(n16961), .ZN(n16970) );
  INV_X1 U20116 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18904) );
  NOR3_X1 U20117 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18904), .A3(n16966), 
        .ZN(n16965) );
  AOI211_X1 U20118 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16963), .A(n16962), .B(
        n17091), .ZN(n16964) );
  AOI211_X1 U20119 ( .C1(n17078), .C2(P3_EBX_REG_10__SCAN_IN), .A(n16965), .B(
        n16964), .ZN(n16969) );
  NOR2_X1 U20120 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16966), .ZN(n16979) );
  AOI21_X1 U20121 ( .B1(n16967), .B2(n17067), .A(n17079), .ZN(n16984) );
  INV_X1 U20122 ( .A(n16984), .ZN(n16993) );
  OAI21_X1 U20123 ( .B1(n16979), .B2(n16993), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16968) );
  NAND4_X1 U20124 ( .A1(n16970), .A2(n16969), .A3(n18345), .A4(n16968), .ZN(
        P3_U2661) );
  INV_X1 U20125 ( .A(n16971), .ZN(n16974) );
  OAI21_X1 U20126 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16988), .A(
        n16972), .ZN(n17920) );
  NAND2_X1 U20127 ( .A1(n16937), .A2(n17070), .ZN(n16999) );
  NOR3_X1 U20128 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17936), .A3(
        n16999), .ZN(n16973) );
  AOI21_X1 U20129 ( .B1(n16974), .B2(n17920), .A(n16973), .ZN(n16975) );
  OAI22_X1 U20130 ( .A1(n16975), .A2(n18866), .B1(n17920), .B2(n17060), .ZN(
        n16976) );
  AOI211_X1 U20131 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17043), .A(
        n9828), .B(n16976), .ZN(n16983) );
  AOI21_X1 U20132 ( .B1(n17056), .B2(n16978), .A(n17078), .ZN(n16977) );
  INV_X1 U20133 ( .A(n16977), .ZN(n16981) );
  NOR2_X1 U20134 ( .A1(n16978), .A2(n17091), .ZN(n16992) );
  AOI221_X1 U20135 ( .B1(n16981), .B2(P3_EBX_REG_9__SCAN_IN), .C1(n16992), 
        .C2(n16980), .A(n16979), .ZN(n16982) );
  OAI211_X1 U20136 ( .C1(n16984), .C2(n18904), .A(n16983), .B(n16982), .ZN(
        P3_U2662) );
  NOR2_X1 U20137 ( .A1(n16985), .A2(n17084), .ZN(n16986) );
  AOI22_X1 U20138 ( .A1(n16987), .A2(n16986), .B1(P3_EBX_REG_8__SCAN_IN), .B2(
        n17078), .ZN(n16996) );
  AOI21_X1 U20139 ( .B1(n17940), .B2(n16998), .A(n16988), .ZN(n17942) );
  INV_X1 U20140 ( .A(n16937), .ZN(n17935) );
  INV_X1 U20141 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17958) );
  NOR2_X1 U20142 ( .A1(n17935), .A2(n17958), .ZN(n17937) );
  AOI21_X1 U20143 ( .B1(n17937), .B2(n17070), .A(n17047), .ZN(n16989) );
  INV_X1 U20144 ( .A(n16989), .ZN(n17001) );
  XNOR2_X1 U20145 ( .A(n17942), .B(n17001), .ZN(n16990) );
  AOI22_X1 U20146 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17043), .B1(
        n17069), .B2(n16990), .ZN(n16995) );
  NAND2_X1 U20147 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17003), .ZN(n16991) );
  AOI22_X1 U20148 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16993), .B1(n16992), 
        .B2(n16991), .ZN(n16994) );
  NAND4_X1 U20149 ( .A1(n16996), .A2(n16995), .A3(n16994), .A4(n18345), .ZN(
        P3_U2663) );
  NOR3_X1 U20150 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17084), .A3(n16997), .ZN(
        n17008) );
  NOR2_X1 U20151 ( .A1(n18027), .A2(n17960), .ZN(n17027) );
  INV_X1 U20152 ( .A(n17027), .ZN(n17011) );
  NOR2_X1 U20153 ( .A1(n17974), .A2(n17011), .ZN(n17010) );
  OAI21_X1 U20154 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17010), .A(
        n16998), .ZN(n17954) );
  INV_X1 U20155 ( .A(n16999), .ZN(n17012) );
  OAI21_X1 U20156 ( .B1(n17012), .B2(n17954), .A(n17069), .ZN(n17000) );
  AOI22_X1 U20157 ( .A1(n17954), .A2(n17001), .B1(n17060), .B2(n17000), .ZN(
        n17007) );
  OAI21_X1 U20158 ( .B1(n17002), .B2(n17084), .A(n17094), .ZN(n17024) );
  INV_X1 U20159 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18898) );
  AND3_X1 U20160 ( .A1(n18898), .A2(n17067), .A3(n17002), .ZN(n17016) );
  OAI21_X1 U20161 ( .B1(n17024), .B2(n17016), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n17005) );
  OAI211_X1 U20162 ( .C1(n17014), .C2(n17362), .A(n17056), .B(n17003), .ZN(
        n17004) );
  OAI211_X1 U20163 ( .C1(n17080), .C2(n17958), .A(n17005), .B(n17004), .ZN(
        n17006) );
  NOR4_X1 U20164 ( .A1(n9828), .A2(n17008), .A3(n17007), .A4(n17006), .ZN(
        n17009) );
  OAI21_X1 U20165 ( .B1(n17362), .B2(n17090), .A(n17009), .ZN(P3_U2664) );
  AOI21_X1 U20166 ( .B1(n17974), .B2(n17011), .A(n17010), .ZN(n17971) );
  NOR3_X1 U20167 ( .A1(n17971), .A2(n17012), .A3(n17081), .ZN(n17013) );
  AOI211_X1 U20168 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17078), .A(n9828), .B(
        n17013), .ZN(n17021) );
  AOI211_X1 U20169 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17025), .A(n17014), .B(
        n17091), .ZN(n17015) );
  AOI211_X1 U20170 ( .C1(n17043), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17016), .B(n17015), .ZN(n17020) );
  NAND2_X1 U20171 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17024), .ZN(n17019) );
  INV_X1 U20172 ( .A(n17017), .ZN(n17076) );
  OAI211_X1 U20173 ( .C1(n17027), .C2(n17047), .A(n17971), .B(n17076), .ZN(
        n17018) );
  NAND4_X1 U20174 ( .A1(n17021), .A2(n17020), .A3(n17019), .A4(n17018), .ZN(
        P3_U2665) );
  NAND2_X1 U20175 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17066) );
  NOR2_X1 U20176 ( .A1(n17084), .A2(n17066), .ZN(n17049) );
  NAND2_X1 U20177 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n17049), .ZN(n17045) );
  OAI21_X1 U20178 ( .B1(n18894), .B2(n17045), .A(n18896), .ZN(n17023) );
  INV_X1 U20179 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17028) );
  OAI22_X1 U20180 ( .A1(n17028), .A2(n17080), .B1(n17026), .B2(n17090), .ZN(
        n17022) );
  AOI21_X1 U20181 ( .B1(n17024), .B2(n17023), .A(n17022), .ZN(n17032) );
  OAI211_X1 U20182 ( .C1(n17034), .C2(n17026), .A(n17056), .B(n17025), .ZN(
        n17031) );
  NAND2_X1 U20183 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17978), .ZN(
        n17035) );
  AOI21_X1 U20184 ( .B1(n17028), .B2(n17035), .A(n17027), .ZN(n17984) );
  AOI21_X1 U20185 ( .B1(n17978), .B2(n17070), .A(n17047), .ZN(n17036) );
  AOI21_X1 U20186 ( .B1(n17984), .B2(n17036), .A(n18866), .ZN(n17029) );
  OAI21_X1 U20187 ( .B1(n17984), .B2(n17036), .A(n17029), .ZN(n17030) );
  NAND4_X1 U20188 ( .A1(n17032), .A2(n18345), .A3(n17031), .A4(n17030), .ZN(
        P3_U2666) );
  AOI21_X1 U20189 ( .B1(n17067), .B2(n17033), .A(n17079), .ZN(n17051) );
  AOI211_X1 U20190 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17055), .A(n17034), .B(
        n17091), .ZN(n17042) );
  NOR2_X1 U20191 ( .A1(n18027), .A2(n17992), .ZN(n17046) );
  OAI21_X1 U20192 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17046), .A(
        n17035), .ZN(n17995) );
  NOR2_X1 U20193 ( .A1(n18366), .A2(n19026), .ZN(n17077) );
  NOR2_X1 U20194 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17992), .ZN(
        n17998) );
  AOI22_X1 U20195 ( .A1(n17070), .A2(n17998), .B1(n17036), .B2(n17995), .ZN(
        n17038) );
  OAI22_X1 U20196 ( .A1(n17038), .A2(n18866), .B1(n17037), .B2(n17090), .ZN(
        n17039) );
  AOI221_X1 U20197 ( .B1(n17340), .B2(n17077), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n17077), .A(n17039), .ZN(
        n17040) );
  OAI211_X1 U20198 ( .C1(n17995), .C2(n17060), .A(n17040), .B(n18345), .ZN(
        n17041) );
  AOI211_X1 U20199 ( .C1(n17043), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n17042), .B(n17041), .ZN(n17044) );
  OAI221_X1 U20200 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17045), .C1(n18894), 
        .C2(n17051), .A(n17044), .ZN(P3_U2667) );
  NAND2_X1 U20201 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n17063), .ZN(
        n18798) );
  AOI21_X1 U20202 ( .B1(n18969), .B2(n18798), .A(n17340), .ZN(n18966) );
  INV_X1 U20203 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17050) );
  NAND2_X1 U20204 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17059) );
  AOI21_X1 U20205 ( .B1(n17050), .B2(n17059), .A(n17046), .ZN(n18009) );
  AOI21_X1 U20206 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17070), .A(
        n17047), .ZN(n17068) );
  OAI21_X1 U20207 ( .B1(n18009), .B2(n17068), .A(n17069), .ZN(n17048) );
  AOI21_X1 U20208 ( .B1(n18009), .B2(n17068), .A(n17048), .ZN(n17054) );
  NOR2_X1 U20209 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n17049), .ZN(n17052) );
  OAI22_X1 U20210 ( .A1(n17052), .A2(n17051), .B1(n17050), .B2(n17080), .ZN(
        n17053) );
  AOI211_X1 U20211 ( .C1(n18966), .C2(n17077), .A(n17054), .B(n17053), .ZN(
        n17058) );
  OAI211_X1 U20212 ( .C1(n17062), .C2(n17374), .A(n17056), .B(n17055), .ZN(
        n17057) );
  OAI211_X1 U20213 ( .C1(n17090), .C2(n17374), .A(n17058), .B(n17057), .ZN(
        P3_U2668) );
  INV_X1 U20214 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18890) );
  OAI21_X1 U20215 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17059), .ZN(n18017) );
  OAI22_X1 U20216 ( .A1(n18890), .A2(n17094), .B1(n18017), .B2(n17060), .ZN(
        n17061) );
  INV_X1 U20217 ( .A(n17061), .ZN(n17074) );
  INV_X1 U20218 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17396) );
  INV_X1 U20219 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17390) );
  NAND2_X1 U20220 ( .A1(n17396), .A2(n17390), .ZN(n17083) );
  AOI211_X1 U20221 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17083), .A(n17062), .B(
        n17091), .ZN(n17065) );
  INV_X1 U20222 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18020) );
  INV_X1 U20223 ( .A(n18799), .ZN(n17075) );
  NOR2_X1 U20224 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n17075), .ZN(
        n18805) );
  AOI21_X1 U20225 ( .B1(n17063), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18805), .ZN(n18975) );
  INV_X1 U20226 ( .A(n18975), .ZN(n18821) );
  INV_X1 U20227 ( .A(n17077), .ZN(n17097) );
  OAI22_X1 U20228 ( .A1(n18020), .A2(n17080), .B1(n18821), .B2(n17097), .ZN(
        n17064) );
  AOI211_X1 U20229 ( .C1(n17078), .C2(P3_EBX_REG_2__SCAN_IN), .A(n17065), .B(
        n17064), .ZN(n17073) );
  OAI211_X1 U20230 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17067), .B(n17066), .ZN(n17072) );
  OAI211_X1 U20231 ( .C1(n17070), .C2(n18017), .A(n17069), .B(n17068), .ZN(
        n17071) );
  NAND4_X1 U20232 ( .A1(n17074), .A2(n17073), .A3(n17072), .A4(n17071), .ZN(
        P3_U2669) );
  AOI21_X1 U20233 ( .B1(n18986), .B2(n18994), .A(n17075), .ZN(n18983) );
  AOI22_X1 U20234 ( .A1(n17077), .A2(n18983), .B1(n17076), .B2(n18027), .ZN(
        n17089) );
  AOI22_X1 U20235 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17079), .B1(
        P3_EBX_REG_1__SCAN_IN), .B2(n17078), .ZN(n17088) );
  OAI21_X1 U20236 ( .B1(n17082), .B2(n17081), .A(n17080), .ZN(n17086) );
  NAND2_X1 U20237 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17383) );
  NAND2_X1 U20238 ( .A1(n17083), .A2(n17383), .ZN(n17392) );
  OAI22_X1 U20239 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17084), .B1(n17091), 
        .B2(n17392), .ZN(n17085) );
  AOI21_X1 U20240 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17086), .A(
        n17085), .ZN(n17087) );
  NAND3_X1 U20241 ( .A1(n17089), .A2(n17088), .A3(n17087), .ZN(P3_U2670) );
  NAND2_X1 U20242 ( .A1(n17091), .A2(n17090), .ZN(n17093) );
  AOI22_X1 U20243 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17093), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17092), .ZN(n17096) );
  NAND3_X1 U20244 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18967), .A3(
        n17094), .ZN(n17095) );
  OAI211_X1 U20245 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17097), .A(
        n17096), .B(n17095), .ZN(P3_U2671) );
  NOR3_X1 U20246 ( .A1(n17100), .A2(n17099), .A3(n17098), .ZN(n17135) );
  INV_X1 U20247 ( .A(n17217), .ZN(n17101) );
  NAND2_X1 U20248 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17101), .ZN(n17180) );
  NOR4_X1 U20249 ( .A1(n17138), .A2(n17102), .A3(n17192), .A4(n17180), .ZN(
        n17103) );
  NAND4_X1 U20250 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n17135), .A4(n17103), .ZN(n17106) );
  NOR2_X1 U20251 ( .A1(n17107), .A2(n17106), .ZN(n17134) );
  NAND2_X1 U20252 ( .A1(n17388), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17105) );
  NAND2_X1 U20253 ( .A1(n17134), .A2(n17367), .ZN(n17104) );
  OAI22_X1 U20254 ( .A1(n17134), .A2(n17105), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17104), .ZN(P3_U2672) );
  NAND2_X1 U20255 ( .A1(n17107), .A2(n17106), .ZN(n17108) );
  NAND2_X1 U20256 ( .A1(n17108), .A2(n17388), .ZN(n17133) );
  AOI22_X1 U20257 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9814), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20258 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17340), .ZN(n17111) );
  AOI22_X1 U20259 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20260 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17109) );
  NAND4_X1 U20261 ( .A1(n17112), .A2(n17111), .A3(n17110), .A4(n17109), .ZN(
        n17119) );
  AOI22_X1 U20262 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10358), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17117) );
  AOI22_X1 U20263 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17167), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17116) );
  AOI22_X1 U20264 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17325), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17326), .ZN(n17115) );
  AOI22_X1 U20265 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n9821), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17113), .ZN(n17114) );
  NAND4_X1 U20266 ( .A1(n17117), .A2(n17116), .A3(n17115), .A4(n17114), .ZN(
        n17118) );
  NOR2_X1 U20267 ( .A1(n17119), .A2(n17118), .ZN(n17132) );
  AOI22_X1 U20268 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10358), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20269 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20270 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17120) );
  OAI21_X1 U20271 ( .B1(n17121), .B2(n17369), .A(n17120), .ZN(n17128) );
  AOI22_X1 U20272 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20273 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17125) );
  AOI22_X1 U20274 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17124) );
  AOI22_X1 U20275 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17123) );
  NAND4_X1 U20276 ( .A1(n17126), .A2(n17125), .A3(n17124), .A4(n17123), .ZN(
        n17127) );
  AOI211_X1 U20277 ( .C1(n17224), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17128), .B(n17127), .ZN(n17129) );
  NAND3_X1 U20278 ( .A1(n17131), .A2(n17130), .A3(n17129), .ZN(n17409) );
  NAND2_X1 U20279 ( .A1(n17410), .A2(n17409), .ZN(n17408) );
  XNOR2_X1 U20280 ( .A(n17132), .B(n17408), .ZN(n17407) );
  OAI22_X1 U20281 ( .A1(n17134), .A2(n17133), .B1(n17407), .B2(n17388), .ZN(
        P3_U2673) );
  INV_X1 U20282 ( .A(n17154), .ZN(n17157) );
  NAND2_X1 U20283 ( .A1(n17157), .A2(n17135), .ZN(n17139) );
  OAI211_X1 U20284 ( .C1(n17410), .C2(n17409), .A(n17394), .B(n17408), .ZN(
        n17136) );
  OAI221_X1 U20285 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n17139), .C1(n17138), 
        .C2(n17137), .A(n17136), .ZN(P3_U2674) );
  AOI21_X1 U20286 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17388), .A(n17140), .ZN(
        n17143) );
  OAI21_X1 U20287 ( .B1(n17145), .B2(n17142), .A(n17141), .ZN(n17424) );
  OAI22_X1 U20288 ( .A1(n17144), .A2(n17143), .B1(n17388), .B2(n17424), .ZN(
        P3_U2676) );
  NAND2_X1 U20289 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17157), .ZN(n17149) );
  AOI21_X1 U20290 ( .B1(n17146), .B2(n17150), .A(n17145), .ZN(n17425) );
  AOI22_X1 U20291 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17147), .B1(n17394), 
        .B2(n17425), .ZN(n17148) );
  OAI21_X1 U20292 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17149), .A(n17148), .ZN(
        P3_U2677) );
  OAI21_X1 U20293 ( .B1(n17152), .B2(n17151), .A(n17150), .ZN(n17433) );
  NAND3_X1 U20294 ( .A1(n17154), .A2(P3_EBX_REG_25__SCAN_IN), .A3(n17388), 
        .ZN(n17153) );
  OAI221_X1 U20295 ( .B1(n17154), .B2(P3_EBX_REG_25__SCAN_IN), .C1(n17388), 
        .C2(n17433), .A(n17153), .ZN(P3_U2678) );
  AOI21_X1 U20296 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17388), .A(n17163), .ZN(
        n17156) );
  XNOR2_X1 U20297 ( .A(n17155), .B(n17159), .ZN(n17438) );
  OAI22_X1 U20298 ( .A1(n17157), .A2(n17156), .B1(n17388), .B2(n17438), .ZN(
        P3_U2679) );
  INV_X1 U20299 ( .A(n17158), .ZN(n17179) );
  AOI21_X1 U20300 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17388), .A(n17179), .ZN(
        n17162) );
  OAI21_X1 U20301 ( .B1(n17161), .B2(n17160), .A(n17159), .ZN(n17443) );
  OAI22_X1 U20302 ( .A1(n17163), .A2(n17162), .B1(n17388), .B2(n17443), .ZN(
        P3_U2680) );
  AOI21_X1 U20303 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17388), .A(n17164), .ZN(
        n17178) );
  AOI22_X1 U20304 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17176) );
  AOI22_X1 U20305 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20306 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17165) );
  OAI21_X1 U20307 ( .B1(n17166), .B2(n17369), .A(n17165), .ZN(n17173) );
  AOI22_X1 U20308 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17171) );
  AOI22_X1 U20309 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17170) );
  AOI22_X1 U20310 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U20311 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17168) );
  NAND4_X1 U20312 ( .A1(n17171), .A2(n17170), .A3(n17169), .A4(n17168), .ZN(
        n17172) );
  AOI211_X1 U20313 ( .C1(n9821), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n17173), .B(n17172), .ZN(n17174) );
  NAND3_X1 U20314 ( .A1(n17176), .A2(n17175), .A3(n17174), .ZN(n17444) );
  INV_X1 U20315 ( .A(n17444), .ZN(n17177) );
  OAI22_X1 U20316 ( .A1(n17179), .A2(n17178), .B1(n17177), .B2(n17388), .ZN(
        P3_U2681) );
  NAND2_X1 U20317 ( .A1(n17388), .A2(n17180), .ZN(n17205) );
  AOI22_X1 U20318 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U20319 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U20320 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17182) );
  AOI22_X1 U20321 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17181) );
  NAND4_X1 U20322 ( .A1(n17184), .A2(n17183), .A3(n17182), .A4(n17181), .ZN(
        n17190) );
  AOI22_X1 U20323 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17188) );
  AOI22_X1 U20324 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U20325 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17186) );
  AOI22_X1 U20326 ( .A1(n9814), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17185) );
  NAND4_X1 U20327 ( .A1(n17188), .A2(n17187), .A3(n17186), .A4(n17185), .ZN(
        n17189) );
  NOR2_X1 U20328 ( .A1(n17190), .A2(n17189), .ZN(n17452) );
  OR2_X1 U20329 ( .A1(n17452), .A2(n17388), .ZN(n17191) );
  OAI221_X1 U20330 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17193), .C1(n17192), 
        .C2(n17205), .A(n17191), .ZN(P3_U2682) );
  AOI22_X1 U20331 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20332 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U20333 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17195) );
  AOI22_X1 U20334 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17194) );
  NAND4_X1 U20335 ( .A1(n17197), .A2(n17196), .A3(n17195), .A4(n17194), .ZN(
        n17203) );
  AOI22_X1 U20336 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17201) );
  AOI22_X1 U20337 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17200) );
  AOI22_X1 U20338 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17199) );
  AOI22_X1 U20339 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17198) );
  NAND4_X1 U20340 ( .A1(n17201), .A2(n17200), .A3(n17199), .A4(n17198), .ZN(
        n17202) );
  NOR2_X1 U20341 ( .A1(n17203), .A2(n17202), .ZN(n17459) );
  NOR2_X1 U20342 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17204), .ZN(n17206) );
  OAI22_X1 U20343 ( .A1(n17459), .A2(n17388), .B1(n17206), .B2(n17205), .ZN(
        P3_U2683) );
  AOI22_X1 U20344 ( .A1(n9814), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20345 ( .A1(n10358), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20346 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20347 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17207) );
  NAND4_X1 U20348 ( .A1(n17210), .A2(n17209), .A3(n17208), .A4(n17207), .ZN(
        n17216) );
  AOI22_X1 U20349 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U20350 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17213) );
  AOI22_X1 U20351 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20352 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17211) );
  NAND4_X1 U20353 ( .A1(n17214), .A2(n17213), .A3(n17212), .A4(n17211), .ZN(
        n17215) );
  NOR2_X1 U20354 ( .A1(n17216), .A2(n17215), .ZN(n17464) );
  OAI21_X1 U20355 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17232), .A(n17217), .ZN(
        n17218) );
  AOI22_X1 U20356 ( .A1(n17394), .A2(n17464), .B1(n17218), .B2(n17388), .ZN(
        P3_U2684) );
  NOR2_X1 U20357 ( .A1(n18402), .A2(n17219), .ZN(n17244) );
  AOI21_X1 U20358 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17388), .A(n17244), .ZN(
        n17231) );
  AOI22_X1 U20359 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20360 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20361 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20362 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17220) );
  NAND4_X1 U20363 ( .A1(n17223), .A2(n17222), .A3(n17221), .A4(n17220), .ZN(
        n17230) );
  AOI22_X1 U20364 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20365 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U20366 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20367 ( .A1(n17347), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17225) );
  NAND4_X1 U20368 ( .A1(n17228), .A2(n17227), .A3(n17226), .A4(n17225), .ZN(
        n17229) );
  NOR2_X1 U20369 ( .A1(n17230), .A2(n17229), .ZN(n17468) );
  OAI22_X1 U20370 ( .A1(n17232), .A2(n17231), .B1(n17468), .B2(n17388), .ZN(
        P3_U2685) );
  AOI22_X1 U20371 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10356), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20372 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U20373 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17234) );
  AOI22_X1 U20374 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17233) );
  NAND4_X1 U20375 ( .A1(n17236), .A2(n17235), .A3(n17234), .A4(n17233), .ZN(
        n17242) );
  AOI22_X1 U20376 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17240) );
  AOI22_X1 U20377 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17239) );
  AOI22_X1 U20378 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U20379 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17237) );
  NAND4_X1 U20380 ( .A1(n17240), .A2(n17239), .A3(n17238), .A4(n17237), .ZN(
        n17241) );
  NOR2_X1 U20381 ( .A1(n17242), .A2(n17241), .ZN(n17474) );
  AND2_X1 U20382 ( .A1(n17367), .A2(n17258), .ZN(n17271) );
  AOI22_X1 U20383 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17388), .B1(n17255), 
        .B2(n17271), .ZN(n17243) );
  OAI22_X1 U20384 ( .A1(n17474), .A2(n17388), .B1(n17244), .B2(n17243), .ZN(
        P3_U2686) );
  AOI22_X1 U20385 ( .A1(n10378), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U20386 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20387 ( .A1(n16071), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17246) );
  AOI22_X1 U20388 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17245) );
  NAND4_X1 U20389 ( .A1(n17248), .A2(n17247), .A3(n17246), .A4(n17245), .ZN(
        n17254) );
  AOI22_X1 U20390 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U20391 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17251) );
  AOI22_X1 U20392 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10358), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17250) );
  AOI22_X1 U20393 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17249) );
  NAND4_X1 U20394 ( .A1(n17252), .A2(n17251), .A3(n17250), .A4(n17249), .ZN(
        n17253) );
  NOR2_X1 U20395 ( .A1(n17254), .A2(n17253), .ZN(n17481) );
  AND2_X1 U20396 ( .A1(n17255), .A2(n17258), .ZN(n17257) );
  AND3_X1 U20397 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n17271), .ZN(n17270) );
  AOI21_X1 U20398 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17388), .A(n17270), .ZN(
        n17256) );
  OAI22_X1 U20399 ( .A1(n17481), .A2(n17388), .B1(n17257), .B2(n17256), .ZN(
        P3_U2687) );
  AND2_X1 U20400 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17258), .ZN(n17284) );
  OAI21_X1 U20401 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17284), .A(n17388), .ZN(
        n17269) );
  AOI22_X1 U20402 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n9813), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17347), .ZN(n17262) );
  AOI22_X1 U20403 ( .A1(n10378), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17325), .ZN(n17261) );
  AOI22_X1 U20404 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9821), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17326), .ZN(n17260) );
  AOI22_X1 U20405 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17259) );
  NAND4_X1 U20406 ( .A1(n17262), .A2(n17261), .A3(n17260), .A4(n17259), .ZN(
        n17268) );
  AOI22_X1 U20407 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17266) );
  AOI22_X1 U20408 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n17331), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17341), .ZN(n17265) );
  AOI22_X1 U20409 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17340), .ZN(n17264) );
  AOI22_X1 U20410 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n9830), .B1(n9833), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17263) );
  NAND4_X1 U20411 ( .A1(n17266), .A2(n17265), .A3(n17264), .A4(n17263), .ZN(
        n17267) );
  NOR2_X1 U20412 ( .A1(n17268), .A2(n17267), .ZN(n17485) );
  OAI22_X1 U20413 ( .A1(n17270), .A2(n17269), .B1(n17485), .B2(n17388), .ZN(
        P3_U2688) );
  OAI21_X1 U20414 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17271), .A(n17388), .ZN(
        n17283) );
  AOI22_X1 U20415 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20416 ( .A1(n10378), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17280) );
  INV_X1 U20417 ( .A(n17325), .ZN(n17345) );
  AOI22_X1 U20418 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17272) );
  OAI21_X1 U20419 ( .B1(n17345), .B2(n17369), .A(n17272), .ZN(n17278) );
  AOI22_X1 U20420 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U20421 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17275) );
  AOI22_X1 U20422 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U20423 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17273) );
  NAND4_X1 U20424 ( .A1(n17276), .A2(n17275), .A3(n17274), .A4(n17273), .ZN(
        n17277) );
  AOI211_X1 U20425 ( .C1(n17167), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n17278), .B(n17277), .ZN(n17279) );
  NAND3_X1 U20426 ( .A1(n17281), .A2(n17280), .A3(n17279), .ZN(n17491) );
  INV_X1 U20427 ( .A(n17491), .ZN(n17282) );
  OAI22_X1 U20428 ( .A1(n17284), .A2(n17283), .B1(n17282), .B2(n17388), .ZN(
        P3_U2689) );
  AOI22_X1 U20429 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17288) );
  AOI22_X1 U20430 ( .A1(n9814), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20431 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20432 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17285) );
  NAND4_X1 U20433 ( .A1(n17288), .A2(n17287), .A3(n17286), .A4(n17285), .ZN(
        n17294) );
  AOI22_X1 U20434 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U20435 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U20436 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10358), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17290) );
  AOI22_X1 U20437 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17289) );
  NAND4_X1 U20438 ( .A1(n17292), .A2(n17291), .A3(n17290), .A4(n17289), .ZN(
        n17293) );
  NOR2_X1 U20439 ( .A1(n17294), .A2(n17293), .ZN(n17500) );
  OAI211_X1 U20440 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17311), .A(n17295), .B(
        n17388), .ZN(n17296) );
  OAI21_X1 U20441 ( .B1(n17500), .B2(n17388), .A(n17296), .ZN(P3_U2691) );
  AOI21_X1 U20442 ( .B1(n17297), .B2(n17322), .A(n17394), .ZN(n17298) );
  INV_X1 U20443 ( .A(n17298), .ZN(n17310) );
  AOI22_X1 U20444 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17299), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17303) );
  AOI22_X1 U20445 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17302) );
  AOI22_X1 U20446 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U20447 ( .A1(n17325), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17300) );
  NAND4_X1 U20448 ( .A1(n17303), .A2(n17302), .A3(n17301), .A4(n17300), .ZN(
        n17309) );
  AOI22_X1 U20449 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17331), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17307) );
  AOI22_X1 U20450 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9813), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17306) );
  AOI22_X1 U20451 ( .A1(n10358), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17305) );
  AOI22_X1 U20452 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17304) );
  NAND4_X1 U20453 ( .A1(n17307), .A2(n17306), .A3(n17305), .A4(n17304), .ZN(
        n17308) );
  NOR2_X1 U20454 ( .A1(n17309), .A2(n17308), .ZN(n17505) );
  OAI22_X1 U20455 ( .A1(n17311), .A2(n17310), .B1(n17505), .B2(n17388), .ZN(
        P3_U2692) );
  AOI22_X1 U20456 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10358), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17315) );
  AOI22_X1 U20457 ( .A1(n9833), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U20458 ( .A1(n17122), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17113), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17313) );
  AOI22_X1 U20459 ( .A1(n9821), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17312) );
  NAND4_X1 U20460 ( .A1(n17315), .A2(n17314), .A3(n17313), .A4(n17312), .ZN(
        n17321) );
  AOI22_X1 U20461 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17319) );
  AOI22_X1 U20462 ( .A1(n17224), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17318) );
  AOI22_X1 U20463 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17341), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17317) );
  AOI22_X1 U20464 ( .A1(n10378), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17316) );
  NAND4_X1 U20465 ( .A1(n17319), .A2(n17318), .A3(n17317), .A4(n17316), .ZN(
        n17320) );
  NOR2_X1 U20466 ( .A1(n17321), .A2(n17320), .ZN(n17512) );
  OAI21_X1 U20467 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17339), .A(n17322), .ZN(
        n17323) );
  AOI22_X1 U20468 ( .A1(n17394), .A2(n17512), .B1(n17323), .B2(n17388), .ZN(
        P3_U2693) );
  INV_X1 U20469 ( .A(n17324), .ZN(n17360) );
  OAI21_X1 U20470 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17360), .A(n17388), .ZN(
        n17338) );
  AOI22_X1 U20471 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U20472 ( .A1(n17340), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20473 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17325), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U20474 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17326), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17327) );
  NAND4_X1 U20475 ( .A1(n17330), .A2(n17329), .A3(n17328), .A4(n17327), .ZN(
        n17337) );
  AOI22_X1 U20476 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17335) );
  AOI22_X1 U20477 ( .A1(n17331), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9814), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U20478 ( .A1(n10378), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10358), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17333) );
  AOI22_X1 U20479 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17224), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17332) );
  NAND4_X1 U20480 ( .A1(n17335), .A2(n17334), .A3(n17333), .A4(n17332), .ZN(
        n17336) );
  NOR2_X1 U20481 ( .A1(n17337), .A2(n17336), .ZN(n17515) );
  OAI22_X1 U20482 ( .A1(n17339), .A2(n17338), .B1(n17515), .B2(n17388), .ZN(
        P3_U2694) );
  AOI22_X1 U20483 ( .A1(n17367), .A2(n17366), .B1(P3_EBX_REG_8__SCAN_IN), .B2(
        n17388), .ZN(n17359) );
  AOI22_X1 U20484 ( .A1(n9835), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9833), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U20485 ( .A1(n17341), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17340), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17356) );
  AOI22_X1 U20486 ( .A1(n17342), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9821), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17343) );
  OAI21_X1 U20487 ( .B1(n17345), .B2(n17344), .A(n17343), .ZN(n17354) );
  AOI22_X1 U20488 ( .A1(n9832), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10356), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U20489 ( .A1(n17346), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17351) );
  AOI22_X1 U20490 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17347), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17350) );
  AOI22_X1 U20491 ( .A1(n10378), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17348), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17349) );
  NAND4_X1 U20492 ( .A1(n17352), .A2(n17351), .A3(n17350), .A4(n17349), .ZN(
        n17353) );
  AOI211_X1 U20493 ( .C1(n17167), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n17354), .B(n17353), .ZN(n17355) );
  NAND3_X1 U20494 ( .A1(n17357), .A2(n17356), .A3(n17355), .ZN(n17519) );
  INV_X1 U20495 ( .A(n17519), .ZN(n17358) );
  OAI22_X1 U20496 ( .A1(n17360), .A2(n17359), .B1(n17358), .B2(n17388), .ZN(
        P3_U2695) );
  AOI21_X1 U20497 ( .B1(n17362), .B2(n17361), .A(n17394), .ZN(n17363) );
  INV_X1 U20498 ( .A(n17363), .ZN(n17365) );
  OAI22_X1 U20499 ( .A1(n17366), .A2(n17365), .B1(n17364), .B2(n17388), .ZN(
        P3_U2696) );
  NAND3_X1 U20500 ( .A1(n17367), .A2(P3_EBX_REG_5__SCAN_IN), .A3(n17377), .ZN(
        n17370) );
  NAND3_X1 U20501 ( .A1(n17370), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17388), .ZN(
        n17368) );
  OAI221_X1 U20502 ( .B1(n17370), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17388), 
        .C2(n17369), .A(n17368), .ZN(P3_U2697) );
  OAI211_X1 U20503 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17377), .A(n17370), .B(
        n17388), .ZN(n17371) );
  OAI21_X1 U20504 ( .B1(n17388), .B2(n17372), .A(n17371), .ZN(P3_U2698) );
  NOR2_X1 U20505 ( .A1(n17373), .A2(n17391), .ZN(n17378) );
  INV_X1 U20506 ( .A(n17378), .ZN(n17384) );
  NOR2_X1 U20507 ( .A1(n17374), .A2(n17384), .ZN(n17381) );
  AOI21_X1 U20508 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17388), .A(n17381), .ZN(
        n17376) );
  INV_X1 U20509 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17375) );
  OAI22_X1 U20510 ( .A1(n17377), .A2(n17376), .B1(n17375), .B2(n17388), .ZN(
        P3_U2699) );
  AOI21_X1 U20511 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17388), .A(n17378), .ZN(
        n17380) );
  OAI22_X1 U20512 ( .A1(n17381), .A2(n17380), .B1(n17379), .B2(n17388), .ZN(
        P3_U2700) );
  NOR2_X1 U20513 ( .A1(n17383), .A2(n17382), .ZN(n17385) );
  OAI21_X1 U20514 ( .B1(n17385), .B2(P3_EBX_REG_2__SCAN_IN), .A(n17384), .ZN(
        n17386) );
  AOI22_X1 U20515 ( .A1(n17394), .A2(n17387), .B1(n17386), .B2(n17388), .ZN(
        P3_U2701) );
  OAI222_X1 U20516 ( .A1(n17392), .A2(n17391), .B1(n17390), .B2(n17397), .C1(
        n17389), .C2(n17388), .ZN(P3_U2702) );
  AOI22_X1 U20517 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17394), .B1(
        n17393), .B2(n17396), .ZN(n17395) );
  OAI21_X1 U20518 ( .B1(n17397), .B2(n17396), .A(n17395), .ZN(P3_U2703) );
  INV_X1 U20519 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17621) );
  INV_X1 U20520 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17617) );
  INV_X1 U20521 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17613) );
  INV_X1 U20522 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17607) );
  INV_X1 U20523 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17660) );
  INV_X1 U20524 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17639) );
  INV_X1 U20525 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17637) );
  INV_X1 U20526 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17635) );
  INV_X1 U20527 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17633) );
  NOR4_X1 U20528 ( .A1(n17639), .A2(n17637), .A3(n17635), .A4(n17633), .ZN(
        n17398) );
  NAND3_X1 U20529 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(n17398), .ZN(n17482) );
  INV_X1 U20530 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17656) );
  INV_X1 U20531 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17643) );
  NAND2_X1 U20532 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n17495) );
  NOR2_X1 U20533 ( .A1(n17643), .A2(n17495), .ZN(n17399) );
  NAND4_X1 U20534 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(n17399), .ZN(n17490) );
  NOR2_X1 U20535 ( .A1(n17656), .A2(n17490), .ZN(n17483) );
  NAND2_X1 U20536 ( .A1(n17521), .A2(n17483), .ZN(n17484) );
  INV_X1 U20537 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17605) );
  INV_X1 U20538 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17603) );
  NOR2_X1 U20539 ( .A1(n17605), .A2(n17603), .ZN(n17400) );
  NAND4_X1 U20540 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n17400), .ZN(n17450) );
  NOR3_X2 U20541 ( .A1(n17607), .A2(n17477), .A3(n17450), .ZN(n17440) );
  NAND2_X1 U20542 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17440), .ZN(n17439) );
  NOR2_X2 U20543 ( .A1(n18402), .A2(n17439), .ZN(n17435) );
  NOR2_X2 U20544 ( .A1(n17613), .A2(n17434), .ZN(n17429) );
  NOR2_X2 U20545 ( .A1(n17621), .A2(n17417), .ZN(n17411) );
  NAND2_X1 U20546 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17411), .ZN(n17404) );
  NAND3_X1 U20547 ( .A1(n17549), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n17404), 
        .ZN(n17403) );
  NAND2_X1 U20548 ( .A1(n18397), .A2(n17513), .ZN(n17451) );
  NAND2_X1 U20549 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17475), .ZN(n17402) );
  OAI211_X1 U20550 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n17404), .A(n17403), .B(
        n17402), .ZN(P3_U2704) );
  NOR2_X2 U20551 ( .A1(n18392), .A2(n17549), .ZN(n17476) );
  AOI22_X1 U20552 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17476), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17475), .ZN(n17406) );
  OAI211_X1 U20553 ( .C1(n17411), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17549), .B(
        n17404), .ZN(n17405) );
  OAI211_X1 U20554 ( .C1(n17407), .C2(n17536), .A(n17406), .B(n17405), .ZN(
        P3_U2705) );
  OAI21_X1 U20555 ( .B1(n17410), .B2(n17409), .A(n17408), .ZN(n17415) );
  AOI22_X1 U20556 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17476), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17475), .ZN(n17414) );
  AOI211_X1 U20557 ( .C1(n17621), .C2(n17417), .A(n17411), .B(n17513), .ZN(
        n17412) );
  INV_X1 U20558 ( .A(n17412), .ZN(n17413) );
  OAI211_X1 U20559 ( .C1(n17415), .C2(n17536), .A(n17414), .B(n17413), .ZN(
        P3_U2706) );
  INV_X1 U20560 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19372) );
  AOI22_X1 U20561 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17476), .B1(n17546), .B2(
        n17416), .ZN(n17419) );
  OAI211_X1 U20562 ( .C1(n17420), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17549), .B(
        n17417), .ZN(n17418) );
  OAI211_X1 U20563 ( .C1(n17451), .C2(n19372), .A(n17419), .B(n17418), .ZN(
        P3_U2707) );
  AOI22_X1 U20564 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17476), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17475), .ZN(n17423) );
  AOI211_X1 U20565 ( .C1(n17617), .C2(n17426), .A(n17420), .B(n17513), .ZN(
        n17421) );
  INV_X1 U20566 ( .A(n17421), .ZN(n17422) );
  OAI211_X1 U20567 ( .C1(n17424), .C2(n17536), .A(n17423), .B(n17422), .ZN(
        P3_U2708) );
  INV_X1 U20568 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18380) );
  AOI22_X1 U20569 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17476), .B1(n17546), .B2(
        n17425), .ZN(n17428) );
  OAI211_X1 U20570 ( .C1(n17429), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17549), .B(
        n17426), .ZN(n17427) );
  OAI211_X1 U20571 ( .C1(n17451), .C2(n18380), .A(n17428), .B(n17427), .ZN(
        P3_U2709) );
  AOI22_X1 U20572 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17476), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17475), .ZN(n17432) );
  AOI211_X1 U20573 ( .C1(n17613), .C2(n17434), .A(n17429), .B(n17513), .ZN(
        n17430) );
  INV_X1 U20574 ( .A(n17430), .ZN(n17431) );
  OAI211_X1 U20575 ( .C1(n17433), .C2(n17536), .A(n17432), .B(n17431), .ZN(
        P3_U2710) );
  AOI22_X1 U20576 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17476), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17475), .ZN(n17437) );
  OAI211_X1 U20577 ( .C1(n17435), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17549), .B(
        n17434), .ZN(n17436) );
  OAI211_X1 U20578 ( .C1(n17438), .C2(n17536), .A(n17437), .B(n17436), .ZN(
        P3_U2711) );
  AOI22_X1 U20579 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17476), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17475), .ZN(n17442) );
  OAI211_X1 U20580 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17440), .A(n17549), .B(
        n17439), .ZN(n17441) );
  OAI211_X1 U20581 ( .C1(n17443), .C2(n17536), .A(n17442), .B(n17441), .ZN(
        P3_U2712) );
  NOR2_X1 U20582 ( .A1(n18402), .A2(n17477), .ZN(n17471) );
  NAND2_X1 U20583 ( .A1(n17471), .A2(n17607), .ZN(n17449) );
  AOI22_X1 U20584 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17475), .B1(n17546), .B2(
        n17444), .ZN(n17448) );
  INV_X1 U20585 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17601) );
  INV_X1 U20586 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17597) );
  NAND2_X1 U20587 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17469), .ZN(n17465) );
  NAND2_X1 U20588 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17460), .ZN(n17456) );
  NAND2_X1 U20589 ( .A1(n17549), .A2(n17456), .ZN(n17455) );
  OAI21_X1 U20590 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17445), .A(n17455), .ZN(
        n17446) );
  AOI22_X1 U20591 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17476), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17446), .ZN(n17447) );
  OAI211_X1 U20592 ( .C1(n17450), .C2(n17449), .A(n17448), .B(n17447), .ZN(
        P3_U2713) );
  INV_X1 U20593 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n19378) );
  OAI22_X1 U20594 ( .A1(n17452), .A2(n17536), .B1(n19378), .B2(n17451), .ZN(
        n17453) );
  AOI21_X1 U20595 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17476), .A(n17453), .ZN(
        n17454) );
  OAI221_X1 U20596 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17456), .C1(n17605), 
        .C2(n17455), .A(n17454), .ZN(P3_U2714) );
  AOI22_X1 U20597 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17476), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17475), .ZN(n17458) );
  OAI211_X1 U20598 ( .C1(n17460), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17549), .B(
        n17456), .ZN(n17457) );
  OAI211_X1 U20599 ( .C1(n17459), .C2(n17536), .A(n17458), .B(n17457), .ZN(
        P3_U2715) );
  AOI22_X1 U20600 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17476), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17475), .ZN(n17463) );
  AOI211_X1 U20601 ( .C1(n17601), .C2(n17465), .A(n17460), .B(n17513), .ZN(
        n17461) );
  INV_X1 U20602 ( .A(n17461), .ZN(n17462) );
  OAI211_X1 U20603 ( .C1(n17464), .C2(n17536), .A(n17463), .B(n17462), .ZN(
        P3_U2716) );
  AOI22_X1 U20604 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17476), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17475), .ZN(n17467) );
  OAI211_X1 U20605 ( .C1(n17469), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17549), .B(
        n17465), .ZN(n17466) );
  OAI211_X1 U20606 ( .C1(n17468), .C2(n17536), .A(n17467), .B(n17466), .ZN(
        P3_U2717) );
  AOI22_X1 U20607 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17476), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17475), .ZN(n17473) );
  INV_X1 U20608 ( .A(n17469), .ZN(n17470) );
  OAI211_X1 U20609 ( .C1(n17471), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17549), .B(
        n17470), .ZN(n17472) );
  OAI211_X1 U20610 ( .C1(n17474), .C2(n17536), .A(n17473), .B(n17472), .ZN(
        P3_U2718) );
  AOI22_X1 U20611 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17476), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17475), .ZN(n17480) );
  OAI211_X1 U20612 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17478), .A(n17549), .B(
        n17477), .ZN(n17479) );
  OAI211_X1 U20613 ( .C1(n17481), .C2(n17536), .A(n17480), .B(n17479), .ZN(
        P3_U2719) );
  NOR3_X1 U20614 ( .A1(n18402), .A2(n17548), .A3(n17482), .ZN(n17526) );
  NAND2_X1 U20615 ( .A1(n17483), .A2(n17526), .ZN(n17488) );
  NAND2_X1 U20616 ( .A1(n17549), .A2(n17484), .ZN(n17493) );
  INV_X1 U20617 ( .A(n17485), .ZN(n17486) );
  AOI22_X1 U20618 ( .A1(n17546), .A2(n17486), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n17547), .ZN(n17487) );
  OAI221_X1 U20619 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17488), .C1(n17660), 
        .C2(n17493), .A(n17487), .ZN(P3_U2720) );
  INV_X1 U20620 ( .A(n17526), .ZN(n17489) );
  NOR2_X1 U20621 ( .A1(n17490), .A2(n17489), .ZN(n17498) );
  INV_X1 U20622 ( .A(n17498), .ZN(n17494) );
  AOI22_X1 U20623 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17547), .B1(n17546), .B2(
        n17491), .ZN(n17492) );
  OAI221_X1 U20624 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17494), .C1(n17656), 
        .C2(n17493), .A(n17492), .ZN(P3_U2721) );
  INV_X1 U20625 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17499) );
  INV_X1 U20626 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17645) );
  NAND2_X1 U20627 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17526), .ZN(n17520) );
  NOR2_X1 U20628 ( .A1(n17645), .A2(n17520), .ZN(n17517) );
  NAND2_X1 U20629 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17517), .ZN(n17509) );
  NOR2_X1 U20630 ( .A1(n17495), .A2(n17509), .ZN(n17502) );
  AOI21_X1 U20631 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17549), .A(n17502), .ZN(
        n17497) );
  OAI222_X1 U20632 ( .A1(n17539), .A2(n17499), .B1(n17498), .B2(n17497), .C1(
        n17536), .C2(n17496), .ZN(P3_U2722) );
  INV_X1 U20633 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17503) );
  INV_X1 U20634 ( .A(n17509), .ZN(n17504) );
  AOI22_X1 U20635 ( .A1(n17504), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n17549), .ZN(n17501) );
  OAI222_X1 U20636 ( .A1(n17539), .A2(n17503), .B1(n17502), .B2(n17501), .C1(
        n17536), .C2(n17500), .ZN(P3_U2723) );
  INV_X1 U20637 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17508) );
  INV_X1 U20638 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17649) );
  NOR2_X1 U20639 ( .A1(n17649), .A2(n17509), .ZN(n17507) );
  AOI21_X1 U20640 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17549), .A(n17504), .ZN(
        n17506) );
  OAI222_X1 U20641 ( .A1(n17539), .A2(n17508), .B1(n17507), .B2(n17506), .C1(
        n17536), .C2(n17505), .ZN(P3_U2724) );
  OAI211_X1 U20642 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17517), .A(n17549), .B(
        n17509), .ZN(n17511) );
  NAND2_X1 U20643 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17547), .ZN(n17510) );
  OAI211_X1 U20644 ( .C1(n17512), .C2(n17536), .A(n17511), .B(n17510), .ZN(
        P3_U2725) );
  INV_X1 U20645 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17518) );
  OAI21_X1 U20646 ( .B1(n17645), .B2(n17513), .A(n17520), .ZN(n17514) );
  INV_X1 U20647 ( .A(n17514), .ZN(n17516) );
  OAI222_X1 U20648 ( .A1(n17539), .A2(n17518), .B1(n17517), .B2(n17516), .C1(
        n17536), .C2(n17515), .ZN(P3_U2726) );
  AOI22_X1 U20649 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17547), .B1(n17546), .B2(
        n17519), .ZN(n17523) );
  OAI211_X1 U20650 ( .C1(n17521), .C2(P3_EAX_REG_8__SCAN_IN), .A(n17549), .B(
        n17520), .ZN(n17522) );
  NAND2_X1 U20651 ( .A1(n17523), .A2(n17522), .ZN(P3_U2727) );
  INV_X1 U20652 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17631) );
  INV_X1 U20653 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17629) );
  OR3_X1 U20654 ( .A1(n18402), .A2(n17548), .A3(n17629), .ZN(n17542) );
  NOR2_X1 U20655 ( .A1(n17631), .A2(n17542), .ZN(n17534) );
  AND2_X1 U20656 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17534), .ZN(n17538) );
  NAND2_X1 U20657 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17538), .ZN(n17527) );
  NOR2_X1 U20658 ( .A1(n17637), .A2(n17527), .ZN(n17530) );
  AOI21_X1 U20659 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17549), .A(n17530), .ZN(
        n17525) );
  OAI222_X1 U20660 ( .A1(n17539), .A2(n18404), .B1(n17526), .B2(n17525), .C1(
        n17536), .C2(n17524), .ZN(P3_U2728) );
  INV_X1 U20661 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18398) );
  INV_X1 U20662 ( .A(n17527), .ZN(n17533) );
  AOI21_X1 U20663 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17549), .A(n17533), .ZN(
        n17529) );
  OAI222_X1 U20664 ( .A1(n18398), .A2(n17539), .B1(n17530), .B2(n17529), .C1(
        n17536), .C2(n17528), .ZN(P3_U2729) );
  INV_X1 U20665 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18393) );
  AOI21_X1 U20666 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17549), .A(n17538), .ZN(
        n17532) );
  OAI222_X1 U20667 ( .A1(n18393), .A2(n17539), .B1(n17533), .B2(n17532), .C1(
        n17536), .C2(n17531), .ZN(P3_U2730) );
  INV_X1 U20668 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18388) );
  AOI21_X1 U20669 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17549), .A(n17534), .ZN(
        n17537) );
  OAI222_X1 U20670 ( .A1(n18388), .A2(n17539), .B1(n17538), .B2(n17537), .C1(
        n17536), .C2(n17535), .ZN(P3_U2731) );
  NAND2_X1 U20671 ( .A1(n17549), .A2(n17542), .ZN(n17545) );
  AOI22_X1 U20672 ( .A1(n17547), .A2(BUF2_REG_3__SCAN_IN), .B1(n17546), .B2(
        n17540), .ZN(n17541) );
  OAI221_X1 U20673 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17542), .C1(n17631), 
        .C2(n17545), .A(n17541), .ZN(P3_U2732) );
  AOI22_X1 U20674 ( .A1(n17547), .A2(BUF2_REG_2__SCAN_IN), .B1(n17546), .B2(
        n17543), .ZN(n17544) );
  OAI221_X1 U20675 ( .B1(n17545), .B2(n17548), .C1(n17545), .C2(n17629), .A(
        n17544), .ZN(P3_U2733) );
  AOI22_X1 U20676 ( .A1(n17547), .A2(BUF2_REG_1__SCAN_IN), .B1(n17546), .B2(
        n9812), .ZN(n17552) );
  OAI211_X1 U20677 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17550), .A(n17549), .B(
        n17548), .ZN(n17551) );
  NAND2_X1 U20678 ( .A1(n17552), .A2(n17551), .ZN(P3_U2734) );
  NOR2_X1 U20679 ( .A1(n18972), .A2(n18870), .ZN(n19011) );
  AND2_X1 U20680 ( .A1(n17567), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20681 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17623) );
  NAND2_X1 U20682 ( .A1(n17554), .A2(n18366), .ZN(n17571) );
  AOI22_X1 U20683 ( .A1(n19011), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17587), .ZN(n17555) );
  OAI21_X1 U20684 ( .B1(n17623), .B2(n17571), .A(n17555), .ZN(P3_U2737) );
  AOI22_X1 U20685 ( .A1(n19011), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17556) );
  OAI21_X1 U20686 ( .B1(n17621), .B2(n17571), .A(n17556), .ZN(P3_U2738) );
  INV_X1 U20687 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17619) );
  AOI22_X1 U20688 ( .A1(n19011), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17567), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17557) );
  OAI21_X1 U20689 ( .B1(n17619), .B2(n17571), .A(n17557), .ZN(P3_U2739) );
  AOI22_X1 U20690 ( .A1(n19011), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17567), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17558) );
  OAI21_X1 U20691 ( .B1(n17617), .B2(n17571), .A(n17558), .ZN(P3_U2740) );
  INV_X1 U20692 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17615) );
  AOI22_X1 U20693 ( .A1(n19011), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17559) );
  OAI21_X1 U20694 ( .B1(n17615), .B2(n17571), .A(n17559), .ZN(P3_U2741) );
  AOI22_X1 U20695 ( .A1(n19011), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17567), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17560) );
  OAI21_X1 U20696 ( .B1(n17613), .B2(n17571), .A(n17560), .ZN(P3_U2742) );
  INV_X1 U20697 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17611) );
  AOI22_X1 U20698 ( .A1(n19011), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17567), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17561) );
  OAI21_X1 U20699 ( .B1(n17611), .B2(n17571), .A(n17561), .ZN(P3_U2743) );
  INV_X1 U20700 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17609) );
  AOI22_X1 U20701 ( .A1(n17588), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17567), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17562) );
  OAI21_X1 U20702 ( .B1(n17609), .B2(n17571), .A(n17562), .ZN(P3_U2744) );
  AOI22_X1 U20703 ( .A1(n17588), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17567), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17563) );
  OAI21_X1 U20704 ( .B1(n17607), .B2(n17571), .A(n17563), .ZN(P3_U2745) );
  AOI22_X1 U20705 ( .A1(n17588), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17567), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17564) );
  OAI21_X1 U20706 ( .B1(n17605), .B2(n17571), .A(n17564), .ZN(P3_U2746) );
  AOI22_X1 U20707 ( .A1(n17588), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17567), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17565) );
  OAI21_X1 U20708 ( .B1(n17603), .B2(n17571), .A(n17565), .ZN(P3_U2747) );
  AOI22_X1 U20709 ( .A1(n17588), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17567), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17566) );
  OAI21_X1 U20710 ( .B1(n17601), .B2(n17571), .A(n17566), .ZN(P3_U2748) );
  INV_X1 U20711 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17599) );
  AOI22_X1 U20712 ( .A1(n17588), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17567), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17568) );
  OAI21_X1 U20713 ( .B1(n17599), .B2(n17571), .A(n17568), .ZN(P3_U2749) );
  AOI22_X1 U20714 ( .A1(n17588), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17569) );
  OAI21_X1 U20715 ( .B1(n17597), .B2(n17571), .A(n17569), .ZN(P3_U2750) );
  INV_X1 U20716 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17595) );
  AOI22_X1 U20717 ( .A1(n17588), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17570) );
  OAI21_X1 U20718 ( .B1(n17595), .B2(n17571), .A(n17570), .ZN(P3_U2751) );
  AOI22_X1 U20719 ( .A1(n17588), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17572) );
  OAI21_X1 U20720 ( .B1(n17660), .B2(n17590), .A(n17572), .ZN(P3_U2752) );
  AOI22_X1 U20721 ( .A1(n17588), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17573) );
  OAI21_X1 U20722 ( .B1(n17656), .B2(n17590), .A(n17573), .ZN(P3_U2753) );
  INV_X1 U20723 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17653) );
  AOI22_X1 U20724 ( .A1(n17588), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17574) );
  OAI21_X1 U20725 ( .B1(n17653), .B2(n17590), .A(n17574), .ZN(P3_U2754) );
  INV_X1 U20726 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17651) );
  AOI22_X1 U20727 ( .A1(n17588), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17575) );
  OAI21_X1 U20728 ( .B1(n17651), .B2(n17590), .A(n17575), .ZN(P3_U2755) );
  AOI22_X1 U20729 ( .A1(n17588), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17576) );
  OAI21_X1 U20730 ( .B1(n17649), .B2(n17590), .A(n17576), .ZN(P3_U2756) );
  INV_X1 U20731 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17647) );
  AOI22_X1 U20732 ( .A1(n17588), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17577) );
  OAI21_X1 U20733 ( .B1(n17647), .B2(n17590), .A(n17577), .ZN(P3_U2757) );
  AOI22_X1 U20734 ( .A1(n17588), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17578) );
  OAI21_X1 U20735 ( .B1(n17645), .B2(n17590), .A(n17578), .ZN(P3_U2758) );
  AOI22_X1 U20736 ( .A1(n17588), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17579) );
  OAI21_X1 U20737 ( .B1(n17643), .B2(n17590), .A(n17579), .ZN(P3_U2759) );
  AOI22_X1 U20738 ( .A1(n17588), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17580) );
  OAI21_X1 U20739 ( .B1(n17639), .B2(n17590), .A(n17580), .ZN(P3_U2760) );
  AOI22_X1 U20740 ( .A1(n17588), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17581) );
  OAI21_X1 U20741 ( .B1(n17637), .B2(n17590), .A(n17581), .ZN(P3_U2761) );
  AOI22_X1 U20742 ( .A1(n17588), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17582) );
  OAI21_X1 U20743 ( .B1(n17635), .B2(n17590), .A(n17582), .ZN(P3_U2762) );
  AOI22_X1 U20744 ( .A1(n17588), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17583) );
  OAI21_X1 U20745 ( .B1(n17633), .B2(n17590), .A(n17583), .ZN(P3_U2763) );
  AOI22_X1 U20746 ( .A1(n17588), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17584) );
  OAI21_X1 U20747 ( .B1(n17631), .B2(n17590), .A(n17584), .ZN(P3_U2764) );
  AOI22_X1 U20748 ( .A1(n17588), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17585) );
  OAI21_X1 U20749 ( .B1(n17629), .B2(n17590), .A(n17585), .ZN(P3_U2765) );
  INV_X1 U20750 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17627) );
  AOI22_X1 U20751 ( .A1(n17588), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17586) );
  OAI21_X1 U20752 ( .B1(n17627), .B2(n17590), .A(n17586), .ZN(P3_U2766) );
  AOI22_X1 U20753 ( .A1(n17588), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17587), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17589) );
  OAI21_X1 U20754 ( .B1(n17625), .B2(n17590), .A(n17589), .ZN(P3_U2767) );
  NAND2_X1 U20755 ( .A1(n18848), .A2(n18375), .ZN(n17592) );
  NOR2_X1 U20756 ( .A1(n17592), .A2(n17591), .ZN(n17640) );
  OAI211_X1 U20757 ( .C1(n19014), .C2(n19015), .A(n18848), .B(n17593), .ZN(
        n17654) );
  AOI22_X1 U20758 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17640), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17657), .ZN(n17594) );
  OAI21_X1 U20759 ( .B1(n17595), .B2(n17642), .A(n17594), .ZN(P3_U2768) );
  AOI22_X1 U20760 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17640), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17657), .ZN(n17596) );
  OAI21_X1 U20761 ( .B1(n17597), .B2(n17642), .A(n17596), .ZN(P3_U2769) );
  AOI22_X1 U20762 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17640), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17657), .ZN(n17598) );
  OAI21_X1 U20763 ( .B1(n17599), .B2(n17642), .A(n17598), .ZN(P3_U2770) );
  AOI22_X1 U20764 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17640), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17657), .ZN(n17600) );
  OAI21_X1 U20765 ( .B1(n17601), .B2(n17642), .A(n17600), .ZN(P3_U2771) );
  AOI22_X1 U20766 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17640), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17657), .ZN(n17602) );
  OAI21_X1 U20767 ( .B1(n17603), .B2(n17642), .A(n17602), .ZN(P3_U2772) );
  AOI22_X1 U20768 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17640), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17657), .ZN(n17604) );
  OAI21_X1 U20769 ( .B1(n17605), .B2(n17642), .A(n17604), .ZN(P3_U2773) );
  AOI22_X1 U20770 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17640), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17657), .ZN(n17606) );
  OAI21_X1 U20771 ( .B1(n17607), .B2(n17642), .A(n17606), .ZN(P3_U2774) );
  AOI22_X1 U20772 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17640), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17654), .ZN(n17608) );
  OAI21_X1 U20773 ( .B1(n17609), .B2(n17642), .A(n17608), .ZN(P3_U2775) );
  AOI22_X1 U20774 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17640), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17654), .ZN(n17610) );
  OAI21_X1 U20775 ( .B1(n17611), .B2(n17642), .A(n17610), .ZN(P3_U2776) );
  AOI22_X1 U20776 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17640), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17654), .ZN(n17612) );
  OAI21_X1 U20777 ( .B1(n17613), .B2(n17642), .A(n17612), .ZN(P3_U2777) );
  AOI22_X1 U20778 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17658), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17654), .ZN(n17614) );
  OAI21_X1 U20779 ( .B1(n17615), .B2(n17642), .A(n17614), .ZN(P3_U2778) );
  AOI22_X1 U20780 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17658), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17654), .ZN(n17616) );
  OAI21_X1 U20781 ( .B1(n17617), .B2(n17642), .A(n17616), .ZN(P3_U2779) );
  AOI22_X1 U20782 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17658), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17657), .ZN(n17618) );
  OAI21_X1 U20783 ( .B1(n17619), .B2(n17642), .A(n17618), .ZN(P3_U2780) );
  AOI22_X1 U20784 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17658), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17657), .ZN(n17620) );
  OAI21_X1 U20785 ( .B1(n17621), .B2(n17642), .A(n17620), .ZN(P3_U2781) );
  AOI22_X1 U20786 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17658), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17657), .ZN(n17622) );
  OAI21_X1 U20787 ( .B1(n17623), .B2(n17642), .A(n17622), .ZN(P3_U2782) );
  AOI22_X1 U20788 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17657), .ZN(n17624) );
  OAI21_X1 U20789 ( .B1(n17625), .B2(n17642), .A(n17624), .ZN(P3_U2783) );
  AOI22_X1 U20790 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17657), .ZN(n17626) );
  OAI21_X1 U20791 ( .B1(n17627), .B2(n17642), .A(n17626), .ZN(P3_U2784) );
  AOI22_X1 U20792 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17657), .ZN(n17628) );
  OAI21_X1 U20793 ( .B1(n17629), .B2(n17642), .A(n17628), .ZN(P3_U2785) );
  AOI22_X1 U20794 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17657), .ZN(n17630) );
  OAI21_X1 U20795 ( .B1(n17631), .B2(n17642), .A(n17630), .ZN(P3_U2786) );
  AOI22_X1 U20796 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17657), .ZN(n17632) );
  OAI21_X1 U20797 ( .B1(n17633), .B2(n17642), .A(n17632), .ZN(P3_U2787) );
  AOI22_X1 U20798 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17657), .ZN(n17634) );
  OAI21_X1 U20799 ( .B1(n17635), .B2(n17642), .A(n17634), .ZN(P3_U2788) );
  AOI22_X1 U20800 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17657), .ZN(n17636) );
  OAI21_X1 U20801 ( .B1(n17637), .B2(n17642), .A(n17636), .ZN(P3_U2789) );
  AOI22_X1 U20802 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17657), .ZN(n17638) );
  OAI21_X1 U20803 ( .B1(n17639), .B2(n17642), .A(n17638), .ZN(P3_U2790) );
  AOI22_X1 U20804 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17640), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17657), .ZN(n17641) );
  OAI21_X1 U20805 ( .B1(n17643), .B2(n17642), .A(n17641), .ZN(P3_U2791) );
  AOI22_X1 U20806 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17654), .ZN(n17644) );
  OAI21_X1 U20807 ( .B1(n17645), .B2(n17642), .A(n17644), .ZN(P3_U2792) );
  AOI22_X1 U20808 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17654), .ZN(n17646) );
  OAI21_X1 U20809 ( .B1(n17647), .B2(n17642), .A(n17646), .ZN(P3_U2793) );
  AOI22_X1 U20810 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17654), .ZN(n17648) );
  OAI21_X1 U20811 ( .B1(n17649), .B2(n17642), .A(n17648), .ZN(P3_U2794) );
  AOI22_X1 U20812 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17654), .ZN(n17650) );
  OAI21_X1 U20813 ( .B1(n17651), .B2(n17642), .A(n17650), .ZN(P3_U2795) );
  AOI22_X1 U20814 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17657), .ZN(n17652) );
  OAI21_X1 U20815 ( .B1(n17653), .B2(n17642), .A(n17652), .ZN(P3_U2796) );
  AOI22_X1 U20816 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17654), .ZN(n17655) );
  OAI21_X1 U20817 ( .B1(n17656), .B2(n17642), .A(n17655), .ZN(P3_U2797) );
  AOI22_X1 U20818 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17658), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17657), .ZN(n17659) );
  OAI21_X1 U20819 ( .B1(n17660), .B2(n17642), .A(n17659), .ZN(P3_U2798) );
  NAND2_X1 U20820 ( .A1(n17662), .A2(n17661), .ZN(n17679) );
  NAND2_X1 U20821 ( .A1(n18037), .A2(n17836), .ZN(n17740) );
  NOR2_X1 U20822 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17663), .ZN(
        n17675) );
  AOI211_X1 U20823 ( .C1(n17666), .C2(n17665), .A(n17664), .B(n17946), .ZN(
        n17674) );
  AND3_X1 U20824 ( .A1(n10071), .A2(n17791), .A3(n17667), .ZN(n17689) );
  INV_X1 U20825 ( .A(n17993), .ZN(n17749) );
  OAI21_X1 U20826 ( .B1(n17667), .B2(n17749), .A(n18032), .ZN(n17668) );
  AOI21_X1 U20827 ( .B1(n17862), .B2(n17669), .A(n17668), .ZN(n17694) );
  OAI21_X1 U20828 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17776), .A(
        n17694), .ZN(n17690) );
  OAI21_X1 U20829 ( .B1(n17689), .B2(n17690), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17671) );
  OAI211_X1 U20830 ( .C1(n17870), .C2(n17672), .A(n17671), .B(n17670), .ZN(
        n17673) );
  AOI211_X1 U20831 ( .C1(n17675), .C2(n17791), .A(n17674), .B(n17673), .ZN(
        n17678) );
  NAND2_X1 U20832 ( .A1(n17901), .A2(n18036), .ZN(n17784) );
  AOI22_X1 U20833 ( .A1(n17943), .A2(n18043), .B1(n18026), .B2(n18045), .ZN(
        n17699) );
  NAND2_X1 U20834 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17699), .ZN(
        n17676) );
  NAND3_X1 U20835 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17784), .A3(
        n17676), .ZN(n17677) );
  OAI211_X1 U20836 ( .C1(n17679), .C2(n17740), .A(n17678), .B(n17677), .ZN(
        P3_U2802) );
  NAND2_X1 U20837 ( .A1(n17681), .A2(n17680), .ZN(n17682) );
  XOR2_X1 U20838 ( .A(n17932), .B(n17682), .Z(n18056) );
  NAND2_X1 U20839 ( .A1(n17683), .A2(n17836), .ZN(n17687) );
  AOI22_X1 U20840 ( .A1(n9828), .A2(P3_REIP_REG_27__SCAN_IN), .B1(n17890), 
        .B2(n17684), .ZN(n17685) );
  OAI221_X1 U20841 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17687), 
        .C1(n17686), .C2(n17699), .A(n17685), .ZN(n17688) );
  AOI211_X1 U20842 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17690), .A(
        n17689), .B(n17688), .ZN(n17691) );
  OAI21_X1 U20843 ( .B1(n18056), .B2(n17946), .A(n17691), .ZN(P3_U2803) );
  AOI21_X1 U20844 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17693), .A(
        n17692), .ZN(n18063) );
  INV_X1 U20845 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18938) );
  NOR2_X1 U20846 ( .A1(n18345), .A2(n18938), .ZN(n18058) );
  INV_X2 U20847 ( .A(n18384), .ZN(n18708) );
  AOI221_X1 U20848 ( .B1(n17696), .B2(n17695), .C1(n18708), .C2(n17695), .A(
        n17694), .ZN(n17704) );
  INV_X1 U20849 ( .A(n17697), .ZN(n17698) );
  AOI21_X1 U20850 ( .B1(n17870), .B2(n17776), .A(n17698), .ZN(n17703) );
  NOR2_X1 U20851 ( .A1(n18057), .A2(n17740), .ZN(n17701) );
  INV_X1 U20852 ( .A(n17699), .ZN(n17700) );
  MUX2_X1 U20853 ( .A(n17701), .B(n17700), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17702) );
  NOR4_X1 U20854 ( .A1(n18058), .A2(n17704), .A3(n17703), .A4(n17702), .ZN(
        n17705) );
  OAI21_X1 U20855 ( .B1(n18063), .B2(n17946), .A(n17705), .ZN(P3_U2804) );
  NAND2_X1 U20856 ( .A1(n18168), .A2(n17712), .ZN(n17706) );
  XOR2_X1 U20857 ( .A(n17706), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18077) );
  NOR2_X1 U20858 ( .A1(n17718), .A2(n18708), .ZN(n17731) );
  AOI211_X1 U20859 ( .C1(n17862), .C2(n17707), .A(n17731), .B(n18021), .ZN(
        n17746) );
  OAI21_X1 U20860 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17776), .A(
        n17746), .ZN(n17719) );
  NOR2_X1 U20861 ( .A1(n18345), .A2(n18936), .ZN(n18072) );
  AND2_X1 U20862 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17710) );
  OAI211_X1 U20863 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17718), .B(n17791), .ZN(n17709) );
  OAI22_X1 U20864 ( .A1(n17710), .A2(n17709), .B1(n17708), .B2(n17870), .ZN(
        n17711) );
  AOI211_X1 U20865 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17719), .A(
        n18072), .B(n17711), .ZN(n17717) );
  NAND2_X1 U20866 ( .A1(n17712), .A2(n18169), .ZN(n17713) );
  XOR2_X1 U20867 ( .A(n17713), .B(n18069), .Z(n18074) );
  AOI21_X1 U20868 ( .B1(n9825), .B2(n17932), .A(n17714), .ZN(n17715) );
  XOR2_X1 U20869 ( .A(n17715), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18073) );
  AOI22_X1 U20870 ( .A1(n17943), .A2(n18074), .B1(n17926), .B2(n18073), .ZN(
        n17716) );
  OAI211_X1 U20871 ( .C1(n18036), .C2(n18077), .A(n17717), .B(n17716), .ZN(
        P3_U2805) );
  OAI22_X1 U20872 ( .A1(n18169), .A2(n17901), .B1(n18168), .B2(n18036), .ZN(
        n17835) );
  AOI21_X1 U20873 ( .B1(n17836), .B2(n18064), .A(n17835), .ZN(n17739) );
  NAND2_X1 U20874 ( .A1(n17718), .A2(n17791), .ZN(n17722) );
  INV_X1 U20875 ( .A(n17719), .ZN(n17720) );
  NAND2_X1 U20876 ( .A1(n9828), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18088) );
  OAI221_X1 U20877 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17722), .C1(
        n17721), .C2(n17720), .A(n18088), .ZN(n17727) );
  AOI21_X1 U20878 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17724), .A(
        n17723), .ZN(n18090) );
  NOR2_X1 U20879 ( .A1(n18091), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18086) );
  INV_X1 U20880 ( .A(n18086), .ZN(n17725) );
  OAI22_X1 U20881 ( .A1(n18090), .A2(n17946), .B1(n17740), .B2(n17725), .ZN(
        n17726) );
  AOI211_X1 U20882 ( .C1(n17890), .C2(n17728), .A(n17727), .B(n17726), .ZN(
        n17729) );
  OAI21_X1 U20883 ( .B1(n17739), .B2(n18083), .A(n17729), .ZN(P3_U2806) );
  INV_X1 U20884 ( .A(n17730), .ZN(n17732) );
  AOI22_X1 U20885 ( .A1(n9828), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17732), 
        .B2(n17731), .ZN(n17744) );
  AOI22_X1 U20886 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17932), .B1(
        n17734), .B2(n17753), .ZN(n17735) );
  NAND2_X1 U20887 ( .A1(n17733), .A2(n17735), .ZN(n17736) );
  XOR2_X1 U20888 ( .A(n17736), .B(n18091), .Z(n18095) );
  INV_X1 U20889 ( .A(n17737), .ZN(n17738) );
  AOI21_X1 U20890 ( .B1(n17870), .B2(n17776), .A(n17738), .ZN(n17742) );
  AOI21_X1 U20891 ( .B1(n18091), .B2(n17740), .A(n17739), .ZN(n17741) );
  AOI211_X1 U20892 ( .C1(n17926), .C2(n18095), .A(n17742), .B(n17741), .ZN(
        n17743) );
  OAI211_X1 U20893 ( .C1(n17746), .C2(n17745), .A(n17744), .B(n17743), .ZN(
        P3_U2807) );
  NAND2_X1 U20894 ( .A1(n17862), .A2(n17747), .ZN(n17748) );
  OAI211_X1 U20895 ( .C1(n9967), .C2(n17749), .A(n18032), .B(n17748), .ZN(
        n17780) );
  AOI21_X1 U20896 ( .B1(n17750), .B2(n17777), .A(n17780), .ZN(n17763) );
  NOR2_X1 U20897 ( .A1(n18345), .A2(n18930), .ZN(n18111) );
  NAND2_X1 U20898 ( .A1(n9967), .A2(n17791), .ZN(n17765) );
  AOI221_X1 U20899 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17764), .C2(n17762), .A(
        n17765), .ZN(n17751) );
  AOI211_X1 U20900 ( .C1(n17752), .C2(n17890), .A(n18111), .B(n17751), .ZN(
        n17761) );
  INV_X1 U20901 ( .A(n17753), .ZN(n17754) );
  OAI221_X1 U20902 ( .B1(n17754), .B2(n18107), .C1(n17754), .C2(n10466), .A(
        n17733), .ZN(n17755) );
  XOR2_X1 U20903 ( .A(n18114), .B(n17755), .Z(n18112) );
  NOR2_X1 U20904 ( .A1(n18097), .A2(n17756), .ZN(n17758) );
  AOI21_X1 U20905 ( .B1(n18097), .B2(n17784), .A(n17835), .ZN(n17775) );
  INV_X1 U20906 ( .A(n17775), .ZN(n17757) );
  MUX2_X1 U20907 ( .A(n17758), .B(n17757), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17759) );
  AOI21_X1 U20908 ( .B1(n17926), .B2(n18112), .A(n17759), .ZN(n17760) );
  OAI211_X1 U20909 ( .C1(n17763), .C2(n17762), .A(n17761), .B(n17760), .ZN(
        P3_U2808) );
  NAND2_X1 U20910 ( .A1(n9828), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18124) );
  OAI221_X1 U20911 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17765), .C1(
        n17764), .C2(n17763), .A(n18124), .ZN(n17772) );
  NOR3_X1 U20912 ( .A1(n17932), .A2(n17814), .A3(n17766), .ZN(n17788) );
  INV_X1 U20913 ( .A(n17767), .ZN(n17810) );
  AOI22_X1 U20914 ( .A1(n18120), .A2(n17788), .B1(n17810), .B2(n17768), .ZN(
        n17769) );
  XOR2_X1 U20915 ( .A(n17769), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(
        n18115) );
  NAND2_X1 U20916 ( .A1(n18120), .A2(n18116), .ZN(n18126) );
  NAND2_X1 U20917 ( .A1(n17770), .A2(n17836), .ZN(n17802) );
  OAI22_X1 U20918 ( .A1(n18115), .A2(n17946), .B1(n18126), .B2(n17802), .ZN(
        n17771) );
  AOI211_X1 U20919 ( .C1(n17890), .C2(n17773), .A(n17772), .B(n17771), .ZN(
        n17774) );
  OAI21_X1 U20920 ( .B1(n17775), .B2(n18116), .A(n17774), .ZN(P3_U2809) );
  OAI21_X1 U20921 ( .B1(n17778), .B2(n18708), .A(n17777), .ZN(n17779) );
  AOI22_X1 U20922 ( .A1(n17781), .A2(n17815), .B1(n17780), .B2(n17779), .ZN(
        n17787) );
  OAI221_X1 U20923 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17809), 
        .C1(n17801), .C2(n17788), .A(n17733), .ZN(n17782) );
  XOR2_X1 U20924 ( .A(n18098), .B(n17782), .Z(n18127) );
  NOR2_X1 U20925 ( .A1(n17783), .A2(n17801), .ZN(n18128) );
  INV_X1 U20926 ( .A(n18128), .ZN(n18099) );
  AOI21_X1 U20927 ( .B1(n17784), .B2(n18099), .A(n17835), .ZN(n17800) );
  NAND2_X1 U20928 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18098), .ZN(
        n18133) );
  OAI22_X1 U20929 ( .A1(n17800), .A2(n18098), .B1(n17802), .B2(n18133), .ZN(
        n17785) );
  AOI21_X1 U20930 ( .B1(n17926), .B2(n18127), .A(n17785), .ZN(n17786) );
  OAI211_X1 U20931 ( .C1(n18345), .C2(n18926), .A(n17787), .B(n17786), .ZN(
        P3_U2810) );
  AOI21_X1 U20932 ( .B1(n17809), .B2(n17810), .A(n17788), .ZN(n17789) );
  XOR2_X1 U20933 ( .A(n17801), .B(n17789), .Z(n18134) );
  NOR2_X1 U20934 ( .A1(n17807), .A2(n17790), .ZN(n17797) );
  OAI211_X1 U20935 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17792), .B(n17791), .ZN(n17796) );
  INV_X1 U20936 ( .A(n17919), .ZN(n18028) );
  OAI21_X1 U20937 ( .B1(n18021), .B2(n17803), .A(n18028), .ZN(n17816) );
  OAI21_X1 U20938 ( .B1(n17793), .B2(n18870), .A(n17816), .ZN(n17806) );
  AOI22_X1 U20939 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17806), .B1(
        n17890), .B2(n17794), .ZN(n17795) );
  NAND2_X1 U20940 ( .A1(n9828), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18136) );
  OAI211_X1 U20941 ( .C1(n17797), .C2(n17796), .A(n17795), .B(n18136), .ZN(
        n17798) );
  AOI21_X1 U20942 ( .B1(n17926), .B2(n18134), .A(n17798), .ZN(n17799) );
  OAI221_X1 U20943 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17802), 
        .C1(n17801), .C2(n17800), .A(n17799), .ZN(P3_U2811) );
  AOI21_X1 U20944 ( .B1(n17836), .B2(n18102), .A(n17835), .ZN(n17825) );
  NOR2_X1 U20945 ( .A1(n17865), .A2(n17803), .ZN(n17808) );
  OAI22_X1 U20946 ( .A1(n18345), .A2(n18922), .B1(n17870), .B2(n17804), .ZN(
        n17805) );
  AOI221_X1 U20947 ( .B1(n17808), .B2(n17807), .C1(n17806), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17805), .ZN(n17813) );
  AOI21_X1 U20948 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17826), .A(
        n17809), .ZN(n17811) );
  XOR2_X1 U20949 ( .A(n17811), .B(n17810), .Z(n18149) );
  NOR2_X1 U20950 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18102), .ZN(
        n18148) );
  AOI22_X1 U20951 ( .A1(n17926), .A2(n18149), .B1(n17836), .B2(n18148), .ZN(
        n17812) );
  OAI211_X1 U20952 ( .C1(n17825), .C2(n17814), .A(n17813), .B(n17812), .ZN(
        P3_U2812) );
  NAND2_X1 U20953 ( .A1(n9828), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18156) );
  INV_X1 U20954 ( .A(n18156), .ZN(n17819) );
  AOI221_X1 U20955 ( .B1(n10603), .B2(n17817), .C1(n18708), .C2(n17817), .A(
        n17816), .ZN(n17818) );
  AOI211_X1 U20956 ( .C1(n17820), .C2(n17815), .A(n17819), .B(n17818), .ZN(
        n17824) );
  OAI21_X1 U20957 ( .B1(n17822), .B2(n18145), .A(n17821), .ZN(n18153) );
  NOR2_X1 U20958 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18162), .ZN(
        n18152) );
  AOI22_X1 U20959 ( .A1(n17926), .A2(n18153), .B1(n17836), .B2(n18152), .ZN(
        n17823) );
  OAI211_X1 U20960 ( .C1(n17825), .C2(n18145), .A(n17824), .B(n17823), .ZN(
        P3_U2813) );
  NAND4_X1 U20961 ( .A1(n17826), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A4(n10452), .ZN(n17924) );
  OAI22_X1 U20962 ( .A1(n17826), .A2(n10466), .B1(n17924), .B2(n18147), .ZN(
        n17827) );
  XOR2_X1 U20963 ( .A(n18162), .B(n17827), .Z(n18167) );
  AOI21_X1 U20964 ( .B1(n17993), .B2(n10021), .A(n18021), .ZN(n17851) );
  OAI21_X1 U20965 ( .B1(n17828), .B2(n18870), .A(n17851), .ZN(n17840) );
  AOI22_X1 U20966 ( .A1(n9828), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17840), .ZN(n17832) );
  NOR3_X1 U20967 ( .A1(n17865), .A2(n17829), .A3(n17866), .ZN(n17842) );
  OAI211_X1 U20968 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17842), .B(n17830), .ZN(n17831) );
  OAI211_X1 U20969 ( .C1(n17870), .C2(n17833), .A(n17832), .B(n17831), .ZN(
        n17834) );
  AOI221_X1 U20970 ( .B1(n17836), .B2(n18162), .C1(n17835), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n17834), .ZN(n17837) );
  OAI21_X1 U20971 ( .B1(n18167), .B2(n17946), .A(n17837), .ZN(P3_U2814) );
  AND2_X1 U20972 ( .A1(n18170), .A2(n10455), .ZN(n17848) );
  OR2_X1 U20973 ( .A1(n17901), .A2(n18169), .ZN(n17847) );
  NAND2_X1 U20974 ( .A1(n9828), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18178) );
  OAI21_X1 U20975 ( .B1(n17870), .B2(n17838), .A(n18178), .ZN(n17839) );
  AOI221_X1 U20976 ( .B1(n17842), .B2(n17841), .C1(n17840), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17839), .ZN(n17846) );
  NOR2_X1 U20977 ( .A1(n18230), .A2(n17924), .ZN(n17905) );
  NAND2_X1 U20978 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17905), .ZN(
        n17878) );
  NOR2_X1 U20979 ( .A1(n10456), .A2(n17878), .ZN(n17857) );
  NAND2_X1 U20980 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n9874), .ZN(
        n17856) );
  OAI221_X1 U20981 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17858), 
        .C1(n18190), .C2(n17857), .A(n17856), .ZN(n17843) );
  XOR2_X1 U20982 ( .A(n10455), .B(n17843), .Z(n18177) );
  NOR2_X1 U20983 ( .A1(n18168), .A2(n18036), .ZN(n17844) );
  OAI21_X1 U20984 ( .B1(n17854), .B2(n18172), .A(n10455), .ZN(n18175) );
  AOI22_X1 U20985 ( .A1(n17926), .A2(n18177), .B1(n17844), .B2(n18175), .ZN(
        n17845) );
  OAI211_X1 U20986 ( .C1(n17848), .C2(n17847), .A(n17846), .B(n17845), .ZN(
        P3_U2815) );
  OAI21_X1 U20987 ( .B1(n17849), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18170), .ZN(n18198) );
  NOR2_X1 U20988 ( .A1(n17866), .A2(n18708), .ZN(n17897) );
  AOI21_X1 U20989 ( .B1(n17867), .B2(n17897), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17850) );
  OAI22_X1 U20990 ( .A1(n17851), .A2(n17850), .B1(n18345), .B2(n18915), .ZN(
        n17852) );
  AOI21_X1 U20991 ( .B1(n17853), .B2(n17815), .A(n17852), .ZN(n17861) );
  NAND2_X1 U20992 ( .A1(n18184), .A2(n18224), .ZN(n18205) );
  NOR2_X1 U20993 ( .A1(n17854), .A2(n18172), .ZN(n17855) );
  AOI221_X1 U20994 ( .B1(n9874), .B2(n18190), .C1(n18205), .C2(n18190), .A(
        n17855), .ZN(n18195) );
  OAI21_X1 U20995 ( .B1(n17858), .B2(n17857), .A(n17856), .ZN(n17859) );
  XOR2_X1 U20996 ( .A(n17859), .B(n18190), .Z(n18194) );
  AOI22_X1 U20997 ( .A1(n18026), .A2(n18195), .B1(n17926), .B2(n18194), .ZN(
        n17860) );
  OAI211_X1 U20998 ( .C1(n17901), .C2(n18198), .A(n17861), .B(n17860), .ZN(
        P3_U2816) );
  AOI22_X1 U20999 ( .A1(n17943), .A2(n18200), .B1(n18026), .B2(n18205), .ZN(
        n17884) );
  AOI21_X1 U21000 ( .B1(n17993), .B2(n17866), .A(n17862), .ZN(n17863) );
  OAI21_X1 U21001 ( .B1(n17864), .B2(n17863), .A(n18032), .ZN(n17880) );
  OR2_X1 U21002 ( .A1(n17866), .A2(n17865), .ZN(n17883) );
  AOI211_X1 U21003 ( .C1(n17882), .C2(n17868), .A(n17867), .B(n17883), .ZN(
        n17872) );
  OAI22_X1 U21004 ( .A1(n18345), .A2(n18912), .B1(n17870), .B2(n17869), .ZN(
        n17871) );
  AOI211_X1 U21005 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17880), .A(
        n17872), .B(n17871), .ZN(n17876) );
  AOI22_X1 U21006 ( .A1(n18184), .A2(n17909), .B1(n17932), .B2(n10456), .ZN(
        n17873) );
  AOI21_X1 U21007 ( .B1(n17877), .B2(n17932), .A(n17873), .ZN(n17874) );
  XOR2_X1 U21008 ( .A(n17874), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18209) );
  AND2_X1 U21009 ( .A1(n9874), .A2(n18184), .ZN(n18208) );
  AOI22_X1 U21010 ( .A1(n17926), .A2(n18209), .B1(n18208), .B2(n17900), .ZN(
        n17875) );
  OAI211_X1 U21011 ( .C1(n17884), .C2(n9874), .A(n17876), .B(n17875), .ZN(
        P3_U2817) );
  NAND2_X1 U21012 ( .A1(n17878), .A2(n17877), .ZN(n17879) );
  XOR2_X1 U21013 ( .A(n17879), .B(n10456), .Z(n18221) );
  INV_X1 U21014 ( .A(n17880), .ZN(n17881) );
  NAND2_X1 U21015 ( .A1(n9828), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18219) );
  OAI221_X1 U21016 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17883), .C1(
        n17882), .C2(n17881), .A(n18219), .ZN(n17888) );
  NOR2_X1 U21017 ( .A1(n17930), .A2(n18201), .ZN(n17886) );
  INV_X1 U21018 ( .A(n17884), .ZN(n17885) );
  MUX2_X1 U21019 ( .A(n17886), .B(n17885), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n17887) );
  AOI211_X1 U21020 ( .C1(n17890), .C2(n17889), .A(n17888), .B(n17887), .ZN(
        n17891) );
  OAI21_X1 U21021 ( .B1(n18221), .B2(n17946), .A(n17891), .ZN(P3_U2818) );
  NOR2_X1 U21022 ( .A1(n17905), .A2(n17892), .ZN(n17893) );
  XOR2_X1 U21023 ( .A(n17893), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18235) );
  NOR2_X1 U21024 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18230), .ZN(
        n18222) );
  NOR2_X1 U21025 ( .A1(n18345), .A2(n18908), .ZN(n17899) );
  NAND3_X1 U21026 ( .A1(n16937), .A2(n17894), .A3(n18738), .ZN(n17923) );
  NOR2_X1 U21027 ( .A1(n17911), .A2(n17923), .ZN(n17910) );
  AOI21_X1 U21028 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18028), .A(
        n17910), .ZN(n17896) );
  OAI22_X1 U21029 ( .A1(n17897), .A2(n17896), .B1(n18018), .B2(n17895), .ZN(
        n17898) );
  AOI211_X1 U21030 ( .C1(n18222), .C2(n17900), .A(n17899), .B(n17898), .ZN(
        n17903) );
  AND2_X1 U21031 ( .A1(n18230), .A2(n17900), .ZN(n17915) );
  OAI22_X1 U21032 ( .A1(n18227), .A2(n17901), .B1(n18036), .B2(n18224), .ZN(
        n17927) );
  OAI21_X1 U21033 ( .B1(n17915), .B2(n17927), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17902) );
  OAI211_X1 U21034 ( .C1(n18235), .C2(n17946), .A(n17903), .B(n17902), .ZN(
        P3_U2819) );
  NAND3_X1 U21035 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17932), .A3(
        n10173), .ZN(n17908) );
  OAI221_X1 U21036 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17904), .C1(
        n10173), .C2(n17924), .A(n10174), .ZN(n17907) );
  INV_X1 U21037 ( .A(n17905), .ZN(n17906) );
  OAI211_X1 U21038 ( .C1(n17909), .C2(n17908), .A(n17907), .B(n17906), .ZN(
        n18244) );
  AOI211_X1 U21039 ( .C1(n17923), .C2(n17911), .A(n17919), .B(n17910), .ZN(
        n17912) );
  INV_X1 U21040 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18906) );
  NOR2_X1 U21041 ( .A1(n18345), .A2(n18906), .ZN(n18241) );
  AOI211_X1 U21042 ( .C1(n17913), .C2(n17815), .A(n17912), .B(n18241), .ZN(
        n17917) );
  NAND2_X1 U21043 ( .A1(n10173), .A2(n10174), .ZN(n17914) );
  AOI22_X1 U21044 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17927), .B1(
        n17915), .B2(n17914), .ZN(n17916) );
  OAI211_X1 U21045 ( .C1(n17946), .C2(n18244), .A(n17917), .B(n17916), .ZN(
        P3_U2820) );
  NAND2_X1 U21046 ( .A1(n16937), .A2(n18738), .ZN(n17951) );
  OAI22_X1 U21047 ( .A1(n17919), .A2(n17918), .B1(n17936), .B2(n17951), .ZN(
        n17922) );
  OAI22_X1 U21048 ( .A1(n18018), .A2(n17920), .B1(n18345), .B2(n18904), .ZN(
        n17921) );
  AOI21_X1 U21049 ( .B1(n17923), .B2(n17922), .A(n17921), .ZN(n17929) );
  NAND2_X1 U21050 ( .A1(n17924), .A2(n17904), .ZN(n17925) );
  XOR2_X1 U21051 ( .A(n17925), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18249) );
  AOI22_X1 U21052 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17927), .B1(
        n17926), .B2(n18249), .ZN(n17928) );
  OAI211_X1 U21053 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17930), .A(
        n17929), .B(n17928), .ZN(P3_U2821) );
  OAI21_X1 U21054 ( .B1(n18267), .B2(n17932), .A(n17931), .ZN(n18270) );
  AOI21_X1 U21055 ( .B1(n17934), .B2(n18263), .A(n17933), .ZN(n18265) );
  AOI21_X1 U21056 ( .B1(n17993), .B2(n17935), .A(n18021), .ZN(n17959) );
  OAI211_X1 U21057 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17937), .A(
        n18384), .B(n17936), .ZN(n17939) );
  INV_X1 U21058 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18903) );
  NOR2_X1 U21059 ( .A1(n18345), .A2(n18903), .ZN(n18261) );
  INV_X1 U21060 ( .A(n18261), .ZN(n17938) );
  OAI211_X1 U21061 ( .C1(n17959), .C2(n17940), .A(n17939), .B(n17938), .ZN(
        n17941) );
  AOI21_X1 U21062 ( .B1(n18026), .B2(n18265), .A(n17941), .ZN(n17945) );
  AOI22_X1 U21063 ( .A1(n17943), .A2(n18267), .B1(n17942), .B2(n17815), .ZN(
        n17944) );
  OAI211_X1 U21064 ( .C1(n17946), .C2(n18270), .A(n17945), .B(n17944), .ZN(
        P3_U2822) );
  OAI21_X1 U21065 ( .B1(n17949), .B2(n17948), .A(n17947), .ZN(n17950) );
  XOR2_X1 U21066 ( .A(n17950), .B(n18280), .Z(n18277) );
  OAI22_X1 U21067 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17951), .B1(
        n18345), .B2(n18900), .ZN(n17956) );
  OAI21_X1 U21068 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17953), .A(
        n17952), .ZN(n18273) );
  OAI22_X1 U21069 ( .A1(n18018), .A2(n17954), .B1(n18035), .B2(n18273), .ZN(
        n17955) );
  AOI211_X1 U21070 ( .C1(n18026), .C2(n18277), .A(n17956), .B(n17955), .ZN(
        n17957) );
  OAI21_X1 U21071 ( .B1(n17959), .B2(n17958), .A(n17957), .ZN(P3_U2823) );
  OAI21_X1 U21072 ( .B1(n18708), .B2(n17960), .A(n18028), .ZN(n17981) );
  OR2_X1 U21073 ( .A1(n17960), .A2(n18708), .ZN(n17964) );
  OAI21_X1 U21074 ( .B1(n17963), .B2(n17962), .A(n17961), .ZN(n18288) );
  OAI22_X1 U21075 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17964), .B1(
        n18035), .B2(n18288), .ZN(n17965) );
  AOI21_X1 U21076 ( .B1(n9828), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17965), .ZN(
        n17973) );
  AOI22_X1 U21077 ( .A1(n17968), .A2(n17975), .B1(n17967), .B2(n17966), .ZN(
        n17969) );
  XOR2_X1 U21078 ( .A(n17970), .B(n17969), .Z(n18281) );
  AOI22_X1 U21079 ( .A1(n18026), .A2(n18281), .B1(n17971), .B2(n17815), .ZN(
        n17972) );
  OAI211_X1 U21080 ( .C1(n17974), .C2(n17981), .A(n17973), .B(n17972), .ZN(
        P3_U2824) );
  OAI21_X1 U21081 ( .B1(n17977), .B2(n17976), .A(n17975), .ZN(n18295) );
  AOI21_X1 U21082 ( .B1(n17978), .B2(n18032), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17982) );
  OAI21_X1 U21083 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17980), .A(
        n17979), .ZN(n18289) );
  OAI22_X1 U21084 ( .A1(n17982), .A2(n17981), .B1(n18035), .B2(n18289), .ZN(
        n17983) );
  AOI21_X1 U21085 ( .B1(n17984), .B2(n17815), .A(n17983), .ZN(n17985) );
  NAND2_X1 U21086 ( .A1(n9828), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18293) );
  OAI211_X1 U21087 ( .C1(n18036), .C2(n18295), .A(n17985), .B(n18293), .ZN(
        P3_U2825) );
  OAI21_X1 U21088 ( .B1(n17988), .B2(n17987), .A(n17986), .ZN(n18298) );
  OAI21_X1 U21089 ( .B1(n17991), .B2(n17990), .A(n17989), .ZN(n18304) );
  OAI22_X1 U21090 ( .A1(n18036), .A2(n18304), .B1(n18345), .B2(n18894), .ZN(
        n17997) );
  AOI21_X1 U21091 ( .B1(n17993), .B2(n17992), .A(n18021), .ZN(n18006) );
  OAI22_X1 U21092 ( .A1(n18018), .A2(n17995), .B1(n17994), .B2(n18006), .ZN(
        n17996) );
  AOI211_X1 U21093 ( .C1(n18384), .C2(n17998), .A(n17997), .B(n17996), .ZN(
        n17999) );
  OAI21_X1 U21094 ( .B1(n18035), .B2(n18298), .A(n17999), .ZN(P3_U2826) );
  OAI21_X1 U21095 ( .B1(n18002), .B2(n18001), .A(n18000), .ZN(n18307) );
  AOI21_X1 U21096 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18032), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18007) );
  OAI21_X1 U21097 ( .B1(n18005), .B2(n18004), .A(n18003), .ZN(n18313) );
  OAI22_X1 U21098 ( .A1(n18007), .A2(n18006), .B1(n18035), .B2(n18313), .ZN(
        n18008) );
  AOI21_X1 U21099 ( .B1(n18009), .B2(n17815), .A(n18008), .ZN(n18010) );
  NAND2_X1 U21100 ( .A1(n9828), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18311) );
  OAI211_X1 U21101 ( .C1(n18036), .C2(n18307), .A(n18010), .B(n18311), .ZN(
        P3_U2827) );
  OAI21_X1 U21102 ( .B1(n18013), .B2(n18012), .A(n18011), .ZN(n18323) );
  OAI21_X1 U21103 ( .B1(n18016), .B2(n18015), .A(n18014), .ZN(n18322) );
  OAI22_X1 U21104 ( .A1(n18018), .A2(n18017), .B1(n18035), .B2(n18322), .ZN(
        n18019) );
  AOI221_X1 U21105 ( .B1(n18021), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18738), .C2(n18020), .A(n18019), .ZN(n18022) );
  NAND2_X1 U21106 ( .A1(n9828), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18327) );
  OAI211_X1 U21107 ( .C1(n18036), .C2(n18323), .A(n18022), .B(n18327), .ZN(
        P3_U2828) );
  OAI21_X1 U21108 ( .B1(n9890), .B2(n18024), .A(n18023), .ZN(n18342) );
  NAND2_X1 U21109 ( .A1(n18991), .A2(n18031), .ZN(n18025) );
  XNOR2_X1 U21110 ( .A(n18025), .B(n18024), .ZN(n18338) );
  AOI22_X1 U21111 ( .A1(n18026), .A2(n18338), .B1(n9828), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18030) );
  AOI22_X1 U21112 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18028), .B1(
        n17815), .B2(n18027), .ZN(n18029) );
  OAI211_X1 U21113 ( .C1(n18035), .C2(n18342), .A(n18030), .B(n18029), .ZN(
        P3_U2829) );
  AOI21_X1 U21114 ( .B1(n18031), .B2(n18991), .A(n9890), .ZN(n18353) );
  INV_X1 U21115 ( .A(n18353), .ZN(n18351) );
  NAND3_X1 U21116 ( .A1(n18972), .A2(n18870), .A3(n18032), .ZN(n18033) );
  AOI22_X1 U21117 ( .A1(n9828), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18033), .ZN(n18034) );
  OAI221_X1 U21118 ( .B1(n18353), .B2(n18036), .C1(n18351), .C2(n18035), .A(
        n18034), .ZN(P3_U2830) );
  NAND2_X1 U21119 ( .A1(n18345), .A2(n18344), .ZN(n18330) );
  NAND2_X1 U21120 ( .A1(n18037), .A2(n18106), .ZN(n18092) );
  NOR2_X1 U21121 ( .A1(n18038), .A2(n18092), .ZN(n18052) );
  NAND2_X1 U21122 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18041) );
  NOR2_X1 U21123 ( .A1(n18812), .A2(n18817), .ZN(n18314) );
  INV_X1 U21124 ( .A(n18314), .ZN(n18144) );
  AOI21_X1 U21125 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18809), .A(
        n18039), .ZN(n18104) );
  NOR2_X1 U21126 ( .A1(n18104), .A2(n18097), .ZN(n18040) );
  AOI21_X1 U21127 ( .B1(n18159), .B2(n18040), .A(n18314), .ZN(n18080) );
  AOI21_X1 U21128 ( .B1(n18041), .B2(n18144), .A(n18080), .ZN(n18065) );
  AOI22_X1 U21129 ( .A1(n18812), .A2(n18069), .B1(n18817), .B2(n18042), .ZN(
        n18048) );
  AOI22_X1 U21130 ( .A1(n18790), .A2(n18045), .B1(n18044), .B2(n18043), .ZN(
        n18047) );
  NAND4_X1 U21131 ( .A1(n18065), .A2(n18048), .A3(n18047), .A4(n18046), .ZN(
        n18060) );
  AOI21_X1 U21132 ( .B1(n18812), .B2(n18049), .A(n18060), .ZN(n18050) );
  INV_X1 U21133 ( .A(n18050), .ZN(n18051) );
  MUX2_X1 U21134 ( .A(n18052), .B(n18051), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n18053) );
  AOI22_X1 U21135 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18334), .B1(
        n18326), .B2(n18053), .ZN(n18055) );
  NAND2_X1 U21136 ( .A1(n9828), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18054) );
  OAI211_X1 U21137 ( .C1(n18056), .C2(n18271), .A(n18055), .B(n18054), .ZN(
        P3_U2835) );
  NOR2_X1 U21138 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18057), .ZN(
        n18059) );
  AOI21_X1 U21139 ( .B1(n18059), .B2(n18087), .A(n18058), .ZN(n18062) );
  OAI211_X1 U21140 ( .C1(n18344), .C2(n18060), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n18345), .ZN(n18061) );
  OAI211_X1 U21141 ( .C1(n18063), .C2(n18271), .A(n18062), .B(n18061), .ZN(
        P3_U2836) );
  NOR2_X1 U21142 ( .A1(n18064), .A2(n18101), .ZN(n18082) );
  OAI221_X1 U21143 ( .B1(n18804), .B2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), 
        .C1(n18804), .C2(n18082), .A(n18065), .ZN(n18066) );
  OAI21_X1 U21144 ( .B1(n18069), .B2(n18066), .A(n18326), .ZN(n18067) );
  AOI221_X1 U21145 ( .B1(n18070), .B2(n18069), .C1(n18068), .C2(n18069), .A(
        n18067), .ZN(n18071) );
  AOI211_X1 U21146 ( .C1(n18334), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18072), .B(n18071), .ZN(n18076) );
  AOI22_X1 U21147 ( .A1(n18266), .A2(n18074), .B1(n18250), .B2(n18073), .ZN(
        n18075) );
  OAI211_X1 U21148 ( .C1(n18352), .C2(n18077), .A(n18076), .B(n18075), .ZN(
        P3_U2837) );
  NAND2_X1 U21149 ( .A1(n18225), .A2(n18226), .ZN(n18229) );
  INV_X1 U21150 ( .A(n18229), .ZN(n18142) );
  NOR2_X1 U21151 ( .A1(n18078), .A2(n18142), .ZN(n18079) );
  OAI22_X1 U21152 ( .A1(n18169), .A2(n18226), .B1(n18168), .B2(n18225), .ZN(
        n18158) );
  NOR4_X1 U21153 ( .A1(n18334), .A2(n18080), .A3(n18079), .A4(n18158), .ZN(
        n18084) );
  NOR2_X1 U21154 ( .A1(n18822), .A2(n18091), .ZN(n18081) );
  AOI221_X1 U21155 ( .B1(n18082), .B2(n18084), .C1(n18081), .C2(n18084), .A(
        n9828), .ZN(n18094) );
  AOI21_X1 U21156 ( .B1(n18297), .B2(n18084), .A(n18083), .ZN(n18085) );
  AOI22_X1 U21157 ( .A1(n18087), .A2(n18086), .B1(n18094), .B2(n18085), .ZN(
        n18089) );
  OAI211_X1 U21158 ( .C1(n18090), .C2(n18271), .A(n18089), .B(n18088), .ZN(
        P3_U2838) );
  OAI21_X1 U21159 ( .B1(n18334), .B2(n18092), .A(n18091), .ZN(n18093) );
  AOI22_X1 U21160 ( .A1(n18250), .A2(n18095), .B1(n18094), .B2(n18093), .ZN(
        n18096) );
  OAI21_X1 U21161 ( .B1(n18345), .B2(n18933), .A(n18096), .ZN(P3_U2839) );
  AOI22_X1 U21162 ( .A1(n18812), .A2(n18098), .B1(n18097), .B2(n18229), .ZN(
        n18119) );
  AOI221_X1 U21163 ( .B1(n18100), .B2(n18812), .C1(n18099), .C2(n18812), .A(
        n18158), .ZN(n18103) );
  OAI21_X1 U21164 ( .B1(n18102), .B2(n18101), .A(n18822), .ZN(n18140) );
  OAI211_X1 U21165 ( .C1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n18804), .A(
        n18103), .B(n18140), .ZN(n18117) );
  AOI211_X1 U21166 ( .C1(n18202), .C2(n18105), .A(n18104), .B(n18117), .ZN(
        n18109) );
  AOI21_X1 U21167 ( .B1(n18107), .B2(n18106), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18108) );
  AOI211_X1 U21168 ( .C1(n18119), .C2(n18109), .A(n18108), .B(n18344), .ZN(
        n18110) );
  AOI211_X1 U21169 ( .C1(n18112), .C2(n18250), .A(n18111), .B(n18110), .ZN(
        n18113) );
  OAI21_X1 U21170 ( .B1(n18114), .B2(n18330), .A(n18113), .ZN(P3_U2840) );
  INV_X1 U21171 ( .A(n18115), .ZN(n18123) );
  NOR2_X1 U21172 ( .A1(n9828), .A2(n18116), .ZN(n18122) );
  NOR2_X1 U21173 ( .A1(n18822), .A2(n18817), .ZN(n18333) );
  AOI211_X1 U21174 ( .C1(n18817), .C2(n18118), .A(n18344), .B(n18117), .ZN(
        n18129) );
  OAI211_X1 U21175 ( .C1(n18120), .C2(n18333), .A(n18129), .B(n18119), .ZN(
        n18121) );
  AOI22_X1 U21176 ( .A1(n18250), .A2(n18123), .B1(n18122), .B2(n18121), .ZN(
        n18125) );
  OAI211_X1 U21177 ( .C1(n18126), .C2(n18138), .A(n18125), .B(n18124), .ZN(
        P3_U2841) );
  AOI22_X1 U21178 ( .A1(n9828), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18250), 
        .B2(n18127), .ZN(n18132) );
  AOI221_X1 U21179 ( .B1(n18142), .B2(n18129), .C1(n18128), .C2(n18129), .A(
        n9828), .ZN(n18135) );
  NOR3_X1 U21180 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18333), .A3(
        n18354), .ZN(n18130) );
  OAI21_X1 U21181 ( .B1(n18135), .B2(n18130), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18131) );
  OAI211_X1 U21182 ( .C1(n18133), .C2(n18138), .A(n18132), .B(n18131), .ZN(
        P3_U2842) );
  AOI22_X1 U21183 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18135), .B1(
        n18250), .B2(n18134), .ZN(n18137) );
  OAI211_X1 U21184 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18138), .A(
        n18137), .B(n18136), .ZN(P3_U2843) );
  NAND2_X1 U21185 ( .A1(n18817), .A2(n18991), .ZN(n18315) );
  NAND3_X1 U21186 ( .A1(n18159), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18315), .ZN(n18139) );
  AOI211_X1 U21187 ( .C1(n18144), .C2(n18139), .A(n18344), .B(n18158), .ZN(
        n18141) );
  OAI211_X1 U21188 ( .C1(n18143), .C2(n18142), .A(n18141), .B(n18140), .ZN(
        n18154) );
  OAI221_X1 U21189 ( .B1(n18154), .B2(n18145), .C1(n18154), .C2(n18144), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18151) );
  NOR2_X1 U21190 ( .A1(n18329), .A2(n18973), .ZN(n18257) );
  AOI22_X1 U21191 ( .A1(n18822), .A2(n18321), .B1(n18257), .B2(n18318), .ZN(
        n18306) );
  NOR2_X1 U21192 ( .A1(n18306), .A2(n18254), .ZN(n18272) );
  NAND3_X1 U21193 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n18272), .ZN(n18189) );
  NAND2_X1 U21194 ( .A1(n18146), .A2(n18189), .ZN(n18213) );
  NAND2_X1 U21195 ( .A1(n18326), .A2(n18213), .ZN(n18253) );
  NOR2_X1 U21196 ( .A1(n18147), .A2(n18253), .ZN(n18163) );
  AOI22_X1 U21197 ( .A1(n18250), .A2(n18149), .B1(n18148), .B2(n18163), .ZN(
        n18150) );
  OAI221_X1 U21198 ( .B1(n9828), .B2(n18151), .C1(n18345), .C2(n18922), .A(
        n18150), .ZN(P3_U2844) );
  AOI22_X1 U21199 ( .A1(n18250), .A2(n18153), .B1(n18163), .B2(n18152), .ZN(
        n18157) );
  NAND3_X1 U21200 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18345), .A3(
        n18154), .ZN(n18155) );
  NAND3_X1 U21201 ( .A1(n18157), .A2(n18156), .A3(n18155), .ZN(P3_U2845) );
  NOR2_X1 U21202 ( .A1(n18344), .A2(n18158), .ZN(n18161) );
  AOI22_X1 U21203 ( .A1(n18809), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18159), .ZN(n18160) );
  OAI22_X1 U21204 ( .A1(n18802), .A2(n18182), .B1(n18181), .B2(n18804), .ZN(
        n18223) );
  AOI211_X1 U21205 ( .C1(n18202), .C2(n18172), .A(n18160), .B(n18223), .ZN(
        n18171) );
  AOI221_X1 U21206 ( .B1(n18297), .B2(n18161), .C1(n18171), .C2(n18161), .A(
        n9828), .ZN(n18164) );
  AOI22_X1 U21207 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18164), .B1(
        n18163), .B2(n18162), .ZN(n18166) );
  NAND2_X1 U21208 ( .A1(n9828), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n18165) );
  OAI211_X1 U21209 ( .C1(n18167), .C2(n18271), .A(n18166), .B(n18165), .ZN(
        P3_U2846) );
  NOR2_X1 U21210 ( .A1(n18168), .A2(n18225), .ZN(n18176) );
  AOI211_X1 U21211 ( .C1(n18170), .C2(n10455), .A(n18169), .B(n18226), .ZN(
        n18174) );
  AOI221_X1 U21212 ( .B1(n18172), .B2(n10455), .C1(n18189), .C2(n10455), .A(
        n18171), .ZN(n18173) );
  AOI211_X1 U21213 ( .C1(n18176), .C2(n18175), .A(n18174), .B(n18173), .ZN(
        n18180) );
  AOI22_X1 U21214 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18334), .B1(
        n18250), .B2(n18177), .ZN(n18179) );
  OAI211_X1 U21215 ( .C1(n18180), .C2(n18344), .A(n18179), .B(n18178), .ZN(
        P3_U2847) );
  NOR2_X1 U21216 ( .A1(n18345), .A2(n18915), .ZN(n18193) );
  OAI221_X1 U21217 ( .B1(n18804), .B2(n18184), .C1(n18804), .C2(n18181), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18187) );
  INV_X1 U21218 ( .A(n18182), .ZN(n18183) );
  OAI21_X1 U21219 ( .B1(n18191), .B2(n18183), .A(n18812), .ZN(n18185) );
  NOR2_X1 U21220 ( .A1(n18991), .A2(n18183), .ZN(n18245) );
  NAND2_X1 U21221 ( .A1(n18184), .A2(n18245), .ZN(n18212) );
  NAND2_X1 U21222 ( .A1(n18817), .A2(n18212), .ZN(n18206) );
  OAI211_X1 U21223 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18333), .A(
        n18185), .B(n18206), .ZN(n18186) );
  OAI21_X1 U21224 ( .B1(n18187), .B2(n18186), .A(n18326), .ZN(n18188) );
  AOI221_X1 U21225 ( .B1(n18191), .B2(n18190), .C1(n18189), .C2(n18190), .A(
        n18188), .ZN(n18192) );
  AOI211_X1 U21226 ( .C1(n18334), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18193), .B(n18192), .ZN(n18197) );
  AOI22_X1 U21227 ( .A1(n18339), .A2(n18195), .B1(n18250), .B2(n18194), .ZN(
        n18196) );
  OAI211_X1 U21228 ( .C1(n18199), .C2(n18198), .A(n18197), .B(n18196), .ZN(
        P3_U2848) );
  INV_X1 U21229 ( .A(n18202), .ZN(n18237) );
  INV_X1 U21230 ( .A(n18200), .ZN(n18203) );
  NAND2_X1 U21231 ( .A1(n18202), .A2(n18201), .ZN(n18231) );
  OAI21_X1 U21232 ( .B1(n18203), .B2(n18226), .A(n18231), .ZN(n18204) );
  AOI211_X1 U21233 ( .C1(n18790), .C2(n18205), .A(n18223), .B(n18204), .ZN(
        n18217) );
  OAI211_X1 U21234 ( .C1(n18237), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18217), .B(n18206), .ZN(n18207) );
  OAI21_X1 U21235 ( .B1(n18344), .B2(n18207), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18211) );
  INV_X1 U21236 ( .A(n18253), .ZN(n18239) );
  AOI22_X1 U21237 ( .A1(n18250), .A2(n18209), .B1(n18239), .B2(n18208), .ZN(
        n18210) );
  OAI221_X1 U21238 ( .B1(n9828), .B2(n18211), .C1(n18345), .C2(n18912), .A(
        n18210), .ZN(P3_U2849) );
  OAI21_X1 U21239 ( .B1(n10456), .B2(n18817), .A(n18212), .ZN(n18216) );
  AOI21_X1 U21240 ( .B1(n18214), .B2(n18213), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18215) );
  AOI211_X1 U21241 ( .C1(n18217), .C2(n18216), .A(n18215), .B(n18344), .ZN(
        n18218) );
  AOI21_X1 U21242 ( .B1(n18334), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18218), .ZN(n18220) );
  OAI211_X1 U21243 ( .C1(n18221), .C2(n18271), .A(n18220), .B(n18219), .ZN(
        P3_U2850) );
  AOI22_X1 U21244 ( .A1(n9828), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18239), 
        .B2(n18222), .ZN(n18234) );
  NOR2_X1 U21245 ( .A1(n18344), .A2(n18223), .ZN(n18246) );
  OAI221_X1 U21246 ( .B1(n18809), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18809), .C2(n18245), .A(n18246), .ZN(n18228) );
  OAI22_X1 U21247 ( .A1(n18227), .A2(n18226), .B1(n18225), .B2(n18224), .ZN(
        n18247) );
  AOI211_X1 U21248 ( .C1(n18230), .C2(n18229), .A(n18228), .B(n18247), .ZN(
        n18236) );
  OAI211_X1 U21249 ( .C1(n18809), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18236), .B(n18231), .ZN(n18232) );
  NAND3_X1 U21250 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18345), .A3(
        n18232), .ZN(n18233) );
  OAI211_X1 U21251 ( .C1(n18235), .C2(n18271), .A(n18234), .B(n18233), .ZN(
        P3_U2851) );
  AOI221_X1 U21252 ( .B1(n18237), .B2(n18236), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18236), .A(n9828), .ZN(n18240) );
  NOR2_X1 U21253 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n10173), .ZN(
        n18238) );
  AOI22_X1 U21254 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18240), .B1(
        n18239), .B2(n18238), .ZN(n18243) );
  INV_X1 U21255 ( .A(n18241), .ZN(n18242) );
  OAI211_X1 U21256 ( .C1(n18271), .C2(n18244), .A(n18243), .B(n18242), .ZN(
        P3_U2852) );
  AOI22_X1 U21257 ( .A1(n18809), .A2(n18246), .B1(n18326), .B2(n18245), .ZN(
        n18248) );
  OAI21_X1 U21258 ( .B1(n18248), .B2(n18247), .A(n18345), .ZN(n18252) );
  AOI22_X1 U21259 ( .A1(n9828), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18250), .B2(
        n18249), .ZN(n18251) );
  OAI221_X1 U21260 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18253), .C1(
        n10173), .C2(n18252), .A(n18251), .ZN(P3_U2853) );
  NOR4_X1 U21261 ( .A1(n18306), .A2(n18344), .A3(n18280), .A4(n18254), .ZN(
        n18264) );
  NAND2_X1 U21262 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18258) );
  AOI21_X1 U21263 ( .B1(n18822), .B2(n18255), .A(n18308), .ZN(n18256) );
  OAI211_X1 U21264 ( .C1(n18257), .C2(n18314), .A(n18256), .B(n18315), .ZN(
        n18296) );
  OAI21_X1 U21265 ( .B1(n18258), .B2(n18296), .A(n18260), .ZN(n18282) );
  OAI21_X1 U21266 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18344), .A(
        n18282), .ZN(n18259) );
  AOI21_X1 U21267 ( .B1(n18260), .B2(n18284), .A(n18259), .ZN(n18275) );
  OAI21_X1 U21268 ( .B1(n18297), .B2(n18275), .A(n18330), .ZN(n18262) );
  AOI221_X1 U21269 ( .B1(n18264), .B2(n18263), .C1(n18262), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18261), .ZN(n18269) );
  AOI22_X1 U21270 ( .A1(n18267), .A2(n18266), .B1(n18339), .B2(n18265), .ZN(
        n18268) );
  OAI211_X1 U21271 ( .C1(n18271), .C2(n18270), .A(n18269), .B(n18268), .ZN(
        P3_U2854) );
  NOR2_X1 U21272 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18272), .ZN(
        n18274) );
  OAI22_X1 U21273 ( .A1(n18275), .A2(n18274), .B1(n18350), .B2(n18273), .ZN(
        n18276) );
  AOI21_X1 U21274 ( .B1(n18339), .B2(n18277), .A(n18276), .ZN(n18279) );
  NAND2_X1 U21275 ( .A1(n9828), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n18278) );
  OAI211_X1 U21276 ( .C1(n18330), .C2(n18280), .A(n18279), .B(n18278), .ZN(
        P3_U2855) );
  AOI22_X1 U21277 ( .A1(n9828), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18339), .B2(
        n18281), .ZN(n18287) );
  NAND2_X1 U21278 ( .A1(n18330), .A2(n18282), .ZN(n18292) );
  NOR3_X1 U21279 ( .A1(n18306), .A2(n18283), .A3(n18344), .ZN(n18285) );
  AOI22_X1 U21280 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18292), .B1(
        n18285), .B2(n18284), .ZN(n18286) );
  OAI211_X1 U21281 ( .C1(n18350), .C2(n18288), .A(n18287), .B(n18286), .ZN(
        P3_U2856) );
  NOR3_X1 U21282 ( .A1(n18306), .A2(n18344), .A3(n18308), .ZN(n18302) );
  NAND2_X1 U21283 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18302), .ZN(
        n18290) );
  OAI22_X1 U21284 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18290), .B1(
        n18289), .B2(n18350), .ZN(n18291) );
  AOI21_X1 U21285 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18292), .A(
        n18291), .ZN(n18294) );
  OAI211_X1 U21286 ( .C1(n18352), .C2(n18295), .A(n18294), .B(n18293), .ZN(
        P3_U2857) );
  INV_X1 U21287 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18301) );
  NAND2_X1 U21288 ( .A1(n18326), .A2(n18296), .ZN(n18305) );
  OAI21_X1 U21289 ( .B1(n18297), .B2(n18305), .A(n18330), .ZN(n18300) );
  OAI22_X1 U21290 ( .A1(n18345), .A2(n18894), .B1(n18350), .B2(n18298), .ZN(
        n18299) );
  AOI221_X1 U21291 ( .B1(n18302), .B2(n18301), .C1(n18300), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18299), .ZN(n18303) );
  OAI21_X1 U21292 ( .B1(n18352), .B2(n18304), .A(n18303), .ZN(P3_U2858) );
  AOI21_X1 U21293 ( .B1(n18306), .B2(n18308), .A(n18305), .ZN(n18310) );
  OAI22_X1 U21294 ( .A1(n18308), .A2(n18330), .B1(n18352), .B2(n18307), .ZN(
        n18309) );
  NOR2_X1 U21295 ( .A1(n18310), .A2(n18309), .ZN(n18312) );
  OAI211_X1 U21296 ( .C1(n18313), .C2(n18350), .A(n18312), .B(n18311), .ZN(
        P3_U2859) );
  AOI21_X1 U21297 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18315), .A(
        n18314), .ZN(n18317) );
  NOR2_X1 U21298 ( .A1(n18973), .A2(n18991), .ZN(n18316) );
  OAI221_X1 U21299 ( .B1(n18317), .B2(n18822), .C1(n18317), .C2(n18316), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18320) );
  NAND3_X1 U21300 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18318), .A3(
        n18329), .ZN(n18319) );
  OAI211_X1 U21301 ( .C1(n18321), .C2(n18804), .A(n18320), .B(n18319), .ZN(
        n18325) );
  OAI22_X1 U21302 ( .A1(n18352), .A2(n18323), .B1(n18350), .B2(n18322), .ZN(
        n18324) );
  AOI21_X1 U21303 ( .B1(n18326), .B2(n18325), .A(n18324), .ZN(n18328) );
  OAI211_X1 U21304 ( .C1(n18330), .C2(n18329), .A(n18328), .B(n18327), .ZN(
        P3_U2860) );
  NOR2_X1 U21305 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18812), .ZN(
        n18332) );
  NOR2_X1 U21306 ( .A1(n18332), .A2(n18331), .ZN(n18336) );
  NOR3_X1 U21307 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18333), .A3(
        n18344), .ZN(n18346) );
  NOR2_X1 U21308 ( .A1(n18334), .A2(n18346), .ZN(n18343) );
  INV_X1 U21309 ( .A(n18343), .ZN(n18335) );
  MUX2_X1 U21310 ( .A(n18336), .B(n18335), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n18337) );
  AOI21_X1 U21311 ( .B1(n18339), .B2(n18338), .A(n18337), .ZN(n18341) );
  NAND2_X1 U21312 ( .A1(n9828), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18340) );
  OAI211_X1 U21313 ( .C1(n18342), .C2(n18350), .A(n18341), .B(n18340), .ZN(
        P3_U2861) );
  OAI21_X1 U21314 ( .B1(n18802), .B2(n18344), .A(n18343), .ZN(n18348) );
  INV_X1 U21315 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19002) );
  NOR2_X1 U21316 ( .A1(n18345), .A2(n19002), .ZN(n18347) );
  AOI211_X1 U21317 ( .C1(n18348), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18347), .B(n18346), .ZN(n18349) );
  OAI221_X1 U21318 ( .B1(n18353), .B2(n18352), .C1(n18351), .C2(n18350), .A(
        n18349), .ZN(P3_U2862) );
  AOI211_X1 U21319 ( .C1(n18356), .C2(n18355), .A(n18354), .B(n18972), .ZN(
        n18851) );
  OAI21_X1 U21320 ( .B1(n18851), .B2(n18411), .A(n18362), .ZN(n18357) );
  OAI221_X1 U21321 ( .B1(n18368), .B2(n19008), .C1(n18368), .C2(n18362), .A(
        n18357), .ZN(P3_U2863) );
  INV_X1 U21322 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18836) );
  NAND2_X1 U21323 ( .A1(n18836), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18540) );
  NAND2_X1 U21324 ( .A1(n18367), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18635) );
  INV_X1 U21325 ( .A(n18635), .ZN(n18637) );
  NAND2_X1 U21326 ( .A1(n18358), .A2(n18637), .ZN(n18659) );
  AND2_X1 U21327 ( .A1(n18540), .A2(n18659), .ZN(n18360) );
  OAI22_X1 U21328 ( .A1(n18361), .A2(n18836), .B1(n18360), .B2(n18359), .ZN(
        P3_U2866) );
  NOR2_X1 U21329 ( .A1(n18363), .A2(n18362), .ZN(P3_U2867) );
  NOR2_X1 U21330 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18814) );
  NAND2_X1 U21331 ( .A1(n18367), .A2(n18836), .ZN(n18496) );
  INV_X1 U21332 ( .A(n18496), .ZN(n18454) );
  NAND2_X1 U21333 ( .A1(n18814), .A2(n18454), .ZN(n18410) );
  NOR2_X1 U21334 ( .A1(n18365), .A2(n18364), .ZN(n18403) );
  NAND2_X1 U21335 ( .A1(n18403), .A2(n18366), .ZN(n18742) );
  AND2_X1 U21336 ( .A1(n18662), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18733) );
  INV_X1 U21337 ( .A(n18732), .ZN(n18860) );
  NAND2_X1 U21338 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18634) );
  INV_X1 U21339 ( .A(n18634), .ZN(n18813) );
  NOR2_X1 U21340 ( .A1(n18367), .A2(n18836), .ZN(n18369) );
  NAND2_X1 U21341 ( .A1(n18813), .A2(n18369), .ZN(n18789) );
  INV_X1 U21342 ( .A(n18789), .ZN(n18449) );
  INV_X1 U21343 ( .A(n18410), .ZN(n18469) );
  NOR2_X1 U21344 ( .A1(n18449), .A2(n18469), .ZN(n18431) );
  NOR2_X1 U21345 ( .A1(n18860), .A2(n18431), .ZN(n18405) );
  AND2_X1 U21346 ( .A1(n18738), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18734) );
  NOR2_X1 U21347 ( .A1(n18636), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18610) );
  NAND2_X1 U21348 ( .A1(n18369), .A2(n18610), .ZN(n18731) );
  INV_X1 U21349 ( .A(n18731), .ZN(n18711) );
  AOI22_X1 U21350 ( .A1(n18733), .A2(n18405), .B1(n18734), .B2(n18711), .ZN(
        n18374) );
  AOI21_X1 U21351 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18431), .ZN(n18370) );
  NOR2_X1 U21352 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18368), .ZN(
        n18586) );
  NOR2_X1 U21353 ( .A1(n18610), .A2(n18586), .ZN(n18660) );
  INV_X1 U21354 ( .A(n18369), .ZN(n18371) );
  NOR2_X1 U21355 ( .A1(n18660), .A2(n18371), .ZN(n18705) );
  AOI22_X1 U21356 ( .A1(n18662), .A2(n18370), .B1(n18738), .B2(n18705), .ZN(
        n18407) );
  NOR2_X1 U21357 ( .A1(n18371), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18737) );
  NAND2_X1 U21358 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18737), .ZN(
        n18704) );
  INV_X1 U21359 ( .A(n18704), .ZN(n18784) );
  INV_X1 U21360 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18372) );
  NOR2_X2 U21361 ( .A1(n18372), .A2(n18708), .ZN(n18739) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18407), .B1(
        n18784), .B2(n18739), .ZN(n18373) );
  OAI211_X1 U21363 ( .C1(n18410), .C2(n18742), .A(n18374), .B(n18373), .ZN(
        P3_U2868) );
  NAND2_X1 U21364 ( .A1(n18403), .A2(n18375), .ZN(n18748) );
  INV_X1 U21365 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18376) );
  NOR2_X2 U21366 ( .A1(n18376), .A2(n18708), .ZN(n18745) );
  AND2_X1 U21367 ( .A1(n18662), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18743) );
  AOI22_X1 U21368 ( .A1(n18784), .A2(n18745), .B1(n18405), .B2(n18743), .ZN(
        n18378) );
  AND2_X1 U21369 ( .A1(n18738), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18744) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18407), .B1(
        n18711), .B2(n18744), .ZN(n18377) );
  OAI211_X1 U21371 ( .C1(n18410), .C2(n18748), .A(n18378), .B(n18377), .ZN(
        P3_U2869) );
  NAND2_X1 U21372 ( .A1(n18403), .A2(n18379), .ZN(n18754) );
  NOR2_X2 U21373 ( .A1(n18380), .A2(n18708), .ZN(n18751) );
  AND2_X1 U21374 ( .A1(n18662), .A2(BUF2_REG_2__SCAN_IN), .ZN(n18749) );
  AOI22_X1 U21375 ( .A1(n18784), .A2(n18751), .B1(n18405), .B2(n18749), .ZN(
        n18382) );
  AND2_X1 U21376 ( .A1(n18738), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18750) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18407), .B1(
        n18711), .B2(n18750), .ZN(n18381) );
  OAI211_X1 U21378 ( .C1(n18410), .C2(n18754), .A(n18382), .B(n18381), .ZN(
        P3_U2870) );
  NAND2_X1 U21379 ( .A1(n18403), .A2(n18383), .ZN(n18760) );
  AND2_X1 U21380 ( .A1(n18662), .A2(BUF2_REG_3__SCAN_IN), .ZN(n18755) );
  AND2_X1 U21381 ( .A1(n18384), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18757) );
  AOI22_X1 U21382 ( .A1(n18405), .A2(n18755), .B1(n18711), .B2(n18757), .ZN(
        n18386) );
  INV_X1 U21383 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n19367) );
  NOR2_X2 U21384 ( .A1(n19367), .A2(n18708), .ZN(n18756) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18407), .B1(
        n18784), .B2(n18756), .ZN(n18385) );
  OAI211_X1 U21386 ( .C1(n18410), .C2(n18760), .A(n18386), .B(n18385), .ZN(
        P3_U2871) );
  NAND2_X1 U21387 ( .A1(n18403), .A2(n18387), .ZN(n18766) );
  NOR2_X2 U21388 ( .A1(n18707), .A2(n18388), .ZN(n18761) );
  INV_X1 U21389 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18389) );
  NOR2_X2 U21390 ( .A1(n18708), .A2(n18389), .ZN(n18762) );
  AOI22_X1 U21391 ( .A1(n18405), .A2(n18761), .B1(n18711), .B2(n18762), .ZN(
        n18391) );
  NOR2_X2 U21392 ( .A1(n19372), .A2(n18708), .ZN(n18763) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18407), .B1(
        n18784), .B2(n18763), .ZN(n18390) );
  OAI211_X1 U21394 ( .C1(n18410), .C2(n18766), .A(n18391), .B(n18390), .ZN(
        P3_U2872) );
  NAND2_X1 U21395 ( .A1(n18403), .A2(n18392), .ZN(n18772) );
  NOR2_X2 U21396 ( .A1(n18707), .A2(n18393), .ZN(n18767) );
  NOR2_X2 U21397 ( .A1(n18708), .A2(n19378), .ZN(n18769) );
  AOI22_X1 U21398 ( .A1(n18405), .A2(n18767), .B1(n18711), .B2(n18769), .ZN(
        n18396) );
  INV_X1 U21399 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18394) );
  NOR2_X2 U21400 ( .A1(n18394), .A2(n18708), .ZN(n18768) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18407), .B1(
        n18784), .B2(n18768), .ZN(n18395) );
  OAI211_X1 U21402 ( .C1(n18410), .C2(n18772), .A(n18396), .B(n18395), .ZN(
        P3_U2873) );
  NAND2_X1 U21403 ( .A1(n18403), .A2(n18397), .ZN(n18778) );
  NOR2_X2 U21404 ( .A1(n18707), .A2(n18398), .ZN(n18773) );
  AND2_X1 U21405 ( .A1(n18738), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18775) );
  AOI22_X1 U21406 ( .A1(n18405), .A2(n18773), .B1(n18711), .B2(n18775), .ZN(
        n18401) );
  INV_X1 U21407 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18399) );
  NOR2_X2 U21408 ( .A1(n18399), .A2(n18708), .ZN(n18774) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18407), .B1(
        n18784), .B2(n18774), .ZN(n18400) );
  OAI211_X1 U21410 ( .C1(n18410), .C2(n18778), .A(n18401), .B(n18400), .ZN(
        P3_U2874) );
  NAND2_X1 U21411 ( .A1(n18403), .A2(n18402), .ZN(n18788) );
  NOR2_X2 U21412 ( .A1(n18404), .A2(n18707), .ZN(n18780) );
  AND2_X1 U21413 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18738), .ZN(n18783) );
  AOI22_X1 U21414 ( .A1(n18405), .A2(n18780), .B1(n18711), .B2(n18783), .ZN(
        n18409) );
  NOR2_X2 U21415 ( .A1(n18708), .A2(n18406), .ZN(n18782) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18407), .B1(
        n18784), .B2(n18782), .ZN(n18408) );
  OAI211_X1 U21417 ( .C1(n18410), .C2(n18788), .A(n18409), .B(n18408), .ZN(
        P3_U2875) );
  NAND2_X1 U21418 ( .A1(n18454), .A2(n18586), .ZN(n18430) );
  NAND2_X1 U21419 ( .A1(n18636), .A2(n18732), .ZN(n18587) );
  NOR2_X1 U21420 ( .A1(n18496), .A2(n18587), .ZN(n18426) );
  AOI22_X1 U21421 ( .A1(n18739), .A2(n18711), .B1(n18733), .B2(n18426), .ZN(
        n18413) );
  NOR2_X1 U21422 ( .A1(n18836), .A2(n18588), .ZN(n18735) );
  NOR2_X1 U21423 ( .A1(n18707), .A2(n18411), .ZN(n18736) );
  INV_X1 U21424 ( .A(n18736), .ZN(n18453) );
  NOR2_X1 U21425 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18453), .ZN(
        n18497) );
  AOI22_X1 U21426 ( .A1(n18738), .A2(n18735), .B1(n18454), .B2(n18497), .ZN(
        n18427) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18427), .B1(
        n18449), .B2(n18734), .ZN(n18412) );
  OAI211_X1 U21428 ( .C1(n18742), .C2(n18430), .A(n18413), .B(n18412), .ZN(
        P3_U2876) );
  AOI22_X1 U21429 ( .A1(n18711), .A2(n18745), .B1(n18743), .B2(n18426), .ZN(
        n18415) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18427), .B1(
        n18449), .B2(n18744), .ZN(n18414) );
  OAI211_X1 U21431 ( .C1(n18748), .C2(n18430), .A(n18415), .B(n18414), .ZN(
        P3_U2877) );
  AOI22_X1 U21432 ( .A1(n18449), .A2(n18750), .B1(n18749), .B2(n18426), .ZN(
        n18417) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18427), .B1(
        n18711), .B2(n18751), .ZN(n18416) );
  OAI211_X1 U21434 ( .C1(n18754), .C2(n18430), .A(n18417), .B(n18416), .ZN(
        P3_U2878) );
  AOI22_X1 U21435 ( .A1(n18711), .A2(n18756), .B1(n18755), .B2(n18426), .ZN(
        n18419) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18427), .B1(
        n18449), .B2(n18757), .ZN(n18418) );
  OAI211_X1 U21437 ( .C1(n18760), .C2(n18430), .A(n18419), .B(n18418), .ZN(
        P3_U2879) );
  AOI22_X1 U21438 ( .A1(n18711), .A2(n18763), .B1(n18761), .B2(n18426), .ZN(
        n18421) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18427), .B1(
        n18449), .B2(n18762), .ZN(n18420) );
  OAI211_X1 U21440 ( .C1(n18766), .C2(n18430), .A(n18421), .B(n18420), .ZN(
        P3_U2880) );
  AOI22_X1 U21441 ( .A1(n18711), .A2(n18768), .B1(n18767), .B2(n18426), .ZN(
        n18423) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18427), .B1(
        n18449), .B2(n18769), .ZN(n18422) );
  OAI211_X1 U21443 ( .C1(n18772), .C2(n18430), .A(n18423), .B(n18422), .ZN(
        P3_U2881) );
  AOI22_X1 U21444 ( .A1(n18449), .A2(n18775), .B1(n18773), .B2(n18426), .ZN(
        n18425) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18427), .B1(
        n18711), .B2(n18774), .ZN(n18424) );
  OAI211_X1 U21446 ( .C1(n18778), .C2(n18430), .A(n18425), .B(n18424), .ZN(
        P3_U2882) );
  AOI22_X1 U21447 ( .A1(n18711), .A2(n18782), .B1(n18780), .B2(n18426), .ZN(
        n18429) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18427), .B1(
        n18449), .B2(n18783), .ZN(n18428) );
  OAI211_X1 U21449 ( .C1(n18788), .C2(n18430), .A(n18429), .B(n18428), .ZN(
        P3_U2883) );
  NAND2_X1 U21450 ( .A1(n18454), .A2(n18610), .ZN(n18452) );
  INV_X1 U21451 ( .A(n18430), .ZN(n18491) );
  INV_X1 U21452 ( .A(n18452), .ZN(n18514) );
  NOR2_X1 U21453 ( .A1(n18491), .A2(n18514), .ZN(n18474) );
  NOR2_X1 U21454 ( .A1(n18860), .A2(n18474), .ZN(n18447) );
  AOI22_X1 U21455 ( .A1(n18469), .A2(n18734), .B1(n18733), .B2(n18447), .ZN(
        n18434) );
  OAI21_X1 U21456 ( .B1(n18431), .B2(n18611), .A(n18474), .ZN(n18432) );
  OAI211_X1 U21457 ( .C1(n18514), .C2(n18963), .A(n18662), .B(n18432), .ZN(
        n18448) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18448), .B1(
        n18739), .B2(n18449), .ZN(n18433) );
  OAI211_X1 U21459 ( .C1(n18742), .C2(n18452), .A(n18434), .B(n18433), .ZN(
        P3_U2884) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18448), .B1(
        n18743), .B2(n18447), .ZN(n18436) );
  AOI22_X1 U21461 ( .A1(n18449), .A2(n18745), .B1(n18469), .B2(n18744), .ZN(
        n18435) );
  OAI211_X1 U21462 ( .C1(n18748), .C2(n18452), .A(n18436), .B(n18435), .ZN(
        P3_U2885) );
  AOI22_X1 U21463 ( .A1(n18449), .A2(n18751), .B1(n18749), .B2(n18447), .ZN(
        n18438) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18448), .B1(
        n18469), .B2(n18750), .ZN(n18437) );
  OAI211_X1 U21465 ( .C1(n18754), .C2(n18452), .A(n18438), .B(n18437), .ZN(
        P3_U2886) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18448), .B1(
        n18755), .B2(n18447), .ZN(n18440) );
  AOI22_X1 U21467 ( .A1(n18449), .A2(n18756), .B1(n18469), .B2(n18757), .ZN(
        n18439) );
  OAI211_X1 U21468 ( .C1(n18760), .C2(n18452), .A(n18440), .B(n18439), .ZN(
        P3_U2887) );
  AOI22_X1 U21469 ( .A1(n18469), .A2(n18762), .B1(n18761), .B2(n18447), .ZN(
        n18442) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18448), .B1(
        n18449), .B2(n18763), .ZN(n18441) );
  OAI211_X1 U21471 ( .C1(n18766), .C2(n18452), .A(n18442), .B(n18441), .ZN(
        P3_U2888) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18448), .B1(
        n18767), .B2(n18447), .ZN(n18444) );
  AOI22_X1 U21473 ( .A1(n18449), .A2(n18768), .B1(n18469), .B2(n18769), .ZN(
        n18443) );
  OAI211_X1 U21474 ( .C1(n18772), .C2(n18452), .A(n18444), .B(n18443), .ZN(
        P3_U2889) );
  AOI22_X1 U21475 ( .A1(n18469), .A2(n18775), .B1(n18773), .B2(n18447), .ZN(
        n18446) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18448), .B1(
        n18449), .B2(n18774), .ZN(n18445) );
  OAI211_X1 U21477 ( .C1(n18778), .C2(n18452), .A(n18446), .B(n18445), .ZN(
        P3_U2890) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18448), .B1(
        n18780), .B2(n18447), .ZN(n18451) );
  AOI22_X1 U21479 ( .A1(n18449), .A2(n18782), .B1(n18469), .B2(n18783), .ZN(
        n18450) );
  OAI211_X1 U21480 ( .C1(n18788), .C2(n18452), .A(n18451), .B(n18450), .ZN(
        P3_U2891) );
  NOR2_X2 U21481 ( .A1(n18634), .A2(n18496), .ZN(n18535) );
  INV_X1 U21482 ( .A(n18535), .ZN(n18473) );
  AOI22_X1 U21483 ( .A1(n18739), .A2(n18469), .B1(n18733), .B2(n10031), .ZN(
        n18456) );
  AOI21_X1 U21484 ( .B1(n18636), .B2(n18611), .A(n18453), .ZN(n18542) );
  NAND2_X1 U21485 ( .A1(n18454), .A2(n18542), .ZN(n18470) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18470), .B1(
        n18734), .B2(n18491), .ZN(n18455) );
  OAI211_X1 U21487 ( .C1(n18742), .C2(n18473), .A(n18456), .B(n18455), .ZN(
        P3_U2892) );
  AOI22_X1 U21488 ( .A1(n18469), .A2(n18745), .B1(n18743), .B2(n10031), .ZN(
        n18458) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18470), .B1(
        n18744), .B2(n18491), .ZN(n18457) );
  OAI211_X1 U21490 ( .C1(n18748), .C2(n18473), .A(n18458), .B(n18457), .ZN(
        P3_U2893) );
  AOI22_X1 U21491 ( .A1(n18469), .A2(n18751), .B1(n18749), .B2(n10031), .ZN(
        n18460) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18470), .B1(
        n18750), .B2(n18491), .ZN(n18459) );
  OAI211_X1 U21493 ( .C1(n18754), .C2(n18473), .A(n18460), .B(n18459), .ZN(
        P3_U2894) );
  AOI22_X1 U21494 ( .A1(n18469), .A2(n18756), .B1(n18755), .B2(n10031), .ZN(
        n18462) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18470), .B1(
        n18757), .B2(n18491), .ZN(n18461) );
  OAI211_X1 U21496 ( .C1(n18760), .C2(n18473), .A(n18462), .B(n18461), .ZN(
        P3_U2895) );
  AOI22_X1 U21497 ( .A1(n18469), .A2(n18763), .B1(n18761), .B2(n10031), .ZN(
        n18464) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18470), .B1(
        n18762), .B2(n18491), .ZN(n18463) );
  OAI211_X1 U21499 ( .C1(n18766), .C2(n18473), .A(n18464), .B(n18463), .ZN(
        P3_U2896) );
  AOI22_X1 U21500 ( .A1(n18769), .A2(n18491), .B1(n18767), .B2(n10031), .ZN(
        n18466) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18470), .B1(
        n18469), .B2(n18768), .ZN(n18465) );
  OAI211_X1 U21502 ( .C1(n18772), .C2(n18473), .A(n18466), .B(n18465), .ZN(
        P3_U2897) );
  AOI22_X1 U21503 ( .A1(n18773), .A2(n10031), .B1(n18775), .B2(n18491), .ZN(
        n18468) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18470), .B1(
        n18469), .B2(n18774), .ZN(n18467) );
  OAI211_X1 U21505 ( .C1(n18778), .C2(n18473), .A(n18468), .B(n18467), .ZN(
        P3_U2898) );
  AOI22_X1 U21506 ( .A1(n18783), .A2(n18491), .B1(n18780), .B2(n10031), .ZN(
        n18472) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18470), .B1(
        n18469), .B2(n18782), .ZN(n18471) );
  OAI211_X1 U21508 ( .C1(n18788), .C2(n18473), .A(n18472), .B(n18471), .ZN(
        P3_U2899) );
  INV_X1 U21509 ( .A(n18540), .ZN(n18541) );
  NAND2_X1 U21510 ( .A1(n18814), .A2(n18541), .ZN(n18495) );
  INV_X1 U21511 ( .A(n18495), .ZN(n18559) );
  NOR2_X1 U21512 ( .A1(n18535), .A2(n18559), .ZN(n18518) );
  NOR2_X1 U21513 ( .A1(n18860), .A2(n18518), .ZN(n18490) );
  AOI22_X1 U21514 ( .A1(n18739), .A2(n18491), .B1(n18733), .B2(n18490), .ZN(
        n18477) );
  OAI22_X1 U21515 ( .A1(n18474), .A2(n18708), .B1(n18518), .B2(n18707), .ZN(
        n18475) );
  OAI21_X1 U21516 ( .B1(n18559), .B2(n18963), .A(n18475), .ZN(n18492) );
  AOI22_X1 U21517 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18492), .B1(
        n18734), .B2(n18514), .ZN(n18476) );
  OAI211_X1 U21518 ( .C1(n18742), .C2(n18495), .A(n18477), .B(n18476), .ZN(
        P3_U2900) );
  AOI22_X1 U21519 ( .A1(n18745), .A2(n18491), .B1(n18743), .B2(n18490), .ZN(
        n18479) );
  AOI22_X1 U21520 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18492), .B1(
        n18744), .B2(n18514), .ZN(n18478) );
  OAI211_X1 U21521 ( .C1(n18748), .C2(n18495), .A(n18479), .B(n18478), .ZN(
        P3_U2901) );
  AOI22_X1 U21522 ( .A1(n18749), .A2(n18490), .B1(n18751), .B2(n18491), .ZN(
        n18481) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18492), .B1(
        n18750), .B2(n18514), .ZN(n18480) );
  OAI211_X1 U21524 ( .C1(n18754), .C2(n18495), .A(n18481), .B(n18480), .ZN(
        P3_U2902) );
  AOI22_X1 U21525 ( .A1(n18756), .A2(n18491), .B1(n18755), .B2(n18490), .ZN(
        n18483) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18492), .B1(
        n18757), .B2(n18514), .ZN(n18482) );
  OAI211_X1 U21527 ( .C1(n18760), .C2(n18495), .A(n18483), .B(n18482), .ZN(
        P3_U2903) );
  AOI22_X1 U21528 ( .A1(n18761), .A2(n18490), .B1(n18762), .B2(n18514), .ZN(
        n18485) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18492), .B1(
        n18763), .B2(n18491), .ZN(n18484) );
  OAI211_X1 U21530 ( .C1(n18766), .C2(n18495), .A(n18485), .B(n18484), .ZN(
        P3_U2904) );
  AOI22_X1 U21531 ( .A1(n18768), .A2(n18491), .B1(n18767), .B2(n18490), .ZN(
        n18487) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18492), .B1(
        n18769), .B2(n18514), .ZN(n18486) );
  OAI211_X1 U21533 ( .C1(n18772), .C2(n18495), .A(n18487), .B(n18486), .ZN(
        P3_U2905) );
  AOI22_X1 U21534 ( .A1(n18773), .A2(n18490), .B1(n18775), .B2(n18514), .ZN(
        n18489) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18492), .B1(
        n18774), .B2(n18491), .ZN(n18488) );
  OAI211_X1 U21536 ( .C1(n18778), .C2(n18495), .A(n18489), .B(n18488), .ZN(
        P3_U2906) );
  AOI22_X1 U21537 ( .A1(n18783), .A2(n18514), .B1(n18780), .B2(n18490), .ZN(
        n18494) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18492), .B1(
        n18782), .B2(n18491), .ZN(n18493) );
  OAI211_X1 U21539 ( .C1(n18788), .C2(n18495), .A(n18494), .B(n18493), .ZN(
        P3_U2907) );
  NAND2_X1 U21540 ( .A1(n18586), .A2(n18541), .ZN(n18543) );
  NOR2_X1 U21541 ( .A1(n18587), .A2(n18540), .ZN(n18513) );
  AOI22_X1 U21542 ( .A1(n18739), .A2(n18514), .B1(n18733), .B2(n18513), .ZN(
        n18500) );
  NOR2_X1 U21543 ( .A1(n18636), .A2(n18496), .ZN(n18498) );
  AOI22_X1 U21544 ( .A1(n18738), .A2(n18498), .B1(n18497), .B2(n18541), .ZN(
        n18515) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18515), .B1(
        n18734), .B2(n18535), .ZN(n18499) );
  OAI211_X1 U21546 ( .C1(n18742), .C2(n18543), .A(n18500), .B(n18499), .ZN(
        P3_U2908) );
  AOI22_X1 U21547 ( .A1(n18745), .A2(n18514), .B1(n18743), .B2(n18513), .ZN(
        n18502) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18515), .B1(
        n18744), .B2(n18535), .ZN(n18501) );
  OAI211_X1 U21549 ( .C1(n18748), .C2(n18543), .A(n18502), .B(n18501), .ZN(
        P3_U2909) );
  AOI22_X1 U21550 ( .A1(n18750), .A2(n18535), .B1(n18749), .B2(n18513), .ZN(
        n18504) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18515), .B1(
        n18751), .B2(n18514), .ZN(n18503) );
  OAI211_X1 U21552 ( .C1(n18754), .C2(n18543), .A(n18504), .B(n18503), .ZN(
        P3_U2910) );
  AOI22_X1 U21553 ( .A1(n18756), .A2(n18514), .B1(n18755), .B2(n18513), .ZN(
        n18506) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18515), .B1(
        n18757), .B2(n18535), .ZN(n18505) );
  OAI211_X1 U21555 ( .C1(n18760), .C2(n18543), .A(n18506), .B(n18505), .ZN(
        P3_U2911) );
  AOI22_X1 U21556 ( .A1(n18761), .A2(n18513), .B1(n18762), .B2(n18535), .ZN(
        n18508) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18515), .B1(
        n18763), .B2(n18514), .ZN(n18507) );
  OAI211_X1 U21558 ( .C1(n18766), .C2(n18543), .A(n18508), .B(n18507), .ZN(
        P3_U2912) );
  AOI22_X1 U21559 ( .A1(n18769), .A2(n18535), .B1(n18767), .B2(n18513), .ZN(
        n18510) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18515), .B1(
        n18768), .B2(n18514), .ZN(n18509) );
  OAI211_X1 U21561 ( .C1(n18772), .C2(n18543), .A(n18510), .B(n18509), .ZN(
        P3_U2913) );
  AOI22_X1 U21562 ( .A1(n18773), .A2(n18513), .B1(n18775), .B2(n18535), .ZN(
        n18512) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18515), .B1(
        n18774), .B2(n18514), .ZN(n18511) );
  OAI211_X1 U21564 ( .C1(n18778), .C2(n18543), .A(n18512), .B(n18511), .ZN(
        P3_U2914) );
  AOI22_X1 U21565 ( .A1(n18782), .A2(n18514), .B1(n18780), .B2(n18513), .ZN(
        n18517) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18515), .B1(
        n18783), .B2(n18535), .ZN(n18516) );
  OAI211_X1 U21567 ( .C1(n18788), .C2(n18543), .A(n18517), .B(n18516), .ZN(
        P3_U2915) );
  NAND2_X1 U21568 ( .A1(n18610), .A2(n18541), .ZN(n18539) );
  AOI21_X1 U21569 ( .B1(n18543), .B2(n18539), .A(n18860), .ZN(n18534) );
  AOI22_X1 U21570 ( .A1(n18733), .A2(n18534), .B1(n18734), .B2(n18559), .ZN(
        n18521) );
  INV_X1 U21571 ( .A(n18539), .ZN(n18606) );
  AOI221_X1 U21572 ( .B1(n18518), .B2(n18543), .C1(n18611), .C2(n18543), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18519) );
  OAI21_X1 U21573 ( .B1(n18606), .B2(n18519), .A(n18662), .ZN(n18536) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18536), .B1(
        n18739), .B2(n18535), .ZN(n18520) );
  OAI211_X1 U21575 ( .C1(n18742), .C2(n18539), .A(n18521), .B(n18520), .ZN(
        P3_U2916) );
  AOI22_X1 U21576 ( .A1(n18745), .A2(n18535), .B1(n18743), .B2(n18534), .ZN(
        n18523) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18536), .B1(
        n18744), .B2(n18559), .ZN(n18522) );
  OAI211_X1 U21578 ( .C1(n18748), .C2(n18539), .A(n18523), .B(n18522), .ZN(
        P3_U2917) );
  AOI22_X1 U21579 ( .A1(n18750), .A2(n18559), .B1(n18749), .B2(n18534), .ZN(
        n18525) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18536), .B1(
        n18751), .B2(n18535), .ZN(n18524) );
  OAI211_X1 U21581 ( .C1(n18754), .C2(n18539), .A(n18525), .B(n18524), .ZN(
        P3_U2918) );
  AOI22_X1 U21582 ( .A1(n18756), .A2(n18535), .B1(n18755), .B2(n18534), .ZN(
        n18527) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18536), .B1(
        n18757), .B2(n18559), .ZN(n18526) );
  OAI211_X1 U21584 ( .C1(n18760), .C2(n18539), .A(n18527), .B(n18526), .ZN(
        P3_U2919) );
  AOI22_X1 U21585 ( .A1(n18763), .A2(n18535), .B1(n18761), .B2(n18534), .ZN(
        n18529) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18536), .B1(
        n18762), .B2(n18559), .ZN(n18528) );
  OAI211_X1 U21587 ( .C1(n18766), .C2(n18539), .A(n18529), .B(n18528), .ZN(
        P3_U2920) );
  AOI22_X1 U21588 ( .A1(n18768), .A2(n18535), .B1(n18767), .B2(n18534), .ZN(
        n18531) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18536), .B1(
        n18769), .B2(n18559), .ZN(n18530) );
  OAI211_X1 U21590 ( .C1(n18772), .C2(n18539), .A(n18531), .B(n18530), .ZN(
        P3_U2921) );
  AOI22_X1 U21591 ( .A1(n18773), .A2(n18534), .B1(n18775), .B2(n18559), .ZN(
        n18533) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18536), .B1(
        n18774), .B2(n18535), .ZN(n18532) );
  OAI211_X1 U21593 ( .C1(n18778), .C2(n18539), .A(n18533), .B(n18532), .ZN(
        P3_U2922) );
  AOI22_X1 U21594 ( .A1(n18783), .A2(n18559), .B1(n18780), .B2(n18534), .ZN(
        n18538) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18536), .B1(
        n18782), .B2(n18535), .ZN(n18537) );
  OAI211_X1 U21596 ( .C1(n18788), .C2(n18539), .A(n18538), .B(n18537), .ZN(
        P3_U2923) );
  NOR2_X2 U21597 ( .A1(n18634), .A2(n18540), .ZN(n18629) );
  INV_X1 U21598 ( .A(n18629), .ZN(n18563) );
  AOI22_X1 U21599 ( .A1(n18739), .A2(n18559), .B1(n18733), .B2(n18558), .ZN(
        n18545) );
  NAND2_X1 U21600 ( .A1(n18542), .A2(n18541), .ZN(n18560) );
  INV_X1 U21601 ( .A(n18543), .ZN(n18581) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18560), .B1(
        n18734), .B2(n18581), .ZN(n18544) );
  OAI211_X1 U21603 ( .C1(n18742), .C2(n18563), .A(n18545), .B(n18544), .ZN(
        P3_U2924) );
  AOI22_X1 U21604 ( .A1(n18745), .A2(n18559), .B1(n18743), .B2(n18558), .ZN(
        n18547) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18560), .B1(
        n18744), .B2(n18581), .ZN(n18546) );
  OAI211_X1 U21606 ( .C1(n18748), .C2(n18563), .A(n18547), .B(n18546), .ZN(
        P3_U2925) );
  AOI22_X1 U21607 ( .A1(n18750), .A2(n18581), .B1(n18749), .B2(n18558), .ZN(
        n18549) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18560), .B1(
        n18751), .B2(n18559), .ZN(n18548) );
  OAI211_X1 U21609 ( .C1(n18754), .C2(n18563), .A(n18549), .B(n18548), .ZN(
        P3_U2926) );
  AOI22_X1 U21610 ( .A1(n18757), .A2(n18581), .B1(n18755), .B2(n18558), .ZN(
        n18551) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18560), .B1(
        n18756), .B2(n18559), .ZN(n18550) );
  OAI211_X1 U21612 ( .C1(n18760), .C2(n18563), .A(n18551), .B(n18550), .ZN(
        P3_U2927) );
  AOI22_X1 U21613 ( .A1(n18763), .A2(n18559), .B1(n18761), .B2(n18558), .ZN(
        n18553) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18560), .B1(
        n18762), .B2(n18581), .ZN(n18552) );
  OAI211_X1 U21615 ( .C1(n18766), .C2(n18563), .A(n18553), .B(n18552), .ZN(
        P3_U2928) );
  AOI22_X1 U21616 ( .A1(n18769), .A2(n18581), .B1(n18767), .B2(n18558), .ZN(
        n18555) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18560), .B1(
        n18768), .B2(n18559), .ZN(n18554) );
  OAI211_X1 U21618 ( .C1(n18772), .C2(n18563), .A(n18555), .B(n18554), .ZN(
        P3_U2929) );
  AOI22_X1 U21619 ( .A1(n18773), .A2(n18558), .B1(n18775), .B2(n18581), .ZN(
        n18557) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18560), .B1(
        n18774), .B2(n18559), .ZN(n18556) );
  OAI211_X1 U21621 ( .C1(n18778), .C2(n18563), .A(n18557), .B(n18556), .ZN(
        P3_U2930) );
  AOI22_X1 U21622 ( .A1(n18783), .A2(n18581), .B1(n18780), .B2(n18558), .ZN(
        n18562) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18560), .B1(
        n18782), .B2(n18559), .ZN(n18561) );
  OAI211_X1 U21624 ( .C1(n18788), .C2(n18563), .A(n18562), .B(n18561), .ZN(
        P3_U2931) );
  NAND2_X1 U21625 ( .A1(n18814), .A2(n18637), .ZN(n18585) );
  INV_X1 U21626 ( .A(n18585), .ZN(n18654) );
  NOR2_X1 U21627 ( .A1(n18629), .A2(n18654), .ZN(n18612) );
  NOR2_X1 U21628 ( .A1(n18860), .A2(n18612), .ZN(n18580) );
  AOI22_X1 U21629 ( .A1(n18739), .A2(n18581), .B1(n18733), .B2(n18580), .ZN(
        n18567) );
  NOR2_X1 U21630 ( .A1(n18581), .A2(n18606), .ZN(n18564) );
  OAI21_X1 U21631 ( .B1(n18564), .B2(n18611), .A(n18612), .ZN(n18565) );
  OAI211_X1 U21632 ( .C1(n18654), .C2(n18963), .A(n18662), .B(n18565), .ZN(
        n18582) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18582), .B1(
        n18734), .B2(n18606), .ZN(n18566) );
  OAI211_X1 U21634 ( .C1(n18742), .C2(n18585), .A(n18567), .B(n18566), .ZN(
        P3_U2932) );
  AOI22_X1 U21635 ( .A1(n18745), .A2(n18581), .B1(n18743), .B2(n18580), .ZN(
        n18569) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18582), .B1(
        n18744), .B2(n18606), .ZN(n18568) );
  OAI211_X1 U21637 ( .C1(n18748), .C2(n18585), .A(n18569), .B(n18568), .ZN(
        P3_U2933) );
  AOI22_X1 U21638 ( .A1(n18749), .A2(n18580), .B1(n18751), .B2(n18581), .ZN(
        n18571) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18582), .B1(
        n18750), .B2(n18606), .ZN(n18570) );
  OAI211_X1 U21640 ( .C1(n18754), .C2(n18585), .A(n18571), .B(n18570), .ZN(
        P3_U2934) );
  AOI22_X1 U21641 ( .A1(n18757), .A2(n18606), .B1(n18755), .B2(n18580), .ZN(
        n18573) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18582), .B1(
        n18756), .B2(n18581), .ZN(n18572) );
  OAI211_X1 U21643 ( .C1(n18760), .C2(n18585), .A(n18573), .B(n18572), .ZN(
        P3_U2935) );
  AOI22_X1 U21644 ( .A1(n18761), .A2(n18580), .B1(n18762), .B2(n18606), .ZN(
        n18575) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18582), .B1(
        n18763), .B2(n18581), .ZN(n18574) );
  OAI211_X1 U21646 ( .C1(n18766), .C2(n18585), .A(n18575), .B(n18574), .ZN(
        P3_U2936) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18582), .B1(
        n18767), .B2(n18580), .ZN(n18577) );
  AOI22_X1 U21648 ( .A1(n18768), .A2(n18581), .B1(n18769), .B2(n18606), .ZN(
        n18576) );
  OAI211_X1 U21649 ( .C1(n18772), .C2(n18585), .A(n18577), .B(n18576), .ZN(
        P3_U2937) );
  AOI22_X1 U21650 ( .A1(n18774), .A2(n18581), .B1(n18773), .B2(n18580), .ZN(
        n18579) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18582), .B1(
        n18775), .B2(n18606), .ZN(n18578) );
  OAI211_X1 U21652 ( .C1(n18778), .C2(n18585), .A(n18579), .B(n18578), .ZN(
        P3_U2938) );
  AOI22_X1 U21653 ( .A1(n18782), .A2(n18581), .B1(n18780), .B2(n18580), .ZN(
        n18584) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18582), .B1(
        n18783), .B2(n18606), .ZN(n18583) );
  OAI211_X1 U21655 ( .C1(n18788), .C2(n18585), .A(n18584), .B(n18583), .ZN(
        P3_U2939) );
  NAND2_X1 U21656 ( .A1(n18586), .A2(n18637), .ZN(n18638) );
  NOR2_X1 U21657 ( .A1(n18587), .A2(n18635), .ZN(n18605) );
  AOI22_X1 U21658 ( .A1(n18739), .A2(n18606), .B1(n18733), .B2(n18605), .ZN(
        n18592) );
  NOR2_X1 U21659 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18588), .ZN(
        n18590) );
  NOR2_X1 U21660 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18635), .ZN(
        n18589) );
  AOI22_X1 U21661 ( .A1(n18738), .A2(n18590), .B1(n18736), .B2(n18589), .ZN(
        n18607) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18607), .B1(
        n18734), .B2(n18629), .ZN(n18591) );
  OAI211_X1 U21663 ( .C1(n18742), .C2(n18638), .A(n18592), .B(n18591), .ZN(
        P3_U2940) );
  AOI22_X1 U21664 ( .A1(n18744), .A2(n18629), .B1(n18743), .B2(n18605), .ZN(
        n18594) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18607), .B1(
        n18745), .B2(n18606), .ZN(n18593) );
  OAI211_X1 U21666 ( .C1(n18748), .C2(n18638), .A(n18594), .B(n18593), .ZN(
        P3_U2941) );
  AOI22_X1 U21667 ( .A1(n18749), .A2(n18605), .B1(n18751), .B2(n18606), .ZN(
        n18596) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18607), .B1(
        n18750), .B2(n18629), .ZN(n18595) );
  OAI211_X1 U21669 ( .C1(n18754), .C2(n18638), .A(n18596), .B(n18595), .ZN(
        P3_U2942) );
  AOI22_X1 U21670 ( .A1(n18757), .A2(n18629), .B1(n18755), .B2(n18605), .ZN(
        n18598) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18607), .B1(
        n18756), .B2(n18606), .ZN(n18597) );
  OAI211_X1 U21672 ( .C1(n18760), .C2(n18638), .A(n18598), .B(n18597), .ZN(
        P3_U2943) );
  AOI22_X1 U21673 ( .A1(n18763), .A2(n18606), .B1(n18761), .B2(n18605), .ZN(
        n18600) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18607), .B1(
        n18762), .B2(n18629), .ZN(n18599) );
  OAI211_X1 U21675 ( .C1(n18766), .C2(n18638), .A(n18600), .B(n18599), .ZN(
        P3_U2944) );
  AOI22_X1 U21676 ( .A1(n18769), .A2(n18629), .B1(n18767), .B2(n18605), .ZN(
        n18602) );
  AOI22_X1 U21677 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18607), .B1(
        n18768), .B2(n18606), .ZN(n18601) );
  OAI211_X1 U21678 ( .C1(n18772), .C2(n18638), .A(n18602), .B(n18601), .ZN(
        P3_U2945) );
  AOI22_X1 U21679 ( .A1(n18773), .A2(n18605), .B1(n18775), .B2(n18629), .ZN(
        n18604) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18607), .B1(
        n18774), .B2(n18606), .ZN(n18603) );
  OAI211_X1 U21681 ( .C1(n18778), .C2(n18638), .A(n18604), .B(n18603), .ZN(
        P3_U2946) );
  AOI22_X1 U21682 ( .A1(n18782), .A2(n18606), .B1(n18780), .B2(n18605), .ZN(
        n18609) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18607), .B1(
        n18783), .B2(n18629), .ZN(n18608) );
  OAI211_X1 U21684 ( .C1(n18788), .C2(n18638), .A(n18609), .B(n18608), .ZN(
        P3_U2947) );
  NAND2_X1 U21685 ( .A1(n18610), .A2(n18637), .ZN(n18633) );
  AOI22_X1 U21686 ( .A1(n18739), .A2(n18629), .B1(n18733), .B2(n18628), .ZN(
        n18615) );
  INV_X1 U21687 ( .A(n18633), .ZN(n18700) );
  AOI221_X1 U21688 ( .B1(n18612), .B2(n18638), .C1(n18611), .C2(n18638), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18613) );
  OAI21_X1 U21689 ( .B1(n18700), .B2(n18613), .A(n18662), .ZN(n18630) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18630), .B1(
        n18734), .B2(n18654), .ZN(n18614) );
  OAI211_X1 U21691 ( .C1(n18742), .C2(n18633), .A(n18615), .B(n18614), .ZN(
        P3_U2948) );
  AOI22_X1 U21692 ( .A1(n18744), .A2(n18654), .B1(n18743), .B2(n18628), .ZN(
        n18617) );
  AOI22_X1 U21693 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18630), .B1(
        n18745), .B2(n18629), .ZN(n18616) );
  OAI211_X1 U21694 ( .C1(n18748), .C2(n18633), .A(n18617), .B(n18616), .ZN(
        P3_U2949) );
  AOI22_X1 U21695 ( .A1(n18749), .A2(n18628), .B1(n18751), .B2(n18629), .ZN(
        n18619) );
  AOI22_X1 U21696 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18630), .B1(
        n18750), .B2(n18654), .ZN(n18618) );
  OAI211_X1 U21697 ( .C1(n18754), .C2(n18633), .A(n18619), .B(n18618), .ZN(
        P3_U2950) );
  AOI22_X1 U21698 ( .A1(n18757), .A2(n18654), .B1(n18755), .B2(n18628), .ZN(
        n18621) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18630), .B1(
        n18756), .B2(n18629), .ZN(n18620) );
  OAI211_X1 U21700 ( .C1(n18760), .C2(n18633), .A(n18621), .B(n18620), .ZN(
        P3_U2951) );
  AOI22_X1 U21701 ( .A1(n18763), .A2(n18629), .B1(n18761), .B2(n18628), .ZN(
        n18623) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18630), .B1(
        n18762), .B2(n18654), .ZN(n18622) );
  OAI211_X1 U21703 ( .C1(n18766), .C2(n18633), .A(n18623), .B(n18622), .ZN(
        P3_U2952) );
  AOI22_X1 U21704 ( .A1(n18768), .A2(n18629), .B1(n18767), .B2(n18628), .ZN(
        n18625) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18630), .B1(
        n18769), .B2(n18654), .ZN(n18624) );
  OAI211_X1 U21706 ( .C1(n18772), .C2(n18633), .A(n18625), .B(n18624), .ZN(
        P3_U2953) );
  AOI22_X1 U21707 ( .A1(n18773), .A2(n18628), .B1(n18775), .B2(n18654), .ZN(
        n18627) );
  AOI22_X1 U21708 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18630), .B1(
        n18774), .B2(n18629), .ZN(n18626) );
  OAI211_X1 U21709 ( .C1(n18778), .C2(n18633), .A(n18627), .B(n18626), .ZN(
        P3_U2954) );
  AOI22_X1 U21710 ( .A1(n18782), .A2(n18629), .B1(n18780), .B2(n18628), .ZN(
        n18632) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18630), .B1(
        n18783), .B2(n18654), .ZN(n18631) );
  OAI211_X1 U21712 ( .C1(n18788), .C2(n18633), .A(n18632), .B(n18631), .ZN(
        P3_U2955) );
  NOR2_X2 U21713 ( .A1(n18634), .A2(n18635), .ZN(n18727) );
  INV_X1 U21714 ( .A(n18727), .ZN(n18658) );
  NOR2_X1 U21715 ( .A1(n18636), .A2(n18635), .ZN(n18684) );
  AND2_X1 U21716 ( .A1(n18732), .A2(n18684), .ZN(n18653) );
  AOI22_X1 U21717 ( .A1(n18739), .A2(n18654), .B1(n18733), .B2(n18653), .ZN(
        n18640) );
  OAI211_X1 U21718 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18738), .A(
        n18736), .B(n18637), .ZN(n18655) );
  INV_X1 U21719 ( .A(n18638), .ZN(n18678) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18655), .B1(
        n18734), .B2(n18678), .ZN(n18639) );
  OAI211_X1 U21721 ( .C1(n18742), .C2(n18658), .A(n18640), .B(n18639), .ZN(
        P3_U2956) );
  AOI22_X1 U21722 ( .A1(n18744), .A2(n18678), .B1(n18743), .B2(n18653), .ZN(
        n18642) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18655), .B1(
        n18745), .B2(n18654), .ZN(n18641) );
  OAI211_X1 U21724 ( .C1(n18748), .C2(n18658), .A(n18642), .B(n18641), .ZN(
        P3_U2957) );
  AOI22_X1 U21725 ( .A1(n18749), .A2(n18653), .B1(n18751), .B2(n18654), .ZN(
        n18644) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18655), .B1(
        n18750), .B2(n18678), .ZN(n18643) );
  OAI211_X1 U21727 ( .C1(n18754), .C2(n18658), .A(n18644), .B(n18643), .ZN(
        P3_U2958) );
  AOI22_X1 U21728 ( .A1(n18757), .A2(n18678), .B1(n18755), .B2(n18653), .ZN(
        n18646) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18655), .B1(
        n18756), .B2(n18654), .ZN(n18645) );
  OAI211_X1 U21730 ( .C1(n18760), .C2(n18658), .A(n18646), .B(n18645), .ZN(
        P3_U2959) );
  AOI22_X1 U21731 ( .A1(n18763), .A2(n18654), .B1(n18761), .B2(n18653), .ZN(
        n18648) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18655), .B1(
        n18762), .B2(n18678), .ZN(n18647) );
  OAI211_X1 U21733 ( .C1(n18766), .C2(n18658), .A(n18648), .B(n18647), .ZN(
        P3_U2960) );
  AOI22_X1 U21734 ( .A1(n18769), .A2(n18678), .B1(n18767), .B2(n18653), .ZN(
        n18650) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18655), .B1(
        n18768), .B2(n18654), .ZN(n18649) );
  OAI211_X1 U21736 ( .C1(n18772), .C2(n18658), .A(n18650), .B(n18649), .ZN(
        P3_U2961) );
  AOI22_X1 U21737 ( .A1(n18773), .A2(n18653), .B1(n18775), .B2(n18678), .ZN(
        n18652) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18655), .B1(
        n18774), .B2(n18654), .ZN(n18651) );
  OAI211_X1 U21739 ( .C1(n18778), .C2(n18658), .A(n18652), .B(n18651), .ZN(
        P3_U2962) );
  AOI22_X1 U21740 ( .A1(n18782), .A2(n18654), .B1(n18780), .B2(n18653), .ZN(
        n18657) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18655), .B1(
        n18783), .B2(n18678), .ZN(n18656) );
  OAI211_X1 U21742 ( .C1(n18788), .C2(n18658), .A(n18657), .B(n18656), .ZN(
        P3_U2963) );
  INV_X1 U21743 ( .A(n18737), .ZN(n18683) );
  NOR2_X2 U21744 ( .A1(n18683), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18781) );
  INV_X1 U21745 ( .A(n18781), .ZN(n18682) );
  NOR2_X1 U21746 ( .A1(n18727), .A2(n18781), .ZN(n18709) );
  OAI21_X1 U21747 ( .B1(n18660), .B2(n18659), .A(n18709), .ZN(n18661) );
  OAI211_X1 U21748 ( .C1(n18781), .C2(n18963), .A(n18662), .B(n18661), .ZN(
        n18679) );
  NOR2_X1 U21749 ( .A1(n18860), .A2(n18709), .ZN(n18677) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18679), .B1(
        n18733), .B2(n18677), .ZN(n18664) );
  AOI22_X1 U21751 ( .A1(n18739), .A2(n18678), .B1(n18734), .B2(n18700), .ZN(
        n18663) );
  OAI211_X1 U21752 ( .C1(n18742), .C2(n18682), .A(n18664), .B(n18663), .ZN(
        P3_U2964) );
  AOI22_X1 U21753 ( .A1(n18745), .A2(n18678), .B1(n18743), .B2(n18677), .ZN(
        n18666) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18679), .B1(
        n18744), .B2(n18700), .ZN(n18665) );
  OAI211_X1 U21755 ( .C1(n18748), .C2(n18682), .A(n18666), .B(n18665), .ZN(
        P3_U2965) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18679), .B1(
        n18749), .B2(n18677), .ZN(n18668) );
  AOI22_X1 U21757 ( .A1(n18750), .A2(n18700), .B1(n18751), .B2(n18678), .ZN(
        n18667) );
  OAI211_X1 U21758 ( .C1(n18754), .C2(n18682), .A(n18668), .B(n18667), .ZN(
        P3_U2966) );
  AOI22_X1 U21759 ( .A1(n18756), .A2(n18678), .B1(n18755), .B2(n18677), .ZN(
        n18670) );
  AOI22_X1 U21760 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18679), .B1(
        n18757), .B2(n18700), .ZN(n18669) );
  OAI211_X1 U21761 ( .C1(n18760), .C2(n18682), .A(n18670), .B(n18669), .ZN(
        P3_U2967) );
  AOI22_X1 U21762 ( .A1(n18763), .A2(n18678), .B1(n18761), .B2(n18677), .ZN(
        n18672) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18679), .B1(
        n18762), .B2(n18700), .ZN(n18671) );
  OAI211_X1 U21764 ( .C1(n18766), .C2(n18682), .A(n18672), .B(n18671), .ZN(
        P3_U2968) );
  AOI22_X1 U21765 ( .A1(n18769), .A2(n18700), .B1(n18767), .B2(n18677), .ZN(
        n18674) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18679), .B1(
        n18768), .B2(n18678), .ZN(n18673) );
  OAI211_X1 U21767 ( .C1(n18772), .C2(n18682), .A(n18674), .B(n18673), .ZN(
        P3_U2969) );
  AOI22_X1 U21768 ( .A1(n18773), .A2(n18677), .B1(n18775), .B2(n18700), .ZN(
        n18676) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18679), .B1(
        n18774), .B2(n18678), .ZN(n18675) );
  OAI211_X1 U21770 ( .C1(n18778), .C2(n18682), .A(n18676), .B(n18675), .ZN(
        P3_U2970) );
  AOI22_X1 U21771 ( .A1(n18782), .A2(n18678), .B1(n18780), .B2(n18677), .ZN(
        n18681) );
  AOI22_X1 U21772 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18679), .B1(
        n18783), .B2(n18700), .ZN(n18680) );
  OAI211_X1 U21773 ( .C1(n18788), .C2(n18682), .A(n18681), .B(n18680), .ZN(
        P3_U2971) );
  NOR2_X1 U21774 ( .A1(n18860), .A2(n18683), .ZN(n18699) );
  AOI22_X1 U21775 ( .A1(n18733), .A2(n18699), .B1(n18734), .B2(n18727), .ZN(
        n18686) );
  AOI22_X1 U21776 ( .A1(n18738), .A2(n18684), .B1(n18737), .B2(n18736), .ZN(
        n18701) );
  AOI22_X1 U21777 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18701), .B1(
        n18739), .B2(n18700), .ZN(n18685) );
  OAI211_X1 U21778 ( .C1(n18704), .C2(n18742), .A(n18686), .B(n18685), .ZN(
        P3_U2972) );
  AOI22_X1 U21779 ( .A1(n18745), .A2(n18700), .B1(n18743), .B2(n18699), .ZN(
        n18688) );
  AOI22_X1 U21780 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18701), .B1(
        n18744), .B2(n18727), .ZN(n18687) );
  OAI211_X1 U21781 ( .C1(n18704), .C2(n18748), .A(n18688), .B(n18687), .ZN(
        P3_U2973) );
  AOI22_X1 U21782 ( .A1(n18750), .A2(n18727), .B1(n18749), .B2(n18699), .ZN(
        n18690) );
  AOI22_X1 U21783 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18701), .B1(
        n18751), .B2(n18700), .ZN(n18689) );
  OAI211_X1 U21784 ( .C1(n18704), .C2(n18754), .A(n18690), .B(n18689), .ZN(
        P3_U2974) );
  AOI22_X1 U21785 ( .A1(n18756), .A2(n18700), .B1(n18755), .B2(n18699), .ZN(
        n18692) );
  AOI22_X1 U21786 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18701), .B1(
        n18757), .B2(n18727), .ZN(n18691) );
  OAI211_X1 U21787 ( .C1(n18704), .C2(n18760), .A(n18692), .B(n18691), .ZN(
        P3_U2975) );
  AOI22_X1 U21788 ( .A1(n18763), .A2(n18700), .B1(n18761), .B2(n18699), .ZN(
        n18694) );
  AOI22_X1 U21789 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18701), .B1(
        n18762), .B2(n18727), .ZN(n18693) );
  OAI211_X1 U21790 ( .C1(n18704), .C2(n18766), .A(n18694), .B(n18693), .ZN(
        P3_U2976) );
  AOI22_X1 U21791 ( .A1(n18769), .A2(n18727), .B1(n18767), .B2(n18699), .ZN(
        n18696) );
  AOI22_X1 U21792 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18701), .B1(
        n18768), .B2(n18700), .ZN(n18695) );
  OAI211_X1 U21793 ( .C1(n18704), .C2(n18772), .A(n18696), .B(n18695), .ZN(
        P3_U2977) );
  AOI22_X1 U21794 ( .A1(n18774), .A2(n18700), .B1(n18773), .B2(n18699), .ZN(
        n18698) );
  AOI22_X1 U21795 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18701), .B1(
        n18775), .B2(n18727), .ZN(n18697) );
  OAI211_X1 U21796 ( .C1(n18704), .C2(n18778), .A(n18698), .B(n18697), .ZN(
        P3_U2978) );
  AOI22_X1 U21797 ( .A1(n18783), .A2(n18727), .B1(n18780), .B2(n18699), .ZN(
        n18703) );
  AOI22_X1 U21798 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18701), .B1(
        n18782), .B2(n18700), .ZN(n18702) );
  OAI211_X1 U21799 ( .C1(n18704), .C2(n18788), .A(n18703), .B(n18702), .ZN(
        P3_U2979) );
  INV_X1 U21800 ( .A(n18705), .ZN(n18706) );
  NOR2_X1 U21801 ( .A1(n18860), .A2(n18706), .ZN(n18726) );
  AOI22_X1 U21802 ( .A1(n18739), .A2(n18727), .B1(n18733), .B2(n18726), .ZN(
        n18713) );
  OAI22_X1 U21803 ( .A1(n18709), .A2(n18708), .B1(n18707), .B2(n18706), .ZN(
        n18710) );
  OAI21_X1 U21804 ( .B1(n18711), .B2(n18963), .A(n18710), .ZN(n18728) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18728), .B1(
        n18734), .B2(n18781), .ZN(n18712) );
  OAI211_X1 U21806 ( .C1(n18742), .C2(n18731), .A(n18713), .B(n18712), .ZN(
        P3_U2980) );
  AOI22_X1 U21807 ( .A1(n18744), .A2(n18781), .B1(n18743), .B2(n18726), .ZN(
        n18715) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18728), .B1(
        n18745), .B2(n18727), .ZN(n18714) );
  OAI211_X1 U21809 ( .C1(n18731), .C2(n18748), .A(n18715), .B(n18714), .ZN(
        P3_U2981) );
  AOI22_X1 U21810 ( .A1(n18749), .A2(n18726), .B1(n18751), .B2(n18727), .ZN(
        n18717) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18728), .B1(
        n18750), .B2(n18781), .ZN(n18716) );
  OAI211_X1 U21812 ( .C1(n18731), .C2(n18754), .A(n18717), .B(n18716), .ZN(
        P3_U2982) );
  AOI22_X1 U21813 ( .A1(n18757), .A2(n18781), .B1(n18755), .B2(n18726), .ZN(
        n18719) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18728), .B1(
        n18756), .B2(n18727), .ZN(n18718) );
  OAI211_X1 U21815 ( .C1(n18731), .C2(n18760), .A(n18719), .B(n18718), .ZN(
        P3_U2983) );
  AOI22_X1 U21816 ( .A1(n18763), .A2(n18727), .B1(n18761), .B2(n18726), .ZN(
        n18721) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18728), .B1(
        n18762), .B2(n18781), .ZN(n18720) );
  OAI211_X1 U21818 ( .C1(n18731), .C2(n18766), .A(n18721), .B(n18720), .ZN(
        P3_U2984) );
  AOI22_X1 U21819 ( .A1(n18769), .A2(n18781), .B1(n18767), .B2(n18726), .ZN(
        n18723) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18728), .B1(
        n18768), .B2(n18727), .ZN(n18722) );
  OAI211_X1 U21821 ( .C1(n18731), .C2(n18772), .A(n18723), .B(n18722), .ZN(
        P3_U2985) );
  AOI22_X1 U21822 ( .A1(n18773), .A2(n18726), .B1(n18775), .B2(n18781), .ZN(
        n18725) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18728), .B1(
        n18774), .B2(n18727), .ZN(n18724) );
  OAI211_X1 U21824 ( .C1(n18731), .C2(n18778), .A(n18725), .B(n18724), .ZN(
        P3_U2986) );
  AOI22_X1 U21825 ( .A1(n18782), .A2(n18727), .B1(n18780), .B2(n18726), .ZN(
        n18730) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18728), .B1(
        n18783), .B2(n18781), .ZN(n18729) );
  OAI211_X1 U21827 ( .C1(n18731), .C2(n18788), .A(n18730), .B(n18729), .ZN(
        P3_U2987) );
  AND2_X1 U21828 ( .A1(n18732), .A2(n18735), .ZN(n18779) );
  AOI22_X1 U21829 ( .A1(n18784), .A2(n18734), .B1(n18733), .B2(n18779), .ZN(
        n18741) );
  AOI22_X1 U21830 ( .A1(n18738), .A2(n18737), .B1(n18736), .B2(n18735), .ZN(
        n18785) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18785), .B1(
        n18739), .B2(n18781), .ZN(n18740) );
  OAI211_X1 U21832 ( .C1(n18789), .C2(n18742), .A(n18741), .B(n18740), .ZN(
        P3_U2988) );
  AOI22_X1 U21833 ( .A1(n18784), .A2(n18744), .B1(n18743), .B2(n18779), .ZN(
        n18747) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18785), .B1(
        n18745), .B2(n18781), .ZN(n18746) );
  OAI211_X1 U21835 ( .C1(n18789), .C2(n18748), .A(n18747), .B(n18746), .ZN(
        P3_U2989) );
  AOI22_X1 U21836 ( .A1(n18784), .A2(n18750), .B1(n18749), .B2(n18779), .ZN(
        n18753) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18785), .B1(
        n18751), .B2(n18781), .ZN(n18752) );
  OAI211_X1 U21838 ( .C1(n18789), .C2(n18754), .A(n18753), .B(n18752), .ZN(
        P3_U2990) );
  AOI22_X1 U21839 ( .A1(n18756), .A2(n18781), .B1(n18755), .B2(n18779), .ZN(
        n18759) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18785), .B1(
        n18784), .B2(n18757), .ZN(n18758) );
  OAI211_X1 U21841 ( .C1(n18789), .C2(n18760), .A(n18759), .B(n18758), .ZN(
        P3_U2991) );
  AOI22_X1 U21842 ( .A1(n18784), .A2(n18762), .B1(n18761), .B2(n18779), .ZN(
        n18765) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18785), .B1(
        n18763), .B2(n18781), .ZN(n18764) );
  OAI211_X1 U21844 ( .C1(n18789), .C2(n18766), .A(n18765), .B(n18764), .ZN(
        P3_U2992) );
  AOI22_X1 U21845 ( .A1(n18768), .A2(n18781), .B1(n18767), .B2(n18779), .ZN(
        n18771) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18785), .B1(
        n18784), .B2(n18769), .ZN(n18770) );
  OAI211_X1 U21847 ( .C1(n18789), .C2(n18772), .A(n18771), .B(n18770), .ZN(
        P3_U2993) );
  AOI22_X1 U21848 ( .A1(n18774), .A2(n18781), .B1(n18773), .B2(n18779), .ZN(
        n18777) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18785), .B1(
        n18784), .B2(n18775), .ZN(n18776) );
  OAI211_X1 U21850 ( .C1(n18789), .C2(n18778), .A(n18777), .B(n18776), .ZN(
        P3_U2994) );
  AOI22_X1 U21851 ( .A1(n18782), .A2(n18781), .B1(n18780), .B2(n18779), .ZN(
        n18787) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18785), .B1(
        n18784), .B2(n18783), .ZN(n18786) );
  OAI211_X1 U21853 ( .C1(n18789), .C2(n18788), .A(n18787), .B(n18786), .ZN(
        P3_U2995) );
  NOR2_X1 U21854 ( .A1(n18822), .A2(n18790), .ZN(n18796) );
  AOI21_X1 U21855 ( .B1(n18793), .B2(n18792), .A(n18791), .ZN(n18794) );
  OAI22_X1 U21856 ( .A1(n18797), .A2(n18796), .B1(n18795), .B2(n18794), .ZN(
        n19007) );
  INV_X1 U21857 ( .A(n18798), .ZN(n18801) );
  AOI22_X1 U21858 ( .A1(n18979), .A2(n18799), .B1(n18825), .B2(n18812), .ZN(
        n18800) );
  OAI21_X1 U21859 ( .B1(n18819), .B2(n18801), .A(n18800), .ZN(n18968) );
  NOR2_X1 U21860 ( .A1(n18969), .A2(n18968), .ZN(n18807) );
  NAND2_X1 U21861 ( .A1(n18802), .A2(n18994), .ZN(n18810) );
  INV_X1 U21862 ( .A(n18810), .ZN(n18803) );
  OAI22_X1 U21863 ( .A1(n18805), .A2(n18804), .B1(n18803), .B2(n18825), .ZN(
        n18964) );
  AOI21_X1 U21864 ( .B1(n18964), .B2(n18832), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18806) );
  AOI21_X1 U21865 ( .B1(n18832), .B2(n18807), .A(n18806), .ZN(n18839) );
  NAND2_X1 U21866 ( .A1(n18809), .A2(n18808), .ZN(n18811) );
  AOI22_X1 U21867 ( .A1(n18983), .A2(n18811), .B1(n18986), .B2(n18810), .ZN(
        n18980) );
  AOI22_X1 U21868 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18812), .B1(
        n18811), .B2(n18994), .ZN(n18987) );
  AOI222_X1 U21869 ( .A1(n18980), .A2(n18987), .B1(n18980), .B2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C1(n18987), .C2(n18813), .ZN(
        n18815) );
  AOI21_X1 U21870 ( .B1(n18815), .B2(n18832), .A(n18814), .ZN(n18834) );
  AOI21_X1 U21871 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18817), .A(
        n18816), .ZN(n18831) );
  INV_X1 U21872 ( .A(n18818), .ZN(n18824) );
  OAI21_X1 U21873 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18820), .A(
        n18819), .ZN(n18823) );
  AOI22_X1 U21874 ( .A1(n18824), .A2(n18823), .B1(n18822), .B2(n18821), .ZN(
        n18829) );
  NAND3_X1 U21875 ( .A1(n18827), .A2(n18826), .A3(n18825), .ZN(n18828) );
  OAI211_X1 U21876 ( .C1(n18831), .C2(n18830), .A(n18829), .B(n18828), .ZN(
        n18977) );
  AOI22_X1 U21877 ( .A1(n18846), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18977), .B2(n18832), .ZN(n18835) );
  OR2_X1 U21878 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18835), .ZN(
        n18833) );
  AOI221_X1 U21879 ( .B1(n18834), .B2(n18833), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n18835), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18838) );
  OAI21_X1 U21880 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18835), .ZN(n18837) );
  AOI222_X1 U21881 ( .A1(n18839), .A2(n18838), .B1(n18839), .B2(n18837), .C1(
        n18838), .C2(n18836), .ZN(n18843) );
  OAI21_X1 U21882 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18840), .ZN(n18842) );
  NAND4_X1 U21883 ( .A1(n18844), .A2(n18843), .A3(n18842), .A4(n18841), .ZN(
        n18845) );
  AOI211_X1 U21884 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18846), .A(
        n19007), .B(n18845), .ZN(n18857) );
  AOI22_X1 U21885 ( .A1(n18988), .A2(n19018), .B1(n18858), .B2(n19011), .ZN(
        n18847) );
  INV_X1 U21886 ( .A(n18847), .ZN(n18853) );
  NAND2_X1 U21887 ( .A1(n19014), .A2(n18848), .ZN(n18849) );
  OAI211_X1 U21888 ( .C1(n18850), .C2(n18849), .A(n19009), .B(n18857), .ZN(
        n18962) );
  OAI21_X1 U21889 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19015), .A(n18962), 
        .ZN(n18861) );
  NOR2_X1 U21890 ( .A1(n18851), .A2(n18861), .ZN(n18852) );
  MUX2_X1 U21891 ( .A(n18853), .B(n18852), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18855) );
  OAI211_X1 U21892 ( .C1(n18857), .C2(n18856), .A(n18855), .B(n18854), .ZN(
        P3_U2996) );
  NAND2_X1 U21893 ( .A1(n18858), .A2(n19011), .ZN(n18865) );
  NOR4_X1 U21894 ( .A1(n18859), .A2(n18972), .A3(n19015), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18868) );
  INV_X1 U21895 ( .A(n18868), .ZN(n18864) );
  OR3_X1 U21896 ( .A1(n18862), .A2(n18861), .A3(n18860), .ZN(n18863) );
  NAND4_X1 U21897 ( .A1(n18866), .A2(n18865), .A3(n18864), .A4(n18863), .ZN(
        P3_U2997) );
  OAI21_X1 U21898 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18867), .ZN(n18869) );
  AOI21_X1 U21899 ( .B1(n18870), .B2(n18869), .A(n18868), .ZN(P3_U2998) );
  AND2_X1 U21900 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18871), .ZN(
        P3_U2999) );
  AND2_X1 U21901 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18871), .ZN(
        P3_U3000) );
  INV_X1 U21902 ( .A(n18960), .ZN(n18872) );
  AND2_X1 U21903 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18872), .ZN(
        P3_U3001) );
  AND2_X1 U21904 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18871), .ZN(
        P3_U3002) );
  AND2_X1 U21905 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18872), .ZN(
        P3_U3003) );
  AND2_X1 U21906 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18871), .ZN(
        P3_U3004) );
  AND2_X1 U21907 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18872), .ZN(
        P3_U3005) );
  AND2_X1 U21908 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18871), .ZN(
        P3_U3006) );
  AND2_X1 U21909 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18872), .ZN(
        P3_U3007) );
  AND2_X1 U21910 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18871), .ZN(
        P3_U3008) );
  AND2_X1 U21911 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18871), .ZN(
        P3_U3009) );
  AND2_X1 U21912 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18872), .ZN(
        P3_U3010) );
  AND2_X1 U21913 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18872), .ZN(
        P3_U3011) );
  AND2_X1 U21914 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18872), .ZN(
        P3_U3012) );
  AND2_X1 U21915 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18872), .ZN(
        P3_U3013) );
  AND2_X1 U21916 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18872), .ZN(
        P3_U3014) );
  AND2_X1 U21917 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18871), .ZN(
        P3_U3015) );
  AND2_X1 U21918 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18871), .ZN(
        P3_U3016) );
  AND2_X1 U21919 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18871), .ZN(
        P3_U3017) );
  AND2_X1 U21920 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18871), .ZN(
        P3_U3018) );
  AND2_X1 U21921 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18871), .ZN(
        P3_U3019) );
  AND2_X1 U21922 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18871), .ZN(
        P3_U3020) );
  AND2_X1 U21923 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18872), .ZN(P3_U3021) );
  AND2_X1 U21924 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18872), .ZN(P3_U3022) );
  AND2_X1 U21925 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18872), .ZN(P3_U3023) );
  AND2_X1 U21926 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18872), .ZN(P3_U3024) );
  AND2_X1 U21927 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18872), .ZN(P3_U3025) );
  AND2_X1 U21928 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18872), .ZN(P3_U3026) );
  AND2_X1 U21929 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18872), .ZN(P3_U3027) );
  AND2_X1 U21930 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18872), .ZN(P3_U3028) );
  NOR2_X1 U21931 ( .A1(n19015), .A2(n18873), .ZN(n18880) );
  INV_X1 U21932 ( .A(n18880), .ZN(n18882) );
  OAI21_X1 U21933 ( .B1(n18874), .B2(n21248), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18876) );
  INV_X1 U21934 ( .A(NA), .ZN(n21254) );
  NOR3_X1 U21935 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .A3(n21254), .ZN(n18875) );
  AOI21_X1 U21936 ( .B1(n19023), .B2(n18876), .A(n18875), .ZN(n18877) );
  OAI221_X1 U21937 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(P3_STATE_REG_0__SCAN_IN), .C1(P3_STATE_REG_2__SCAN_IN), .C2(n18882), .A(n18877), .ZN(P3_U3029) );
  NAND2_X1 U21938 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n18881) );
  AOI22_X1 U21939 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18881), .B1(HOLD), 
        .B2(n18878), .ZN(n18879) );
  OAI211_X1 U21940 ( .C1(n18879), .C2(n18886), .A(n18882), .B(n19012), .ZN(
        P3_U3030) );
  AOI221_X1 U21941 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18886), .C1(n21254), 
        .C2(n18886), .A(n18880), .ZN(n18887) );
  INV_X1 U21942 ( .A(n18881), .ZN(n18884) );
  OAI22_X1 U21943 ( .A1(NA), .A2(n18882), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18883) );
  OAI22_X1 U21944 ( .A1(n18884), .A2(n18883), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18885) );
  OAI22_X1 U21945 ( .A1(n18887), .A2(n18888), .B1(n18886), .B2(n18885), .ZN(
        P3_U3031) );
  OAI222_X1 U21946 ( .A1(n18996), .A2(n18944), .B1(n18889), .B2(n18955), .C1(
        n18890), .C2(n18947), .ZN(P3_U3032) );
  INV_X1 U21947 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18892) );
  OAI222_X1 U21948 ( .A1(n18947), .A2(n18892), .B1(n18891), .B2(n18955), .C1(
        n18890), .C2(n18951), .ZN(P3_U3033) );
  OAI222_X1 U21949 ( .A1(n18947), .A2(n18894), .B1(n18893), .B2(n18955), .C1(
        n18892), .C2(n18944), .ZN(P3_U3034) );
  OAI222_X1 U21950 ( .A1(n18947), .A2(n18896), .B1(n18895), .B2(n18955), .C1(
        n18894), .C2(n18944), .ZN(P3_U3035) );
  OAI222_X1 U21951 ( .A1(n18947), .A2(n18898), .B1(n18897), .B2(n18955), .C1(
        n18896), .C2(n18944), .ZN(P3_U3036) );
  OAI222_X1 U21952 ( .A1(n18947), .A2(n18900), .B1(n18899), .B2(n18955), .C1(
        n18898), .C2(n18944), .ZN(P3_U3037) );
  OAI222_X1 U21953 ( .A1(n18947), .A2(n18903), .B1(n18901), .B2(n18955), .C1(
        n18900), .C2(n18944), .ZN(P3_U3038) );
  OAI222_X1 U21954 ( .A1(n18903), .A2(n18944), .B1(n18902), .B2(n18955), .C1(
        n18904), .C2(n18947), .ZN(P3_U3039) );
  OAI222_X1 U21955 ( .A1(n18947), .A2(n18906), .B1(n18905), .B2(n18955), .C1(
        n18904), .C2(n18944), .ZN(P3_U3040) );
  OAI222_X1 U21956 ( .A1(n18947), .A2(n18908), .B1(n18907), .B2(n18955), .C1(
        n18906), .C2(n18944), .ZN(P3_U3041) );
  OAI222_X1 U21957 ( .A1(n18947), .A2(n18910), .B1(n18909), .B2(n18955), .C1(
        n18908), .C2(n18944), .ZN(P3_U3042) );
  OAI222_X1 U21958 ( .A1(n18947), .A2(n18912), .B1(n18911), .B2(n18955), .C1(
        n18910), .C2(n18944), .ZN(P3_U3043) );
  OAI222_X1 U21959 ( .A1(n18947), .A2(n18915), .B1(n18913), .B2(n18955), .C1(
        n18912), .C2(n18951), .ZN(P3_U3044) );
  OAI222_X1 U21960 ( .A1(n18915), .A2(n18944), .B1(n18914), .B2(n18955), .C1(
        n18916), .C2(n18947), .ZN(P3_U3045) );
  OAI222_X1 U21961 ( .A1(n18947), .A2(n18918), .B1(n18917), .B2(n18955), .C1(
        n18916), .C2(n18951), .ZN(P3_U3046) );
  OAI222_X1 U21962 ( .A1(n18947), .A2(n18921), .B1(n18919), .B2(n18955), .C1(
        n18918), .C2(n18951), .ZN(P3_U3047) );
  OAI222_X1 U21963 ( .A1(n18921), .A2(n18944), .B1(n18920), .B2(n18955), .C1(
        n18922), .C2(n18947), .ZN(P3_U3048) );
  INV_X1 U21964 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18924) );
  OAI222_X1 U21965 ( .A1(n18947), .A2(n18924), .B1(n18923), .B2(n18955), .C1(
        n18922), .C2(n18951), .ZN(P3_U3049) );
  OAI222_X1 U21966 ( .A1(n18947), .A2(n18926), .B1(n18925), .B2(n18955), .C1(
        n18924), .C2(n18951), .ZN(P3_U3050) );
  OAI222_X1 U21967 ( .A1(n18947), .A2(n18928), .B1(n18927), .B2(n18955), .C1(
        n18926), .C2(n18951), .ZN(P3_U3051) );
  OAI222_X1 U21968 ( .A1(n18947), .A2(n18930), .B1(n18929), .B2(n18955), .C1(
        n18928), .C2(n18951), .ZN(P3_U3052) );
  OAI222_X1 U21969 ( .A1(n18947), .A2(n18933), .B1(n18931), .B2(n18955), .C1(
        n18930), .C2(n18944), .ZN(P3_U3053) );
  OAI222_X1 U21970 ( .A1(n18933), .A2(n18944), .B1(n18932), .B2(n18955), .C1(
        n18934), .C2(n18947), .ZN(P3_U3054) );
  OAI222_X1 U21971 ( .A1(n18947), .A2(n18936), .B1(n18935), .B2(n18955), .C1(
        n18934), .C2(n18951), .ZN(P3_U3055) );
  OAI222_X1 U21972 ( .A1(n18947), .A2(n18938), .B1(n18937), .B2(n18955), .C1(
        n18936), .C2(n18944), .ZN(P3_U3056) );
  OAI222_X1 U21973 ( .A1(n18947), .A2(n18940), .B1(n18939), .B2(n18955), .C1(
        n18938), .C2(n18944), .ZN(P3_U3057) );
  OAI222_X1 U21974 ( .A1(n18947), .A2(n18943), .B1(n18941), .B2(n18955), .C1(
        n18940), .C2(n18944), .ZN(P3_U3058) );
  OAI222_X1 U21975 ( .A1(n18943), .A2(n18944), .B1(n18942), .B2(n18955), .C1(
        n18945), .C2(n18947), .ZN(P3_U3059) );
  OAI222_X1 U21976 ( .A1(n18947), .A2(n18950), .B1(n18946), .B2(n18955), .C1(
        n18945), .C2(n18944), .ZN(P3_U3060) );
  INV_X1 U21977 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18949) );
  OAI222_X1 U21978 ( .A1(n18951), .A2(n18950), .B1(n18949), .B2(n18955), .C1(
        n18948), .C2(n18947), .ZN(P3_U3061) );
  OAI22_X1 U21979 ( .A1(n19023), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18955), .ZN(n18952) );
  INV_X1 U21980 ( .A(n18952), .ZN(P3_U3274) );
  OAI22_X1 U21981 ( .A1(n19023), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18955), .ZN(n18953) );
  INV_X1 U21982 ( .A(n18953), .ZN(P3_U3275) );
  OAI22_X1 U21983 ( .A1(n19023), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18955), .ZN(n18954) );
  INV_X1 U21984 ( .A(n18954), .ZN(P3_U3276) );
  OAI22_X1 U21985 ( .A1(n19023), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18955), .ZN(n18956) );
  INV_X1 U21986 ( .A(n18956), .ZN(P3_U3277) );
  OAI21_X1 U21987 ( .B1(n18960), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18958), 
        .ZN(n18957) );
  INV_X1 U21988 ( .A(n18957), .ZN(P3_U3280) );
  OAI21_X1 U21989 ( .B1(n18960), .B2(n18959), .A(n18958), .ZN(P3_U3281) );
  OAI221_X1 U21990 ( .B1(n18963), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18963), 
        .C2(n18962), .A(n18961), .ZN(P3_U3282) );
  NOR2_X1 U21991 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18967), .ZN(
        n18965) );
  AOI22_X1 U21992 ( .A1(n18988), .A2(n18966), .B1(n18965), .B2(n18964), .ZN(
        n18971) );
  INV_X1 U21993 ( .A(n18967), .ZN(n18990) );
  AOI21_X1 U21994 ( .B1(n18990), .B2(n18968), .A(n18995), .ZN(n18970) );
  OAI22_X1 U21995 ( .A1(n18995), .A2(n18971), .B1(n18970), .B2(n18969), .ZN(
        P3_U3285) );
  NOR2_X1 U21996 ( .A1(n18972), .A2(n18991), .ZN(n18981) );
  OAI22_X1 U21997 ( .A1(n18974), .A2(n18973), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18982) );
  INV_X1 U21998 ( .A(n18982), .ZN(n18976) );
  AOI222_X1 U21999 ( .A1(n18977), .A2(n18990), .B1(n18981), .B2(n18976), .C1(
        n18988), .C2(n18975), .ZN(n18978) );
  AOI22_X1 U22000 ( .A1(n18995), .A2(n18979), .B1(n18978), .B2(n18992), .ZN(
        P3_U3288) );
  INV_X1 U22001 ( .A(n18980), .ZN(n18984) );
  AOI222_X1 U22002 ( .A1(n18984), .A2(n18990), .B1(n18988), .B2(n18983), .C1(
        n18982), .C2(n18981), .ZN(n18985) );
  AOI22_X1 U22003 ( .A1(n18995), .A2(n18986), .B1(n18985), .B2(n18992), .ZN(
        P3_U3289) );
  INV_X1 U22004 ( .A(n18987), .ZN(n18989) );
  AOI222_X1 U22005 ( .A1(n18991), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18990), 
        .B2(n18989), .C1(n18994), .C2(n18988), .ZN(n18993) );
  AOI22_X1 U22006 ( .A1(n18995), .A2(n18994), .B1(n18993), .B2(n18992), .ZN(
        P3_U3290) );
  AOI21_X1 U22007 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18997) );
  AOI22_X1 U22008 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18997), .B2(n18996), .ZN(n18999) );
  INV_X1 U22009 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18998) );
  AOI22_X1 U22010 ( .A1(n19000), .A2(n18999), .B1(n18998), .B2(n19003), .ZN(
        P3_U3292) );
  INV_X1 U22011 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19004) );
  NOR2_X1 U22012 ( .A1(n19003), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19001) );
  AOI22_X1 U22013 ( .A1(n19004), .A2(n19003), .B1(n19002), .B2(n19001), .ZN(
        P3_U3293) );
  INV_X1 U22014 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19005) );
  AOI22_X1 U22015 ( .A1(n18955), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19005), 
        .B2(n19023), .ZN(P3_U3294) );
  MUX2_X1 U22016 ( .A(P3_MORE_REG_SCAN_IN), .B(n19007), .S(n19006), .Z(
        P3_U3295) );
  OAI21_X1 U22017 ( .B1(n19009), .B2(n19008), .A(n19026), .ZN(n19010) );
  AOI21_X1 U22018 ( .B1(n19011), .B2(n19015), .A(n19010), .ZN(n19022) );
  AOI21_X1 U22019 ( .B1(n19014), .B2(n19013), .A(n19012), .ZN(n19016) );
  OAI211_X1 U22020 ( .C1(n19017), .C2(n19016), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19015), .ZN(n19019) );
  AOI21_X1 U22021 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19019), .A(n19018), 
        .ZN(n19021) );
  NAND2_X1 U22022 ( .A1(n19022), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19020) );
  OAI21_X1 U22023 ( .B1(n19022), .B2(n19021), .A(n19020), .ZN(P3_U3296) );
  MUX2_X1 U22024 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .B(P3_M_IO_N_REG_SCAN_IN), 
        .S(n19023), .Z(P3_U3297) );
  OAI21_X1 U22025 ( .B1(n19027), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n19026), 
        .ZN(n19024) );
  OAI21_X1 U22026 ( .B1(n19026), .B2(n19025), .A(n19024), .ZN(P3_U3298) );
  OAI21_X1 U22027 ( .B1(n19027), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n19026), 
        .ZN(n19029) );
  NAND2_X1 U22028 ( .A1(n19029), .A2(n19028), .ZN(P3_U3299) );
  INV_X1 U22029 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19917) );
  NAND2_X1 U22030 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19917), .ZN(n19908) );
  INV_X1 U22031 ( .A(n19908), .ZN(n19030) );
  NOR2_X1 U22032 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19904) );
  AOI21_X1 U22033 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19030), .A(n19904), 
        .ZN(n19899) );
  INV_X1 U22034 ( .A(n19899), .ZN(n19983) );
  AOI21_X1 U22035 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19983), .ZN(n19031) );
  INV_X1 U22036 ( .A(n19031), .ZN(P2_U2815) );
  NOR2_X1 U22037 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19032), .ZN(n19893) );
  AOI22_X1 U22038 ( .A1(n19033), .A2(n19893), .B1(P2_CODEFETCH_REG_SCAN_IN), 
        .B2(n20043), .ZN(n19034) );
  INV_X1 U22039 ( .A(n19034), .ZN(P2_U2816) );
  AOI21_X1 U22040 ( .B1(n19900), .B2(n19917), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19035) );
  AOI22_X1 U22041 ( .A1(n20050), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19035), 
        .B2(n20051), .ZN(P2_U2817) );
  INV_X1 U22042 ( .A(BS16), .ZN(n21075) );
  INV_X1 U22043 ( .A(n19983), .ZN(n19980) );
  AOI21_X1 U22044 ( .B1(n19910), .B2(n21075), .A(n19980), .ZN(n19978) );
  INV_X1 U22045 ( .A(n19978), .ZN(n19981) );
  OAI21_X1 U22046 ( .B1(n19983), .B2(n19629), .A(n19981), .ZN(P2_U2818) );
  NOR4_X1 U22047 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19039) );
  NOR4_X1 U22048 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19038) );
  NOR4_X1 U22049 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19037) );
  NOR4_X1 U22050 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19036) );
  NAND4_X1 U22051 ( .A1(n19039), .A2(n19038), .A3(n19037), .A4(n19036), .ZN(
        n19045) );
  NOR4_X1 U22052 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19043) );
  AOI211_X1 U22053 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19042) );
  NOR4_X1 U22054 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19041) );
  NOR4_X1 U22055 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19040) );
  NAND4_X1 U22056 ( .A1(n19043), .A2(n19042), .A3(n19041), .A4(n19040), .ZN(
        n19044) );
  NOR2_X1 U22057 ( .A1(n19045), .A2(n19044), .ZN(n19055) );
  INV_X1 U22058 ( .A(n19055), .ZN(n19053) );
  NOR2_X1 U22059 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19053), .ZN(n19048) );
  INV_X1 U22060 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19219) );
  INV_X1 U22061 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19046) );
  AOI22_X1 U22062 ( .A1(n19048), .A2(n19219), .B1(n19053), .B2(n19046), .ZN(
        P2_U2820) );
  INV_X1 U22063 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19982) );
  INV_X1 U22064 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19979) );
  NAND3_X1 U22065 ( .A1(n19219), .A2(n19982), .A3(n19979), .ZN(n19052) );
  INV_X1 U22066 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19047) );
  AOI22_X1 U22067 ( .A1(n19048), .A2(n19052), .B1(n19053), .B2(n19047), .ZN(
        P2_U2821) );
  NAND2_X1 U22068 ( .A1(n19048), .A2(n19982), .ZN(n19051) );
  OAI21_X1 U22069 ( .B1(n19219), .B2(n10734), .A(n19055), .ZN(n19049) );
  OAI21_X1 U22070 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19055), .A(n19049), 
        .ZN(n19050) );
  OAI221_X1 U22071 ( .B1(n19051), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19051), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19050), .ZN(P2_U2822) );
  INV_X1 U22072 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19054) );
  OAI221_X1 U22073 ( .B1(n19055), .B2(n19054), .C1(n19053), .C2(n19052), .A(
        n19051), .ZN(P2_U2823) );
  INV_X1 U22074 ( .A(n19228), .ZN(n19107) );
  NOR2_X1 U22075 ( .A1(n19056), .A2(n19202), .ZN(n19061) );
  AOI22_X1 U22076 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19199), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n19168), .ZN(n19058) );
  NAND2_X1 U22077 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19229), .ZN(
        n19057) );
  OAI211_X1 U22078 ( .C1(n19214), .C2(n19059), .A(n19058), .B(n19057), .ZN(
        n19060) );
  AOI211_X1 U22079 ( .C1(n19062), .C2(n19110), .A(n19061), .B(n19060), .ZN(
        n19067) );
  INV_X1 U22080 ( .A(n19063), .ZN(n19064) );
  OAI21_X1 U22081 ( .B1(n19065), .B2(n19068), .A(n19064), .ZN(n19066) );
  OAI211_X1 U22082 ( .C1(n19068), .C2(n19107), .A(n19067), .B(n19066), .ZN(
        P2_U2835) );
  NAND2_X1 U22083 ( .A1(n10206), .A2(n19069), .ZN(n19070) );
  XOR2_X1 U22084 ( .A(n19071), .B(n19070), .Z(n19080) );
  AOI22_X1 U22085 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19229), .B1(
        P2_EBX_REG_19__SCAN_IN), .B2(n19168), .ZN(n19072) );
  OAI21_X1 U22086 ( .B1(n19073), .B2(n19217), .A(n19072), .ZN(n19074) );
  AOI211_X1 U22087 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n19199), .A(n19172), 
        .B(n19074), .ZN(n19079) );
  INV_X1 U22088 ( .A(n19075), .ZN(n19077) );
  AOI22_X1 U22089 ( .A1(n19077), .A2(n19223), .B1(n19076), .B2(n19200), .ZN(
        n19078) );
  OAI211_X1 U22090 ( .C1(n19895), .C2(n19080), .A(n19079), .B(n19078), .ZN(
        P2_U2836) );
  OAI21_X1 U22091 ( .B1(n19948), .B2(n19220), .A(n19181), .ZN(n19084) );
  OAI22_X1 U22092 ( .A1(n19082), .A2(n19217), .B1(n19081), .B2(n19215), .ZN(
        n19083) );
  AOI211_X1 U22093 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19229), .A(
        n19084), .B(n19083), .ZN(n19091) );
  NOR2_X1 U22094 ( .A1(n19206), .A2(n19094), .ZN(n19086) );
  XNOR2_X1 U22095 ( .A(n19086), .B(n19085), .ZN(n19089) );
  INV_X1 U22096 ( .A(n19087), .ZN(n19088) );
  AOI22_X1 U22097 ( .A1(n19089), .A2(n19191), .B1(n19223), .B2(n19088), .ZN(
        n19090) );
  OAI211_X1 U22098 ( .C1(n19092), .C2(n19214), .A(n19091), .B(n19090), .ZN(
        P2_U2837) );
  AOI211_X1 U22099 ( .C1(n19096), .C2(n19095), .A(n19094), .B(n19093), .ZN(
        n19102) );
  NAND2_X1 U22100 ( .A1(n19097), .A2(n19110), .ZN(n19100) );
  AOI22_X1 U22101 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19229), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19168), .ZN(n19099) );
  NAND2_X1 U22102 ( .A1(n19199), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n19098) );
  NAND4_X1 U22103 ( .A1(n19100), .A2(n19099), .A3(n19181), .A4(n19098), .ZN(
        n19101) );
  NOR2_X1 U22104 ( .A1(n19102), .A2(n19101), .ZN(n19106) );
  AOI22_X1 U22105 ( .A1(n19104), .A2(n19223), .B1(n19103), .B2(n19200), .ZN(
        n19105) );
  OAI211_X1 U22106 ( .C1(n19108), .C2(n19107), .A(n19106), .B(n19105), .ZN(
        P2_U2838) );
  INV_X1 U22107 ( .A(n19109), .ZN(n19111) );
  AOI22_X1 U22108 ( .A1(n19111), .A2(n19110), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19229), .ZN(n19112) );
  OAI211_X1 U22109 ( .C1(n19944), .C2(n19220), .A(n19112), .B(n19181), .ZN(
        n19113) );
  AOI21_X1 U22110 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n19168), .A(n19113), .ZN(
        n19120) );
  NOR2_X1 U22111 ( .A1(n19206), .A2(n19114), .ZN(n19116) );
  XNOR2_X1 U22112 ( .A(n19116), .B(n19115), .ZN(n19118) );
  AOI22_X1 U22113 ( .A1(n19118), .A2(n19191), .B1(n19117), .B2(n19223), .ZN(
        n19119) );
  OAI211_X1 U22114 ( .C1(n19121), .C2(n19214), .A(n19120), .B(n19119), .ZN(
        P2_U2839) );
  NAND2_X1 U22115 ( .A1(n10206), .A2(n19122), .ZN(n19123) );
  XOR2_X1 U22116 ( .A(n19124), .B(n19123), .Z(n19131) );
  AOI22_X1 U22117 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19229), .B1(
        P2_EBX_REG_15__SCAN_IN), .B2(n19168), .ZN(n19125) );
  OAI21_X1 U22118 ( .B1(n19126), .B2(n19217), .A(n19125), .ZN(n19127) );
  AOI211_X1 U22119 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19199), .A(n19172), 
        .B(n19127), .ZN(n19130) );
  AOI22_X1 U22120 ( .A1(n19128), .A2(n19223), .B1(n19200), .B2(n19238), .ZN(
        n19129) );
  OAI211_X1 U22121 ( .C1(n19895), .C2(n19131), .A(n19130), .B(n19129), .ZN(
        P2_U2840) );
  NOR2_X1 U22122 ( .A1(n19206), .A2(n19132), .ZN(n19134) );
  XOR2_X1 U22123 ( .A(n19134), .B(n19133), .Z(n19142) );
  AOI22_X1 U22124 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19229), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19168), .ZN(n19135) );
  OAI21_X1 U22125 ( .B1(n19136), .B2(n19217), .A(n19135), .ZN(n19137) );
  AOI211_X1 U22126 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19199), .A(n19328), 
        .B(n19137), .ZN(n19141) );
  AOI22_X1 U22127 ( .A1(n19139), .A2(n19223), .B1(n19200), .B2(n19138), .ZN(
        n19140) );
  OAI211_X1 U22128 ( .C1(n19895), .C2(n19142), .A(n19141), .B(n19140), .ZN(
        P2_U2841) );
  AOI22_X1 U22129 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19229), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n19168), .ZN(n19143) );
  OAI21_X1 U22130 ( .B1(n19144), .B2(n19217), .A(n19143), .ZN(n19145) );
  AOI211_X1 U22131 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19199), .A(n19328), 
        .B(n19145), .ZN(n19153) );
  NOR2_X1 U22132 ( .A1(n19206), .A2(n19146), .ZN(n19148) );
  XNOR2_X1 U22133 ( .A(n19148), .B(n19147), .ZN(n19151) );
  INV_X1 U22134 ( .A(n19149), .ZN(n19150) );
  AOI22_X1 U22135 ( .A1(n19151), .A2(n19191), .B1(n19223), .B2(n19150), .ZN(
        n19152) );
  OAI211_X1 U22136 ( .C1(n19154), .C2(n19214), .A(n19153), .B(n19152), .ZN(
        P2_U2843) );
  OAI22_X1 U22137 ( .A1(n19156), .A2(n19217), .B1(n19155), .B2(n10223), .ZN(
        n19157) );
  INV_X1 U22138 ( .A(n19157), .ZN(n19158) );
  OAI211_X1 U22139 ( .C1(n19933), .C2(n19220), .A(n19158), .B(n19181), .ZN(
        n19159) );
  AOI21_X1 U22140 ( .B1(P2_EBX_REG_10__SCAN_IN), .B2(n19168), .A(n19159), .ZN(
        n19166) );
  NOR2_X1 U22141 ( .A1(n19206), .A2(n19160), .ZN(n19162) );
  XNOR2_X1 U22142 ( .A(n19162), .B(n19161), .ZN(n19164) );
  AOI22_X1 U22143 ( .A1(n19164), .A2(n19191), .B1(n19223), .B2(n19163), .ZN(
        n19165) );
  OAI211_X1 U22144 ( .C1(n19167), .C2(n19214), .A(n19166), .B(n19165), .ZN(
        P2_U2845) );
  AOI22_X1 U22145 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19229), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19168), .ZN(n19169) );
  OAI21_X1 U22146 ( .B1(n19170), .B2(n19217), .A(n19169), .ZN(n19171) );
  AOI211_X1 U22147 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19199), .A(n19172), .B(
        n19171), .ZN(n19179) );
  NOR2_X1 U22148 ( .A1(n19206), .A2(n19173), .ZN(n19175) );
  XNOR2_X1 U22149 ( .A(n19175), .B(n19174), .ZN(n19177) );
  AOI22_X1 U22150 ( .A1(n19177), .A2(n19191), .B1(n19223), .B2(n19176), .ZN(
        n19178) );
  OAI211_X1 U22151 ( .C1(n19180), .C2(n19214), .A(n19179), .B(n19178), .ZN(
        P2_U2847) );
  OAI21_X1 U22152 ( .B1(n19926), .B2(n19220), .A(n19181), .ZN(n19185) );
  INV_X1 U22153 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19182) );
  OAI22_X1 U22154 ( .A1(n19183), .A2(n19217), .B1(n19215), .B2(n19182), .ZN(
        n19184) );
  AOI211_X1 U22155 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19229), .A(
        n19185), .B(n19184), .ZN(n19194) );
  NOR2_X1 U22156 ( .A1(n19206), .A2(n19186), .ZN(n19188) );
  XNOR2_X1 U22157 ( .A(n19188), .B(n19187), .ZN(n19192) );
  INV_X1 U22158 ( .A(n19189), .ZN(n19190) );
  AOI22_X1 U22159 ( .A1(n19192), .A2(n19191), .B1(n19223), .B2(n19190), .ZN(
        n19193) );
  OAI211_X1 U22160 ( .C1(n19214), .C2(n19195), .A(n19194), .B(n19193), .ZN(
        P2_U2849) );
  OAI22_X1 U22161 ( .A1(n19197), .A2(n19217), .B1(n19196), .B2(n19215), .ZN(
        n19198) );
  AOI211_X1 U22162 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19199), .A(n19328), .B(
        n19198), .ZN(n19213) );
  AOI22_X1 U22163 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19229), .B1(
        n19200), .B2(n19260), .ZN(n19212) );
  OAI22_X1 U22164 ( .A1(n19262), .A2(n19203), .B1(n19202), .B2(n19201), .ZN(
        n19204) );
  INV_X1 U22165 ( .A(n19204), .ZN(n19211) );
  INV_X1 U22166 ( .A(n19340), .ZN(n19209) );
  NOR2_X1 U22167 ( .A1(n19206), .A2(n19205), .ZN(n19208) );
  AOI21_X1 U22168 ( .B1(n19209), .B2(n19208), .A(n19895), .ZN(n19207) );
  OAI21_X1 U22169 ( .B1(n19209), .B2(n19208), .A(n19207), .ZN(n19210) );
  NAND4_X1 U22170 ( .A1(n19213), .A2(n19212), .A3(n19211), .A4(n19210), .ZN(
        P2_U2851) );
  OAI22_X1 U22171 ( .A1(n19215), .A2(n11136), .B1(n19214), .B2(n19254), .ZN(
        n19222) );
  INV_X1 U22172 ( .A(n19216), .ZN(n19218) );
  OAI22_X1 U22173 ( .A1(n19220), .A2(n19219), .B1(n19218), .B2(n19217), .ZN(
        n19221) );
  AOI22_X1 U22174 ( .A1(n20017), .A2(n19227), .B1(n19226), .B2(n19225), .ZN(
        n19231) );
  OAI21_X1 U22175 ( .B1(n19229), .B2(n19228), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19230) );
  NAND3_X1 U22176 ( .A1(n19232), .A2(n19231), .A3(n19230), .ZN(P2_U2855) );
  AOI22_X1 U22177 ( .A1(n19234), .A2(n19285), .B1(n19233), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19237) );
  AOI22_X1 U22178 ( .A1(n19235), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19284), .ZN(n19236) );
  NAND2_X1 U22179 ( .A1(n19237), .A2(n19236), .ZN(P2_U2888) );
  INV_X1 U22180 ( .A(n19252), .ZN(n19247) );
  AOI22_X1 U22181 ( .A1(n19247), .A2(n19238), .B1(P2_EAX_REG_15__SCAN_IN), 
        .B2(n19284), .ZN(n19239) );
  OAI21_X1 U22182 ( .B1(n19291), .B2(n19240), .A(n19239), .ZN(P2_U2904) );
  INV_X1 U22183 ( .A(n19291), .ZN(n19242) );
  AOI22_X1 U22184 ( .A1(n19242), .A2(n19241), .B1(P2_EAX_REG_13__SCAN_IN), 
        .B2(n19284), .ZN(n19243) );
  OAI21_X1 U22185 ( .B1(n19252), .B2(n19244), .A(n19243), .ZN(P2_U2906) );
  INV_X1 U22186 ( .A(n19245), .ZN(n19392) );
  AOI22_X1 U22187 ( .A1(n19247), .A2(n19246), .B1(P2_EAX_REG_7__SCAN_IN), .B2(
        n19284), .ZN(n19248) );
  OAI21_X1 U22188 ( .B1(n19392), .B2(n19291), .A(n19248), .ZN(P2_U2912) );
  INV_X1 U22189 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19249) );
  OAI22_X1 U22190 ( .A1(n19252), .A2(n19251), .B1(n19250), .B2(n19249), .ZN(
        n19253) );
  INV_X1 U22191 ( .A(n19253), .ZN(n19259) );
  XOR2_X1 U22192 ( .A(n19266), .B(n19988), .Z(n19269) );
  INV_X1 U22193 ( .A(n19998), .ZN(n19255) );
  XNOR2_X1 U22194 ( .A(n19998), .B(n20000), .ZN(n19275) );
  XOR2_X1 U22195 ( .A(n20003), .B(n19986), .Z(n19280) );
  INV_X1 U22196 ( .A(n19254), .ZN(n19288) );
  NAND2_X1 U22197 ( .A1(n20017), .A2(n19288), .ZN(n19287) );
  NAND2_X1 U22198 ( .A1(n19280), .A2(n19287), .ZN(n19279) );
  OAI21_X1 U22199 ( .B1(n20003), .B2(n19986), .A(n19279), .ZN(n19274) );
  NAND2_X1 U22200 ( .A1(n19275), .A2(n19274), .ZN(n19273) );
  OAI21_X1 U22201 ( .B1(n20000), .B2(n19255), .A(n19273), .ZN(n19268) );
  NAND2_X1 U22202 ( .A1(n19269), .A2(n19268), .ZN(n19267) );
  NAND2_X1 U22203 ( .A1(n19988), .A2(n19266), .ZN(n19256) );
  AOI21_X1 U22204 ( .B1(n19267), .B2(n19256), .A(n19260), .ZN(n19261) );
  OR3_X1 U22205 ( .A1(n19261), .A2(n19262), .A3(n19257), .ZN(n19258) );
  OAI211_X1 U22206 ( .C1(n19381), .C2(n19291), .A(n19259), .B(n19258), .ZN(
        P2_U2914) );
  AOI22_X1 U22207 ( .A1(n19285), .A2(n19260), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19284), .ZN(n19265) );
  XOR2_X1 U22208 ( .A(n19262), .B(n19261), .Z(n19263) );
  NAND2_X1 U22209 ( .A1(n19263), .A2(n19286), .ZN(n19264) );
  OAI211_X1 U22210 ( .C1(n19374), .C2(n19291), .A(n19265), .B(n19264), .ZN(
        P2_U2915) );
  INV_X1 U22211 ( .A(n19266), .ZN(n19991) );
  AOI22_X1 U22212 ( .A1(n19285), .A2(n19991), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19284), .ZN(n19272) );
  OAI21_X1 U22213 ( .B1(n19269), .B2(n19268), .A(n19267), .ZN(n19270) );
  NAND2_X1 U22214 ( .A1(n19270), .A2(n19286), .ZN(n19271) );
  OAI211_X1 U22215 ( .C1(n19368), .C2(n19291), .A(n19272), .B(n19271), .ZN(
        P2_U2916) );
  AOI22_X1 U22216 ( .A1(n20000), .A2(n19285), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19284), .ZN(n19278) );
  OAI21_X1 U22217 ( .B1(n19275), .B2(n19274), .A(n19273), .ZN(n19276) );
  NAND2_X1 U22218 ( .A1(n19276), .A2(n19286), .ZN(n19277) );
  OAI211_X1 U22219 ( .C1(n19362), .C2(n19291), .A(n19278), .B(n19277), .ZN(
        P2_U2917) );
  AOI22_X1 U22220 ( .A1(n19285), .A2(n20003), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19284), .ZN(n19283) );
  OAI21_X1 U22221 ( .B1(n19280), .B2(n19287), .A(n19279), .ZN(n19281) );
  NAND2_X1 U22222 ( .A1(n19281), .A2(n19286), .ZN(n19282) );
  OAI211_X1 U22223 ( .C1(n19357), .C2(n19291), .A(n19283), .B(n19282), .ZN(
        P2_U2918) );
  AOI22_X1 U22224 ( .A1(n19285), .A2(n19288), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19284), .ZN(n19290) );
  OAI211_X1 U22225 ( .C1(n20017), .C2(n19288), .A(n19287), .B(n19286), .ZN(
        n19289) );
  OAI211_X1 U22226 ( .C1(n19292), .C2(n19291), .A(n19290), .B(n19289), .ZN(
        P2_U2919) );
  AND2_X1 U22227 ( .A1(n19312), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  INV_X1 U22228 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19295) );
  AOI22_X1 U22229 ( .A1(n20047), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19294) );
  OAI21_X1 U22230 ( .B1(n19295), .B2(n19326), .A(n19294), .ZN(P2_U2936) );
  AOI22_X1 U22231 ( .A1(n20047), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19296) );
  OAI21_X1 U22232 ( .B1(n19297), .B2(n19326), .A(n19296), .ZN(P2_U2937) );
  AOI22_X1 U22233 ( .A1(n20047), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19298) );
  OAI21_X1 U22234 ( .B1(n19299), .B2(n19326), .A(n19298), .ZN(P2_U2938) );
  AOI22_X1 U22235 ( .A1(n20047), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19300) );
  OAI21_X1 U22236 ( .B1(n19301), .B2(n19326), .A(n19300), .ZN(P2_U2939) );
  AOI22_X1 U22237 ( .A1(n20047), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19312), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19302) );
  OAI21_X1 U22238 ( .B1(n19303), .B2(n19326), .A(n19302), .ZN(P2_U2940) );
  AOI22_X1 U22239 ( .A1(n20047), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19312), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19304) );
  OAI21_X1 U22240 ( .B1(n19305), .B2(n19326), .A(n19304), .ZN(P2_U2941) );
  AOI22_X1 U22241 ( .A1(n20047), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19312), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19306) );
  OAI21_X1 U22242 ( .B1(n19307), .B2(n19326), .A(n19306), .ZN(P2_U2942) );
  AOI22_X1 U22243 ( .A1(n20047), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19312), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19308) );
  OAI21_X1 U22244 ( .B1(n19309), .B2(n19326), .A(n19308), .ZN(P2_U2943) );
  INV_X1 U22245 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19311) );
  AOI22_X1 U22246 ( .A1(n20047), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19312), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19310) );
  OAI21_X1 U22247 ( .B1(n19311), .B2(n19326), .A(n19310), .ZN(P2_U2944) );
  AOI22_X1 U22248 ( .A1(n20047), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19312), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19313) );
  OAI21_X1 U22249 ( .B1(n19314), .B2(n19326), .A(n19313), .ZN(P2_U2945) );
  AOI22_X1 U22250 ( .A1(n20047), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19315) );
  OAI21_X1 U22251 ( .B1(n19249), .B2(n19326), .A(n19315), .ZN(P2_U2946) );
  INV_X1 U22252 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19317) );
  AOI22_X1 U22253 ( .A1(n20047), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19316) );
  OAI21_X1 U22254 ( .B1(n19317), .B2(n19326), .A(n19316), .ZN(P2_U2947) );
  INV_X1 U22255 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19319) );
  AOI22_X1 U22256 ( .A1(n20047), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19318) );
  OAI21_X1 U22257 ( .B1(n19319), .B2(n19326), .A(n19318), .ZN(P2_U2948) );
  INV_X1 U22258 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19321) );
  AOI22_X1 U22259 ( .A1(n20047), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19320) );
  OAI21_X1 U22260 ( .B1(n19321), .B2(n19326), .A(n19320), .ZN(P2_U2949) );
  INV_X1 U22261 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19323) );
  AOI22_X1 U22262 ( .A1(n20047), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19322) );
  OAI21_X1 U22263 ( .B1(n19323), .B2(n19326), .A(n19322), .ZN(P2_U2950) );
  INV_X1 U22264 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19327) );
  AOI22_X1 U22265 ( .A1(n20047), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19324), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19325) );
  OAI21_X1 U22266 ( .B1(n19327), .B2(n19326), .A(n19325), .ZN(P2_U2951) );
  AOI22_X1 U22267 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19329), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19328), .ZN(n19339) );
  INV_X1 U22268 ( .A(n19330), .ZN(n19334) );
  OAI22_X1 U22269 ( .A1(n19334), .A2(n19333), .B1(n19332), .B2(n19331), .ZN(
        n19335) );
  AOI21_X1 U22270 ( .B1(n19337), .B2(n19336), .A(n19335), .ZN(n19338) );
  OAI211_X1 U22271 ( .C1(n19341), .C2(n19340), .A(n19339), .B(n19338), .ZN(
        P2_U3010) );
  NOR2_X2 U22272 ( .A1(n19759), .A2(n19788), .ZN(n19885) );
  NOR3_X2 U22273 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19455), .ZN(n19391) );
  AOI22_X1 U22274 ( .A1(n19840), .A2(n19885), .B1(n19832), .B2(n19391), .ZN(
        n19355) );
  OAI21_X1 U22275 ( .B1(n19885), .B2(n19413), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19344) );
  NAND2_X1 U22276 ( .A1(n19344), .A2(n19990), .ZN(n19353) );
  INV_X1 U22277 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19995) );
  NOR2_X1 U22278 ( .A1(n19345), .A2(n19995), .ZN(n19880) );
  NOR2_X1 U22279 ( .A1(n19880), .A2(n19391), .ZN(n19352) );
  INV_X1 U22280 ( .A(n19352), .ZN(n19349) );
  INV_X1 U22281 ( .A(n19391), .ZN(n19346) );
  OAI211_X1 U22282 ( .C1(n19347), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19346), 
        .B(n19599), .ZN(n19348) );
  OAI211_X1 U22283 ( .C1(n19353), .C2(n19349), .A(n19833), .B(n19348), .ZN(
        n19394) );
  OAI21_X1 U22284 ( .B1(n19350), .B2(n19391), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19351) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19394), .B1(
        n14132), .B2(n19393), .ZN(n19354) );
  OAI211_X1 U22286 ( .C1(n19843), .C2(n19424), .A(n19355), .B(n19354), .ZN(
        P2_U3048) );
  AOI22_X1 U22287 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19389), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19388), .ZN(n19767) );
  AOI22_X1 U22288 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19389), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19388), .ZN(n19848) );
  NOR2_X2 U22289 ( .A1(n19356), .A2(n19390), .ZN(n19844) );
  AOI22_X1 U22290 ( .A1(n19764), .A2(n19885), .B1(n19844), .B2(n19391), .ZN(
        n19360) );
  AOI22_X1 U22291 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19394), .B1(
        n19358), .B2(n19393), .ZN(n19359) );
  OAI211_X1 U22292 ( .C1(n19767), .C2(n19424), .A(n19360), .B(n19359), .ZN(
        P2_U3049) );
  AOI22_X1 U22293 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19389), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19388), .ZN(n19771) );
  AOI22_X1 U22294 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19388), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19389), .ZN(n19853) );
  INV_X1 U22295 ( .A(n19853), .ZN(n19768) );
  NOR2_X2 U22296 ( .A1(n19361), .A2(n19390), .ZN(n19849) );
  AOI22_X1 U22297 ( .A1(n19768), .A2(n19885), .B1(n19849), .B2(n19391), .ZN(
        n19365) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19394), .B1(
        n19363), .B2(n19393), .ZN(n19364) );
  OAI211_X1 U22299 ( .C1(n19771), .C2(n19424), .A(n19365), .B(n19364), .ZN(
        P2_U3050) );
  AOI22_X2 U22300 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19389), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19388), .ZN(n19859) );
  OAI22_X2 U22301 ( .A1(n19367), .A2(n19377), .B1(n19366), .B2(n19379), .ZN(
        n19856) );
  NOR2_X2 U22302 ( .A1(n9819), .A2(n19390), .ZN(n19854) );
  AOI22_X1 U22303 ( .A1(n19856), .A2(n19885), .B1(n19854), .B2(n19391), .ZN(
        n19370) );
  NOR2_X2 U22304 ( .A1(n19368), .A2(n19792), .ZN(n19855) );
  AOI22_X1 U22305 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19394), .B1(
        n19855), .B2(n19393), .ZN(n19369) );
  OAI211_X1 U22306 ( .C1(n19859), .C2(n19424), .A(n19370), .B(n19369), .ZN(
        P2_U3051) );
  AOI22_X1 U22307 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19389), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19388), .ZN(n19812) );
  OAI22_X1 U22308 ( .A1(n19372), .A2(n19377), .B1(n19371), .B2(n19379), .ZN(
        n19809) );
  AOI22_X1 U22309 ( .A1(n19809), .A2(n19885), .B1(n19860), .B2(n19391), .ZN(
        n19376) );
  NOR2_X2 U22310 ( .A1(n19374), .A2(n19792), .ZN(n19861) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19394), .B1(
        n19861), .B2(n19393), .ZN(n19375) );
  OAI211_X1 U22312 ( .C1(n19812), .C2(n19424), .A(n19376), .B(n19375), .ZN(
        P2_U3052) );
  OAI22_X1 U22313 ( .A1(n19380), .A2(n19379), .B1(n19378), .B2(n19377), .ZN(
        n19776) );
  AOI22_X1 U22314 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19389), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19388), .ZN(n19780) );
  NOR2_X2 U22315 ( .A1(n14575), .A2(n19390), .ZN(n19866) );
  AOI22_X1 U22316 ( .A1(n19868), .A2(n19885), .B1(n19866), .B2(n19391), .ZN(
        n19383) );
  NOR2_X2 U22317 ( .A1(n19381), .A2(n19792), .ZN(n19867) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19394), .B1(
        n19867), .B2(n19393), .ZN(n19382) );
  OAI211_X1 U22319 ( .C1(n19871), .C2(n19424), .A(n19383), .B(n19382), .ZN(
        P2_U3053) );
  AOI22_X1 U22320 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19389), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19388), .ZN(n19819) );
  NOR2_X2 U22321 ( .A1(n19384), .A2(n19390), .ZN(n19872) );
  AOI22_X1 U22322 ( .A1(n19874), .A2(n19885), .B1(n19872), .B2(n19391), .ZN(
        n19387) );
  NOR2_X2 U22323 ( .A1(n19385), .A2(n19792), .ZN(n19873) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19394), .B1(
        n19873), .B2(n19393), .ZN(n19386) );
  OAI211_X1 U22325 ( .C1(n19879), .C2(n19424), .A(n19387), .B(n19386), .ZN(
        P2_U3054) );
  AOI22_X1 U22326 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19389), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19388), .ZN(n19890) );
  NOR2_X2 U22327 ( .A1(n11511), .A2(n19390), .ZN(n19881) );
  AOI22_X1 U22328 ( .A1(n19822), .A2(n19885), .B1(n19881), .B2(n19391), .ZN(
        n19396) );
  NOR2_X2 U22329 ( .A1(n19392), .A2(n19792), .ZN(n19882) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19394), .B1(
        n19882), .B2(n19393), .ZN(n19395) );
  OAI211_X1 U22331 ( .C1(n19827), .C2(n19424), .A(n19396), .B(n19395), .ZN(
        P2_U3055) );
  NAND2_X1 U22332 ( .A1(n19457), .A2(n20011), .ZN(n19400) );
  NOR2_X1 U22333 ( .A1(n19634), .A2(n19455), .ZN(n19419) );
  NOR3_X1 U22334 ( .A1(n19397), .A2(n19419), .A3(n20039), .ZN(n19399) );
  AOI211_X2 U22335 ( .C1(n19400), .C2(n20039), .A(n19398), .B(n19399), .ZN(
        n19420) );
  AOI22_X1 U22336 ( .A1(n19420), .A2(n14132), .B1(n19832), .B2(n19419), .ZN(
        n19404) );
  NAND2_X1 U22337 ( .A1(n19574), .A2(n19639), .ZN(n19401) );
  AOI21_X1 U22338 ( .B1(n19401), .B2(n19400), .A(n19399), .ZN(n19402) );
  OAI211_X1 U22339 ( .C1(n19419), .C2(n20012), .A(n19402), .B(n19833), .ZN(
        n19421) );
  NAND2_X1 U22340 ( .A1(n19639), .A2(n19578), .ZN(n19416) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19421), .B1(
        n19450), .B2(n19760), .ZN(n19403) );
  OAI211_X1 U22342 ( .C1(n19763), .C2(n19424), .A(n19404), .B(n19403), .ZN(
        P2_U3056) );
  AOI22_X1 U22343 ( .A1(n19420), .A2(n19358), .B1(n19844), .B2(n19419), .ZN(
        n19406) );
  INV_X1 U22344 ( .A(n19767), .ZN(n19845) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19421), .B1(
        n19450), .B2(n19845), .ZN(n19405) );
  OAI211_X1 U22346 ( .C1(n19848), .C2(n19424), .A(n19406), .B(n19405), .ZN(
        P2_U3057) );
  AOI22_X1 U22347 ( .A1(n19420), .A2(n19363), .B1(n19849), .B2(n19419), .ZN(
        n19408) );
  INV_X1 U22348 ( .A(n19771), .ZN(n19850) );
  AOI22_X1 U22349 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19421), .B1(
        n19450), .B2(n19850), .ZN(n19407) );
  OAI211_X1 U22350 ( .C1(n19853), .C2(n19424), .A(n19408), .B(n19407), .ZN(
        P2_U3058) );
  AOI22_X1 U22351 ( .A1(n19420), .A2(n19855), .B1(n19854), .B2(n19419), .ZN(
        n19410) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19421), .B1(
        n19413), .B2(n19856), .ZN(n19409) );
  OAI211_X1 U22353 ( .C1(n19859), .C2(n19416), .A(n19410), .B(n19409), .ZN(
        P2_U3059) );
  AOI22_X1 U22354 ( .A1(n19420), .A2(n19861), .B1(n19860), .B2(n19419), .ZN(
        n19412) );
  INV_X1 U22355 ( .A(n19812), .ZN(n19862) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19421), .B1(
        n19450), .B2(n19862), .ZN(n19411) );
  OAI211_X1 U22357 ( .C1(n19865), .C2(n19424), .A(n19412), .B(n19411), .ZN(
        P2_U3060) );
  AOI22_X1 U22358 ( .A1(n19420), .A2(n19867), .B1(n19866), .B2(n19419), .ZN(
        n19415) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19421), .B1(
        n19413), .B2(n19868), .ZN(n19414) );
  OAI211_X1 U22360 ( .C1(n19871), .C2(n19416), .A(n19415), .B(n19414), .ZN(
        P2_U3061) );
  AOI22_X1 U22361 ( .A1(n19420), .A2(n19873), .B1(n19872), .B2(n19419), .ZN(
        n19418) );
  INV_X1 U22362 ( .A(n19879), .ZN(n19815) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19421), .B1(
        n19450), .B2(n19815), .ZN(n19417) );
  OAI211_X1 U22364 ( .C1(n19819), .C2(n19424), .A(n19418), .B(n19417), .ZN(
        P2_U3062) );
  AOI22_X1 U22365 ( .A1(n19420), .A2(n19882), .B1(n19881), .B2(n19419), .ZN(
        n19423) );
  INV_X1 U22366 ( .A(n19827), .ZN(n19884) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19421), .B1(
        n19450), .B2(n19884), .ZN(n19422) );
  OAI211_X1 U22368 ( .C1(n19890), .C2(n19424), .A(n19423), .B(n19422), .ZN(
        P2_U3063) );
  NOR2_X1 U22369 ( .A1(n19670), .A2(n19455), .ZN(n19448) );
  OAI21_X1 U22370 ( .B1(n19425), .B2(n19448), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19426) );
  NAND2_X1 U22371 ( .A1(n19457), .A2(n19669), .ZN(n19429) );
  NAND2_X1 U22372 ( .A1(n19426), .A2(n19429), .ZN(n19449) );
  AOI22_X1 U22373 ( .A1(n19449), .A2(n14132), .B1(n19832), .B2(n19448), .ZN(
        n19435) );
  INV_X1 U22374 ( .A(n19448), .ZN(n19427) );
  OAI21_X1 U22375 ( .B1(n19428), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19427), 
        .ZN(n19432) );
  OAI21_X1 U22376 ( .B1(n19483), .B2(n19450), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19430) );
  NAND2_X1 U22377 ( .A1(n19430), .A2(n19429), .ZN(n19431) );
  MUX2_X1 U22378 ( .A(n19432), .B(n19431), .S(n19990), .Z(n19433) );
  NAND2_X1 U22379 ( .A1(n19433), .A2(n19833), .ZN(n19451) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19451), .B1(
        n19450), .B2(n19840), .ZN(n19434) );
  OAI211_X1 U22381 ( .C1(n19843), .C2(n19479), .A(n19435), .B(n19434), .ZN(
        P2_U3064) );
  AOI22_X1 U22382 ( .A1(n19449), .A2(n19358), .B1(n19844), .B2(n19448), .ZN(
        n19437) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19451), .B1(
        n19450), .B2(n19764), .ZN(n19436) );
  OAI211_X1 U22384 ( .C1(n19767), .C2(n19479), .A(n19437), .B(n19436), .ZN(
        P2_U3065) );
  AOI22_X1 U22385 ( .A1(n19449), .A2(n19363), .B1(n19849), .B2(n19448), .ZN(
        n19439) );
  AOI22_X1 U22386 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19451), .B1(
        n19450), .B2(n19768), .ZN(n19438) );
  OAI211_X1 U22387 ( .C1(n19771), .C2(n19479), .A(n19439), .B(n19438), .ZN(
        P2_U3066) );
  AOI22_X1 U22388 ( .A1(n19449), .A2(n19855), .B1(n19854), .B2(n19448), .ZN(
        n19441) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19451), .B1(
        n19450), .B2(n19856), .ZN(n19440) );
  OAI211_X1 U22390 ( .C1(n19859), .C2(n19479), .A(n19441), .B(n19440), .ZN(
        P2_U3067) );
  AOI22_X1 U22391 ( .A1(n19449), .A2(n19861), .B1(n10033), .B2(n19448), .ZN(
        n19443) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19451), .B1(
        n19450), .B2(n19809), .ZN(n19442) );
  OAI211_X1 U22393 ( .C1(n19812), .C2(n19479), .A(n19443), .B(n19442), .ZN(
        P2_U3068) );
  AOI22_X1 U22394 ( .A1(n19449), .A2(n19867), .B1(n19866), .B2(n19448), .ZN(
        n19445) );
  AOI22_X1 U22395 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19451), .B1(
        n19450), .B2(n19868), .ZN(n19444) );
  OAI211_X1 U22396 ( .C1(n19871), .C2(n19479), .A(n19445), .B(n19444), .ZN(
        P2_U3069) );
  AOI22_X1 U22397 ( .A1(n19449), .A2(n19873), .B1(n19872), .B2(n19448), .ZN(
        n19447) );
  AOI22_X1 U22398 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19451), .B1(
        n19450), .B2(n19874), .ZN(n19446) );
  OAI211_X1 U22399 ( .C1(n19879), .C2(n19479), .A(n19447), .B(n19446), .ZN(
        P2_U3070) );
  AOI22_X1 U22400 ( .A1(n19449), .A2(n19882), .B1(n19881), .B2(n19448), .ZN(
        n19453) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19451), .B1(
        n19450), .B2(n19822), .ZN(n19452) );
  OAI211_X1 U22402 ( .C1(n19827), .C2(n19479), .A(n19453), .B(n19452), .ZN(
        P2_U3071) );
  NOR2_X1 U22403 ( .A1(n19455), .A2(n19454), .ZN(n19482) );
  AOI22_X1 U22404 ( .A1(n19840), .A2(n19483), .B1(n19832), .B2(n19482), .ZN(
        n19468) );
  INV_X1 U22405 ( .A(n19482), .ZN(n19456) );
  OAI21_X1 U22406 ( .B1(n10945), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19456), 
        .ZN(n19459) );
  NAND2_X1 U22407 ( .A1(n19574), .A2(n19984), .ZN(n19463) );
  NAND2_X1 U22408 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19457), .ZN(
        n19461) );
  NAND2_X1 U22409 ( .A1(n19463), .A2(n19461), .ZN(n19458) );
  MUX2_X1 U22410 ( .A(n19459), .B(n19458), .S(n19990), .Z(n19460) );
  NAND2_X1 U22411 ( .A1(n19460), .A2(n19833), .ZN(n19485) );
  INV_X1 U22412 ( .A(n19461), .ZN(n19462) );
  NAND3_X1 U22413 ( .A1(n19463), .A2(n19990), .A3(n19462), .ZN(n19466) );
  OAI21_X1 U22414 ( .B1(n19464), .B2(n19482), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19465) );
  NAND2_X1 U22415 ( .A1(n19466), .A2(n19465), .ZN(n19484) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19485), .B1(
        n14132), .B2(n19484), .ZN(n19467) );
  OAI211_X1 U22417 ( .C1(n19843), .C2(n19491), .A(n19468), .B(n19467), .ZN(
        P2_U3072) );
  AOI22_X1 U22418 ( .A1(n19845), .A2(n19513), .B1(n19482), .B2(n19844), .ZN(
        n19470) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19485), .B1(
        n19358), .B2(n19484), .ZN(n19469) );
  OAI211_X1 U22420 ( .C1(n19848), .C2(n19479), .A(n19470), .B(n19469), .ZN(
        P2_U3073) );
  AOI22_X1 U22421 ( .A1(n19768), .A2(n19483), .B1(n19482), .B2(n19849), .ZN(
        n19472) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19485), .B1(
        n19363), .B2(n19484), .ZN(n19471) );
  OAI211_X1 U22423 ( .C1(n19771), .C2(n19491), .A(n19472), .B(n19471), .ZN(
        P2_U3074) );
  AOI22_X1 U22424 ( .A1(n19856), .A2(n19483), .B1(n19482), .B2(n19854), .ZN(
        n19474) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19485), .B1(
        n19855), .B2(n19484), .ZN(n19473) );
  OAI211_X1 U22426 ( .C1(n19859), .C2(n19491), .A(n19474), .B(n19473), .ZN(
        P2_U3075) );
  AOI22_X1 U22427 ( .A1(n19809), .A2(n19483), .B1(n19482), .B2(n19860), .ZN(
        n19476) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19485), .B1(
        n19861), .B2(n19484), .ZN(n19475) );
  OAI211_X1 U22429 ( .C1(n19812), .C2(n19491), .A(n19476), .B(n19475), .ZN(
        P2_U3076) );
  AOI22_X1 U22430 ( .A1(n19776), .A2(n19513), .B1(n19482), .B2(n19866), .ZN(
        n19478) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19485), .B1(
        n19867), .B2(n19484), .ZN(n19477) );
  OAI211_X1 U22432 ( .C1(n19780), .C2(n19479), .A(n19478), .B(n19477), .ZN(
        P2_U3077) );
  AOI22_X1 U22433 ( .A1(n19874), .A2(n19483), .B1(n19482), .B2(n19872), .ZN(
        n19481) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19485), .B1(
        n19873), .B2(n19484), .ZN(n19480) );
  OAI211_X1 U22435 ( .C1(n19879), .C2(n19491), .A(n19481), .B(n19480), .ZN(
        P2_U3078) );
  AOI22_X1 U22436 ( .A1(n19822), .A2(n19483), .B1(n19482), .B2(n19881), .ZN(
        n19487) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19485), .B1(
        n19882), .B2(n19484), .ZN(n19486) );
  OAI211_X1 U22438 ( .C1(n19827), .C2(n19491), .A(n19487), .B(n19486), .ZN(
        P2_U3079) );
  NAND3_X1 U22439 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19995), .A3(
        n20011), .ZN(n19521) );
  NOR2_X1 U22440 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19521), .ZN(
        n19511) );
  NOR3_X1 U22441 ( .A1(n19488), .A2(n19511), .A3(n20039), .ZN(n19492) );
  NOR2_X1 U22442 ( .A1(n19489), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19496) );
  AOI21_X1 U22443 ( .B1(n20012), .B2(n19496), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19490) );
  NOR2_X1 U22444 ( .A1(n19492), .A2(n19490), .ZN(n19512) );
  AOI22_X1 U22445 ( .A1(n19512), .A2(n14132), .B1(n19832), .B2(n19511), .ZN(
        n19498) );
  AOI21_X1 U22446 ( .B1(n19491), .B2(n19537), .A(n19629), .ZN(n19495) );
  INV_X1 U22447 ( .A(n19511), .ZN(n19493) );
  AOI211_X1 U22448 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19493), .A(n19792), 
        .B(n19492), .ZN(n19494) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19840), .ZN(n19497) );
  OAI211_X1 U22450 ( .C1(n19843), .C2(n19537), .A(n19498), .B(n19497), .ZN(
        P2_U3080) );
  AOI22_X1 U22451 ( .A1(n19512), .A2(n19358), .B1(n19844), .B2(n19511), .ZN(
        n19500) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19764), .ZN(n19499) );
  OAI211_X1 U22453 ( .C1(n19767), .C2(n19537), .A(n19500), .B(n19499), .ZN(
        P2_U3081) );
  AOI22_X1 U22454 ( .A1(n19512), .A2(n19363), .B1(n19849), .B2(n19511), .ZN(
        n19502) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19768), .ZN(n19501) );
  OAI211_X1 U22456 ( .C1(n19771), .C2(n19537), .A(n19502), .B(n19501), .ZN(
        P2_U3082) );
  AOI22_X1 U22457 ( .A1(n19512), .A2(n19855), .B1(n19854), .B2(n19511), .ZN(
        n19504) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19856), .ZN(n19503) );
  OAI211_X1 U22459 ( .C1(n19859), .C2(n19537), .A(n19504), .B(n19503), .ZN(
        P2_U3083) );
  AOI22_X1 U22460 ( .A1(n19512), .A2(n19861), .B1(n10033), .B2(n19511), .ZN(
        n19506) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19809), .ZN(n19505) );
  OAI211_X1 U22462 ( .C1(n19812), .C2(n19537), .A(n19506), .B(n19505), .ZN(
        P2_U3084) );
  AOI22_X1 U22463 ( .A1(n19512), .A2(n19867), .B1(n19866), .B2(n19511), .ZN(
        n19508) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19868), .ZN(n19507) );
  OAI211_X1 U22465 ( .C1(n19871), .C2(n19537), .A(n19508), .B(n19507), .ZN(
        P2_U3085) );
  AOI22_X1 U22466 ( .A1(n19512), .A2(n19873), .B1(n19872), .B2(n19511), .ZN(
        n19510) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19874), .ZN(n19509) );
  OAI211_X1 U22468 ( .C1(n19879), .C2(n19537), .A(n19510), .B(n19509), .ZN(
        P2_U3086) );
  AOI22_X1 U22469 ( .A1(n19512), .A2(n19882), .B1(n19881), .B2(n19511), .ZN(
        n19516) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19514), .B1(
        n19513), .B2(n19822), .ZN(n19515) );
  OAI211_X1 U22471 ( .C1(n19827), .C2(n19537), .A(n19516), .B(n19515), .ZN(
        P2_U3087) );
  NOR2_X1 U22472 ( .A1(n20020), .A2(n19521), .ZN(n19547) );
  AOI22_X1 U22473 ( .A1(n19760), .A2(n19567), .B1(n19832), .B2(n19547), .ZN(
        n19524) );
  AOI21_X1 U22474 ( .B1(n19756), .B2(n19574), .A(n19599), .ZN(n19519) );
  NOR2_X1 U22475 ( .A1(n19517), .A2(n19547), .ZN(n19520) );
  AOI22_X1 U22476 ( .A1(n19519), .A2(n19521), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19520), .ZN(n19518) );
  OAI211_X1 U22477 ( .C1(n19547), .C2(n20012), .A(n19518), .B(n19833), .ZN(
        n19540) );
  INV_X1 U22478 ( .A(n19519), .ZN(n19522) );
  OAI22_X1 U22479 ( .A1(n19522), .A2(n19521), .B1(n19520), .B2(n20039), .ZN(
        n19539) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19540), .B1(
        n14132), .B2(n19539), .ZN(n19523) );
  OAI211_X1 U22481 ( .C1(n19763), .C2(n19537), .A(n19524), .B(n19523), .ZN(
        P2_U3088) );
  INV_X1 U22482 ( .A(n19537), .ZN(n19538) );
  AOI22_X1 U22483 ( .A1(n19764), .A2(n19538), .B1(n19844), .B2(n19547), .ZN(
        n19526) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19540), .B1(
        n19358), .B2(n19539), .ZN(n19525) );
  OAI211_X1 U22485 ( .C1(n19767), .C2(n19564), .A(n19526), .B(n19525), .ZN(
        P2_U3089) );
  AOI22_X1 U22486 ( .A1(n19850), .A2(n19567), .B1(n19547), .B2(n19849), .ZN(
        n19528) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19540), .B1(
        n19363), .B2(n19539), .ZN(n19527) );
  OAI211_X1 U22488 ( .C1(n19853), .C2(n19537), .A(n19528), .B(n19527), .ZN(
        P2_U3090) );
  AOI22_X1 U22489 ( .A1(n19856), .A2(n19538), .B1(n19547), .B2(n19854), .ZN(
        n19530) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19540), .B1(
        n19855), .B2(n19539), .ZN(n19529) );
  OAI211_X1 U22491 ( .C1(n19859), .C2(n19564), .A(n19530), .B(n19529), .ZN(
        P2_U3091) );
  AOI22_X1 U22492 ( .A1(n19862), .A2(n19567), .B1(n19547), .B2(n19860), .ZN(
        n19532) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19540), .B1(
        n19861), .B2(n19539), .ZN(n19531) );
  OAI211_X1 U22494 ( .C1(n19865), .C2(n19537), .A(n19532), .B(n19531), .ZN(
        P2_U3092) );
  AOI22_X1 U22495 ( .A1(n19776), .A2(n19567), .B1(n19547), .B2(n19866), .ZN(
        n19534) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19540), .B1(
        n19867), .B2(n19539), .ZN(n19533) );
  OAI211_X1 U22497 ( .C1(n19780), .C2(n19537), .A(n19534), .B(n19533), .ZN(
        P2_U3093) );
  AOI22_X1 U22498 ( .A1(n19815), .A2(n19567), .B1(n19547), .B2(n19872), .ZN(
        n19536) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19540), .B1(
        n19873), .B2(n19539), .ZN(n19535) );
  OAI211_X1 U22500 ( .C1(n19819), .C2(n19537), .A(n19536), .B(n19535), .ZN(
        P2_U3094) );
  AOI22_X1 U22501 ( .A1(n19822), .A2(n19538), .B1(n19547), .B2(n19881), .ZN(
        n19542) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19540), .B1(
        n19882), .B2(n19539), .ZN(n19541) );
  OAI211_X1 U22503 ( .C1(n19827), .C2(n19564), .A(n19542), .B(n19541), .ZN(
        P2_U3095) );
  INV_X1 U22504 ( .A(n19577), .ZN(n19573) );
  NOR2_X1 U22505 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19573), .ZN(
        n19565) );
  NOR2_X1 U22506 ( .A1(n19547), .A2(n19565), .ZN(n19544) );
  OR2_X1 U22507 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19544), .ZN(n19545) );
  NOR3_X1 U22508 ( .A1(n10957), .A2(n19565), .A3(n20039), .ZN(n19548) );
  AOI21_X1 U22509 ( .B1(n20039), .B2(n19545), .A(n19548), .ZN(n19566) );
  AOI22_X1 U22510 ( .A1(n19566), .A2(n14132), .B1(n19832), .B2(n19565), .ZN(
        n19551) );
  AOI21_X1 U22511 ( .B1(n19564), .B2(n19591), .A(n19629), .ZN(n19546) );
  AOI221_X1 U22512 ( .B1(n20012), .B2(n19547), .C1(n20012), .C2(n19546), .A(
        n19565), .ZN(n19549) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19568), .B1(
        n19567), .B2(n19840), .ZN(n19550) );
  OAI211_X1 U22514 ( .C1(n19843), .C2(n19591), .A(n19551), .B(n19550), .ZN(
        P2_U3096) );
  AOI22_X1 U22515 ( .A1(n19566), .A2(n19358), .B1(n19844), .B2(n19565), .ZN(
        n19553) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19568), .B1(
        n19595), .B2(n19845), .ZN(n19552) );
  OAI211_X1 U22517 ( .C1(n19848), .C2(n19564), .A(n19553), .B(n19552), .ZN(
        P2_U3097) );
  AOI22_X1 U22518 ( .A1(n19566), .A2(n19363), .B1(n19849), .B2(n19565), .ZN(
        n19555) );
  AOI22_X1 U22519 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19568), .B1(
        n19595), .B2(n19850), .ZN(n19554) );
  OAI211_X1 U22520 ( .C1(n19853), .C2(n19564), .A(n19555), .B(n19554), .ZN(
        P2_U3098) );
  AOI22_X1 U22521 ( .A1(n19566), .A2(n19855), .B1(n19854), .B2(n19565), .ZN(
        n19557) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19568), .B1(
        n19567), .B2(n19856), .ZN(n19556) );
  OAI211_X1 U22523 ( .C1(n19859), .C2(n19591), .A(n19557), .B(n19556), .ZN(
        P2_U3099) );
  AOI22_X1 U22524 ( .A1(n19566), .A2(n19861), .B1(n10033), .B2(n19565), .ZN(
        n19559) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19568), .B1(
        n19595), .B2(n19862), .ZN(n19558) );
  OAI211_X1 U22526 ( .C1(n19865), .C2(n19564), .A(n19559), .B(n19558), .ZN(
        P2_U3100) );
  AOI22_X1 U22527 ( .A1(n19566), .A2(n19867), .B1(n19866), .B2(n19565), .ZN(
        n19561) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19568), .B1(
        n19595), .B2(n19776), .ZN(n19560) );
  OAI211_X1 U22529 ( .C1(n19780), .C2(n19564), .A(n19561), .B(n19560), .ZN(
        P2_U3101) );
  AOI22_X1 U22530 ( .A1(n19566), .A2(n19873), .B1(n19872), .B2(n19565), .ZN(
        n19563) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19568), .B1(
        n19595), .B2(n19815), .ZN(n19562) );
  OAI211_X1 U22532 ( .C1(n19819), .C2(n19564), .A(n19563), .B(n19562), .ZN(
        P2_U3102) );
  AOI22_X1 U22533 ( .A1(n19566), .A2(n19882), .B1(n19881), .B2(n19565), .ZN(
        n19570) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19568), .B1(
        n19567), .B2(n19822), .ZN(n19569) );
  OAI211_X1 U22535 ( .C1(n19827), .C2(n19591), .A(n19570), .B(n19569), .ZN(
        P2_U3103) );
  INV_X1 U22536 ( .A(n19602), .ZN(n19605) );
  OAI21_X1 U22537 ( .B1(n19571), .B2(n19605), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19572) );
  OAI21_X1 U22538 ( .B1(n19573), .B2(n19599), .A(n19572), .ZN(n19594) );
  AOI22_X1 U22539 ( .A1(n19594), .A2(n14132), .B1(n19605), .B2(n19832), .ZN(
        n19580) );
  INV_X1 U22540 ( .A(n19574), .ZN(n19575) );
  NOR2_X1 U22541 ( .A1(n19575), .A2(n19788), .ZN(n19989) );
  OAI211_X1 U22542 ( .C1(n10942), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19602), 
        .B(n19599), .ZN(n19576) );
  OAI211_X1 U22543 ( .C1(n19989), .C2(n19577), .A(n19576), .B(n19833), .ZN(
        n19596) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19596), .B1(
        n19624), .B2(n19760), .ZN(n19579) );
  OAI211_X1 U22545 ( .C1(n19763), .C2(n19591), .A(n19580), .B(n19579), .ZN(
        P2_U3104) );
  AOI22_X1 U22546 ( .A1(n19594), .A2(n19358), .B1(n19605), .B2(n19844), .ZN(
        n19582) );
  AOI22_X1 U22547 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19596), .B1(
        n19624), .B2(n19845), .ZN(n19581) );
  OAI211_X1 U22548 ( .C1(n19848), .C2(n19591), .A(n19582), .B(n19581), .ZN(
        P2_U3105) );
  AOI22_X1 U22549 ( .A1(n19594), .A2(n19363), .B1(n19605), .B2(n19849), .ZN(
        n19584) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19596), .B1(
        n19624), .B2(n19850), .ZN(n19583) );
  OAI211_X1 U22551 ( .C1(n19853), .C2(n19591), .A(n19584), .B(n19583), .ZN(
        P2_U3106) );
  AOI22_X1 U22552 ( .A1(n19594), .A2(n19855), .B1(n19605), .B2(n19854), .ZN(
        n19586) );
  AOI22_X1 U22553 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19596), .B1(
        n19595), .B2(n19856), .ZN(n19585) );
  OAI211_X1 U22554 ( .C1(n19859), .C2(n19618), .A(n19586), .B(n19585), .ZN(
        P2_U3107) );
  AOI22_X1 U22555 ( .A1(n19594), .A2(n19861), .B1(n19605), .B2(n19860), .ZN(
        n19588) );
  AOI22_X1 U22556 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19596), .B1(
        n19624), .B2(n19862), .ZN(n19587) );
  OAI211_X1 U22557 ( .C1(n19865), .C2(n19591), .A(n19588), .B(n19587), .ZN(
        P2_U3108) );
  AOI22_X1 U22558 ( .A1(n19594), .A2(n19867), .B1(n19605), .B2(n19866), .ZN(
        n19590) );
  AOI22_X1 U22559 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19596), .B1(
        n19624), .B2(n19776), .ZN(n19589) );
  OAI211_X1 U22560 ( .C1(n19780), .C2(n19591), .A(n19590), .B(n19589), .ZN(
        P2_U3109) );
  AOI22_X1 U22561 ( .A1(n19594), .A2(n19873), .B1(n19605), .B2(n19872), .ZN(
        n19593) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19596), .B1(
        n19595), .B2(n19874), .ZN(n19592) );
  OAI211_X1 U22563 ( .C1(n19879), .C2(n19618), .A(n19593), .B(n19592), .ZN(
        P2_U3110) );
  AOI22_X1 U22564 ( .A1(n19594), .A2(n19882), .B1(n19605), .B2(n19881), .ZN(
        n19598) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19596), .B1(
        n19595), .B2(n19822), .ZN(n19597) );
  OAI211_X1 U22566 ( .C1(n19827), .C2(n19618), .A(n19598), .B(n19597), .ZN(
        P2_U3111) );
  NAND2_X1 U22567 ( .A1(n20002), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19701) );
  OR2_X1 U22568 ( .A1(n19701), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19643) );
  NOR2_X1 U22569 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19643), .ZN(
        n19623) );
  AOI22_X1 U22570 ( .A1(n19840), .A2(n19624), .B1(n19832), .B2(n19623), .ZN(
        n19609) );
  AOI21_X1 U22571 ( .B1(n19667), .B2(n19618), .A(n19629), .ZN(n19600) );
  NOR2_X1 U22572 ( .A1(n19600), .A2(n19599), .ZN(n19604) );
  OAI21_X1 U22573 ( .B1(n10940), .B2(n20039), .A(n20012), .ZN(n19601) );
  AOI21_X1 U22574 ( .B1(n19604), .B2(n19602), .A(n19601), .ZN(n19603) );
  OAI21_X1 U22575 ( .B1(n19605), .B2(n19623), .A(n19604), .ZN(n19607) );
  OAI21_X1 U22576 ( .B1(n10940), .B2(n19623), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19606) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19626), .B1(
        n14132), .B2(n19625), .ZN(n19608) );
  OAI211_X1 U22578 ( .C1(n19843), .C2(n19667), .A(n19609), .B(n19608), .ZN(
        P2_U3112) );
  AOI22_X1 U22579 ( .A1(n19764), .A2(n19624), .B1(n19844), .B2(n19623), .ZN(
        n19611) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19626), .B1(
        n19625), .B2(n19358), .ZN(n19610) );
  OAI211_X1 U22581 ( .C1(n19767), .C2(n19667), .A(n19611), .B(n19610), .ZN(
        P2_U3113) );
  AOI22_X1 U22582 ( .A1(n19768), .A2(n19624), .B1(n19849), .B2(n19623), .ZN(
        n19613) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19626), .B1(
        n19625), .B2(n19363), .ZN(n19612) );
  OAI211_X1 U22584 ( .C1(n19771), .C2(n19667), .A(n19613), .B(n19612), .ZN(
        P2_U3114) );
  AOI22_X1 U22585 ( .A1(n19856), .A2(n19624), .B1(n19854), .B2(n19623), .ZN(
        n19615) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19626), .B1(
        n19625), .B2(n19855), .ZN(n19614) );
  OAI211_X1 U22587 ( .C1(n19859), .C2(n19667), .A(n19615), .B(n19614), .ZN(
        P2_U3115) );
  AOI22_X1 U22588 ( .A1(n19862), .A2(n19655), .B1(n19860), .B2(n19623), .ZN(
        n19617) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19626), .B1(
        n19625), .B2(n19861), .ZN(n19616) );
  OAI211_X1 U22590 ( .C1(n19865), .C2(n19618), .A(n19617), .B(n19616), .ZN(
        P2_U3116) );
  AOI22_X1 U22591 ( .A1(n19868), .A2(n19624), .B1(n19866), .B2(n19623), .ZN(
        n19620) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19626), .B1(
        n19625), .B2(n19867), .ZN(n19619) );
  OAI211_X1 U22593 ( .C1(n19871), .C2(n19667), .A(n19620), .B(n19619), .ZN(
        P2_U3117) );
  AOI22_X1 U22594 ( .A1(n19874), .A2(n19624), .B1(n19872), .B2(n19623), .ZN(
        n19622) );
  AOI22_X1 U22595 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19626), .B1(
        n19625), .B2(n19873), .ZN(n19621) );
  OAI211_X1 U22596 ( .C1(n19879), .C2(n19667), .A(n19622), .B(n19621), .ZN(
        P2_U3118) );
  AOI22_X1 U22597 ( .A1(n19822), .A2(n19624), .B1(n19881), .B2(n19623), .ZN(
        n19628) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19626), .B1(
        n19625), .B2(n19882), .ZN(n19627) );
  OAI211_X1 U22599 ( .C1(n19827), .C2(n19667), .A(n19628), .B(n19627), .ZN(
        P2_U3119) );
  NOR2_X1 U22600 ( .A1(n19988), .A2(n19629), .ZN(n19837) );
  NAND2_X1 U22601 ( .A1(n19837), .A2(n19639), .ZN(n19630) );
  NAND2_X1 U22602 ( .A1(n19630), .A2(n19990), .ZN(n19644) );
  INV_X1 U22603 ( .A(n19643), .ZN(n19631) );
  OR2_X1 U22604 ( .A1(n19644), .A2(n19631), .ZN(n19638) );
  NAND2_X1 U22605 ( .A1(n19632), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19633) );
  NAND2_X1 U22606 ( .A1(n19633), .A2(n20012), .ZN(n19636) );
  NOR2_X1 U22607 ( .A1(n19634), .A2(n19701), .ZN(n19673) );
  INV_X1 U22608 ( .A(n19673), .ZN(n19635) );
  AOI21_X1 U22609 ( .B1(n19636), .B2(n19635), .A(n19792), .ZN(n19637) );
  INV_X1 U22610 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19647) );
  AOI22_X1 U22611 ( .A1(n19760), .A2(n19693), .B1(n19832), .B2(n19673), .ZN(
        n19646) );
  OAI21_X1 U22612 ( .B1(n19641), .B2(n19673), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19642) );
  OAI21_X1 U22613 ( .B1(n19644), .B2(n19643), .A(n19642), .ZN(n19663) );
  AOI22_X1 U22614 ( .A1(n14132), .A2(n19663), .B1(n19655), .B2(n19840), .ZN(
        n19645) );
  OAI211_X1 U22615 ( .C1(n19650), .C2(n19647), .A(n19646), .B(n19645), .ZN(
        P2_U3120) );
  AOI22_X1 U22616 ( .A1(n19764), .A2(n19655), .B1(n19844), .B2(n19673), .ZN(
        n19649) );
  AOI22_X1 U22617 ( .A1(n19358), .A2(n19663), .B1(n19693), .B2(n19845), .ZN(
        n19648) );
  OAI211_X1 U22618 ( .C1(n19650), .C2(n10826), .A(n19649), .B(n19648), .ZN(
        P2_U3121) );
  AOI22_X1 U22619 ( .A1(n19850), .A2(n19693), .B1(n19849), .B2(n19673), .ZN(
        n19652) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19664), .B1(
        n19363), .B2(n19663), .ZN(n19651) );
  OAI211_X1 U22621 ( .C1(n19853), .C2(n19667), .A(n19652), .B(n19651), .ZN(
        P2_U3122) );
  INV_X1 U22622 ( .A(n19693), .ZN(n19658) );
  AOI22_X1 U22623 ( .A1(n19856), .A2(n19655), .B1(n19854), .B2(n19673), .ZN(
        n19654) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19664), .B1(
        n19855), .B2(n19663), .ZN(n19653) );
  OAI211_X1 U22625 ( .C1(n19859), .C2(n19658), .A(n19654), .B(n19653), .ZN(
        P2_U3123) );
  AOI22_X1 U22626 ( .A1(n19809), .A2(n19655), .B1(n19860), .B2(n19673), .ZN(
        n19657) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19664), .B1(
        n19861), .B2(n19663), .ZN(n19656) );
  OAI211_X1 U22628 ( .C1(n19812), .C2(n19658), .A(n19657), .B(n19656), .ZN(
        P2_U3124) );
  AOI22_X1 U22629 ( .A1(n19776), .A2(n19693), .B1(n19866), .B2(n19673), .ZN(
        n19660) );
  AOI22_X1 U22630 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19664), .B1(
        n19867), .B2(n19663), .ZN(n19659) );
  OAI211_X1 U22631 ( .C1(n19780), .C2(n19667), .A(n19660), .B(n19659), .ZN(
        P2_U3125) );
  AOI22_X1 U22632 ( .A1(n19815), .A2(n19693), .B1(n19872), .B2(n19673), .ZN(
        n19662) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19664), .B1(
        n19873), .B2(n19663), .ZN(n19661) );
  OAI211_X1 U22634 ( .C1(n19819), .C2(n19667), .A(n19662), .B(n19661), .ZN(
        P2_U3126) );
  AOI22_X1 U22635 ( .A1(n19884), .A2(n19693), .B1(n19881), .B2(n19673), .ZN(
        n19666) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19664), .B1(
        n19882), .B2(n19663), .ZN(n19665) );
  OAI211_X1 U22637 ( .C1(n19890), .C2(n19667), .A(n19666), .B(n19665), .ZN(
        P2_U3127) );
  INV_X1 U22638 ( .A(n19669), .ZN(n19672) );
  NOR2_X1 U22639 ( .A1(n19670), .A2(n19701), .ZN(n19691) );
  OAI21_X1 U22640 ( .B1(n10992), .B2(n19691), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19671) );
  OAI21_X1 U22641 ( .B1(n19701), .B2(n19672), .A(n19671), .ZN(n19692) );
  AOI22_X1 U22642 ( .A1(n19692), .A2(n14132), .B1(n19832), .B2(n19691), .ZN(
        n19678) );
  AOI221_X1 U22643 ( .B1(n19721), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19693), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19673), .ZN(n19674) );
  AOI211_X1 U22644 ( .C1(n19675), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19674), .ZN(n19676) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n19840), .ZN(n19677) );
  OAI211_X1 U22646 ( .C1(n19843), .C2(n19729), .A(n19678), .B(n19677), .ZN(
        P2_U3128) );
  AOI22_X1 U22647 ( .A1(n19692), .A2(n19358), .B1(n19844), .B2(n19691), .ZN(
        n19680) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n19764), .ZN(n19679) );
  OAI211_X1 U22649 ( .C1(n19767), .C2(n19729), .A(n19680), .B(n19679), .ZN(
        P2_U3129) );
  AOI22_X1 U22650 ( .A1(n19692), .A2(n19363), .B1(n19849), .B2(n19691), .ZN(
        n19682) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n19768), .ZN(n19681) );
  OAI211_X1 U22652 ( .C1(n19771), .C2(n19729), .A(n19682), .B(n19681), .ZN(
        P2_U3130) );
  AOI22_X1 U22653 ( .A1(n19692), .A2(n19855), .B1(n19854), .B2(n19691), .ZN(
        n19684) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n19856), .ZN(n19683) );
  OAI211_X1 U22655 ( .C1(n19859), .C2(n19729), .A(n19684), .B(n19683), .ZN(
        P2_U3131) );
  AOI22_X1 U22656 ( .A1(n19692), .A2(n19861), .B1(n10033), .B2(n19691), .ZN(
        n19686) );
  AOI22_X1 U22657 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n19809), .ZN(n19685) );
  OAI211_X1 U22658 ( .C1(n19812), .C2(n19729), .A(n19686), .B(n19685), .ZN(
        P2_U3132) );
  AOI22_X1 U22659 ( .A1(n19692), .A2(n19867), .B1(n19866), .B2(n19691), .ZN(
        n19688) );
  AOI22_X1 U22660 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n19868), .ZN(n19687) );
  OAI211_X1 U22661 ( .C1(n19871), .C2(n19729), .A(n19688), .B(n19687), .ZN(
        P2_U3133) );
  AOI22_X1 U22662 ( .A1(n19692), .A2(n19873), .B1(n19872), .B2(n19691), .ZN(
        n19690) );
  AOI22_X1 U22663 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n19874), .ZN(n19689) );
  OAI211_X1 U22664 ( .C1(n19879), .C2(n19729), .A(n19690), .B(n19689), .ZN(
        P2_U3134) );
  AOI22_X1 U22665 ( .A1(n19692), .A2(n19882), .B1(n19881), .B2(n19691), .ZN(
        n19696) );
  AOI22_X1 U22666 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19694), .B1(
        n19693), .B2(n19822), .ZN(n19695) );
  OAI211_X1 U22667 ( .C1(n19827), .C2(n19729), .A(n19696), .B(n19695), .ZN(
        P2_U3135) );
  INV_X1 U22668 ( .A(n19701), .ZN(n19697) );
  NAND2_X1 U22669 ( .A1(n19698), .A2(n19697), .ZN(n19704) );
  AND2_X1 U22670 ( .A1(n19704), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19699) );
  NAND2_X1 U22671 ( .A1(n19700), .A2(n19699), .ZN(n19705) );
  NOR2_X1 U22672 ( .A1(n20011), .A2(n19701), .ZN(n19708) );
  INV_X1 U22673 ( .A(n19708), .ZN(n19702) );
  OAI21_X1 U22674 ( .B1(n19702), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20039), 
        .ZN(n19703) );
  AND2_X1 U22675 ( .A1(n19705), .A2(n19703), .ZN(n19725) );
  INV_X1 U22676 ( .A(n19704), .ZN(n19724) );
  AOI22_X1 U22677 ( .A1(n19725), .A2(n14132), .B1(n19832), .B2(n19724), .ZN(
        n19710) );
  OAI211_X1 U22678 ( .C1(n19724), .C2(n20012), .A(n19705), .B(n19833), .ZN(
        n19706) );
  INV_X1 U22679 ( .A(n19706), .ZN(n19707) );
  OAI221_X1 U22680 ( .B1(n19708), .B2(n19984), .C1(n19708), .C2(n19837), .A(
        n19707), .ZN(n19726) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19726), .B1(
        n19742), .B2(n19760), .ZN(n19709) );
  OAI211_X1 U22682 ( .C1(n19763), .C2(n19729), .A(n19710), .B(n19709), .ZN(
        P2_U3136) );
  AOI22_X1 U22683 ( .A1(n19725), .A2(n19358), .B1(n19844), .B2(n19724), .ZN(
        n19712) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19726), .B1(
        n19721), .B2(n19764), .ZN(n19711) );
  OAI211_X1 U22685 ( .C1(n19767), .C2(n19750), .A(n19712), .B(n19711), .ZN(
        P2_U3137) );
  AOI22_X1 U22686 ( .A1(n19725), .A2(n19363), .B1(n19849), .B2(n19724), .ZN(
        n19714) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19726), .B1(
        n19742), .B2(n19850), .ZN(n19713) );
  OAI211_X1 U22688 ( .C1(n19853), .C2(n19729), .A(n19714), .B(n19713), .ZN(
        P2_U3138) );
  AOI22_X1 U22689 ( .A1(n19725), .A2(n19855), .B1(n19854), .B2(n19724), .ZN(
        n19716) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19726), .B1(
        n19721), .B2(n19856), .ZN(n19715) );
  OAI211_X1 U22691 ( .C1(n19859), .C2(n19750), .A(n19716), .B(n19715), .ZN(
        P2_U3139) );
  AOI22_X1 U22692 ( .A1(n19725), .A2(n19861), .B1(n10033), .B2(n19724), .ZN(
        n19718) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19726), .B1(
        n19721), .B2(n19809), .ZN(n19717) );
  OAI211_X1 U22694 ( .C1(n19812), .C2(n19750), .A(n19718), .B(n19717), .ZN(
        P2_U3140) );
  AOI22_X1 U22695 ( .A1(n19725), .A2(n19867), .B1(n19866), .B2(n19724), .ZN(
        n19720) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19726), .B1(
        n19721), .B2(n19868), .ZN(n19719) );
  OAI211_X1 U22697 ( .C1(n19871), .C2(n19750), .A(n19720), .B(n19719), .ZN(
        P2_U3141) );
  AOI22_X1 U22698 ( .A1(n19725), .A2(n19873), .B1(n19872), .B2(n19724), .ZN(
        n19723) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19726), .B1(
        n19721), .B2(n19874), .ZN(n19722) );
  OAI211_X1 U22700 ( .C1(n19879), .C2(n19750), .A(n19723), .B(n19722), .ZN(
        P2_U3142) );
  AOI22_X1 U22701 ( .A1(n19725), .A2(n19882), .B1(n19881), .B2(n19724), .ZN(
        n19728) );
  AOI22_X1 U22702 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19726), .B1(
        n19742), .B2(n19884), .ZN(n19727) );
  OAI211_X1 U22703 ( .C1(n19890), .C2(n19729), .A(n19728), .B(n19727), .ZN(
        P2_U3143) );
  AOI22_X1 U22704 ( .A1(n19746), .A2(n19358), .B1(n19844), .B2(n19745), .ZN(
        n19731) );
  AOI22_X1 U22705 ( .A1(n19742), .A2(n19764), .B1(n19784), .B2(n19845), .ZN(
        n19730) );
  OAI211_X1 U22706 ( .C1(n19733), .C2(n19732), .A(n19731), .B(n19730), .ZN(
        P2_U3145) );
  AOI22_X1 U22707 ( .A1(n19746), .A2(n19363), .B1(n19849), .B2(n19745), .ZN(
        n19735) );
  AOI22_X1 U22708 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19747), .B1(
        n19784), .B2(n19850), .ZN(n19734) );
  OAI211_X1 U22709 ( .C1(n19853), .C2(n19750), .A(n19735), .B(n19734), .ZN(
        P2_U3146) );
  AOI22_X1 U22710 ( .A1(n19746), .A2(n19855), .B1(n19854), .B2(n19745), .ZN(
        n19737) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19747), .B1(
        n19742), .B2(n19856), .ZN(n19736) );
  OAI211_X1 U22712 ( .C1(n19859), .C2(n19779), .A(n19737), .B(n19736), .ZN(
        P2_U3147) );
  AOI22_X1 U22713 ( .A1(n19746), .A2(n19861), .B1(n10033), .B2(n19745), .ZN(
        n19739) );
  AOI22_X1 U22714 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19747), .B1(
        n19784), .B2(n19862), .ZN(n19738) );
  OAI211_X1 U22715 ( .C1(n19865), .C2(n19750), .A(n19739), .B(n19738), .ZN(
        P2_U3148) );
  AOI22_X1 U22716 ( .A1(n19746), .A2(n19867), .B1(n19866), .B2(n19745), .ZN(
        n19741) );
  AOI22_X1 U22717 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19747), .B1(
        n19784), .B2(n19776), .ZN(n19740) );
  OAI211_X1 U22718 ( .C1(n19780), .C2(n19750), .A(n19741), .B(n19740), .ZN(
        P2_U3149) );
  AOI22_X1 U22719 ( .A1(n19746), .A2(n19873), .B1(n19872), .B2(n19745), .ZN(
        n19744) );
  AOI22_X1 U22720 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19747), .B1(
        n19742), .B2(n19874), .ZN(n19743) );
  OAI211_X1 U22721 ( .C1(n19879), .C2(n19779), .A(n19744), .B(n19743), .ZN(
        P2_U3150) );
  AOI22_X1 U22722 ( .A1(n19746), .A2(n19882), .B1(n19881), .B2(n19745), .ZN(
        n19749) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19747), .B1(
        n19784), .B2(n19884), .ZN(n19748) );
  OAI211_X1 U22724 ( .C1(n19890), .C2(n19750), .A(n19749), .B(n19748), .ZN(
        P2_U3151) );
  NOR2_X1 U22725 ( .A1(n20020), .A2(n19751), .ZN(n19791) );
  NOR3_X1 U22726 ( .A1(n10941), .A2(n19791), .A3(n20039), .ZN(n19753) );
  INV_X1 U22727 ( .A(n19751), .ZN(n19757) );
  AOI21_X1 U22728 ( .B1(n20012), .B2(n19757), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19752) );
  NOR2_X1 U22729 ( .A1(n19753), .A2(n19752), .ZN(n19783) );
  AOI22_X1 U22730 ( .A1(n19783), .A2(n14132), .B1(n19832), .B2(n19791), .ZN(
        n19762) );
  INV_X1 U22731 ( .A(n19791), .ZN(n19754) );
  AOI211_X1 U22732 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19754), .A(n19792), 
        .B(n19753), .ZN(n19755) );
  OAI221_X1 U22733 ( .B1(n19757), .B2(n19756), .C1(n19757), .C2(n19837), .A(
        n19755), .ZN(n19785) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19785), .B1(
        n19821), .B2(n19760), .ZN(n19761) );
  OAI211_X1 U22735 ( .C1(n19763), .C2(n19779), .A(n19762), .B(n19761), .ZN(
        P2_U3152) );
  AOI22_X1 U22736 ( .A1(n19783), .A2(n19358), .B1(n19844), .B2(n19791), .ZN(
        n19766) );
  AOI22_X1 U22737 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19785), .B1(
        n19784), .B2(n19764), .ZN(n19765) );
  OAI211_X1 U22738 ( .C1(n19767), .C2(n19818), .A(n19766), .B(n19765), .ZN(
        P2_U3153) );
  AOI22_X1 U22739 ( .A1(n19783), .A2(n19363), .B1(n19849), .B2(n19791), .ZN(
        n19770) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19785), .B1(
        n19784), .B2(n19768), .ZN(n19769) );
  OAI211_X1 U22741 ( .C1(n19771), .C2(n19818), .A(n19770), .B(n19769), .ZN(
        P2_U3154) );
  AOI22_X1 U22742 ( .A1(n19783), .A2(n19855), .B1(n19854), .B2(n19791), .ZN(
        n19773) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19785), .B1(
        n19784), .B2(n19856), .ZN(n19772) );
  OAI211_X1 U22744 ( .C1(n19859), .C2(n19818), .A(n19773), .B(n19772), .ZN(
        P2_U3155) );
  AOI22_X1 U22745 ( .A1(n19783), .A2(n19861), .B1(n10033), .B2(n19791), .ZN(
        n19775) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19785), .B1(
        n19821), .B2(n19862), .ZN(n19774) );
  OAI211_X1 U22747 ( .C1(n19865), .C2(n19779), .A(n19775), .B(n19774), .ZN(
        P2_U3156) );
  AOI22_X1 U22748 ( .A1(n19783), .A2(n19867), .B1(n19866), .B2(n19791), .ZN(
        n19778) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19785), .B1(
        n19821), .B2(n19776), .ZN(n19777) );
  OAI211_X1 U22750 ( .C1(n19780), .C2(n19779), .A(n19778), .B(n19777), .ZN(
        P2_U3157) );
  AOI22_X1 U22751 ( .A1(n19783), .A2(n19873), .B1(n19872), .B2(n19791), .ZN(
        n19782) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19785), .B1(
        n19784), .B2(n19874), .ZN(n19781) );
  OAI211_X1 U22753 ( .C1(n19879), .C2(n19818), .A(n19782), .B(n19781), .ZN(
        P2_U3158) );
  AOI22_X1 U22754 ( .A1(n19783), .A2(n19882), .B1(n19881), .B2(n19791), .ZN(
        n19787) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19785), .B1(
        n19784), .B2(n19822), .ZN(n19786) );
  OAI211_X1 U22756 ( .C1(n19827), .C2(n19818), .A(n19787), .B(n19786), .ZN(
        P2_U3159) );
  NOR3_X1 U22757 ( .A1(n19995), .A2(n20002), .A3(n20011), .ZN(n19839) );
  INV_X1 U22758 ( .A(n19839), .ZN(n19830) );
  NOR2_X1 U22759 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19830), .ZN(
        n19820) );
  AOI22_X1 U22760 ( .A1(n19840), .A2(n19821), .B1(n19832), .B2(n19820), .ZN(
        n19802) );
  OAI21_X1 U22761 ( .B1(n19875), .B2(n19821), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19790) );
  NAND2_X1 U22762 ( .A1(n19790), .A2(n19990), .ZN(n19800) );
  NOR2_X1 U22763 ( .A1(n19820), .A2(n19791), .ZN(n19799) );
  INV_X1 U22764 ( .A(n19799), .ZN(n19796) );
  OAI21_X1 U22765 ( .B1(n19797), .B2(n20039), .A(n20012), .ZN(n19794) );
  INV_X1 U22766 ( .A(n19820), .ZN(n19793) );
  AOI21_X1 U22767 ( .B1(n19794), .B2(n19793), .A(n19792), .ZN(n19795) );
  OAI21_X1 U22768 ( .B1(n19797), .B2(n19820), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19798) );
  AOI22_X1 U22769 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19824), .B1(
        n14132), .B2(n19823), .ZN(n19801) );
  OAI211_X1 U22770 ( .C1(n19843), .C2(n19889), .A(n19802), .B(n19801), .ZN(
        P2_U3160) );
  AOI22_X1 U22771 ( .A1(n19845), .A2(n19875), .B1(n19844), .B2(n19820), .ZN(
        n19804) );
  AOI22_X1 U22772 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19824), .B1(
        n19358), .B2(n19823), .ZN(n19803) );
  OAI211_X1 U22773 ( .C1(n19848), .C2(n19818), .A(n19804), .B(n19803), .ZN(
        P2_U3161) );
  AOI22_X1 U22774 ( .A1(n19850), .A2(n19875), .B1(n19849), .B2(n19820), .ZN(
        n19806) );
  AOI22_X1 U22775 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19824), .B1(
        n19363), .B2(n19823), .ZN(n19805) );
  OAI211_X1 U22776 ( .C1(n19853), .C2(n19818), .A(n19806), .B(n19805), .ZN(
        P2_U3162) );
  AOI22_X1 U22777 ( .A1(n19856), .A2(n19821), .B1(n19854), .B2(n19820), .ZN(
        n19808) );
  AOI22_X1 U22778 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19824), .B1(
        n19855), .B2(n19823), .ZN(n19807) );
  OAI211_X1 U22779 ( .C1(n19859), .C2(n19889), .A(n19808), .B(n19807), .ZN(
        P2_U3163) );
  AOI22_X1 U22780 ( .A1(n19809), .A2(n19821), .B1(n19860), .B2(n19820), .ZN(
        n19811) );
  AOI22_X1 U22781 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19824), .B1(
        n19861), .B2(n19823), .ZN(n19810) );
  OAI211_X1 U22782 ( .C1(n19812), .C2(n19889), .A(n19811), .B(n19810), .ZN(
        P2_U3164) );
  AOI22_X1 U22783 ( .A1(n19868), .A2(n19821), .B1(n19866), .B2(n19820), .ZN(
        n19814) );
  AOI22_X1 U22784 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19824), .B1(
        n19867), .B2(n19823), .ZN(n19813) );
  OAI211_X1 U22785 ( .C1(n19871), .C2(n19889), .A(n19814), .B(n19813), .ZN(
        P2_U3165) );
  AOI22_X1 U22786 ( .A1(n19815), .A2(n19875), .B1(n19872), .B2(n19820), .ZN(
        n19817) );
  AOI22_X1 U22787 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19824), .B1(
        n19873), .B2(n19823), .ZN(n19816) );
  OAI211_X1 U22788 ( .C1(n19819), .C2(n19818), .A(n19817), .B(n19816), .ZN(
        P2_U3166) );
  AOI22_X1 U22789 ( .A1(n19822), .A2(n19821), .B1(n19881), .B2(n19820), .ZN(
        n19826) );
  AOI22_X1 U22790 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19824), .B1(
        n19882), .B2(n19823), .ZN(n19825) );
  OAI211_X1 U22791 ( .C1(n19827), .C2(n19889), .A(n19826), .B(n19825), .ZN(
        P2_U3167) );
  INV_X1 U22792 ( .A(n19885), .ZN(n19878) );
  NOR2_X1 U22793 ( .A1(n19880), .A2(n20039), .ZN(n19828) );
  NAND2_X1 U22794 ( .A1(n19829), .A2(n19828), .ZN(n19834) );
  OAI21_X1 U22795 ( .B1(n19830), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20039), 
        .ZN(n19831) );
  AND2_X1 U22796 ( .A1(n19834), .A2(n19831), .ZN(n19883) );
  AOI22_X1 U22797 ( .A1(n19883), .A2(n14132), .B1(n19832), .B2(n19880), .ZN(
        n19842) );
  OAI211_X1 U22798 ( .C1(n19880), .C2(n20012), .A(n19834), .B(n19833), .ZN(
        n19835) );
  INV_X1 U22799 ( .A(n19835), .ZN(n19836) );
  OAI221_X1 U22800 ( .B1(n19839), .B2(n19838), .C1(n19839), .C2(n19837), .A(
        n19836), .ZN(n19886) );
  AOI22_X1 U22801 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19886), .B1(
        n19875), .B2(n19840), .ZN(n19841) );
  OAI211_X1 U22802 ( .C1(n19843), .C2(n19878), .A(n19842), .B(n19841), .ZN(
        P2_U3168) );
  AOI22_X1 U22803 ( .A1(n19883), .A2(n19358), .B1(n19844), .B2(n19880), .ZN(
        n19847) );
  AOI22_X1 U22804 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19886), .B1(
        n19885), .B2(n19845), .ZN(n19846) );
  OAI211_X1 U22805 ( .C1(n19848), .C2(n19889), .A(n19847), .B(n19846), .ZN(
        P2_U3169) );
  AOI22_X1 U22806 ( .A1(n19883), .A2(n19363), .B1(n19849), .B2(n19880), .ZN(
        n19852) );
  AOI22_X1 U22807 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19886), .B1(
        n19885), .B2(n19850), .ZN(n19851) );
  OAI211_X1 U22808 ( .C1(n19853), .C2(n19889), .A(n19852), .B(n19851), .ZN(
        P2_U3170) );
  AOI22_X1 U22809 ( .A1(n19883), .A2(n19855), .B1(n19854), .B2(n19880), .ZN(
        n19858) );
  AOI22_X1 U22810 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19886), .B1(
        n19875), .B2(n19856), .ZN(n19857) );
  OAI211_X1 U22811 ( .C1(n19859), .C2(n19878), .A(n19858), .B(n19857), .ZN(
        P2_U3171) );
  AOI22_X1 U22812 ( .A1(n19883), .A2(n19861), .B1(n10033), .B2(n19880), .ZN(
        n19864) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19886), .B1(
        n19885), .B2(n19862), .ZN(n19863) );
  OAI211_X1 U22814 ( .C1(n19865), .C2(n19889), .A(n19864), .B(n19863), .ZN(
        P2_U3172) );
  AOI22_X1 U22815 ( .A1(n19883), .A2(n19867), .B1(n19866), .B2(n19880), .ZN(
        n19870) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19886), .B1(
        n19875), .B2(n19868), .ZN(n19869) );
  OAI211_X1 U22817 ( .C1(n19871), .C2(n19878), .A(n19870), .B(n19869), .ZN(
        P2_U3173) );
  AOI22_X1 U22818 ( .A1(n19883), .A2(n19873), .B1(n19872), .B2(n19880), .ZN(
        n19877) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19886), .B1(
        n19875), .B2(n19874), .ZN(n19876) );
  OAI211_X1 U22820 ( .C1(n19879), .C2(n19878), .A(n19877), .B(n19876), .ZN(
        P2_U3174) );
  AOI22_X1 U22821 ( .A1(n19883), .A2(n19882), .B1(n19881), .B2(n19880), .ZN(
        n19888) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19886), .B1(
        n19885), .B2(n19884), .ZN(n19887) );
  OAI211_X1 U22823 ( .C1(n19890), .C2(n19889), .A(n19888), .B(n19887), .ZN(
        P2_U3175) );
  OAI211_X1 U22824 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20046), .A(n19892), 
        .B(n19891), .ZN(n19897) );
  OAI211_X1 U22825 ( .C1(n19894), .C2(n19893), .A(n20040), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19896) );
  OAI211_X1 U22826 ( .C1(n19898), .C2(n19897), .A(n19896), .B(n19895), .ZN(
        P2_U3177) );
  AND2_X1 U22827 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19980), .ZN(
        P2_U3179) );
  AND2_X1 U22828 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19980), .ZN(
        P2_U3180) );
  AND2_X1 U22829 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19980), .ZN(
        P2_U3181) );
  AND2_X1 U22830 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19980), .ZN(
        P2_U3182) );
  AND2_X1 U22831 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19980), .ZN(
        P2_U3183) );
  AND2_X1 U22832 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19899), .ZN(
        P2_U3184) );
  AND2_X1 U22833 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19899), .ZN(
        P2_U3185) );
  AND2_X1 U22834 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19899), .ZN(
        P2_U3186) );
  AND2_X1 U22835 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19899), .ZN(
        P2_U3187) );
  AND2_X1 U22836 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19899), .ZN(
        P2_U3188) );
  AND2_X1 U22837 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19899), .ZN(
        P2_U3189) );
  AND2_X1 U22838 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19899), .ZN(
        P2_U3190) );
  AND2_X1 U22839 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19899), .ZN(
        P2_U3191) );
  AND2_X1 U22840 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19899), .ZN(
        P2_U3192) );
  AND2_X1 U22841 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19899), .ZN(
        P2_U3193) );
  AND2_X1 U22842 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19899), .ZN(
        P2_U3194) );
  AND2_X1 U22843 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19980), .ZN(
        P2_U3195) );
  AND2_X1 U22844 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19980), .ZN(
        P2_U3196) );
  AND2_X1 U22845 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19980), .ZN(
        P2_U3197) );
  AND2_X1 U22846 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19980), .ZN(
        P2_U3198) );
  AND2_X1 U22847 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19980), .ZN(
        P2_U3199) );
  AND2_X1 U22848 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19980), .ZN(
        P2_U3200) );
  AND2_X1 U22849 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19899), .ZN(P2_U3201) );
  AND2_X1 U22850 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19980), .ZN(P2_U3202) );
  AND2_X1 U22851 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19980), .ZN(P2_U3203) );
  AND2_X1 U22852 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19980), .ZN(P2_U3204) );
  AND2_X1 U22853 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19980), .ZN(P2_U3205) );
  AND2_X1 U22854 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19980), .ZN(P2_U3206) );
  AND2_X1 U22855 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19980), .ZN(P2_U3207) );
  AND2_X1 U22856 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19980), .ZN(P2_U3208) );
  NAND2_X1 U22857 ( .A1(n20040), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19909) );
  INV_X1 U22858 ( .A(n19909), .ZN(n19914) );
  INV_X1 U22859 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19901) );
  NOR3_X1 U22860 ( .A1(n19914), .A2(n19901), .A3(n19900), .ZN(n19903) );
  OAI211_X1 U22861 ( .C1(HOLD), .C2(n19901), .A(n20051), .B(n19910), .ZN(
        n19902) );
  NAND2_X1 U22862 ( .A1(NA), .A2(n19904), .ZN(n19912) );
  OAI211_X1 U22863 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n19903), .A(n19902), 
        .B(n19912), .ZN(P2_U3209) );
  NAND2_X1 U22864 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21248), .ZN(n19913) );
  OAI21_X1 U22865 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n19904), .A(n19913), 
        .ZN(n19905) );
  AOI21_X1 U22866 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n19905), .A(n19914), .ZN(n19907) );
  OAI211_X1 U22867 ( .C1(n21248), .C2(n19908), .A(n19907), .B(n19906), .ZN(
        P2_U3210) );
  OAI22_X1 U22868 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19910), .B1(NA), 
        .B2(n19909), .ZN(n19911) );
  OAI211_X1 U22869 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19911), .ZN(n19916) );
  OAI211_X1 U22870 ( .C1(n19914), .C2(n19913), .A(P2_STATE_REG_2__SCAN_IN), 
        .B(n19912), .ZN(n19915) );
  NAND2_X1 U22871 ( .A1(n19916), .A2(n19915), .ZN(P2_U3211) );
  INV_X1 U22872 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19920) );
  OAI222_X1 U22873 ( .A1(n19974), .A2(n19920), .B1(n19918), .B2(n20050), .C1(
        n10734), .C2(n19972), .ZN(P2_U3212) );
  OAI222_X1 U22874 ( .A1(n19972), .A2(n19920), .B1(n19919), .B2(n20050), .C1(
        n14014), .C2(n19974), .ZN(P2_U3213) );
  INV_X1 U22875 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19922) );
  OAI222_X1 U22876 ( .A1(n19972), .A2(n14014), .B1(n19921), .B2(n20050), .C1(
        n19922), .C2(n19974), .ZN(P2_U3214) );
  OAI222_X1 U22877 ( .A1(n19974), .A2(n19924), .B1(n19923), .B2(n20050), .C1(
        n19922), .C2(n19972), .ZN(P2_U3215) );
  OAI222_X1 U22878 ( .A1(n19974), .A2(n19926), .B1(n19925), .B2(n20050), .C1(
        n19924), .C2(n19972), .ZN(P2_U3216) );
  INV_X1 U22879 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19928) );
  OAI222_X1 U22880 ( .A1(n19974), .A2(n19928), .B1(n19927), .B2(n20050), .C1(
        n19926), .C2(n19972), .ZN(P2_U3217) );
  OAI222_X1 U22881 ( .A1(n19974), .A2(n19930), .B1(n19929), .B2(n20050), .C1(
        n19928), .C2(n19972), .ZN(P2_U3218) );
  OAI222_X1 U22882 ( .A1(n19974), .A2(n14114), .B1(n19931), .B2(n20050), .C1(
        n19930), .C2(n19972), .ZN(P2_U3219) );
  OAI222_X1 U22883 ( .A1(n19974), .A2(n19933), .B1(n19932), .B2(n20050), .C1(
        n14114), .C2(n19972), .ZN(P2_U3220) );
  OAI222_X1 U22884 ( .A1(n19974), .A2(n14082), .B1(n19934), .B2(n20050), .C1(
        n19933), .C2(n19972), .ZN(P2_U3221) );
  OAI222_X1 U22885 ( .A1(n19974), .A2(n19936), .B1(n19935), .B2(n20050), .C1(
        n14082), .C2(n19972), .ZN(P2_U3222) );
  OAI222_X1 U22886 ( .A1(n19974), .A2(n19938), .B1(n19937), .B2(n20050), .C1(
        n19936), .C2(n19972), .ZN(P2_U3223) );
  INV_X1 U22887 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19940) );
  OAI222_X1 U22888 ( .A1(n19974), .A2(n19940), .B1(n19939), .B2(n20050), .C1(
        n19938), .C2(n19972), .ZN(P2_U3224) );
  INV_X1 U22889 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19942) );
  OAI222_X1 U22890 ( .A1(n19974), .A2(n19942), .B1(n19941), .B2(n20050), .C1(
        n19940), .C2(n19972), .ZN(P2_U3225) );
  OAI222_X1 U22891 ( .A1(n19974), .A2(n19944), .B1(n19943), .B2(n20050), .C1(
        n19942), .C2(n19972), .ZN(P2_U3226) );
  OAI222_X1 U22892 ( .A1(n19974), .A2(n19946), .B1(n19945), .B2(n20050), .C1(
        n19944), .C2(n19972), .ZN(P2_U3227) );
  OAI222_X1 U22893 ( .A1(n19974), .A2(n19948), .B1(n19947), .B2(n20050), .C1(
        n19946), .C2(n19972), .ZN(P2_U3228) );
  INV_X1 U22894 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19950) );
  OAI222_X1 U22895 ( .A1(n19974), .A2(n19950), .B1(n19949), .B2(n20050), .C1(
        n19948), .C2(n19972), .ZN(P2_U3229) );
  OAI222_X1 U22896 ( .A1(n19974), .A2(n19952), .B1(n19951), .B2(n20050), .C1(
        n19950), .C2(n19972), .ZN(P2_U3230) );
  OAI222_X1 U22897 ( .A1(n19974), .A2(n19954), .B1(n19953), .B2(n20050), .C1(
        n19952), .C2(n19972), .ZN(P2_U3231) );
  OAI222_X1 U22898 ( .A1(n19974), .A2(n19956), .B1(n19955), .B2(n20050), .C1(
        n19954), .C2(n19972), .ZN(P2_U3232) );
  OAI222_X1 U22899 ( .A1(n19974), .A2(n19958), .B1(n19957), .B2(n20050), .C1(
        n19956), .C2(n19972), .ZN(P2_U3233) );
  OAI222_X1 U22900 ( .A1(n19974), .A2(n19960), .B1(n19959), .B2(n20050), .C1(
        n19958), .C2(n19972), .ZN(P2_U3234) );
  INV_X1 U22901 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19962) );
  OAI222_X1 U22902 ( .A1(n19974), .A2(n19962), .B1(n19961), .B2(n20050), .C1(
        n19960), .C2(n19972), .ZN(P2_U3235) );
  OAI222_X1 U22903 ( .A1(n19974), .A2(n19964), .B1(n19963), .B2(n20050), .C1(
        n19962), .C2(n19972), .ZN(P2_U3236) );
  INV_X1 U22904 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19967) );
  OAI222_X1 U22905 ( .A1(n19974), .A2(n19967), .B1(n19965), .B2(n20050), .C1(
        n19964), .C2(n19972), .ZN(P2_U3237) );
  OAI222_X1 U22906 ( .A1(n19972), .A2(n19967), .B1(n19966), .B2(n20050), .C1(
        n19968), .C2(n19974), .ZN(P2_U3238) );
  INV_X1 U22907 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19970) );
  OAI222_X1 U22908 ( .A1(n19974), .A2(n19970), .B1(n19969), .B2(n20050), .C1(
        n19968), .C2(n19972), .ZN(P2_U3239) );
  OAI222_X1 U22909 ( .A1(n19974), .A2(n11723), .B1(n19971), .B2(n20050), .C1(
        n19970), .C2(n19972), .ZN(P2_U3240) );
  INV_X1 U22910 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19973) );
  OAI222_X1 U22911 ( .A1(n19974), .A2(n15361), .B1(n19973), .B2(n20050), .C1(
        n11723), .C2(n19972), .ZN(P2_U3241) );
  OAI22_X1 U22912 ( .A1(n20051), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20050), .ZN(n19975) );
  INV_X1 U22913 ( .A(n19975), .ZN(P2_U3585) );
  MUX2_X1 U22914 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20051), .Z(P2_U3586) );
  OAI22_X1 U22915 ( .A1(n20051), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20050), .ZN(n19976) );
  INV_X1 U22916 ( .A(n19976), .ZN(P2_U3587) );
  OAI22_X1 U22917 ( .A1(n20051), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20050), .ZN(n19977) );
  INV_X1 U22918 ( .A(n19977), .ZN(P2_U3588) );
  AOI21_X1 U22919 ( .B1(n19980), .B2(n19979), .A(n19978), .ZN(P2_U3591) );
  OAI21_X1 U22920 ( .B1(n19983), .B2(n19982), .A(n19981), .ZN(P2_U3592) );
  NAND2_X1 U22921 ( .A1(n19984), .A2(n20004), .ZN(n19996) );
  NAND3_X1 U22922 ( .A1(n19986), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19985), 
        .ZN(n19987) );
  NAND2_X1 U22923 ( .A1(n19987), .A2(n20016), .ZN(n19997) );
  NAND2_X1 U22924 ( .A1(n19996), .A2(n19997), .ZN(n19993) );
  INV_X1 U22925 ( .A(n19988), .ZN(n19992) );
  AOI222_X1 U22926 ( .A1(n19993), .A2(n19992), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19991), .C1(n19990), .C2(n19989), .ZN(n19994) );
  AOI22_X1 U22927 ( .A1(n20021), .A2(n19995), .B1(n19994), .B2(n20018), .ZN(
        P2_U3602) );
  OAI21_X1 U22928 ( .B1(n19998), .B2(n19997), .A(n19996), .ZN(n19999) );
  AOI21_X1 U22929 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20000), .A(n19999), 
        .ZN(n20001) );
  AOI22_X1 U22930 ( .A1(n20021), .A2(n20002), .B1(n20001), .B2(n20018), .ZN(
        P2_U3603) );
  AOI22_X1 U22931 ( .A1(n20007), .A2(n20004), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20003), .ZN(n20010) );
  INV_X1 U22932 ( .A(n20016), .ZN(n20006) );
  AND2_X1 U22933 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20005) );
  NOR3_X1 U22934 ( .A1(n20007), .A2(n20006), .A3(n20005), .ZN(n20008) );
  NOR2_X1 U22935 ( .A1(n20021), .A2(n20008), .ZN(n20009) );
  AOI22_X1 U22936 ( .A1(n20011), .A2(n20021), .B1(n20010), .B2(n20009), .ZN(
        P2_U3604) );
  NOR2_X1 U22937 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20012), .ZN(
        n20015) );
  INV_X1 U22938 ( .A(n20013), .ZN(n20014) );
  AOI211_X1 U22939 ( .C1(n20017), .C2(n20016), .A(n20015), .B(n20014), .ZN(
        n20019) );
  AOI22_X1 U22940 ( .A1(n20021), .A2(n20020), .B1(n20019), .B2(n20018), .ZN(
        P2_U3605) );
  INV_X1 U22941 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20022) );
  AOI22_X1 U22942 ( .A1(n20050), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20022), 
        .B2(n20051), .ZN(P2_U3608) );
  INV_X1 U22943 ( .A(n20023), .ZN(n20031) );
  INV_X1 U22944 ( .A(n20024), .ZN(n20029) );
  NAND3_X1 U22945 ( .A1(n20027), .A2(n20026), .A3(n20025), .ZN(n20028) );
  OAI211_X1 U22946 ( .C1(n20031), .C2(n20030), .A(n20029), .B(n20028), .ZN(
        n20033) );
  MUX2_X1 U22947 ( .A(P2_MORE_REG_SCAN_IN), .B(n20033), .S(n20032), .Z(
        P2_U3609) );
  OAI21_X1 U22948 ( .B1(n20035), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20034), 
        .ZN(n20036) );
  NAND3_X1 U22949 ( .A1(n20037), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20036), 
        .ZN(n20042) );
  OAI21_X1 U22950 ( .B1(n20040), .B2(n20039), .A(n20038), .ZN(n20041) );
  NAND2_X1 U22951 ( .A1(n20042), .A2(n20041), .ZN(n20049) );
  OAI21_X1 U22952 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20044), .A(n20043), 
        .ZN(n20045) );
  AOI21_X1 U22953 ( .B1(n20047), .B2(n20046), .A(n20045), .ZN(n20048) );
  MUX2_X1 U22954 ( .A(n20049), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n20048), 
        .Z(P2_U3610) );
  OAI22_X1 U22955 ( .A1(n20051), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20050), .ZN(n20052) );
  INV_X1 U22956 ( .A(n20052), .ZN(P2_U3611) );
  AOI21_X1 U22957 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20867), .A(n13417), 
        .ZN(n20054) );
  INV_X1 U22958 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21190) );
  INV_X1 U22959 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20858) );
  NOR2_X1 U22960 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20858), .ZN(n20939) );
  AOI21_X1 U22961 ( .B1(n20054), .B2(n21190), .A(n20939), .ZN(P1_U2802) );
  NOR2_X1 U22962 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20055) );
  OAI21_X1 U22963 ( .B1(n20055), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20927), .ZN(
        n20053) );
  OAI21_X1 U22964 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20927), .A(n20053), 
        .ZN(P1_U2804) );
  NOR2_X1 U22965 ( .A1(n20939), .A2(n20054), .ZN(n20912) );
  OAI21_X1 U22966 ( .B1(BS16), .B2(n20055), .A(n20912), .ZN(n20910) );
  OAI21_X1 U22967 ( .B1(n20912), .B2(n21085), .A(n20910), .ZN(P1_U2805) );
  OAI21_X1 U22968 ( .B1(n20058), .B2(n20057), .A(n20056), .ZN(P1_U2806) );
  NOR4_X1 U22969 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20062) );
  NOR4_X1 U22970 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20061) );
  NOR4_X1 U22971 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20060) );
  NOR4_X1 U22972 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20059) );
  NAND4_X1 U22973 ( .A1(n20062), .A2(n20061), .A3(n20060), .A4(n20059), .ZN(
        n20068) );
  NOR4_X1 U22974 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20066) );
  AOI211_X1 U22975 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20065) );
  NOR4_X1 U22976 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20064) );
  NOR4_X1 U22977 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20063) );
  NAND4_X1 U22978 ( .A1(n20066), .A2(n20065), .A3(n20064), .A4(n20063), .ZN(
        n20067) );
  NOR2_X1 U22979 ( .A1(n20068), .A2(n20067), .ZN(n20923) );
  INV_X1 U22980 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21262) );
  NOR3_X1 U22981 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20070) );
  OAI21_X1 U22982 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20070), .A(n20923), .ZN(
        n20069) );
  OAI21_X1 U22983 ( .B1(n20923), .B2(n21262), .A(n20069), .ZN(P1_U2807) );
  INV_X1 U22984 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20911) );
  AOI21_X1 U22985 ( .B1(n13685), .B2(n20911), .A(n20070), .ZN(n20072) );
  INV_X1 U22986 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20071) );
  INV_X1 U22987 ( .A(n20923), .ZN(n20925) );
  AOI22_X1 U22988 ( .A1(n20923), .A2(n20072), .B1(n20071), .B2(n20925), .ZN(
        P1_U2808) );
  OAI21_X1 U22989 ( .B1(n20115), .B2(n20073), .A(n20113), .ZN(n20077) );
  NOR3_X1 U22990 ( .A1(n20075), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n20074), .ZN(
        n20076) );
  AOI211_X1 U22991 ( .C1(n20127), .C2(P1_EBX_REG_9__SCAN_IN), .A(n20077), .B(
        n20076), .ZN(n20078) );
  OAI21_X1 U22992 ( .B1(n20080), .B2(n20079), .A(n20078), .ZN(n20081) );
  AOI21_X1 U22993 ( .B1(n20082), .B2(n20106), .A(n20081), .ZN(n20087) );
  AOI22_X1 U22994 ( .A1(n20085), .A2(n20084), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n20083), .ZN(n20086) );
  NAND2_X1 U22995 ( .A1(n20087), .A2(n20086), .ZN(P1_U2831) );
  INV_X1 U22996 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21095) );
  INV_X1 U22997 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21229) );
  NOR2_X1 U22998 ( .A1(n21095), .A2(n21229), .ZN(n20089) );
  INV_X1 U22999 ( .A(n20089), .ZN(n20088) );
  NOR3_X1 U23000 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20088), .A3(n20120), .ZN(
        n20093) );
  INV_X1 U23001 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20091) );
  AOI21_X1 U23002 ( .B1(n20089), .B2(n20111), .A(n20112), .ZN(n20101) );
  AOI22_X1 U23003 ( .A1(n20101), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20127), 
        .B2(P1_EBX_REG_7__SCAN_IN), .ZN(n20090) );
  OAI211_X1 U23004 ( .C1(n20115), .C2(n20091), .A(n20090), .B(n20113), .ZN(
        n20092) );
  AOI211_X1 U23005 ( .C1(n20094), .C2(n20126), .A(n20093), .B(n20092), .ZN(
        n20097) );
  NAND2_X1 U23006 ( .A1(n20095), .A2(n20106), .ZN(n20096) );
  OAI211_X1 U23007 ( .C1(n20140), .C2(n20098), .A(n20097), .B(n20096), .ZN(
        P1_U2833) );
  NOR2_X1 U23008 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20120), .ZN(n20099) );
  AOI22_X1 U23009 ( .A1(n20126), .A2(n20100), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n20099), .ZN(n20109) );
  NAND2_X1 U23010 ( .A1(n20101), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n20103) );
  AOI21_X1 U23011 ( .B1(n20133), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20132), .ZN(n20102) );
  OAI211_X1 U23012 ( .C1(n20104), .C2(n21296), .A(n20103), .B(n20102), .ZN(
        n20105) );
  AOI21_X1 U23013 ( .B1(n20107), .B2(n20106), .A(n20105), .ZN(n20108) );
  OAI211_X1 U23014 ( .C1(n20110), .C2(n20140), .A(n20109), .B(n20108), .ZN(
        P1_U2834) );
  NOR2_X1 U23015 ( .A1(n20112), .A2(n20111), .ZN(n20137) );
  NAND2_X1 U23016 ( .A1(n20137), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n20119) );
  NAND2_X1 U23017 ( .A1(n20127), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n20114) );
  OAI211_X1 U23018 ( .C1(n12468), .C2(n20115), .A(n20114), .B(n20113), .ZN(
        n20116) );
  AOI21_X1 U23019 ( .B1(n20126), .B2(n20117), .A(n20116), .ZN(n20118) );
  OAI211_X1 U23020 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n20120), .A(n20119), .B(
        n20118), .ZN(n20121) );
  AOI21_X1 U23021 ( .B1(n20122), .B2(n20135), .A(n20121), .ZN(n20123) );
  OAI21_X1 U23022 ( .B1(n20124), .B2(n20140), .A(n20123), .ZN(P1_U2835) );
  INV_X1 U23023 ( .A(n20125), .ZN(n20194) );
  AOI22_X1 U23024 ( .A1(n20127), .A2(P1_EBX_REG_4__SCAN_IN), .B1(n20126), .B2(
        n20194), .ZN(n20128) );
  OAI21_X1 U23025 ( .B1(n20130), .B2(n20129), .A(n20128), .ZN(n20131) );
  AOI211_X1 U23026 ( .C1(n20133), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20132), .B(n20131), .ZN(n20139) );
  OAI21_X1 U23027 ( .B1(n20870), .B2(n20134), .A(n21228), .ZN(n20136) );
  AOI22_X1 U23028 ( .A1(n20137), .A2(n20136), .B1(n20187), .B2(n20135), .ZN(
        n20138) );
  OAI211_X1 U23029 ( .C1(n20192), .C2(n20140), .A(n20139), .B(n20138), .ZN(
        P1_U2836) );
  AOI22_X1 U23030 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20144), .B1(n20163), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20141) );
  OAI21_X1 U23031 ( .B1(n20143), .B2(n20142), .A(n20141), .ZN(P1_U2921) );
  AOI22_X1 U23032 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20145) );
  OAI21_X1 U23033 ( .B1(n14974), .B2(n20166), .A(n20145), .ZN(P1_U2922) );
  AOI22_X1 U23034 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20146) );
  OAI21_X1 U23035 ( .B1(n14977), .B2(n20166), .A(n20146), .ZN(P1_U2923) );
  AOI22_X1 U23036 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20147) );
  OAI21_X1 U23037 ( .B1(n14981), .B2(n20166), .A(n20147), .ZN(P1_U2924) );
  AOI22_X1 U23038 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20148) );
  OAI21_X1 U23039 ( .B1(n14984), .B2(n20166), .A(n20148), .ZN(P1_U2925) );
  INV_X1 U23040 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20150) );
  AOI22_X1 U23041 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20149) );
  OAI21_X1 U23042 ( .B1(n20150), .B2(n20166), .A(n20149), .ZN(P1_U2926) );
  AOI22_X1 U23043 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20151) );
  OAI21_X1 U23044 ( .B1(n14251), .B2(n20166), .A(n20151), .ZN(P1_U2927) );
  AOI22_X1 U23045 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20152) );
  OAI21_X1 U23046 ( .B1(n20153), .B2(n20166), .A(n20152), .ZN(P1_U2928) );
  AOI22_X1 U23047 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20154) );
  OAI21_X1 U23048 ( .B1(n14184), .B2(n20166), .A(n20154), .ZN(P1_U2929) );
  AOI22_X1 U23049 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20155) );
  OAI21_X1 U23050 ( .B1(n20156), .B2(n20166), .A(n20155), .ZN(P1_U2930) );
  AOI22_X1 U23051 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20157) );
  OAI21_X1 U23052 ( .B1(n12471), .B2(n20166), .A(n20157), .ZN(P1_U2931) );
  AOI22_X1 U23053 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20158) );
  OAI21_X1 U23054 ( .B1(n20159), .B2(n20166), .A(n20158), .ZN(P1_U2932) );
  AOI22_X1 U23055 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20160) );
  OAI21_X1 U23056 ( .B1(n12422), .B2(n20166), .A(n20160), .ZN(P1_U2933) );
  AOI22_X1 U23057 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20161) );
  OAI21_X1 U23058 ( .B1(n12368), .B2(n20166), .A(n20161), .ZN(P1_U2934) );
  AOI22_X1 U23059 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20162) );
  OAI21_X1 U23060 ( .B1(n12372), .B2(n20166), .A(n20162), .ZN(P1_U2935) );
  AOI22_X1 U23061 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20164), .B1(n20163), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20165) );
  OAI21_X1 U23062 ( .B1(n20167), .B2(n20166), .A(n20165), .ZN(P1_U2936) );
  AOI22_X1 U23063 ( .A1(n20179), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20178), .ZN(n20169) );
  NAND2_X1 U23064 ( .A1(n20169), .A2(n20168), .ZN(P1_U2961) );
  AOI22_X1 U23065 ( .A1(n20179), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20178), .ZN(n20171) );
  NAND2_X1 U23066 ( .A1(n20171), .A2(n20170), .ZN(P1_U2962) );
  AOI22_X1 U23067 ( .A1(n20179), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20178), .ZN(n20173) );
  NAND2_X1 U23068 ( .A1(n20173), .A2(n20172), .ZN(P1_U2963) );
  AOI22_X1 U23069 ( .A1(n20179), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20178), .ZN(n20175) );
  NAND2_X1 U23070 ( .A1(n20175), .A2(n20174), .ZN(P1_U2964) );
  AOI22_X1 U23071 ( .A1(n20179), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20178), .ZN(n20177) );
  NAND2_X1 U23072 ( .A1(n20177), .A2(n20176), .ZN(P1_U2965) );
  AOI22_X1 U23073 ( .A1(n20179), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20178), .ZN(n20181) );
  NAND2_X1 U23074 ( .A1(n20181), .A2(n20180), .ZN(P1_U2966) );
  AOI22_X1 U23075 ( .A1(n20182), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n10057), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20191) );
  OAI21_X1 U23076 ( .B1(n20183), .B2(n20185), .A(n20184), .ZN(n20186) );
  INV_X1 U23077 ( .A(n20186), .ZN(n20197) );
  AOI22_X1 U23078 ( .A1(n20197), .A2(n20189), .B1(n20188), .B2(n20187), .ZN(
        n20190) );
  OAI211_X1 U23079 ( .C1(n20193), .C2(n20192), .A(n20191), .B(n20190), .ZN(
        P1_U2995) );
  OAI21_X1 U23080 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20202), .ZN(n20200) );
  AOI22_X1 U23081 ( .A1(n20194), .A2(n20205), .B1(n10057), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20199) );
  OAI21_X1 U23082 ( .B1(n20218), .B2(n20196), .A(n20195), .ZN(n20207) );
  AOI22_X1 U23083 ( .A1(n20197), .A2(n20215), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20207), .ZN(n20198) );
  OAI211_X1 U23084 ( .C1(n20201), .C2(n20200), .A(n20199), .B(n20198), .ZN(
        P1_U3027) );
  INV_X1 U23085 ( .A(n20202), .ZN(n20210) );
  AOI21_X1 U23086 ( .B1(n20205), .B2(n20204), .A(n20203), .ZN(n20209) );
  AOI22_X1 U23087 ( .A1(n20207), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20215), .B2(n20206), .ZN(n20208) );
  OAI211_X1 U23088 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20210), .A(
        n20209), .B(n20208), .ZN(P1_U3028) );
  NAND2_X1 U23089 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20211), .ZN(
        n20233) );
  AOI21_X1 U23090 ( .B1(n20214), .B2(n20213), .A(n20212), .ZN(n20231) );
  NAND3_X1 U23091 ( .A1(n20216), .A2(n15152), .A3(n20215), .ZN(n20229) );
  AND2_X1 U23092 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20217) );
  NAND2_X1 U23093 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n20217), .ZN(
        n20219) );
  NAND2_X1 U23094 ( .A1(n20219), .A2(n20218), .ZN(n20220) );
  AND2_X1 U23095 ( .A1(n20221), .A2(n20220), .ZN(n20227) );
  OAI22_X1 U23096 ( .A1(n20225), .A2(n20224), .B1(n20223), .B2(n20222), .ZN(
        n20226) );
  NOR2_X1 U23097 ( .A1(n20227), .A2(n20226), .ZN(n20228) );
  AND2_X1 U23098 ( .A1(n20229), .A2(n20228), .ZN(n20230) );
  OAI221_X1 U23099 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20233), .C1(
        n20232), .C2(n20231), .A(n20230), .ZN(P1_U3029) );
  NOR2_X1 U23100 ( .A1(n16140), .A2(n20234), .ZN(P1_U3032) );
  INV_X1 U23101 ( .A(DATAI_16_), .ZN(n21265) );
  NAND2_X1 U23102 ( .A1(n20235), .A2(n20188), .ZN(n20284) );
  NAND2_X1 U23103 ( .A1(n20188), .A2(n20236), .ZN(n20285) );
  OAI22_X1 U23104 ( .A1(n21265), .A2(n20284), .B1(n20237), .B2(n20285), .ZN(
        n20792) );
  INV_X1 U23105 ( .A(n20792), .ZN(n20736) );
  INV_X1 U23106 ( .A(n13914), .ZN(n20239) );
  INV_X1 U23107 ( .A(n20628), .ZN(n20241) );
  INV_X1 U23108 ( .A(n20285), .ZN(n20287) );
  INV_X1 U23109 ( .A(n20284), .ZN(n20288) );
  AOI22_X1 U23110 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20287), .B1(DATAI_24_), 
        .B2(n20288), .ZN(n20795) );
  INV_X1 U23111 ( .A(n20795), .ZN(n20733) );
  NAND3_X1 U23112 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20932), .A3(n20242), 
        .ZN(n20276) );
  NAND2_X1 U23113 ( .A1(n20289), .A2(n20243), .ZN(n20783) );
  NOR3_X1 U23114 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20302) );
  NAND2_X1 U23115 ( .A1(n20690), .A2(n20302), .ZN(n20248) );
  INV_X1 U23116 ( .A(n20248), .ZN(n20290) );
  AOI22_X1 U23117 ( .A1(n20843), .A2(n20733), .B1(n20725), .B2(n20290), .ZN(
        n20257) );
  INV_X1 U23118 ( .A(n20582), .ZN(n20244) );
  NOR2_X1 U23119 ( .A1(n20244), .A2(n20529), .ZN(n20253) );
  INV_X1 U23120 ( .A(n20245), .ZN(n20252) );
  NAND2_X1 U23121 ( .A1(n20252), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20722) );
  NAND2_X1 U23122 ( .A1(n20308), .A2(n20790), .ZN(n20246) );
  NAND2_X1 U23123 ( .A1(n20790), .A2(n21085), .ZN(n20652) );
  OAI21_X1 U23124 ( .B1(n20246), .B2(n20843), .A(n20652), .ZN(n20251) );
  NAND2_X1 U23125 ( .A1(n10019), .A2(n20528), .ZN(n20254) );
  AOI22_X1 U23126 ( .A1(n20251), .A2(n20254), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20248), .ZN(n20249) );
  OAI211_X1 U23127 ( .C1(n20253), .C2(n20929), .A(n20589), .B(n20249), .ZN(
        n20294) );
  NAND2_X1 U23128 ( .A1(n20250), .A2(n20292), .ZN(n20782) );
  INV_X1 U23129 ( .A(n20251), .ZN(n20255) );
  NOR2_X1 U23130 ( .A1(n20252), .A2(n20929), .ZN(n20584) );
  INV_X1 U23131 ( .A(n20584), .ZN(n20530) );
  INV_X1 U23132 ( .A(n20253), .ZN(n20402) );
  OAI22_X1 U23133 ( .A1(n20255), .A2(n20254), .B1(n20530), .B2(n20402), .ZN(
        n20293) );
  AOI22_X1 U23134 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20294), .B1(
        n20724), .B2(n20293), .ZN(n20256) );
  OAI211_X1 U23135 ( .C1(n20736), .C2(n20308), .A(n20257), .B(n20256), .ZN(
        P1_U3033) );
  INV_X1 U23136 ( .A(DATAI_17_), .ZN(n21072) );
  OAI22_X1 U23137 ( .A1(n20258), .A2(n20285), .B1(n21072), .B2(n20284), .ZN(
        n20798) );
  INV_X1 U23138 ( .A(n20798), .ZN(n20740) );
  AOI22_X1 U23139 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20287), .B1(DATAI_25_), 
        .B2(n20288), .ZN(n20801) );
  INV_X1 U23140 ( .A(n20801), .ZN(n20737) );
  AOI22_X1 U23141 ( .A1(n20843), .A2(n20737), .B1(n20797), .B2(n20290), .ZN(
        n20261) );
  NAND2_X1 U23142 ( .A1(n20259), .A2(n20292), .ZN(n20669) );
  AOI22_X1 U23143 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20294), .B1(
        n20796), .B2(n20293), .ZN(n20260) );
  OAI211_X1 U23144 ( .C1(n20740), .C2(n20308), .A(n20261), .B(n20260), .ZN(
        P1_U3034) );
  INV_X1 U23145 ( .A(DATAI_18_), .ZN(n21024) );
  OAI22_X1 U23146 ( .A1(n20262), .A2(n20285), .B1(n21024), .B2(n20284), .ZN(
        n20805) );
  INV_X1 U23147 ( .A(n20805), .ZN(n20746) );
  AOI22_X1 U23148 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20287), .B1(DATAI_26_), 
        .B2(n20288), .ZN(n20808) );
  INV_X1 U23149 ( .A(n20808), .ZN(n20743) );
  NAND2_X1 U23150 ( .A1(n20289), .A2(n20263), .ZN(n20803) );
  AOI22_X1 U23151 ( .A1(n20843), .A2(n20743), .B1(n20742), .B2(n20290), .ZN(
        n20266) );
  NAND2_X1 U23152 ( .A1(n20264), .A2(n20292), .ZN(n20802) );
  AOI22_X1 U23153 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20294), .B1(
        n20741), .B2(n20293), .ZN(n20265) );
  OAI211_X1 U23154 ( .C1(n20746), .C2(n20308), .A(n20266), .B(n20265), .ZN(
        P1_U3035) );
  INV_X1 U23155 ( .A(DATAI_19_), .ZN(n21251) );
  OAI22_X1 U23156 ( .A1(n20267), .A2(n20285), .B1(n21251), .B2(n20284), .ZN(
        n20812) );
  INV_X1 U23157 ( .A(n20812), .ZN(n20752) );
  AOI22_X1 U23158 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20287), .B1(DATAI_27_), 
        .B2(n20288), .ZN(n20815) );
  INV_X1 U23159 ( .A(n20815), .ZN(n20749) );
  NAND2_X1 U23160 ( .A1(n20289), .A2(n20268), .ZN(n20810) );
  AOI22_X1 U23161 ( .A1(n20843), .A2(n20749), .B1(n20748), .B2(n20290), .ZN(
        n20271) );
  NAND2_X1 U23162 ( .A1(n20269), .A2(n20292), .ZN(n20809) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20294), .B1(
        n20747), .B2(n20293), .ZN(n20270) );
  OAI211_X1 U23164 ( .C1(n20752), .C2(n20308), .A(n20271), .B(n20270), .ZN(
        P1_U3036) );
  OAI22_X1 U23165 ( .A1(n20272), .A2(n20285), .B1(n14950), .B2(n20284), .ZN(
        n20819) );
  INV_X1 U23166 ( .A(n20819), .ZN(n20758) );
  AOI22_X1 U23167 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20287), .B1(DATAI_28_), 
        .B2(n20288), .ZN(n20822) );
  INV_X1 U23168 ( .A(n20822), .ZN(n20755) );
  NAND2_X1 U23169 ( .A1(n20289), .A2(n12301), .ZN(n20817) );
  AOI22_X1 U23170 ( .A1(n20843), .A2(n20755), .B1(n20754), .B2(n20290), .ZN(
        n20275) );
  NAND2_X1 U23171 ( .A1(n20273), .A2(n20292), .ZN(n20816) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20294), .B1(
        n20753), .B2(n20293), .ZN(n20274) );
  OAI211_X1 U23173 ( .C1(n20758), .C2(n20308), .A(n20275), .B(n20274), .ZN(
        P1_U3037) );
  AOI22_X1 U23174 ( .A1(DATAI_21_), .A2(n20288), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20287), .ZN(n20762) );
  AOI22_X1 U23175 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20287), .B1(DATAI_29_), 
        .B2(n20288), .ZN(n20828) );
  INV_X1 U23176 ( .A(n20828), .ZN(n20759) );
  NOR2_X2 U23177 ( .A1(n20276), .A2(n10059), .ZN(n20824) );
  AOI22_X1 U23178 ( .A1(n20843), .A2(n20759), .B1(n20824), .B2(n20290), .ZN(
        n20279) );
  NAND2_X1 U23179 ( .A1(n20277), .A2(n20292), .ZN(n20678) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20294), .B1(
        n20823), .B2(n20293), .ZN(n20278) );
  OAI211_X1 U23181 ( .C1(n20762), .C2(n20308), .A(n20279), .B(n20278), .ZN(
        P1_U3038) );
  INV_X1 U23182 ( .A(DATAI_22_), .ZN(n21014) );
  OAI22_X1 U23183 ( .A1(n20280), .A2(n20285), .B1(n21014), .B2(n20284), .ZN(
        n20834) );
  INV_X1 U23184 ( .A(n20834), .ZN(n20768) );
  AOI22_X1 U23185 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20287), .B1(DATAI_30_), 
        .B2(n20288), .ZN(n20837) );
  INV_X1 U23186 ( .A(n20837), .ZN(n20765) );
  NAND2_X1 U23187 ( .A1(n20289), .A2(n12239), .ZN(n20832) );
  AOI22_X1 U23188 ( .A1(n20843), .A2(n20765), .B1(n20764), .B2(n20290), .ZN(
        n20283) );
  NAND2_X1 U23189 ( .A1(n20281), .A2(n20292), .ZN(n20830) );
  AOI22_X1 U23190 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20294), .B1(
        n20763), .B2(n20293), .ZN(n20282) );
  OAI211_X1 U23191 ( .C1(n20768), .C2(n20308), .A(n20283), .B(n20282), .ZN(
        P1_U3039) );
  INV_X1 U23192 ( .A(DATAI_23_), .ZN(n21089) );
  OAI22_X1 U23193 ( .A1(n20286), .A2(n20285), .B1(n21089), .B2(n20284), .ZN(
        n20842) );
  INV_X1 U23194 ( .A(n20842), .ZN(n20776) );
  AOI22_X1 U23195 ( .A1(DATAI_31_), .A2(n20288), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20287), .ZN(n20848) );
  INV_X1 U23196 ( .A(n20848), .ZN(n20771) );
  NAND2_X1 U23197 ( .A1(n20289), .A2(n13015), .ZN(n20614) );
  AOI22_X1 U23198 ( .A1(n20843), .A2(n20771), .B1(n20840), .B2(n20290), .ZN(
        n20296) );
  AOI22_X1 U23199 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20294), .B1(
        n20839), .B2(n20293), .ZN(n20295) );
  OAI211_X1 U23200 ( .C1(n20776), .C2(n20308), .A(n20296), .B(n20295), .ZN(
        P1_U3040) );
  INV_X1 U23201 ( .A(n20302), .ZN(n20298) );
  NOR2_X1 U23202 ( .A1(n20690), .A2(n20298), .ZN(n20320) );
  INV_X1 U23203 ( .A(n20297), .ZN(n20692) );
  AOI21_X1 U23204 ( .B1(n10019), .B2(n20692), .A(n20320), .ZN(n20300) );
  OAI22_X1 U23205 ( .A1(n20300), .A2(n20779), .B1(n20298), .B2(n20929), .ZN(
        n20319) );
  AOI22_X1 U23206 ( .A1(n20725), .A2(n20320), .B1(n20724), .B2(n20319), .ZN(
        n20304) );
  INV_X1 U23207 ( .A(n20363), .ZN(n20299) );
  NOR2_X1 U23208 ( .A1(n20299), .A2(n20779), .ZN(n20361) );
  INV_X1 U23209 ( .A(n20652), .ZN(n20695) );
  OAI21_X1 U23210 ( .B1(n20361), .B2(n20695), .A(n20300), .ZN(n20301) );
  OAI211_X1 U23211 ( .C1(n20790), .C2(n20302), .A(n20789), .B(n20301), .ZN(
        n20322) );
  AOI22_X1 U23212 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20733), .ZN(n20303) );
  OAI211_X1 U23213 ( .C1(n20736), .C2(n20352), .A(n20304), .B(n20303), .ZN(
        P1_U3041) );
  AOI22_X1 U23214 ( .A1(n20797), .A2(n20320), .B1(n20319), .B2(n20796), .ZN(
        n20307) );
  INV_X1 U23215 ( .A(n20352), .ZN(n20305) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20322), .B1(
        n20305), .B2(n20798), .ZN(n20306) );
  OAI211_X1 U23217 ( .C1(n20801), .C2(n20308), .A(n20307), .B(n20306), .ZN(
        P1_U3042) );
  AOI22_X1 U23218 ( .A1(n20742), .A2(n20320), .B1(n20741), .B2(n20319), .ZN(
        n20310) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20743), .ZN(n20309) );
  OAI211_X1 U23220 ( .C1(n20746), .C2(n20352), .A(n20310), .B(n20309), .ZN(
        P1_U3043) );
  AOI22_X1 U23221 ( .A1(n20748), .A2(n20320), .B1(n20747), .B2(n20319), .ZN(
        n20312) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20749), .ZN(n20311) );
  OAI211_X1 U23223 ( .C1(n20752), .C2(n20352), .A(n20312), .B(n20311), .ZN(
        P1_U3044) );
  AOI22_X1 U23224 ( .A1(n20754), .A2(n20320), .B1(n20753), .B2(n20319), .ZN(
        n20314) );
  AOI22_X1 U23225 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20755), .ZN(n20313) );
  OAI211_X1 U23226 ( .C1(n20758), .C2(n20352), .A(n20314), .B(n20313), .ZN(
        P1_U3045) );
  AOI22_X1 U23227 ( .A1(n20824), .A2(n20320), .B1(n20319), .B2(n20823), .ZN(
        n20316) );
  AOI22_X1 U23228 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20759), .ZN(n20315) );
  OAI211_X1 U23229 ( .C1(n20762), .C2(n20352), .A(n20316), .B(n20315), .ZN(
        P1_U3046) );
  AOI22_X1 U23230 ( .A1(n20764), .A2(n20320), .B1(n20763), .B2(n20319), .ZN(
        n20318) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20765), .ZN(n20317) );
  OAI211_X1 U23232 ( .C1(n20768), .C2(n20352), .A(n20318), .B(n20317), .ZN(
        P1_U3047) );
  AOI22_X1 U23233 ( .A1(n20840), .A2(n20320), .B1(n20839), .B2(n20319), .ZN(
        n20324) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20322), .B1(
        n20321), .B2(n20771), .ZN(n20323) );
  OAI211_X1 U23235 ( .C1(n20776), .C2(n20352), .A(n20324), .B(n20323), .ZN(
        P1_U3048) );
  INV_X1 U23236 ( .A(n20718), .ZN(n20454) );
  NOR3_X1 U23237 ( .A1(n20585), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20365) );
  NAND2_X1 U23238 ( .A1(n20690), .A2(n20365), .ZN(n20351) );
  OAI22_X1 U23239 ( .A1(n20352), .A2(n20795), .B1(n20783), .B2(n20351), .ZN(
        n20325) );
  INV_X1 U23240 ( .A(n20325), .ZN(n20332) );
  AOI21_X1 U23241 ( .B1(n20394), .B2(n20352), .A(n21085), .ZN(n20326) );
  NOR2_X1 U23242 ( .A1(n20326), .A2(n20779), .ZN(n20328) );
  INV_X1 U23243 ( .A(n20528), .ZN(n20727) );
  NAND2_X1 U23244 ( .A1(n10019), .A2(n20727), .ZN(n20329) );
  AOI22_X1 U23245 ( .A1(n20328), .A2(n20329), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20351), .ZN(n20327) );
  OR2_X1 U23246 ( .A1(n20582), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20460) );
  NAND2_X1 U23247 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20460), .ZN(n20457) );
  NAND3_X1 U23248 ( .A1(n20589), .A2(n20327), .A3(n20457), .ZN(n20355) );
  INV_X1 U23249 ( .A(n20328), .ZN(n20330) );
  OAI22_X1 U23250 ( .A1(n20330), .A2(n20329), .B1(n20530), .B2(n20460), .ZN(
        n20354) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20355), .B1(
        n20724), .B2(n20354), .ZN(n20331) );
  OAI211_X1 U23252 ( .C1(n20736), .C2(n20394), .A(n20332), .B(n20331), .ZN(
        P1_U3049) );
  INV_X1 U23253 ( .A(n20394), .ZN(n20390) );
  INV_X1 U23254 ( .A(n20351), .ZN(n20333) );
  AOI22_X1 U23255 ( .A1(n20390), .A2(n20798), .B1(n20797), .B2(n20333), .ZN(
        n20335) );
  AOI22_X1 U23256 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20355), .B1(
        n20796), .B2(n20354), .ZN(n20334) );
  OAI211_X1 U23257 ( .C1(n20801), .C2(n20352), .A(n20335), .B(n20334), .ZN(
        P1_U3050) );
  OAI22_X1 U23258 ( .A1(n20394), .A2(n20746), .B1(n20803), .B2(n20351), .ZN(
        n20336) );
  INV_X1 U23259 ( .A(n20336), .ZN(n20338) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20355), .B1(
        n20741), .B2(n20354), .ZN(n20337) );
  OAI211_X1 U23261 ( .C1(n20808), .C2(n20352), .A(n20338), .B(n20337), .ZN(
        P1_U3051) );
  OAI22_X1 U23262 ( .A1(n20352), .A2(n20815), .B1(n20810), .B2(n20351), .ZN(
        n20339) );
  INV_X1 U23263 ( .A(n20339), .ZN(n20341) );
  AOI22_X1 U23264 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20355), .B1(
        n20747), .B2(n20354), .ZN(n20340) );
  OAI211_X1 U23265 ( .C1(n20752), .C2(n20394), .A(n20341), .B(n20340), .ZN(
        P1_U3052) );
  OAI22_X1 U23266 ( .A1(n20394), .A2(n20758), .B1(n20817), .B2(n20351), .ZN(
        n20342) );
  INV_X1 U23267 ( .A(n20342), .ZN(n20344) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20355), .B1(
        n20753), .B2(n20354), .ZN(n20343) );
  OAI211_X1 U23269 ( .C1(n20822), .C2(n20352), .A(n20344), .B(n20343), .ZN(
        P1_U3053) );
  INV_X1 U23270 ( .A(n20824), .ZN(n20385) );
  OAI22_X1 U23271 ( .A1(n20352), .A2(n20828), .B1(n20385), .B2(n20351), .ZN(
        n20345) );
  INV_X1 U23272 ( .A(n20345), .ZN(n20347) );
  AOI22_X1 U23273 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20355), .B1(
        n20823), .B2(n20354), .ZN(n20346) );
  OAI211_X1 U23274 ( .C1(n20762), .C2(n20394), .A(n20347), .B(n20346), .ZN(
        P1_U3054) );
  OAI22_X1 U23275 ( .A1(n20394), .A2(n20768), .B1(n20832), .B2(n20351), .ZN(
        n20348) );
  INV_X1 U23276 ( .A(n20348), .ZN(n20350) );
  AOI22_X1 U23277 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20355), .B1(
        n20763), .B2(n20354), .ZN(n20349) );
  OAI211_X1 U23278 ( .C1(n20837), .C2(n20352), .A(n20350), .B(n20349), .ZN(
        P1_U3055) );
  OAI22_X1 U23279 ( .A1(n20352), .A2(n20848), .B1(n20614), .B2(n20351), .ZN(
        n20353) );
  INV_X1 U23280 ( .A(n20353), .ZN(n20357) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20355), .B1(
        n20839), .B2(n20354), .ZN(n20356) );
  OAI211_X1 U23282 ( .C1(n20776), .C2(n20394), .A(n20357), .B(n20356), .ZN(
        P1_U3056) );
  AND2_X1 U23283 ( .A1(n20358), .A2(n12378), .ZN(n20777) );
  INV_X1 U23284 ( .A(n20621), .ZN(n20359) );
  NAND2_X1 U23285 ( .A1(n20359), .A2(n20658), .ZN(n20393) );
  INV_X1 U23286 ( .A(n20393), .ZN(n20360) );
  AOI21_X1 U23287 ( .B1(n10019), .B2(n20777), .A(n20360), .ZN(n20368) );
  INV_X1 U23288 ( .A(n20368), .ZN(n20362) );
  AOI22_X1 U23289 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20365), .B1(n20362), 
        .B2(n20367), .ZN(n20399) );
  OAI22_X1 U23290 ( .A1(n20403), .A2(n20736), .B1(n20783), .B2(n20393), .ZN(
        n20364) );
  INV_X1 U23291 ( .A(n20364), .ZN(n20371) );
  INV_X1 U23292 ( .A(n20365), .ZN(n20366) );
  AOI22_X1 U23293 ( .A1(n20368), .A2(n20367), .B1(n20779), .B2(n20366), .ZN(
        n20369) );
  NAND2_X1 U23294 ( .A1(n20789), .A2(n20369), .ZN(n20396) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20396), .B1(
        n20390), .B2(n20733), .ZN(n20370) );
  OAI211_X1 U23296 ( .C1(n20399), .C2(n20782), .A(n20371), .B(n20370), .ZN(
        P1_U3057) );
  INV_X1 U23297 ( .A(n20797), .ZN(n20372) );
  OAI22_X1 U23298 ( .A1(n20394), .A2(n20801), .B1(n20372), .B2(n20393), .ZN(
        n20373) );
  INV_X1 U23299 ( .A(n20373), .ZN(n20375) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20396), .B1(
        n20424), .B2(n20798), .ZN(n20374) );
  OAI211_X1 U23301 ( .C1(n20399), .C2(n20669), .A(n20375), .B(n20374), .ZN(
        P1_U3058) );
  OAI22_X1 U23302 ( .A1(n20394), .A2(n20808), .B1(n20803), .B2(n20393), .ZN(
        n20376) );
  INV_X1 U23303 ( .A(n20376), .ZN(n20378) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20396), .B1(
        n20424), .B2(n20805), .ZN(n20377) );
  OAI211_X1 U23305 ( .C1(n20399), .C2(n20802), .A(n20378), .B(n20377), .ZN(
        P1_U3059) );
  OAI22_X1 U23306 ( .A1(n20394), .A2(n20815), .B1(n20810), .B2(n20393), .ZN(
        n20379) );
  INV_X1 U23307 ( .A(n20379), .ZN(n20381) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20396), .B1(
        n20424), .B2(n20812), .ZN(n20380) );
  OAI211_X1 U23309 ( .C1(n20399), .C2(n20809), .A(n20381), .B(n20380), .ZN(
        P1_U3060) );
  OAI22_X1 U23310 ( .A1(n20403), .A2(n20758), .B1(n20817), .B2(n20393), .ZN(
        n20382) );
  INV_X1 U23311 ( .A(n20382), .ZN(n20384) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20396), .B1(
        n20390), .B2(n20755), .ZN(n20383) );
  OAI211_X1 U23313 ( .C1(n20399), .C2(n20816), .A(n20384), .B(n20383), .ZN(
        P1_U3061) );
  OAI22_X1 U23314 ( .A1(n20394), .A2(n20828), .B1(n20385), .B2(n20393), .ZN(
        n20386) );
  INV_X1 U23315 ( .A(n20386), .ZN(n20388) );
  INV_X1 U23316 ( .A(n20762), .ZN(n20825) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20396), .B1(
        n20424), .B2(n20825), .ZN(n20387) );
  OAI211_X1 U23318 ( .C1(n20399), .C2(n20678), .A(n20388), .B(n20387), .ZN(
        P1_U3062) );
  OAI22_X1 U23319 ( .A1(n20403), .A2(n20768), .B1(n20832), .B2(n20393), .ZN(
        n20389) );
  INV_X1 U23320 ( .A(n20389), .ZN(n20392) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20396), .B1(
        n20390), .B2(n20765), .ZN(n20391) );
  OAI211_X1 U23322 ( .C1(n20399), .C2(n20830), .A(n20392), .B(n20391), .ZN(
        P1_U3063) );
  INV_X1 U23323 ( .A(n20839), .ZN(n20686) );
  OAI22_X1 U23324 ( .A1(n20394), .A2(n20848), .B1(n20614), .B2(n20393), .ZN(
        n20395) );
  INV_X1 U23325 ( .A(n20395), .ZN(n20398) );
  AOI22_X1 U23326 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20396), .B1(
        n20424), .B2(n20842), .ZN(n20397) );
  OAI211_X1 U23327 ( .C1(n20399), .C2(n20686), .A(n20398), .B(n20397), .ZN(
        P1_U3064) );
  NOR3_X1 U23328 ( .A1(n13020), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20432) );
  INV_X1 U23329 ( .A(n20432), .ZN(n20428) );
  NOR2_X1 U23330 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20428), .ZN(
        n20423) );
  NOR2_X1 U23331 ( .A1(n20655), .A2(n20400), .ZN(n20490) );
  NAND3_X1 U23332 ( .A1(n20490), .A2(n20790), .A3(n20528), .ZN(n20401) );
  OAI21_X1 U23333 ( .B1(n20402), .B2(n20722), .A(n20401), .ZN(n20422) );
  AOI22_X1 U23334 ( .A1(n20725), .A2(n20423), .B1(n20724), .B2(n20422), .ZN(
        n20409) );
  AOI21_X1 U23335 ( .B1(n20403), .B2(n20441), .A(n21085), .ZN(n20404) );
  AOI21_X1 U23336 ( .B1(n20490), .B2(n20528), .A(n20404), .ZN(n20405) );
  NOR2_X1 U23337 ( .A1(n20405), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20407) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20733), .ZN(n20408) );
  OAI211_X1 U23339 ( .C1(n20736), .C2(n20441), .A(n20409), .B(n20408), .ZN(
        P1_U3065) );
  AOI22_X1 U23340 ( .A1(n20797), .A2(n20423), .B1(n20796), .B2(n20422), .ZN(
        n20411) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20737), .ZN(n20410) );
  OAI211_X1 U23342 ( .C1(n20740), .C2(n20441), .A(n20411), .B(n20410), .ZN(
        P1_U3066) );
  AOI22_X1 U23343 ( .A1(n20742), .A2(n20423), .B1(n20741), .B2(n20422), .ZN(
        n20413) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20743), .ZN(n20412) );
  OAI211_X1 U23345 ( .C1(n20746), .C2(n20441), .A(n20413), .B(n20412), .ZN(
        P1_U3067) );
  AOI22_X1 U23346 ( .A1(n20748), .A2(n20423), .B1(n20747), .B2(n20422), .ZN(
        n20415) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20749), .ZN(n20414) );
  OAI211_X1 U23348 ( .C1(n20752), .C2(n20441), .A(n20415), .B(n20414), .ZN(
        P1_U3068) );
  AOI22_X1 U23349 ( .A1(n20754), .A2(n20423), .B1(n20753), .B2(n20422), .ZN(
        n20417) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20755), .ZN(n20416) );
  OAI211_X1 U23351 ( .C1(n20758), .C2(n20441), .A(n20417), .B(n20416), .ZN(
        P1_U3069) );
  AOI22_X1 U23352 ( .A1(n20824), .A2(n20423), .B1(n20823), .B2(n20422), .ZN(
        n20419) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20759), .ZN(n20418) );
  OAI211_X1 U23354 ( .C1(n20762), .C2(n20441), .A(n20419), .B(n20418), .ZN(
        P1_U3070) );
  AOI22_X1 U23355 ( .A1(n20764), .A2(n20423), .B1(n20763), .B2(n20422), .ZN(
        n20421) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20765), .ZN(n20420) );
  OAI211_X1 U23357 ( .C1(n20768), .C2(n20441), .A(n20421), .B(n20420), .ZN(
        P1_U3071) );
  AOI22_X1 U23358 ( .A1(n20840), .A2(n20423), .B1(n20839), .B2(n20422), .ZN(
        n20427) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20771), .ZN(n20426) );
  OAI211_X1 U23360 ( .C1(n20776), .C2(n20441), .A(n20427), .B(n20426), .ZN(
        P1_U3072) );
  NOR2_X1 U23361 ( .A1(n20690), .A2(n20428), .ZN(n20449) );
  AOI21_X1 U23362 ( .B1(n20490), .B2(n20692), .A(n20449), .ZN(n20430) );
  OAI22_X1 U23363 ( .A1(n20430), .A2(n20779), .B1(n20428), .B2(n20929), .ZN(
        n20448) );
  AOI22_X1 U23364 ( .A1(n20725), .A2(n20449), .B1(n20724), .B2(n20448), .ZN(
        n20434) );
  NOR2_X1 U23365 ( .A1(n20429), .A2(n20779), .ZN(n20495) );
  OAI21_X1 U23366 ( .B1(n20495), .B2(n20695), .A(n20430), .ZN(n20431) );
  OAI211_X1 U23367 ( .C1(n20790), .C2(n20432), .A(n20789), .B(n20431), .ZN(
        n20451) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20451), .B1(
        n20450), .B2(n20733), .ZN(n20433) );
  OAI211_X1 U23369 ( .C1(n20736), .C2(n20484), .A(n20434), .B(n20433), .ZN(
        P1_U3073) );
  AOI22_X1 U23370 ( .A1(n20797), .A2(n20449), .B1(n20796), .B2(n20448), .ZN(
        n20436) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20451), .B1(
        n20450), .B2(n20737), .ZN(n20435) );
  OAI211_X1 U23372 ( .C1(n20740), .C2(n20484), .A(n20436), .B(n20435), .ZN(
        P1_U3074) );
  AOI22_X1 U23373 ( .A1(n20742), .A2(n20449), .B1(n20741), .B2(n20448), .ZN(
        n20438) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20451), .B1(
        n20450), .B2(n20743), .ZN(n20437) );
  OAI211_X1 U23375 ( .C1(n20746), .C2(n20484), .A(n20438), .B(n20437), .ZN(
        P1_U3075) );
  AOI22_X1 U23376 ( .A1(n20748), .A2(n20449), .B1(n20747), .B2(n20448), .ZN(
        n20440) );
  INV_X1 U23377 ( .A(n20484), .ZN(n20477) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20451), .B1(
        n20477), .B2(n20812), .ZN(n20439) );
  OAI211_X1 U23379 ( .C1(n20815), .C2(n20441), .A(n20440), .B(n20439), .ZN(
        P1_U3076) );
  AOI22_X1 U23380 ( .A1(n20754), .A2(n20449), .B1(n20753), .B2(n20448), .ZN(
        n20443) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20451), .B1(
        n20450), .B2(n20755), .ZN(n20442) );
  OAI211_X1 U23382 ( .C1(n20758), .C2(n20484), .A(n20443), .B(n20442), .ZN(
        P1_U3077) );
  AOI22_X1 U23383 ( .A1(n20824), .A2(n20449), .B1(n20823), .B2(n20448), .ZN(
        n20445) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20451), .B1(
        n20450), .B2(n20759), .ZN(n20444) );
  OAI211_X1 U23385 ( .C1(n20762), .C2(n20484), .A(n20445), .B(n20444), .ZN(
        P1_U3078) );
  AOI22_X1 U23386 ( .A1(n20764), .A2(n20449), .B1(n20763), .B2(n20448), .ZN(
        n20447) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20451), .B1(
        n20450), .B2(n20765), .ZN(n20446) );
  OAI211_X1 U23388 ( .C1(n20768), .C2(n20484), .A(n20447), .B(n20446), .ZN(
        P1_U3079) );
  AOI22_X1 U23389 ( .A1(n20840), .A2(n20449), .B1(n20839), .B2(n20448), .ZN(
        n20453) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20451), .B1(
        n20450), .B2(n20771), .ZN(n20452) );
  OAI211_X1 U23391 ( .C1(n20776), .C2(n20484), .A(n20453), .B(n20452), .ZN(
        P1_U3080) );
  NAND2_X1 U23392 ( .A1(n20690), .A2(n10313), .ZN(n20483) );
  OAI22_X1 U23393 ( .A1(n20484), .A2(n20795), .B1(n20783), .B2(n20483), .ZN(
        n20455) );
  INV_X1 U23394 ( .A(n20455), .ZN(n20464) );
  AOI21_X1 U23395 ( .B1(n20518), .B2(n20484), .A(n21085), .ZN(n20456) );
  NOR2_X1 U23396 ( .A1(n20456), .A2(n20779), .ZN(n20459) );
  NAND2_X1 U23397 ( .A1(n20490), .A2(n20727), .ZN(n20461) );
  AOI22_X1 U23398 ( .A1(n20459), .A2(n20461), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20483), .ZN(n20458) );
  NAND3_X1 U23399 ( .A1(n20730), .A2(n20458), .A3(n20457), .ZN(n20487) );
  INV_X1 U23400 ( .A(n20459), .ZN(n20462) );
  OAI22_X1 U23401 ( .A1(n20462), .A2(n20461), .B1(n20722), .B2(n20460), .ZN(
        n20486) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20487), .B1(
        n20724), .B2(n20486), .ZN(n20463) );
  OAI211_X1 U23403 ( .C1(n20736), .C2(n20518), .A(n20464), .B(n20463), .ZN(
        P1_U3081) );
  INV_X1 U23404 ( .A(n20483), .ZN(n20476) );
  AOI22_X1 U23405 ( .A1(n20477), .A2(n20737), .B1(n20476), .B2(n20797), .ZN(
        n20466) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20487), .B1(
        n20796), .B2(n20486), .ZN(n20465) );
  OAI211_X1 U23407 ( .C1(n20740), .C2(n20518), .A(n20466), .B(n20465), .ZN(
        P1_U3082) );
  OAI22_X1 U23408 ( .A1(n20518), .A2(n20746), .B1(n20483), .B2(n20803), .ZN(
        n20467) );
  INV_X1 U23409 ( .A(n20467), .ZN(n20469) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20487), .B1(
        n20741), .B2(n20486), .ZN(n20468) );
  OAI211_X1 U23411 ( .C1(n20808), .C2(n20484), .A(n20469), .B(n20468), .ZN(
        P1_U3083) );
  OAI22_X1 U23412 ( .A1(n20484), .A2(n20815), .B1(n20483), .B2(n20810), .ZN(
        n20470) );
  INV_X1 U23413 ( .A(n20470), .ZN(n20472) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20487), .B1(
        n20747), .B2(n20486), .ZN(n20471) );
  OAI211_X1 U23415 ( .C1(n20752), .C2(n20518), .A(n20472), .B(n20471), .ZN(
        P1_U3084) );
  OAI22_X1 U23416 ( .A1(n20484), .A2(n20822), .B1(n20483), .B2(n20817), .ZN(
        n20473) );
  INV_X1 U23417 ( .A(n20473), .ZN(n20475) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20487), .B1(
        n20753), .B2(n20486), .ZN(n20474) );
  OAI211_X1 U23419 ( .C1(n20758), .C2(n20518), .A(n20475), .B(n20474), .ZN(
        P1_U3085) );
  AOI22_X1 U23420 ( .A1(n20477), .A2(n20759), .B1(n20476), .B2(n20824), .ZN(
        n20479) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20487), .B1(
        n20823), .B2(n20486), .ZN(n20478) );
  OAI211_X1 U23422 ( .C1(n20762), .C2(n20518), .A(n20479), .B(n20478), .ZN(
        P1_U3086) );
  OAI22_X1 U23423 ( .A1(n20518), .A2(n20768), .B1(n20483), .B2(n20832), .ZN(
        n20480) );
  INV_X1 U23424 ( .A(n20480), .ZN(n20482) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20487), .B1(
        n20763), .B2(n20486), .ZN(n20481) );
  OAI211_X1 U23426 ( .C1(n20837), .C2(n20484), .A(n20482), .B(n20481), .ZN(
        P1_U3087) );
  OAI22_X1 U23427 ( .A1(n20484), .A2(n20848), .B1(n20483), .B2(n20614), .ZN(
        n20485) );
  INV_X1 U23428 ( .A(n20485), .ZN(n20489) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20487), .B1(
        n20839), .B2(n20486), .ZN(n20488) );
  OAI211_X1 U23430 ( .C1(n20776), .C2(n20518), .A(n20489), .B(n20488), .ZN(
        P1_U3088) );
  INV_X1 U23431 ( .A(n20514), .ZN(n20520) );
  AOI21_X1 U23432 ( .B1(n20490), .B2(n20777), .A(n20520), .ZN(n20494) );
  OR2_X1 U23433 ( .A1(n20494), .A2(n20779), .ZN(n20492) );
  NAND2_X1 U23434 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n10313), .ZN(n20491) );
  NAND2_X1 U23435 ( .A1(n20492), .A2(n20491), .ZN(n20519) );
  INV_X1 U23436 ( .A(n20519), .ZN(n20513) );
  OAI22_X1 U23437 ( .A1(n20783), .A2(n20514), .B1(n20513), .B2(n20782), .ZN(
        n20493) );
  INV_X1 U23438 ( .A(n20493), .ZN(n20499) );
  OAI21_X1 U23439 ( .B1(n20787), .B2(n20495), .A(n20494), .ZN(n20496) );
  OAI211_X1 U23440 ( .C1(n10313), .C2(n20790), .A(n20789), .B(n20496), .ZN(
        n20522) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20522), .B1(
        n20551), .B2(n20792), .ZN(n20498) );
  OAI211_X1 U23442 ( .C1(n20795), .C2(n20518), .A(n20499), .B(n20498), .ZN(
        P1_U3089) );
  AOI22_X1 U23443 ( .A1(n20797), .A2(n20520), .B1(n20796), .B2(n20519), .ZN(
        n20501) );
  INV_X1 U23444 ( .A(n20518), .ZN(n20521) );
  AOI22_X1 U23445 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20522), .B1(
        n20521), .B2(n20737), .ZN(n20500) );
  OAI211_X1 U23446 ( .C1(n20740), .C2(n20525), .A(n20501), .B(n20500), .ZN(
        P1_U3090) );
  OAI22_X1 U23447 ( .A1(n20803), .A2(n20514), .B1(n20513), .B2(n20802), .ZN(
        n20502) );
  INV_X1 U23448 ( .A(n20502), .ZN(n20504) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20522), .B1(
        n20521), .B2(n20743), .ZN(n20503) );
  OAI211_X1 U23450 ( .C1(n20746), .C2(n20525), .A(n20504), .B(n20503), .ZN(
        P1_U3091) );
  OAI22_X1 U23451 ( .A1(n20810), .A2(n20514), .B1(n20513), .B2(n20809), .ZN(
        n20505) );
  INV_X1 U23452 ( .A(n20505), .ZN(n20507) );
  AOI22_X1 U23453 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20522), .B1(
        n20551), .B2(n20812), .ZN(n20506) );
  OAI211_X1 U23454 ( .C1(n20815), .C2(n20518), .A(n20507), .B(n20506), .ZN(
        P1_U3092) );
  OAI22_X1 U23455 ( .A1(n20817), .A2(n20514), .B1(n20513), .B2(n20816), .ZN(
        n20508) );
  INV_X1 U23456 ( .A(n20508), .ZN(n20510) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20522), .B1(
        n20551), .B2(n20819), .ZN(n20509) );
  OAI211_X1 U23458 ( .C1(n20822), .C2(n20518), .A(n20510), .B(n20509), .ZN(
        P1_U3093) );
  AOI22_X1 U23459 ( .A1(n20824), .A2(n20520), .B1(n20823), .B2(n20519), .ZN(
        n20512) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20522), .B1(
        n20551), .B2(n20825), .ZN(n20511) );
  OAI211_X1 U23461 ( .C1(n20828), .C2(n20518), .A(n20512), .B(n20511), .ZN(
        P1_U3094) );
  OAI22_X1 U23462 ( .A1(n20832), .A2(n20514), .B1(n20513), .B2(n20830), .ZN(
        n20515) );
  INV_X1 U23463 ( .A(n20515), .ZN(n20517) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20522), .B1(
        n20551), .B2(n20834), .ZN(n20516) );
  OAI211_X1 U23465 ( .C1(n20837), .C2(n20518), .A(n20517), .B(n20516), .ZN(
        P1_U3095) );
  AOI22_X1 U23466 ( .A1(n20520), .A2(n20840), .B1(n20839), .B2(n20519), .ZN(
        n20524) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20522), .B1(
        n20521), .B2(n20771), .ZN(n20523) );
  OAI211_X1 U23468 ( .C1(n20776), .C2(n20525), .A(n20524), .B(n20523), .ZN(
        P1_U3096) );
  NOR3_X1 U23469 ( .A1(n20658), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20558) );
  INV_X1 U23470 ( .A(n20558), .ZN(n20555) );
  NOR2_X1 U23471 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20555), .ZN(
        n20550) );
  AND2_X1 U23472 ( .A1(n20527), .A2(n20655), .ZN(n20622) );
  AOI21_X1 U23473 ( .B1(n20622), .B2(n20528), .A(n20550), .ZN(n20532) );
  AND2_X1 U23474 ( .A1(n20529), .A2(n20582), .ZN(n20656) );
  INV_X1 U23475 ( .A(n20656), .ZN(n20660) );
  OAI22_X1 U23476 ( .A1(n20532), .A2(n20779), .B1(n20660), .B2(n20530), .ZN(
        n20549) );
  AOI22_X1 U23477 ( .A1(n20725), .A2(n20550), .B1(n20724), .B2(n20549), .ZN(
        n20536) );
  INV_X1 U23478 ( .A(n20578), .ZN(n20531) );
  OAI21_X1 U23479 ( .B1(n20531), .B2(n20551), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20533) );
  NAND2_X1 U23480 ( .A1(n20533), .A2(n20532), .ZN(n20534) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20552), .B1(
        n20551), .B2(n20733), .ZN(n20535) );
  OAI211_X1 U23482 ( .C1(n20736), .C2(n20578), .A(n20536), .B(n20535), .ZN(
        P1_U3097) );
  AOI22_X1 U23483 ( .A1(n20797), .A2(n20550), .B1(n20549), .B2(n20796), .ZN(
        n20538) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20552), .B1(
        n20551), .B2(n20737), .ZN(n20537) );
  OAI211_X1 U23485 ( .C1(n20740), .C2(n20578), .A(n20538), .B(n20537), .ZN(
        P1_U3098) );
  AOI22_X1 U23486 ( .A1(n20742), .A2(n20550), .B1(n20741), .B2(n20549), .ZN(
        n20540) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20552), .B1(
        n20551), .B2(n20743), .ZN(n20539) );
  OAI211_X1 U23488 ( .C1(n20746), .C2(n20578), .A(n20540), .B(n20539), .ZN(
        P1_U3099) );
  AOI22_X1 U23489 ( .A1(n20748), .A2(n20550), .B1(n20747), .B2(n20549), .ZN(
        n20542) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20552), .B1(
        n20551), .B2(n20749), .ZN(n20541) );
  OAI211_X1 U23491 ( .C1(n20752), .C2(n20578), .A(n20542), .B(n20541), .ZN(
        P1_U3100) );
  AOI22_X1 U23492 ( .A1(n20754), .A2(n20550), .B1(n20753), .B2(n20549), .ZN(
        n20544) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20552), .B1(
        n20551), .B2(n20755), .ZN(n20543) );
  OAI211_X1 U23494 ( .C1(n20758), .C2(n20578), .A(n20544), .B(n20543), .ZN(
        P1_U3101) );
  AOI22_X1 U23495 ( .A1(n20824), .A2(n20550), .B1(n20549), .B2(n20823), .ZN(
        n20546) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20552), .B1(
        n20551), .B2(n20759), .ZN(n20545) );
  OAI211_X1 U23497 ( .C1(n20762), .C2(n20578), .A(n20546), .B(n20545), .ZN(
        P1_U3102) );
  AOI22_X1 U23498 ( .A1(n20764), .A2(n20550), .B1(n20763), .B2(n20549), .ZN(
        n20548) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20552), .B1(
        n20551), .B2(n20765), .ZN(n20547) );
  OAI211_X1 U23500 ( .C1(n20768), .C2(n20578), .A(n20548), .B(n20547), .ZN(
        P1_U3103) );
  AOI22_X1 U23501 ( .A1(n20840), .A2(n20550), .B1(n20839), .B2(n20549), .ZN(
        n20554) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20552), .B1(
        n20551), .B2(n20771), .ZN(n20553) );
  OAI211_X1 U23503 ( .C1(n20776), .C2(n20578), .A(n20554), .B(n20553), .ZN(
        P1_U3104) );
  NOR2_X1 U23504 ( .A1(n20690), .A2(n20555), .ZN(n20574) );
  AOI21_X1 U23505 ( .B1(n20622), .B2(n20692), .A(n20574), .ZN(n20556) );
  OAI22_X1 U23506 ( .A1(n20556), .A2(n20779), .B1(n20555), .B2(n20929), .ZN(
        n20573) );
  AOI22_X1 U23507 ( .A1(n20725), .A2(n20574), .B1(n20724), .B2(n20573), .ZN(
        n20560) );
  AND2_X1 U23508 ( .A1(n20629), .A2(n20790), .ZN(n20625) );
  OAI21_X1 U23509 ( .B1(n20625), .B2(n20695), .A(n20556), .ZN(n20557) );
  OAI211_X1 U23510 ( .C1(n20790), .C2(n20558), .A(n20789), .B(n20557), .ZN(
        n20575) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20575), .B1(
        n20616), .B2(n20792), .ZN(n20559) );
  OAI211_X1 U23512 ( .C1(n20795), .C2(n20578), .A(n20560), .B(n20559), .ZN(
        P1_U3105) );
  AOI22_X1 U23513 ( .A1(n20797), .A2(n20574), .B1(n20573), .B2(n20796), .ZN(
        n20562) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20575), .B1(
        n20616), .B2(n20798), .ZN(n20561) );
  OAI211_X1 U23515 ( .C1(n20801), .C2(n20578), .A(n20562), .B(n20561), .ZN(
        P1_U3106) );
  AOI22_X1 U23516 ( .A1(n20742), .A2(n20574), .B1(n20741), .B2(n20573), .ZN(
        n20564) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20575), .B1(
        n20616), .B2(n20805), .ZN(n20563) );
  OAI211_X1 U23518 ( .C1(n20808), .C2(n20578), .A(n20564), .B(n20563), .ZN(
        P1_U3107) );
  AOI22_X1 U23519 ( .A1(n20748), .A2(n20574), .B1(n20747), .B2(n20573), .ZN(
        n20566) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20575), .B1(
        n20616), .B2(n20812), .ZN(n20565) );
  OAI211_X1 U23521 ( .C1(n20815), .C2(n20578), .A(n20566), .B(n20565), .ZN(
        P1_U3108) );
  AOI22_X1 U23522 ( .A1(n20754), .A2(n20574), .B1(n20753), .B2(n20573), .ZN(
        n20568) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20575), .B1(
        n20616), .B2(n20819), .ZN(n20567) );
  OAI211_X1 U23524 ( .C1(n20822), .C2(n20578), .A(n20568), .B(n20567), .ZN(
        P1_U3109) );
  AOI22_X1 U23525 ( .A1(n20824), .A2(n20574), .B1(n20573), .B2(n20823), .ZN(
        n20570) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20575), .B1(
        n20616), .B2(n20825), .ZN(n20569) );
  OAI211_X1 U23527 ( .C1(n20828), .C2(n20578), .A(n20570), .B(n20569), .ZN(
        P1_U3110) );
  AOI22_X1 U23528 ( .A1(n20764), .A2(n20574), .B1(n20763), .B2(n20573), .ZN(
        n20572) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20575), .B1(
        n20616), .B2(n20834), .ZN(n20571) );
  OAI211_X1 U23530 ( .C1(n20837), .C2(n20578), .A(n20572), .B(n20571), .ZN(
        P1_U3111) );
  AOI22_X1 U23531 ( .A1(n20840), .A2(n20574), .B1(n20839), .B2(n20573), .ZN(
        n20577) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20575), .B1(
        n20616), .B2(n20842), .ZN(n20576) );
  OAI211_X1 U23533 ( .C1(n20848), .C2(n20578), .A(n20577), .B(n20576), .ZN(
        P1_U3112) );
  INV_X1 U23534 ( .A(n20616), .ZN(n20580) );
  NAND3_X1 U23535 ( .A1(n20580), .A2(n20790), .A3(n20649), .ZN(n20581) );
  NAND2_X1 U23536 ( .A1(n20581), .A2(n20652), .ZN(n20587) );
  AND2_X1 U23537 ( .A1(n20622), .A2(n20727), .ZN(n20591) );
  OR2_X1 U23538 ( .A1(n20582), .A2(n20658), .ZN(n20723) );
  INV_X1 U23539 ( .A(n20723), .ZN(n20583) );
  NOR3_X1 U23540 ( .A1(n20658), .A2(n20585), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20627) );
  INV_X1 U23541 ( .A(n20627), .ZN(n20623) );
  NOR2_X1 U23542 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20623), .ZN(
        n20606) );
  INV_X1 U23543 ( .A(n20606), .ZN(n20613) );
  OAI22_X1 U23544 ( .A1(n20649), .A2(n20736), .B1(n20783), .B2(n20613), .ZN(
        n20586) );
  INV_X1 U23545 ( .A(n20586), .ZN(n20594) );
  INV_X1 U23546 ( .A(n20587), .ZN(n20592) );
  NAND2_X1 U23547 ( .A1(n20723), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20729) );
  OAI21_X1 U23548 ( .B1(n20664), .B2(n20606), .A(n20729), .ZN(n20588) );
  INV_X1 U23549 ( .A(n20588), .ZN(n20590) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20617), .B1(
        n20616), .B2(n20733), .ZN(n20593) );
  OAI211_X1 U23551 ( .C1(n20620), .C2(n20782), .A(n20594), .B(n20593), .ZN(
        P1_U3113) );
  AOI22_X1 U23552 ( .A1(n20616), .A2(n20737), .B1(n20797), .B2(n20606), .ZN(
        n20596) );
  INV_X1 U23553 ( .A(n20649), .ZN(n20607) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20617), .B1(
        n20607), .B2(n20798), .ZN(n20595) );
  OAI211_X1 U23555 ( .C1(n20620), .C2(n20669), .A(n20596), .B(n20595), .ZN(
        P1_U3114) );
  OAI22_X1 U23556 ( .A1(n20649), .A2(n20746), .B1(n20803), .B2(n20613), .ZN(
        n20597) );
  INV_X1 U23557 ( .A(n20597), .ZN(n20599) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20617), .B1(
        n20616), .B2(n20743), .ZN(n20598) );
  OAI211_X1 U23559 ( .C1(n20620), .C2(n20802), .A(n20599), .B(n20598), .ZN(
        P1_U3115) );
  OAI22_X1 U23560 ( .A1(n20649), .A2(n20752), .B1(n20810), .B2(n20613), .ZN(
        n20600) );
  INV_X1 U23561 ( .A(n20600), .ZN(n20602) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20617), .B1(
        n20616), .B2(n20749), .ZN(n20601) );
  OAI211_X1 U23563 ( .C1(n20620), .C2(n20809), .A(n20602), .B(n20601), .ZN(
        P1_U3116) );
  OAI22_X1 U23564 ( .A1(n20649), .A2(n20758), .B1(n20817), .B2(n20613), .ZN(
        n20603) );
  INV_X1 U23565 ( .A(n20603), .ZN(n20605) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20617), .B1(
        n20616), .B2(n20755), .ZN(n20604) );
  OAI211_X1 U23567 ( .C1(n20620), .C2(n20816), .A(n20605), .B(n20604), .ZN(
        P1_U3117) );
  AOI22_X1 U23568 ( .A1(n20616), .A2(n20759), .B1(n20824), .B2(n20606), .ZN(
        n20609) );
  AOI22_X1 U23569 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20617), .B1(
        n20607), .B2(n20825), .ZN(n20608) );
  OAI211_X1 U23570 ( .C1(n20620), .C2(n20678), .A(n20609), .B(n20608), .ZN(
        P1_U3118) );
  OAI22_X1 U23571 ( .A1(n20649), .A2(n20768), .B1(n20832), .B2(n20613), .ZN(
        n20610) );
  INV_X1 U23572 ( .A(n20610), .ZN(n20612) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20617), .B1(
        n20616), .B2(n20765), .ZN(n20611) );
  OAI211_X1 U23574 ( .C1(n20620), .C2(n20830), .A(n20612), .B(n20611), .ZN(
        P1_U3119) );
  OAI22_X1 U23575 ( .A1(n20649), .A2(n20776), .B1(n20614), .B2(n20613), .ZN(
        n20615) );
  INV_X1 U23576 ( .A(n20615), .ZN(n20619) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20617), .B1(
        n20616), .B2(n20771), .ZN(n20618) );
  OAI211_X1 U23578 ( .C1(n20620), .C2(n20686), .A(n20619), .B(n20618), .ZN(
        P1_U3120) );
  NOR2_X1 U23579 ( .A1(n20621), .A2(n20658), .ZN(n20645) );
  AOI21_X1 U23580 ( .B1(n20622), .B2(n20777), .A(n20645), .ZN(n20624) );
  OAI22_X1 U23581 ( .A1(n20624), .A2(n20779), .B1(n20623), .B2(n20929), .ZN(
        n20644) );
  AOI22_X1 U23582 ( .A1(n20725), .A2(n20645), .B1(n20724), .B2(n20644), .ZN(
        n20631) );
  OAI21_X1 U23583 ( .B1(n20787), .B2(n20625), .A(n20624), .ZN(n20626) );
  OAI211_X1 U23584 ( .C1(n20790), .C2(n20627), .A(n20789), .B(n20626), .ZN(
        n20646) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20646), .B1(
        n20682), .B2(n20792), .ZN(n20630) );
  OAI211_X1 U23586 ( .C1(n20795), .C2(n20649), .A(n20631), .B(n20630), .ZN(
        P1_U3121) );
  AOI22_X1 U23587 ( .A1(n20797), .A2(n20645), .B1(n20644), .B2(n20796), .ZN(
        n20633) );
  AOI22_X1 U23588 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20646), .B1(
        n20682), .B2(n20798), .ZN(n20632) );
  OAI211_X1 U23589 ( .C1(n20801), .C2(n20649), .A(n20633), .B(n20632), .ZN(
        P1_U3122) );
  AOI22_X1 U23590 ( .A1(n20742), .A2(n20645), .B1(n20644), .B2(n20741), .ZN(
        n20635) );
  AOI22_X1 U23591 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20646), .B1(
        n20682), .B2(n20805), .ZN(n20634) );
  OAI211_X1 U23592 ( .C1(n20808), .C2(n20649), .A(n20635), .B(n20634), .ZN(
        P1_U3123) );
  AOI22_X1 U23593 ( .A1(n20748), .A2(n20645), .B1(n20644), .B2(n20747), .ZN(
        n20637) );
  AOI22_X1 U23594 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20646), .B1(
        n20682), .B2(n20812), .ZN(n20636) );
  OAI211_X1 U23595 ( .C1(n20815), .C2(n20649), .A(n20637), .B(n20636), .ZN(
        P1_U3124) );
  AOI22_X1 U23596 ( .A1(n20754), .A2(n20645), .B1(n20644), .B2(n20753), .ZN(
        n20639) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20646), .B1(
        n20682), .B2(n20819), .ZN(n20638) );
  OAI211_X1 U23598 ( .C1(n20822), .C2(n20649), .A(n20639), .B(n20638), .ZN(
        P1_U3125) );
  AOI22_X1 U23599 ( .A1(n20824), .A2(n20645), .B1(n20644), .B2(n20823), .ZN(
        n20641) );
  AOI22_X1 U23600 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20646), .B1(
        n20682), .B2(n20825), .ZN(n20640) );
  OAI211_X1 U23601 ( .C1(n20828), .C2(n20649), .A(n20641), .B(n20640), .ZN(
        P1_U3126) );
  AOI22_X1 U23602 ( .A1(n20764), .A2(n20645), .B1(n20644), .B2(n20763), .ZN(
        n20643) );
  AOI22_X1 U23603 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20646), .B1(
        n20682), .B2(n20834), .ZN(n20642) );
  OAI211_X1 U23604 ( .C1(n20837), .C2(n20649), .A(n20643), .B(n20642), .ZN(
        P1_U3127) );
  AOI22_X1 U23605 ( .A1(n20840), .A2(n20645), .B1(n20839), .B2(n20644), .ZN(
        n20648) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20646), .B1(
        n20682), .B2(n20842), .ZN(n20647) );
  OAI211_X1 U23607 ( .C1(n20848), .C2(n20649), .A(n20648), .B(n20647), .ZN(
        P1_U3128) );
  INV_X1 U23608 ( .A(n20682), .ZN(n20650) );
  NAND2_X1 U23609 ( .A1(n20650), .A2(n20790), .ZN(n20653) );
  OAI21_X1 U23610 ( .B1(n20653), .B2(n20714), .A(n20652), .ZN(n20662) );
  OR2_X1 U23611 ( .A1(n20655), .A2(n20654), .ZN(n20691) );
  NOR2_X1 U23612 ( .A1(n20691), .A2(n20727), .ZN(n20659) );
  INV_X1 U23613 ( .A(n20722), .ZN(n20657) );
  NOR3_X1 U23614 ( .A1(n13020), .A2(n20658), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20697) );
  INV_X1 U23615 ( .A(n20697), .ZN(n20693) );
  NOR2_X1 U23616 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20693), .ZN(
        n20681) );
  AOI22_X1 U23617 ( .A1(n20714), .A2(n20792), .B1(n20725), .B2(n20681), .ZN(
        n20666) );
  INV_X1 U23618 ( .A(n20659), .ZN(n20661) );
  AOI22_X1 U23619 ( .A1(n20662), .A2(n20661), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20660), .ZN(n20663) );
  AOI22_X1 U23620 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20733), .ZN(n20665) );
  OAI211_X1 U23621 ( .C1(n20687), .C2(n20782), .A(n20666), .B(n20665), .ZN(
        P1_U3129) );
  AOI22_X1 U23622 ( .A1(n20714), .A2(n20798), .B1(n20797), .B2(n20681), .ZN(
        n20668) );
  AOI22_X1 U23623 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20737), .ZN(n20667) );
  OAI211_X1 U23624 ( .C1(n20687), .C2(n20669), .A(n20668), .B(n20667), .ZN(
        P1_U3130) );
  AOI22_X1 U23625 ( .A1(n20714), .A2(n20805), .B1(n20742), .B2(n20681), .ZN(
        n20671) );
  AOI22_X1 U23626 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20743), .ZN(n20670) );
  OAI211_X1 U23627 ( .C1(n20687), .C2(n20802), .A(n20671), .B(n20670), .ZN(
        P1_U3131) );
  AOI22_X1 U23628 ( .A1(n20714), .A2(n20812), .B1(n20748), .B2(n20681), .ZN(
        n20673) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20749), .ZN(n20672) );
  OAI211_X1 U23630 ( .C1(n20687), .C2(n20809), .A(n20673), .B(n20672), .ZN(
        P1_U3132) );
  AOI22_X1 U23631 ( .A1(n20714), .A2(n20819), .B1(n20754), .B2(n20681), .ZN(
        n20675) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20755), .ZN(n20674) );
  OAI211_X1 U23633 ( .C1(n20687), .C2(n20816), .A(n20675), .B(n20674), .ZN(
        P1_U3133) );
  AOI22_X1 U23634 ( .A1(n20714), .A2(n20825), .B1(n20824), .B2(n20681), .ZN(
        n20677) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20759), .ZN(n20676) );
  OAI211_X1 U23636 ( .C1(n20687), .C2(n20678), .A(n20677), .B(n20676), .ZN(
        P1_U3134) );
  AOI22_X1 U23637 ( .A1(n20714), .A2(n20834), .B1(n20764), .B2(n20681), .ZN(
        n20680) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20765), .ZN(n20679) );
  OAI211_X1 U23639 ( .C1(n20687), .C2(n20830), .A(n20680), .B(n20679), .ZN(
        P1_U3135) );
  AOI22_X1 U23640 ( .A1(n20714), .A2(n20842), .B1(n20840), .B2(n20681), .ZN(
        n20685) );
  AOI22_X1 U23641 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20683), .B1(
        n20682), .B2(n20771), .ZN(n20684) );
  OAI211_X1 U23642 ( .C1(n20687), .C2(n20686), .A(n20685), .B(n20684), .ZN(
        P1_U3136) );
  INV_X1 U23643 ( .A(n20688), .ZN(n20689) );
  NOR2_X1 U23644 ( .A1(n20690), .A2(n20693), .ZN(n20713) );
  AOI21_X1 U23645 ( .B1(n20778), .B2(n20692), .A(n20713), .ZN(n20694) );
  OAI22_X1 U23646 ( .A1(n20694), .A2(n20779), .B1(n20693), .B2(n20929), .ZN(
        n20712) );
  AOI22_X1 U23647 ( .A1(n20725), .A2(n20713), .B1(n20724), .B2(n20712), .ZN(
        n20699) );
  NOR2_X1 U23648 ( .A1(n20719), .A2(n20779), .ZN(n20786) );
  OAI21_X1 U23649 ( .B1(n20786), .B2(n20695), .A(n20694), .ZN(n20696) );
  OAI211_X1 U23650 ( .C1(n20790), .C2(n20697), .A(n20789), .B(n20696), .ZN(
        n20715) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n20733), .ZN(n20698) );
  OAI211_X1 U23652 ( .C1(n20736), .C2(n20732), .A(n20699), .B(n20698), .ZN(
        P1_U3137) );
  AOI22_X1 U23653 ( .A1(n20797), .A2(n20713), .B1(n20796), .B2(n20712), .ZN(
        n20701) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n20737), .ZN(n20700) );
  OAI211_X1 U23655 ( .C1(n20740), .C2(n20732), .A(n20701), .B(n20700), .ZN(
        P1_U3138) );
  AOI22_X1 U23656 ( .A1(n20742), .A2(n20713), .B1(n20741), .B2(n20712), .ZN(
        n20703) );
  AOI22_X1 U23657 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n20743), .ZN(n20702) );
  OAI211_X1 U23658 ( .C1(n20746), .C2(n20732), .A(n20703), .B(n20702), .ZN(
        P1_U3139) );
  AOI22_X1 U23659 ( .A1(n20748), .A2(n20713), .B1(n20747), .B2(n20712), .ZN(
        n20705) );
  AOI22_X1 U23660 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n20749), .ZN(n20704) );
  OAI211_X1 U23661 ( .C1(n20752), .C2(n20732), .A(n20705), .B(n20704), .ZN(
        P1_U3140) );
  AOI22_X1 U23662 ( .A1(n20754), .A2(n20713), .B1(n20753), .B2(n20712), .ZN(
        n20707) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n20755), .ZN(n20706) );
  OAI211_X1 U23664 ( .C1(n20758), .C2(n20732), .A(n20707), .B(n20706), .ZN(
        P1_U3141) );
  AOI22_X1 U23665 ( .A1(n20824), .A2(n20713), .B1(n20823), .B2(n20712), .ZN(
        n20709) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n20759), .ZN(n20708) );
  OAI211_X1 U23667 ( .C1(n20762), .C2(n20732), .A(n20709), .B(n20708), .ZN(
        P1_U3142) );
  AOI22_X1 U23668 ( .A1(n20764), .A2(n20713), .B1(n20763), .B2(n20712), .ZN(
        n20711) );
  AOI22_X1 U23669 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n20765), .ZN(n20710) );
  OAI211_X1 U23670 ( .C1(n20768), .C2(n20732), .A(n20711), .B(n20710), .ZN(
        P1_U3143) );
  AOI22_X1 U23671 ( .A1(n20840), .A2(n20713), .B1(n20839), .B2(n20712), .ZN(
        n20717) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20715), .B1(
        n20714), .B2(n20771), .ZN(n20716) );
  OAI211_X1 U23673 ( .C1(n20776), .C2(n20732), .A(n20717), .B(n20716), .ZN(
        P1_U3144) );
  INV_X1 U23674 ( .A(n20791), .ZN(n20720) );
  NOR2_X1 U23675 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20720), .ZN(
        n20770) );
  NAND3_X1 U23676 ( .A1(n20778), .A2(n20727), .A3(n20790), .ZN(n20721) );
  OAI21_X1 U23677 ( .B1(n20723), .B2(n20722), .A(n20721), .ZN(n20769) );
  AOI22_X1 U23678 ( .A1(n20725), .A2(n20770), .B1(n20724), .B2(n20769), .ZN(
        n20735) );
  AOI21_X1 U23679 ( .B1(n20732), .B2(n20847), .A(n21085), .ZN(n20726) );
  AOI21_X1 U23680 ( .B1(n20778), .B2(n20727), .A(n20726), .ZN(n20728) );
  NOR2_X1 U23681 ( .A1(n20728), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20731) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20773), .B1(
        n20772), .B2(n20733), .ZN(n20734) );
  OAI211_X1 U23683 ( .C1(n20736), .C2(n20847), .A(n20735), .B(n20734), .ZN(
        P1_U3145) );
  AOI22_X1 U23684 ( .A1(n20797), .A2(n20770), .B1(n20796), .B2(n20769), .ZN(
        n20739) );
  AOI22_X1 U23685 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20773), .B1(
        n20772), .B2(n20737), .ZN(n20738) );
  OAI211_X1 U23686 ( .C1(n20740), .C2(n20847), .A(n20739), .B(n20738), .ZN(
        P1_U3146) );
  AOI22_X1 U23687 ( .A1(n20742), .A2(n20770), .B1(n20741), .B2(n20769), .ZN(
        n20745) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20773), .B1(
        n20772), .B2(n20743), .ZN(n20744) );
  OAI211_X1 U23689 ( .C1(n20746), .C2(n20847), .A(n20745), .B(n20744), .ZN(
        P1_U3147) );
  AOI22_X1 U23690 ( .A1(n20748), .A2(n20770), .B1(n20747), .B2(n20769), .ZN(
        n20751) );
  AOI22_X1 U23691 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20773), .B1(
        n20772), .B2(n20749), .ZN(n20750) );
  OAI211_X1 U23692 ( .C1(n20752), .C2(n20847), .A(n20751), .B(n20750), .ZN(
        P1_U3148) );
  AOI22_X1 U23693 ( .A1(n20754), .A2(n20770), .B1(n20753), .B2(n20769), .ZN(
        n20757) );
  AOI22_X1 U23694 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20773), .B1(
        n20772), .B2(n20755), .ZN(n20756) );
  OAI211_X1 U23695 ( .C1(n20758), .C2(n20847), .A(n20757), .B(n20756), .ZN(
        P1_U3149) );
  AOI22_X1 U23696 ( .A1(n20824), .A2(n20770), .B1(n20823), .B2(n20769), .ZN(
        n20761) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20773), .B1(
        n20772), .B2(n20759), .ZN(n20760) );
  OAI211_X1 U23698 ( .C1(n20762), .C2(n20847), .A(n20761), .B(n20760), .ZN(
        P1_U3150) );
  AOI22_X1 U23699 ( .A1(n20764), .A2(n20770), .B1(n20763), .B2(n20769), .ZN(
        n20767) );
  AOI22_X1 U23700 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20773), .B1(
        n20772), .B2(n20765), .ZN(n20766) );
  OAI211_X1 U23701 ( .C1(n20768), .C2(n20847), .A(n20767), .B(n20766), .ZN(
        P1_U3151) );
  AOI22_X1 U23702 ( .A1(n20840), .A2(n20770), .B1(n20839), .B2(n20769), .ZN(
        n20775) );
  AOI22_X1 U23703 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20773), .B1(
        n20772), .B2(n20771), .ZN(n20774) );
  OAI211_X1 U23704 ( .C1(n20776), .C2(n20847), .A(n20775), .B(n20774), .ZN(
        P1_U3152) );
  INV_X1 U23705 ( .A(n20831), .ZN(n20841) );
  AOI21_X1 U23706 ( .B1(n20778), .B2(n20777), .A(n20841), .ZN(n20785) );
  OR2_X1 U23707 ( .A1(n20785), .A2(n20779), .ZN(n20781) );
  NAND2_X1 U23708 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20791), .ZN(n20780) );
  NAND2_X1 U23709 ( .A1(n20781), .A2(n20780), .ZN(n20838) );
  INV_X1 U23710 ( .A(n20838), .ZN(n20829) );
  OAI22_X1 U23711 ( .A1(n20783), .A2(n20831), .B1(n20782), .B2(n20829), .ZN(
        n20784) );
  INV_X1 U23712 ( .A(n20784), .ZN(n20794) );
  OAI21_X1 U23713 ( .B1(n20787), .B2(n20786), .A(n20785), .ZN(n20788) );
  OAI211_X1 U23714 ( .C1(n20791), .C2(n20790), .A(n20789), .B(n20788), .ZN(
        n20844) );
  AOI22_X1 U23715 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20844), .B1(
        n20843), .B2(n20792), .ZN(n20793) );
  OAI211_X1 U23716 ( .C1(n20795), .C2(n20847), .A(n20794), .B(n20793), .ZN(
        P1_U3153) );
  AOI22_X1 U23717 ( .A1(n20797), .A2(n20841), .B1(n20796), .B2(n20838), .ZN(
        n20800) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20844), .B1(
        n20843), .B2(n20798), .ZN(n20799) );
  OAI211_X1 U23719 ( .C1(n20801), .C2(n20847), .A(n20800), .B(n20799), .ZN(
        P1_U3154) );
  OAI22_X1 U23720 ( .A1(n20803), .A2(n20831), .B1(n20802), .B2(n20829), .ZN(
        n20804) );
  INV_X1 U23721 ( .A(n20804), .ZN(n20807) );
  AOI22_X1 U23722 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20844), .B1(
        n20843), .B2(n20805), .ZN(n20806) );
  OAI211_X1 U23723 ( .C1(n20808), .C2(n20847), .A(n20807), .B(n20806), .ZN(
        P1_U3155) );
  OAI22_X1 U23724 ( .A1(n20810), .A2(n20831), .B1(n20809), .B2(n20829), .ZN(
        n20811) );
  INV_X1 U23725 ( .A(n20811), .ZN(n20814) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20844), .B1(
        n20843), .B2(n20812), .ZN(n20813) );
  OAI211_X1 U23727 ( .C1(n20815), .C2(n20847), .A(n20814), .B(n20813), .ZN(
        P1_U3156) );
  OAI22_X1 U23728 ( .A1(n20817), .A2(n20831), .B1(n20816), .B2(n20829), .ZN(
        n20818) );
  INV_X1 U23729 ( .A(n20818), .ZN(n20821) );
  AOI22_X1 U23730 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20844), .B1(
        n20843), .B2(n20819), .ZN(n20820) );
  OAI211_X1 U23731 ( .C1(n20822), .C2(n20847), .A(n20821), .B(n20820), .ZN(
        P1_U3157) );
  AOI22_X1 U23732 ( .A1(n20824), .A2(n20841), .B1(n20823), .B2(n20838), .ZN(
        n20827) );
  AOI22_X1 U23733 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20844), .B1(
        n20843), .B2(n20825), .ZN(n20826) );
  OAI211_X1 U23734 ( .C1(n20828), .C2(n20847), .A(n20827), .B(n20826), .ZN(
        P1_U3158) );
  OAI22_X1 U23735 ( .A1(n20832), .A2(n20831), .B1(n20830), .B2(n20829), .ZN(
        n20833) );
  INV_X1 U23736 ( .A(n20833), .ZN(n20836) );
  AOI22_X1 U23737 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20844), .B1(
        n20843), .B2(n20834), .ZN(n20835) );
  OAI211_X1 U23738 ( .C1(n20837), .C2(n20847), .A(n20836), .B(n20835), .ZN(
        P1_U3159) );
  AOI22_X1 U23739 ( .A1(n20841), .A2(n20840), .B1(n20839), .B2(n20838), .ZN(
        n20846) );
  AOI22_X1 U23740 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20844), .B1(
        n20843), .B2(n20842), .ZN(n20845) );
  OAI211_X1 U23741 ( .C1(n20848), .C2(n20847), .A(n20846), .B(n20845), .ZN(
        P1_U3160) );
  NOR2_X1 U23742 ( .A1(n20932), .A2(n20849), .ZN(n20852) );
  INV_X1 U23743 ( .A(n20850), .ZN(n20851) );
  OAI21_X1 U23744 ( .B1(n20852), .B2(n20929), .A(n20851), .ZN(P1_U3163) );
  INV_X1 U23745 ( .A(n20912), .ZN(n20853) );
  AND2_X1 U23746 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20853), .ZN(
        P1_U3164) );
  AND2_X1 U23747 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20853), .ZN(
        P1_U3165) );
  AND2_X1 U23748 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20853), .ZN(
        P1_U3166) );
  AND2_X1 U23749 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20853), .ZN(
        P1_U3167) );
  AND2_X1 U23750 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20853), .ZN(
        P1_U3168) );
  AND2_X1 U23751 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20853), .ZN(
        P1_U3169) );
  AND2_X1 U23752 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20853), .ZN(
        P1_U3170) );
  AND2_X1 U23753 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20853), .ZN(
        P1_U3171) );
  AND2_X1 U23754 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20853), .ZN(
        P1_U3172) );
  AND2_X1 U23755 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20853), .ZN(
        P1_U3173) );
  AND2_X1 U23756 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20853), .ZN(
        P1_U3174) );
  AND2_X1 U23757 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20853), .ZN(
        P1_U3175) );
  AND2_X1 U23758 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20853), .ZN(
        P1_U3176) );
  AND2_X1 U23759 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20853), .ZN(
        P1_U3177) );
  AND2_X1 U23760 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20853), .ZN(
        P1_U3178) );
  AND2_X1 U23761 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20853), .ZN(
        P1_U3179) );
  AND2_X1 U23762 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20853), .ZN(
        P1_U3180) );
  AND2_X1 U23763 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20853), .ZN(
        P1_U3181) );
  AND2_X1 U23764 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20853), .ZN(
        P1_U3182) );
  AND2_X1 U23765 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20853), .ZN(
        P1_U3183) );
  AND2_X1 U23766 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20853), .ZN(
        P1_U3184) );
  AND2_X1 U23767 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20853), .ZN(
        P1_U3185) );
  AND2_X1 U23768 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20853), .ZN(P1_U3186) );
  AND2_X1 U23769 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20853), .ZN(P1_U3187) );
  AND2_X1 U23770 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20853), .ZN(P1_U3188) );
  AND2_X1 U23771 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20853), .ZN(P1_U3189) );
  AND2_X1 U23772 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20853), .ZN(P1_U3190) );
  AND2_X1 U23773 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20853), .ZN(P1_U3191) );
  AND2_X1 U23774 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20853), .ZN(P1_U3192) );
  AND2_X1 U23775 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20853), .ZN(P1_U3193) );
  NAND2_X1 U23776 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20860), .ZN(n20863) );
  INV_X1 U23777 ( .A(n20863), .ZN(n20857) );
  OAI21_X1 U23778 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21254), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20854) );
  AOI211_X1 U23779 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20855), .B(
        n20854), .ZN(n20856) );
  OAI22_X1 U23780 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20857), .B1(n20939), 
        .B2(n20856), .ZN(P1_U3194) );
  AOI211_X1 U23781 ( .C1(n20859), .C2(n21254), .A(P1_STATE_REG_2__SCAN_IN), 
        .B(n20858), .ZN(n20866) );
  AOI21_X1 U23782 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20867), .A(n21248), .ZN(n20862) );
  INV_X1 U23783 ( .A(n20860), .ZN(n20861) );
  OAI221_X1 U23784 ( .B1(n20862), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20862), .C2(n20861), .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20865) );
  OAI211_X1 U23785 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21254), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20863), .ZN(n20864) );
  OAI21_X1 U23786 ( .B1(n20866), .B2(n20865), .A(n20864), .ZN(P1_U3196) );
  OR2_X1 U23787 ( .A1(n20927), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20895) );
  NOR2_X1 U23788 ( .A1(n20867), .A2(n20927), .ZN(n20903) );
  INV_X1 U23789 ( .A(n20903), .ZN(n20892) );
  INV_X1 U23790 ( .A(n20892), .ZN(n20901) );
  AOI222_X1 U23791 ( .A1(n9829), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20901), .ZN(n20868) );
  INV_X1 U23792 ( .A(n20868), .ZN(P1_U3197) );
  AOI222_X1 U23793 ( .A1(n20901), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n9829), .ZN(n20869) );
  INV_X1 U23794 ( .A(n20869), .ZN(P1_U3198) );
  OAI222_X1 U23795 ( .A1(n20895), .A2(n21228), .B1(n20871), .B2(n20939), .C1(
        n20870), .C2(n20892), .ZN(P1_U3199) );
  AOI222_X1 U23796 ( .A1(n9829), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20901), .ZN(n20872) );
  INV_X1 U23797 ( .A(n20872), .ZN(P1_U3200) );
  AOI222_X1 U23798 ( .A1(n20901), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n9829), .ZN(n20873) );
  INV_X1 U23799 ( .A(n20873), .ZN(P1_U3201) );
  AOI222_X1 U23800 ( .A1(n20901), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n9829), .ZN(n20874) );
  INV_X1 U23801 ( .A(n20874), .ZN(P1_U3202) );
  AOI222_X1 U23802 ( .A1(n20901), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n9829), .ZN(n20875) );
  INV_X1 U23803 ( .A(n20875), .ZN(P1_U3203) );
  AOI222_X1 U23804 ( .A1(n20901), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n9829), .ZN(n20876) );
  INV_X1 U23805 ( .A(n20876), .ZN(P1_U3204) );
  AOI222_X1 U23806 ( .A1(n20901), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n9829), .ZN(n20877) );
  INV_X1 U23807 ( .A(n20877), .ZN(P1_U3205) );
  INV_X1 U23808 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21226) );
  AOI22_X1 U23809 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20927), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n9829), .ZN(n20878) );
  OAI21_X1 U23810 ( .B1(n21226), .B2(n20892), .A(n20878), .ZN(P1_U3206) );
  INV_X1 U23811 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21050) );
  AOI22_X1 U23812 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20927), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20901), .ZN(n20879) );
  OAI21_X1 U23813 ( .B1(n21050), .B2(n20895), .A(n20879), .ZN(P1_U3207) );
  AOI222_X1 U23814 ( .A1(n20901), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n9829), .ZN(n20880) );
  INV_X1 U23815 ( .A(n20880), .ZN(P1_U3208) );
  AOI22_X1 U23816 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20927), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n9829), .ZN(n20881) );
  OAI21_X1 U23817 ( .B1(n20882), .B2(n20892), .A(n20881), .ZN(P1_U3209) );
  AOI22_X1 U23818 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20927), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20903), .ZN(n20883) );
  OAI21_X1 U23819 ( .B1(n21225), .B2(n20895), .A(n20883), .ZN(P1_U3210) );
  AOI222_X1 U23820 ( .A1(n9829), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20901), .ZN(n20884) );
  INV_X1 U23821 ( .A(n20884), .ZN(P1_U3211) );
  AOI222_X1 U23822 ( .A1(n20903), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n9829), .ZN(n20885) );
  INV_X1 U23823 ( .A(n20885), .ZN(P1_U3212) );
  AOI222_X1 U23824 ( .A1(n9829), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20901), .ZN(n20886) );
  INV_X1 U23825 ( .A(n20886), .ZN(P1_U3213) );
  AOI222_X1 U23826 ( .A1(n9829), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20901), .ZN(n20887) );
  INV_X1 U23827 ( .A(n20887), .ZN(P1_U3214) );
  AOI222_X1 U23828 ( .A1(n20903), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n9829), .ZN(n20888) );
  INV_X1 U23829 ( .A(n20888), .ZN(P1_U3215) );
  AOI222_X1 U23830 ( .A1(n20903), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n9829), .ZN(n20889) );
  INV_X1 U23831 ( .A(n20889), .ZN(P1_U3216) );
  AOI222_X1 U23832 ( .A1(n9829), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20901), .ZN(n20890) );
  INV_X1 U23833 ( .A(n20890), .ZN(P1_U3217) );
  AOI22_X1 U23834 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20927), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n9829), .ZN(n20891) );
  OAI21_X1 U23835 ( .B1(n20893), .B2(n20892), .A(n20891), .ZN(P1_U3218) );
  AOI22_X1 U23836 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20927), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20903), .ZN(n20894) );
  OAI21_X1 U23837 ( .B1(n21232), .B2(n20895), .A(n20894), .ZN(P1_U3219) );
  AOI222_X1 U23838 ( .A1(n20903), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n9829), .ZN(n20896) );
  INV_X1 U23839 ( .A(n20896), .ZN(P1_U3220) );
  AOI222_X1 U23840 ( .A1(n20903), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n9829), .ZN(n20897) );
  INV_X1 U23841 ( .A(n20897), .ZN(P1_U3221) );
  AOI222_X1 U23842 ( .A1(n20903), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n9829), .ZN(n20898) );
  INV_X1 U23843 ( .A(n20898), .ZN(P1_U3222) );
  AOI222_X1 U23844 ( .A1(n20901), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n9829), .ZN(n20899) );
  INV_X1 U23845 ( .A(n20899), .ZN(P1_U3223) );
  AOI222_X1 U23846 ( .A1(n20901), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n9829), .ZN(n20900) );
  INV_X1 U23847 ( .A(n20900), .ZN(P1_U3224) );
  AOI222_X1 U23848 ( .A1(n9829), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20901), .ZN(n20902) );
  INV_X1 U23849 ( .A(n20902), .ZN(P1_U3225) );
  AOI222_X1 U23850 ( .A1(n20903), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20927), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n9829), .ZN(n20904) );
  INV_X1 U23851 ( .A(n20904), .ZN(P1_U3226) );
  OAI22_X1 U23852 ( .A1(n20927), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20939), .ZN(n20905) );
  INV_X1 U23853 ( .A(n20905), .ZN(P1_U3458) );
  OAI22_X1 U23854 ( .A1(n20927), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20939), .ZN(n20906) );
  INV_X1 U23855 ( .A(n20906), .ZN(P1_U3459) );
  OAI22_X1 U23856 ( .A1(n20927), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20939), .ZN(n20907) );
  INV_X1 U23857 ( .A(n20907), .ZN(P1_U3460) );
  OAI22_X1 U23858 ( .A1(n20927), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20939), .ZN(n20908) );
  INV_X1 U23859 ( .A(n20908), .ZN(P1_U3461) );
  OAI21_X1 U23860 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20912), .A(n20910), 
        .ZN(n20909) );
  INV_X1 U23861 ( .A(n20909), .ZN(P1_U3464) );
  OAI21_X1 U23862 ( .B1(n20912), .B2(n20911), .A(n20910), .ZN(P1_U3465) );
  INV_X1 U23863 ( .A(n20913), .ZN(n20917) );
  OAI22_X1 U23864 ( .A1(n20917), .A2(n20916), .B1(n20915), .B2(n20914), .ZN(
        n20920) );
  MUX2_X1 U23865 ( .A(n20920), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20918), .Z(P1_U3469) );
  AOI21_X1 U23866 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20921) );
  AOI22_X1 U23867 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20921), .B2(n13685), .ZN(n20922) );
  INV_X1 U23868 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21070) );
  AOI22_X1 U23869 ( .A1(n20923), .A2(n20922), .B1(n21070), .B2(n20925), .ZN(
        P1_U3481) );
  INV_X1 U23870 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20926) );
  INV_X1 U23871 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21087) );
  NOR2_X1 U23872 ( .A1(n20925), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20924) );
  AOI22_X1 U23873 ( .A1(n20926), .A2(n20925), .B1(n21087), .B2(n20924), .ZN(
        P1_U3482) );
  AOI22_X1 U23874 ( .A1(n20939), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21261), 
        .B2(n20927), .ZN(P1_U3483) );
  AOI211_X1 U23875 ( .C1(n20930), .C2(n21085), .A(n20929), .B(n20928), .ZN(
        n20933) );
  OAI21_X1 U23876 ( .B1(n20933), .B2(n20932), .A(n20931), .ZN(n20938) );
  AOI211_X1 U23877 ( .C1(n20164), .C2(n20936), .A(n20935), .B(n20934), .ZN(
        n20937) );
  MUX2_X1 U23878 ( .A(n20938), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20937), 
        .Z(P1_U3485) );
  OAI22_X1 U23879 ( .A1(n20927), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20939), .ZN(n20940) );
  INV_X1 U23880 ( .A(n20940), .ZN(P1_U3486) );
  OAI22_X1 U23881 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(keyinput_g109), .B1(
        keyinput_g12), .B2(DATAI_20_), .ZN(n20941) );
  AOI221_X1 U23882 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(keyinput_g109), .C1(
        DATAI_20_), .C2(keyinput_g12), .A(n20941), .ZN(n20948) );
  OAI22_X1 U23883 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g49), .B1(
        keyinput_g33), .B2(HOLD), .ZN(n20942) );
  AOI221_X1 U23884 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g49), 
        .C1(HOLD), .C2(keyinput_g33), .A(n20942), .ZN(n20947) );
  OAI22_X1 U23885 ( .A1(P1_EBX_REG_0__SCAN_IN), .A2(keyinput_g115), .B1(
        DATAI_25_), .B2(keyinput_g7), .ZN(n20943) );
  AOI221_X1 U23886 ( .B1(P1_EBX_REG_0__SCAN_IN), .B2(keyinput_g115), .C1(
        keyinput_g7), .C2(DATAI_25_), .A(n20943), .ZN(n20946) );
  OAI22_X1 U23887 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(keyinput_g110), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(keyinput_g80), .ZN(n20944) );
  AOI221_X1 U23888 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(keyinput_g110), .C1(
        keyinput_g80), .C2(P1_REIP_REG_3__SCAN_IN), .A(n20944), .ZN(n20945) );
  NAND4_X1 U23889 ( .A1(n20948), .A2(n20947), .A3(n20946), .A4(n20945), .ZN(
        n20976) );
  OAI22_X1 U23890 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(keyinput_g64), .B1(
        keyinput_g18), .B2(DATAI_14_), .ZN(n20949) );
  AOI221_X1 U23891 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(keyinput_g64), .C1(
        DATAI_14_), .C2(keyinput_g18), .A(n20949), .ZN(n20956) );
  OAI22_X1 U23892 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(keyinput_g112), .B1(
        DATAI_6_), .B2(keyinput_g26), .ZN(n20950) );
  AOI221_X1 U23893 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(keyinput_g112), .C1(
        keyinput_g26), .C2(DATAI_6_), .A(n20950), .ZN(n20955) );
  OAI22_X1 U23894 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_g123), .B1(
        keyinput_g38), .B2(P1_READREQUEST_REG_SCAN_IN), .ZN(n20951) );
  AOI221_X1 U23895 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_g123), .C1(
        P1_READREQUEST_REG_SCAN_IN), .C2(keyinput_g38), .A(n20951), .ZN(n20954) );
  OAI22_X1 U23896 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_g88), .B1(
        keyinput_g78), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n20952) );
  AOI221_X1 U23897 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput_g88), .C1(
        P1_REIP_REG_5__SCAN_IN), .C2(keyinput_g78), .A(n20952), .ZN(n20953) );
  NAND4_X1 U23898 ( .A1(n20956), .A2(n20955), .A3(n20954), .A4(n20953), .ZN(
        n20975) );
  OAI22_X1 U23899 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_g60), .B1(
        keyinput_g43), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20957) );
  AOI221_X1 U23900 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .C1(
        P1_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_g43), .A(n20957), .ZN(
        n20964) );
  OAI22_X1 U23901 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(keyinput_g74), .B1(
        keyinput_g69), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n20958) );
  AOI221_X1 U23902 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(keyinput_g74), .C1(
        P1_REIP_REG_14__SCAN_IN), .C2(keyinput_g69), .A(n20958), .ZN(n20963)
         );
  OAI22_X1 U23903 ( .A1(P1_EAX_REG_27__SCAN_IN), .A2(keyinput_g120), .B1(
        keyinput_g58), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n20959) );
  AOI221_X1 U23904 ( .B1(P1_EAX_REG_27__SCAN_IN), .B2(keyinput_g120), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_g58), .A(n20959), .ZN(n20962)
         );
  OAI22_X1 U23905 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(keyinput_g100), .B1(
        DATAI_28_), .B2(keyinput_g4), .ZN(n20960) );
  AOI221_X1 U23906 ( .B1(P1_EBX_REG_15__SCAN_IN), .B2(keyinput_g100), .C1(
        keyinput_g4), .C2(DATAI_28_), .A(n20960), .ZN(n20961) );
  NAND4_X1 U23907 ( .A1(n20964), .A2(n20963), .A3(n20962), .A4(n20961), .ZN(
        n20974) );
  OAI22_X1 U23908 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(keyinput_g68), .B1(
        keyinput_g0), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20965) );
  AOI221_X1 U23909 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(keyinput_g68), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_g0), .A(n20965), .ZN(n20972)
         );
  OAI22_X1 U23910 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(keyinput_g94), .B1(
        DATAI_5_), .B2(keyinput_g27), .ZN(n20966) );
  AOI221_X1 U23911 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(keyinput_g94), .C1(
        keyinput_g27), .C2(DATAI_5_), .A(n20966), .ZN(n20971) );
  OAI22_X1 U23912 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput_g61), .B1(
        keyinput_g25), .B2(DATAI_7_), .ZN(n20967) );
  AOI221_X1 U23913 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_g61), .C1(
        DATAI_7_), .C2(keyinput_g25), .A(n20967), .ZN(n20970) );
  OAI22_X1 U23914 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(keyinput_g103), .B1(
        P1_EBX_REG_11__SCAN_IN), .B2(keyinput_g104), .ZN(n20968) );
  AOI221_X1 U23915 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(keyinput_g103), .C1(
        keyinput_g104), .C2(P1_EBX_REG_11__SCAN_IN), .A(n20968), .ZN(n20969)
         );
  NAND4_X1 U23916 ( .A1(n20972), .A2(n20971), .A3(n20970), .A4(n20969), .ZN(
        n20973) );
  NOR4_X1 U23917 ( .A1(n20976), .A2(n20975), .A3(n20974), .A4(n20973), .ZN(
        n21319) );
  OAI22_X1 U23918 ( .A1(P1_EAX_REG_30__SCAN_IN), .A2(keyinput_g117), .B1(
        keyinput_g48), .B2(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20977) );
  AOI221_X1 U23919 ( .B1(P1_EAX_REG_30__SCAN_IN), .B2(keyinput_g117), .C1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_g48), .A(n20977), .ZN(
        n20984) );
  OAI22_X1 U23920 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(keyinput_g72), .B1(
        keyinput_g5), .B2(DATAI_27_), .ZN(n20978) );
  AOI221_X1 U23921 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(keyinput_g72), .C1(
        DATAI_27_), .C2(keyinput_g5), .A(n20978), .ZN(n20983) );
  OAI22_X1 U23922 ( .A1(DATAI_11_), .A2(keyinput_g21), .B1(
        P1_FLUSH_REG_SCAN_IN), .B2(keyinput_g46), .ZN(n20979) );
  AOI221_X1 U23923 ( .B1(DATAI_11_), .B2(keyinput_g21), .C1(keyinput_g46), 
        .C2(P1_FLUSH_REG_SCAN_IN), .A(n20979), .ZN(n20982) );
  OAI22_X1 U23924 ( .A1(P1_EBX_REG_24__SCAN_IN), .A2(keyinput_g91), .B1(
        P1_EBX_REG_13__SCAN_IN), .B2(keyinput_g102), .ZN(n20980) );
  AOI221_X1 U23925 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(keyinput_g91), .C1(
        keyinput_g102), .C2(P1_EBX_REG_13__SCAN_IN), .A(n20980), .ZN(n20981)
         );
  NAND4_X1 U23926 ( .A1(n20984), .A2(n20983), .A3(n20982), .A4(n20981), .ZN(
        n21113) );
  OAI22_X1 U23927 ( .A1(P1_EAX_REG_23__SCAN_IN), .A2(keyinput_g124), .B1(
        keyinput_g54), .B2(P1_REIP_REG_29__SCAN_IN), .ZN(n20985) );
  AOI221_X1 U23928 ( .B1(P1_EAX_REG_23__SCAN_IN), .B2(keyinput_g124), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_g54), .A(n20985), .ZN(n21010)
         );
  OAI22_X1 U23929 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g51), .ZN(n20986) );
  AOI221_X1 U23930 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        keyinput_g51), .C2(P1_BYTEENABLE_REG_3__SCAN_IN), .A(n20986), .ZN(
        n20989) );
  OAI22_X1 U23931 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(keyinput_g79), .B1(NA), 
        .B2(keyinput_g34), .ZN(n20987) );
  AOI221_X1 U23932 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(keyinput_g79), .C1(
        keyinput_g34), .C2(NA), .A(n20987), .ZN(n20988) );
  OAI211_X1 U23933 ( .C1(n21252), .C2(keyinput_g106), .A(n20989), .B(n20988), 
        .ZN(n20990) );
  AOI21_X1 U23934 ( .B1(n21252), .B2(keyinput_g106), .A(n20990), .ZN(n21009)
         );
  AOI22_X1 U23935 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_g45), .B1(DATAI_8_), 
        .B2(keyinput_g24), .ZN(n20991) );
  OAI221_X1 U23936 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_g45), .C1(DATAI_8_), .C2(keyinput_g24), .A(n20991), .ZN(n20998) );
  AOI22_X1 U23937 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput_g75), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(keyinput_g125), .ZN(n20992) );
  OAI221_X1 U23938 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput_g75), .C1(
        P1_EAX_REG_22__SCAN_IN), .C2(keyinput_g125), .A(n20992), .ZN(n20997)
         );
  AOI22_X1 U23939 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .ZN(n20993) );
  OAI221_X1 U23940 ( .B1(P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_g59), .A(n20993), .ZN(n20996)
         );
  AOI22_X1 U23941 ( .A1(DATAI_2_), .A2(keyinput_g30), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_g56), .ZN(n20994) );
  OAI221_X1 U23942 ( .B1(DATAI_2_), .B2(keyinput_g30), .C1(
        P1_REIP_REG_27__SCAN_IN), .C2(keyinput_g56), .A(n20994), .ZN(n20995)
         );
  NOR4_X1 U23943 ( .A1(n20998), .A2(n20997), .A3(n20996), .A4(n20995), .ZN(
        n21008) );
  AOI22_X1 U23944 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_g65), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(keyinput_g86), .ZN(n20999) );
  OAI221_X1 U23945 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(keyinput_g65), .C1(
        P1_EBX_REG_29__SCAN_IN), .C2(keyinput_g86), .A(n20999), .ZN(n21006) );
  AOI22_X1 U23946 ( .A1(DATAI_21_), .A2(keyinput_g11), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(keyinput_g70), .ZN(n21000) );
  OAI221_X1 U23947 ( .B1(DATAI_21_), .B2(keyinput_g11), .C1(
        P1_REIP_REG_13__SCAN_IN), .C2(keyinput_g70), .A(n21000), .ZN(n21005)
         );
  AOI22_X1 U23948 ( .A1(DATAI_30_), .A2(keyinput_g2), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(keyinput_g127), .ZN(n21001) );
  OAI221_X1 U23949 ( .B1(DATAI_30_), .B2(keyinput_g2), .C1(
        P1_EAX_REG_20__SCAN_IN), .C2(keyinput_g127), .A(n21001), .ZN(n21004)
         );
  AOI22_X1 U23950 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_g63), .B1(
        P1_EBX_REG_16__SCAN_IN), .B2(keyinput_g99), .ZN(n21002) );
  OAI221_X1 U23951 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .C1(
        P1_EBX_REG_16__SCAN_IN), .C2(keyinput_g99), .A(n21002), .ZN(n21003) );
  NOR4_X1 U23952 ( .A1(n21006), .A2(n21005), .A3(n21004), .A4(n21003), .ZN(
        n21007) );
  NAND4_X1 U23953 ( .A1(n21010), .A2(n21009), .A3(n21008), .A4(n21007), .ZN(
        n21112) );
  AOI22_X1 U23954 ( .A1(DATAI_15_), .A2(keyinput_g17), .B1(
        P1_EBX_REG_7__SCAN_IN), .B2(keyinput_g108), .ZN(n21011) );
  OAI221_X1 U23955 ( .B1(DATAI_15_), .B2(keyinput_g17), .C1(
        P1_EBX_REG_7__SCAN_IN), .C2(keyinput_g108), .A(n21011), .ZN(n21019) );
  AOI22_X1 U23956 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(keyinput_g82), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(keyinput_g85), .ZN(n21012) );
  OAI221_X1 U23957 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(keyinput_g82), .C1(
        P1_EBX_REG_30__SCAN_IN), .C2(keyinput_g85), .A(n21012), .ZN(n21018) );
  AOI22_X1 U23958 ( .A1(n21014), .A2(keyinput_g10), .B1(n14932), .B2(
        keyinput_g8), .ZN(n21013) );
  OAI221_X1 U23959 ( .B1(n21014), .B2(keyinput_g10), .C1(n14932), .C2(
        keyinput_g8), .A(n21013), .ZN(n21017) );
  INV_X1 U23960 ( .A(DATAI_0_), .ZN(n21290) );
  AOI22_X1 U23961 ( .A1(n21267), .A2(keyinput_g111), .B1(keyinput_g32), .B2(
        n21290), .ZN(n21015) );
  OAI221_X1 U23962 ( .B1(n21267), .B2(keyinput_g111), .C1(n21290), .C2(
        keyinput_g32), .A(n21015), .ZN(n21016) );
  NOR4_X1 U23963 ( .A1(n21019), .A2(n21018), .A3(n21017), .A4(n21016), .ZN(
        n21058) );
  INV_X1 U23964 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21292) );
  AOI22_X1 U23965 ( .A1(n14851), .A2(keyinput_g93), .B1(keyinput_g76), .B2(
        n21292), .ZN(n21020) );
  OAI221_X1 U23966 ( .B1(n14851), .B2(keyinput_g93), .C1(n21292), .C2(
        keyinput_g76), .A(n21020), .ZN(n21030) );
  INV_X1 U23967 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21231) );
  INV_X1 U23968 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n21196) );
  AOI22_X1 U23969 ( .A1(n21231), .A2(keyinput_g62), .B1(n21196), .B2(
        keyinput_g96), .ZN(n21021) );
  OAI221_X1 U23970 ( .B1(n21231), .B2(keyinput_g62), .C1(n21196), .C2(
        keyinput_g96), .A(n21021), .ZN(n21029) );
  AOI22_X1 U23971 ( .A1(n21024), .A2(keyinput_g14), .B1(n21023), .B2(
        keyinput_g90), .ZN(n21022) );
  OAI221_X1 U23972 ( .B1(n21024), .B2(keyinput_g14), .C1(n21023), .C2(
        keyinput_g90), .A(n21022), .ZN(n21028) );
  INV_X1 U23973 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n21026) );
  AOI22_X1 U23974 ( .A1(n21026), .A2(keyinput_g116), .B1(keyinput_g97), .B2(
        n21289), .ZN(n21025) );
  OAI221_X1 U23975 ( .B1(n21026), .B2(keyinput_g116), .C1(n21289), .C2(
        keyinput_g97), .A(n21025), .ZN(n21027) );
  NOR4_X1 U23976 ( .A1(n21030), .A2(n21029), .A3(n21028), .A4(n21027), .ZN(
        n21057) );
  INV_X1 U23977 ( .A(DATAI_4_), .ZN(n21033) );
  AOI22_X1 U23978 ( .A1(n21033), .A2(keyinput_g28), .B1(n21032), .B2(
        keyinput_g119), .ZN(n21031) );
  OAI221_X1 U23979 ( .B1(n21033), .B2(keyinput_g28), .C1(n21032), .C2(
        keyinput_g119), .A(n21031), .ZN(n21042) );
  INV_X1 U23980 ( .A(DATAI_3_), .ZN(n21277) );
  AOI22_X1 U23981 ( .A1(n21277), .A2(keyinput_g29), .B1(n13954), .B2(
        keyinput_g113), .ZN(n21034) );
  OAI221_X1 U23982 ( .B1(n21277), .B2(keyinput_g29), .C1(n13954), .C2(
        keyinput_g113), .A(n21034), .ZN(n21041) );
  INV_X1 U23983 ( .A(DATAI_1_), .ZN(n21036) );
  AOI22_X1 U23984 ( .A1(n21036), .A2(keyinput_g31), .B1(n21234), .B2(
        keyinput_g121), .ZN(n21035) );
  OAI221_X1 U23985 ( .B1(n21036), .B2(keyinput_g31), .C1(n21234), .C2(
        keyinput_g121), .A(n21035), .ZN(n21040) );
  INV_X1 U23986 ( .A(DATAI_10_), .ZN(n21235) );
  AOI22_X1 U23987 ( .A1(n21038), .A2(keyinput_g89), .B1(keyinput_g22), .B2(
        n21235), .ZN(n21037) );
  OAI221_X1 U23988 ( .B1(n21038), .B2(keyinput_g89), .C1(n21235), .C2(
        keyinput_g22), .A(n21037), .ZN(n21039) );
  NOR4_X1 U23989 ( .A1(n21042), .A2(n21041), .A3(n21040), .A4(n21039), .ZN(
        n21056) );
  AOI22_X1 U23990 ( .A1(n21226), .A2(keyinput_g73), .B1(n21044), .B2(
        keyinput_g126), .ZN(n21043) );
  OAI221_X1 U23991 ( .B1(n21226), .B2(keyinput_g73), .C1(n21044), .C2(
        keyinput_g126), .A(n21043), .ZN(n21054) );
  INV_X1 U23992 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21213) );
  AOI22_X1 U23993 ( .A1(n21046), .A2(keyinput_g118), .B1(keyinput_g53), .B2(
        n21213), .ZN(n21045) );
  OAI221_X1 U23994 ( .B1(n21046), .B2(keyinput_g118), .C1(n21213), .C2(
        keyinput_g53), .A(n21045), .ZN(n21053) );
  INV_X1 U23995 ( .A(DATAI_26_), .ZN(n21279) );
  INV_X1 U23996 ( .A(DATAI_12_), .ZN(n21280) );
  AOI22_X1 U23997 ( .A1(n21279), .A2(keyinput_g6), .B1(n21280), .B2(
        keyinput_g20), .ZN(n21047) );
  OAI221_X1 U23998 ( .B1(n21279), .B2(keyinput_g6), .C1(n21280), .C2(
        keyinput_g20), .A(n21047), .ZN(n21052) );
  INV_X1 U23999 ( .A(READY1), .ZN(n21049) );
  AOI22_X1 U24000 ( .A1(n21050), .A2(keyinput_g71), .B1(n21049), .B2(
        keyinput_g36), .ZN(n21048) );
  OAI221_X1 U24001 ( .B1(n21050), .B2(keyinput_g71), .C1(n21049), .C2(
        keyinput_g36), .A(n21048), .ZN(n21051) );
  NOR4_X1 U24002 ( .A1(n21054), .A2(n21053), .A3(n21052), .A4(n21051), .ZN(
        n21055) );
  NAND4_X1 U24003 ( .A1(n21058), .A2(n21057), .A3(n21056), .A4(n21055), .ZN(
        n21111) );
  AOI22_X1 U24004 ( .A1(n21190), .A2(keyinput_g39), .B1(n14835), .B2(
        keyinput_g107), .ZN(n21059) );
  OAI221_X1 U24005 ( .B1(n21190), .B2(keyinput_g39), .C1(n14835), .C2(
        keyinput_g107), .A(n21059), .ZN(n21068) );
  AOI22_X1 U24006 ( .A1(n21204), .A2(keyinput_g105), .B1(keyinput_g16), .B2(
        n21265), .ZN(n21060) );
  OAI221_X1 U24007 ( .B1(n21204), .B2(keyinput_g105), .C1(n21265), .C2(
        keyinput_g16), .A(n21060), .ZN(n21067) );
  AOI22_X1 U24008 ( .A1(n14996), .A2(keyinput_g55), .B1(n21283), .B2(
        keyinput_g98), .ZN(n21061) );
  OAI221_X1 U24009 ( .B1(n14996), .B2(keyinput_g55), .C1(n21283), .C2(
        keyinput_g98), .A(n21061), .ZN(n21066) );
  INV_X1 U24010 ( .A(DATAI_13_), .ZN(n21064) );
  INV_X1 U24011 ( .A(READY2), .ZN(n21063) );
  AOI22_X1 U24012 ( .A1(n21064), .A2(keyinput_g19), .B1(keyinput_g37), .B2(
        n21063), .ZN(n21062) );
  OAI221_X1 U24013 ( .B1(n21064), .B2(keyinput_g19), .C1(n21063), .C2(
        keyinput_g37), .A(n21062), .ZN(n21065) );
  NOR4_X1 U24014 ( .A1(n21068), .A2(n21067), .A3(n21066), .A4(n21065), .ZN(
        n21109) );
  INV_X1 U24015 ( .A(DATAI_9_), .ZN(n21282) );
  AOI22_X1 U24016 ( .A1(n21282), .A2(keyinput_g23), .B1(keyinput_g50), .B2(
        n21070), .ZN(n21069) );
  OAI221_X1 U24017 ( .B1(n21282), .B2(keyinput_g23), .C1(n21070), .C2(
        keyinput_g50), .A(n21069), .ZN(n21081) );
  AOI22_X1 U24018 ( .A1(n21073), .A2(keyinput_g66), .B1(keyinput_g15), .B2(
        n21072), .ZN(n21071) );
  OAI221_X1 U24019 ( .B1(n21073), .B2(keyinput_g66), .C1(n21072), .C2(
        keyinput_g15), .A(n21071), .ZN(n21080) );
  AOI22_X1 U24020 ( .A1(n21076), .A2(keyinput_g40), .B1(keyinput_g35), .B2(
        n21075), .ZN(n21074) );
  OAI221_X1 U24021 ( .B1(n21076), .B2(keyinput_g40), .C1(n21075), .C2(
        keyinput_g35), .A(n21074), .ZN(n21079) );
  AOI22_X1 U24022 ( .A1(n21216), .A2(keyinput_g92), .B1(n21294), .B2(
        keyinput_g87), .ZN(n21077) );
  OAI221_X1 U24023 ( .B1(n21216), .B2(keyinput_g92), .C1(n21294), .C2(
        keyinput_g87), .A(n21077), .ZN(n21078) );
  NOR4_X1 U24024 ( .A1(n21081), .A2(n21080), .A3(n21079), .A4(n21078), .ZN(
        n21108) );
  AOI22_X1 U24025 ( .A1(n21083), .A2(keyinput_g52), .B1(keyinput_g101), .B2(
        n21255), .ZN(n21082) );
  OAI221_X1 U24026 ( .B1(n21083), .B2(keyinput_g52), .C1(n21255), .C2(
        keyinput_g101), .A(n21082), .ZN(n21093) );
  AOI22_X1 U24027 ( .A1(n14644), .A2(keyinput_g84), .B1(n21085), .B2(
        keyinput_g44), .ZN(n21084) );
  OAI221_X1 U24028 ( .B1(n14644), .B2(keyinput_g84), .C1(n21085), .C2(
        keyinput_g44), .A(n21084), .ZN(n21092) );
  AOI22_X1 U24029 ( .A1(n21087), .A2(keyinput_g83), .B1(n21251), .B2(
        keyinput_g13), .ZN(n21086) );
  OAI221_X1 U24030 ( .B1(n21087), .B2(keyinput_g83), .C1(n21251), .C2(
        keyinput_g13), .A(n21086), .ZN(n21091) );
  AOI22_X1 U24031 ( .A1(n21089), .A2(keyinput_g9), .B1(n21264), .B2(
        keyinput_g122), .ZN(n21088) );
  OAI221_X1 U24032 ( .B1(n21089), .B2(keyinput_g9), .C1(n21264), .C2(
        keyinput_g122), .A(n21088), .ZN(n21090) );
  NOR4_X1 U24033 ( .A1(n21093), .A2(n21092), .A3(n21091), .A4(n21090), .ZN(
        n21107) );
  AOI22_X1 U24034 ( .A1(n21261), .A2(keyinput_g47), .B1(n21095), .B2(
        keyinput_g77), .ZN(n21094) );
  OAI221_X1 U24035 ( .B1(n21261), .B2(keyinput_g47), .C1(n21095), .C2(
        keyinput_g77), .A(n21094), .ZN(n21105) );
  INV_X1 U24036 ( .A(DATAI_31_), .ZN(n21097) );
  AOI22_X1 U24037 ( .A1(n21097), .A2(keyinput_g1), .B1(n21215), .B2(
        keyinput_g95), .ZN(n21096) );
  OAI221_X1 U24038 ( .B1(n21097), .B2(keyinput_g1), .C1(n21215), .C2(
        keyinput_g95), .A(n21096), .ZN(n21104) );
  AOI22_X1 U24039 ( .A1(n21099), .A2(keyinput_g114), .B1(keyinput_g67), .B2(
        n15098), .ZN(n21098) );
  OAI221_X1 U24040 ( .B1(n21099), .B2(keyinput_g114), .C1(n15098), .C2(
        keyinput_g67), .A(n21098), .ZN(n21103) );
  INV_X1 U24041 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21101) );
  AOI22_X1 U24042 ( .A1(n21101), .A2(keyinput_g57), .B1(keyinput_g3), .B2(
        n14909), .ZN(n21100) );
  OAI221_X1 U24043 ( .B1(n21101), .B2(keyinput_g57), .C1(n14909), .C2(
        keyinput_g3), .A(n21100), .ZN(n21102) );
  NOR4_X1 U24044 ( .A1(n21105), .A2(n21104), .A3(n21103), .A4(n21102), .ZN(
        n21106) );
  NAND4_X1 U24045 ( .A1(n21109), .A2(n21108), .A3(n21107), .A4(n21106), .ZN(
        n21110) );
  NOR4_X1 U24046 ( .A1(n21113), .A2(n21112), .A3(n21111), .A4(n21110), .ZN(
        n21318) );
  AOI22_X1 U24047 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(keyinput_f126), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n21114) );
  OAI221_X1 U24048 ( .B1(P1_EAX_REG_21__SCAN_IN), .B2(keyinput_f126), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_f44), .A(n21114), .ZN(n21121)
         );
  AOI22_X1 U24049 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_f60), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(keyinput_f127), .ZN(n21115) );
  OAI221_X1 U24050 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_f60), .C1(
        P1_EAX_REG_20__SCAN_IN), .C2(keyinput_f127), .A(n21115), .ZN(n21120)
         );
  AOI22_X1 U24051 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(keyinput_f66), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(keyinput_f57), .ZN(n21116) );
  OAI221_X1 U24052 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(keyinput_f66), .C1(
        P1_REIP_REG_26__SCAN_IN), .C2(keyinput_f57), .A(n21116), .ZN(n21119)
         );
  AOI22_X1 U24053 ( .A1(keyinput_f42), .A2(P1_D_C_N_REG_SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(keyinput_f119), .ZN(n21117) );
  OAI221_X1 U24054 ( .B1(keyinput_f42), .B2(P1_D_C_N_REG_SCAN_IN), .C1(
        P1_EAX_REG_28__SCAN_IN), .C2(keyinput_f119), .A(n21117), .ZN(n21118)
         );
  NOR4_X1 U24055 ( .A1(n21121), .A2(n21120), .A3(n21119), .A4(n21118), .ZN(
        n21312) );
  AOI22_X1 U24056 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(keyinput_f72), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput_f118), .ZN(n21122) );
  OAI221_X1 U24057 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(keyinput_f72), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput_f118), .A(n21122), .ZN(n21148)
         );
  OAI22_X1 U24058 ( .A1(DATAI_7_), .A2(keyinput_f25), .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_f46), .ZN(n21123) );
  AOI221_X1 U24059 ( .B1(DATAI_7_), .B2(keyinput_f25), .C1(keyinput_f46), .C2(
        P1_FLUSH_REG_SCAN_IN), .A(n21123), .ZN(n21127) );
  AOI22_X1 U24060 ( .A1(DATAI_4_), .A2(keyinput_f28), .B1(READY1), .B2(
        keyinput_f36), .ZN(n21124) );
  OAI221_X1 U24061 ( .B1(DATAI_4_), .B2(keyinput_f28), .C1(READY1), .C2(
        keyinput_f36), .A(n21124), .ZN(n21125) );
  AOI21_X1 U24062 ( .B1(keyinput_f58), .B2(n21128), .A(n21125), .ZN(n21126) );
  OAI211_X1 U24063 ( .C1(keyinput_f58), .C2(n21128), .A(n21127), .B(n21126), 
        .ZN(n21147) );
  OAI22_X1 U24064 ( .A1(P1_EAX_REG_23__SCAN_IN), .A2(keyinput_f124), .B1(
        keyinput_f80), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n21129) );
  AOI221_X1 U24065 ( .B1(P1_EAX_REG_23__SCAN_IN), .B2(keyinput_f124), .C1(
        P1_REIP_REG_3__SCAN_IN), .C2(keyinput_f80), .A(n21129), .ZN(n21136) );
  OAI22_X1 U24066 ( .A1(DATAI_31_), .A2(keyinput_f1), .B1(keyinput_f63), .B2(
        P1_REIP_REG_20__SCAN_IN), .ZN(n21130) );
  AOI221_X1 U24067 ( .B1(DATAI_31_), .B2(keyinput_f1), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_f63), .A(n21130), .ZN(n21135)
         );
  OAI22_X1 U24068 ( .A1(P1_EAX_REG_27__SCAN_IN), .A2(keyinput_f120), .B1(
        keyinput_f10), .B2(DATAI_22_), .ZN(n21131) );
  AOI221_X1 U24069 ( .B1(P1_EAX_REG_27__SCAN_IN), .B2(keyinput_f120), .C1(
        DATAI_22_), .C2(keyinput_f10), .A(n21131), .ZN(n21134) );
  OAI22_X1 U24070 ( .A1(P1_EBX_REG_30__SCAN_IN), .A2(keyinput_f85), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(keyinput_f71), .ZN(n21132) );
  AOI221_X1 U24071 ( .B1(P1_EBX_REG_30__SCAN_IN), .B2(keyinput_f85), .C1(
        keyinput_f71), .C2(P1_REIP_REG_12__SCAN_IN), .A(n21132), .ZN(n21133)
         );
  NAND4_X1 U24072 ( .A1(n21136), .A2(n21135), .A3(n21134), .A4(n21133), .ZN(
        n21146) );
  OAI22_X1 U24073 ( .A1(P1_EBX_REG_25__SCAN_IN), .A2(keyinput_f90), .B1(
        DATAI_29_), .B2(keyinput_f3), .ZN(n21137) );
  AOI221_X1 U24074 ( .B1(P1_EBX_REG_25__SCAN_IN), .B2(keyinput_f90), .C1(
        keyinput_f3), .C2(DATAI_29_), .A(n21137), .ZN(n21144) );
  OAI22_X1 U24075 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_f88), .B1(
        DATAI_27_), .B2(keyinput_f5), .ZN(n21138) );
  AOI221_X1 U24076 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput_f88), .C1(
        keyinput_f5), .C2(DATAI_27_), .A(n21138), .ZN(n21143) );
  OAI22_X1 U24077 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(keyinput_f112), .B1(
        keyinput_f69), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n21139) );
  AOI221_X1 U24078 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(keyinput_f112), .C1(
        P1_REIP_REG_14__SCAN_IN), .C2(keyinput_f69), .A(n21139), .ZN(n21142)
         );
  OAI22_X1 U24079 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(keyinput_f56), .B1(
        keyinput_f37), .B2(READY2), .ZN(n21140) );
  AOI221_X1 U24080 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(keyinput_f56), .C1(
        READY2), .C2(keyinput_f37), .A(n21140), .ZN(n21141) );
  NAND4_X1 U24081 ( .A1(n21144), .A2(n21143), .A3(n21142), .A4(n21141), .ZN(
        n21145) );
  NOR4_X1 U24082 ( .A1(n21148), .A2(n21147), .A3(n21146), .A4(n21145), .ZN(
        n21311) );
  OAI22_X1 U24083 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(keyinput_f114), .B1(
        DATAI_13_), .B2(keyinput_f19), .ZN(n21149) );
  AOI221_X1 U24084 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(keyinput_f114), .C1(
        keyinput_f19), .C2(DATAI_13_), .A(n21149), .ZN(n21156) );
  OAI22_X1 U24085 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(keyinput_f110), .B1(
        keyinput_f65), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n21150) );
  AOI221_X1 U24086 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(keyinput_f110), .C1(
        P1_REIP_REG_18__SCAN_IN), .C2(keyinput_f65), .A(n21150), .ZN(n21155)
         );
  OAI22_X1 U24087 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(keyinput_f100), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_f48), .ZN(n21151) );
  AOI221_X1 U24088 ( .B1(P1_EBX_REG_15__SCAN_IN), .B2(keyinput_f100), .C1(
        keyinput_f48), .C2(P1_BYTEENABLE_REG_0__SCAN_IN), .A(n21151), .ZN(
        n21154) );
  OAI22_X1 U24089 ( .A1(DATAI_24_), .A2(keyinput_f8), .B1(keyinput_f50), .B2(
        P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21152) );
  AOI221_X1 U24090 ( .B1(DATAI_24_), .B2(keyinput_f8), .C1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_f50), .A(n21152), .ZN(
        n21153) );
  NAND4_X1 U24091 ( .A1(n21156), .A2(n21155), .A3(n21154), .A4(n21153), .ZN(
        n21184) );
  OAI22_X1 U24092 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(keyinput_f52), .B1(
        P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f0), .ZN(n21157) );
  AOI221_X1 U24093 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(keyinput_f52), .C1(
        keyinput_f0), .C2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n21157), .ZN(n21164)
         );
  OAI22_X1 U24094 ( .A1(P1_EBX_REG_24__SCAN_IN), .A2(keyinput_f91), .B1(
        P1_EBX_REG_13__SCAN_IN), .B2(keyinput_f102), .ZN(n21158) );
  AOI221_X1 U24095 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(keyinput_f91), .C1(
        keyinput_f102), .C2(P1_EBX_REG_13__SCAN_IN), .A(n21158), .ZN(n21163)
         );
  OAI22_X1 U24096 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput_f61), .B1(
        P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f43), .ZN(n21159) );
  AOI221_X1 U24097 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_f61), .C1(
        keyinput_f43), .C2(P1_REQUESTPENDING_REG_SCAN_IN), .A(n21159), .ZN(
        n21162) );
  OAI22_X1 U24098 ( .A1(P1_EBX_REG_8__SCAN_IN), .A2(keyinput_f107), .B1(
        DATAI_23_), .B2(keyinput_f9), .ZN(n21160) );
  AOI221_X1 U24099 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(keyinput_f107), .C1(
        keyinput_f9), .C2(DATAI_23_), .A(n21160), .ZN(n21161) );
  NAND4_X1 U24100 ( .A1(n21164), .A2(n21163), .A3(n21162), .A4(n21161), .ZN(
        n21183) );
  OAI22_X1 U24101 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(keyinput_f83), .B1(BS16), 
        .B2(keyinput_f35), .ZN(n21165) );
  AOI221_X1 U24102 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(keyinput_f83), .C1(
        keyinput_f35), .C2(BS16), .A(n21165), .ZN(n21172) );
  OAI22_X1 U24103 ( .A1(DATAI_30_), .A2(keyinput_f2), .B1(keyinput_f11), .B2(
        DATAI_21_), .ZN(n21166) );
  AOI221_X1 U24104 ( .B1(DATAI_30_), .B2(keyinput_f2), .C1(DATAI_21_), .C2(
        keyinput_f11), .A(n21166), .ZN(n21171) );
  OAI22_X1 U24105 ( .A1(DATAI_11_), .A2(keyinput_f21), .B1(keyinput_f40), .B2(
        P1_CODEFETCH_REG_SCAN_IN), .ZN(n21167) );
  AOI221_X1 U24106 ( .B1(DATAI_11_), .B2(keyinput_f21), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(keyinput_f40), .A(n21167), .ZN(n21170)
         );
  OAI22_X1 U24107 ( .A1(P1_EAX_REG_30__SCAN_IN), .A2(keyinput_f117), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(keyinput_f70), .ZN(n21168) );
  AOI221_X1 U24108 ( .B1(P1_EAX_REG_30__SCAN_IN), .B2(keyinput_f117), .C1(
        keyinput_f70), .C2(P1_REIP_REG_13__SCAN_IN), .A(n21168), .ZN(n21169)
         );
  NAND4_X1 U24109 ( .A1(n21172), .A2(n21171), .A3(n21170), .A4(n21169), .ZN(
        n21182) );
  OAI22_X1 U24110 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(keyinput_f113), .B1(
        keyinput_f14), .B2(DATAI_18_), .ZN(n21173) );
  AOI221_X1 U24111 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(keyinput_f113), .C1(
        DATAI_18_), .C2(keyinput_f14), .A(n21173), .ZN(n21180) );
  OAI22_X1 U24112 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(keyinput_f116), .B1(
        keyinput_f115), .B2(P1_EBX_REG_0__SCAN_IN), .ZN(n21174) );
  AOI221_X1 U24113 ( .B1(P1_EAX_REG_31__SCAN_IN), .B2(keyinput_f116), .C1(
        P1_EBX_REG_0__SCAN_IN), .C2(keyinput_f115), .A(n21174), .ZN(n21179) );
  OAI22_X1 U24114 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(keyinput_f94), .B1(
        DATAI_1_), .B2(keyinput_f31), .ZN(n21175) );
  AOI221_X1 U24115 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(keyinput_f94), .C1(
        keyinput_f31), .C2(DATAI_1_), .A(n21175), .ZN(n21178) );
  OAI22_X1 U24116 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(keyinput_f125), .B1(
        P1_EBX_REG_26__SCAN_IN), .B2(keyinput_f89), .ZN(n21176) );
  AOI221_X1 U24117 ( .B1(P1_EAX_REG_22__SCAN_IN), .B2(keyinput_f125), .C1(
        keyinput_f89), .C2(P1_EBX_REG_26__SCAN_IN), .A(n21176), .ZN(n21177) );
  NAND4_X1 U24118 ( .A1(n21180), .A2(n21179), .A3(n21178), .A4(n21177), .ZN(
        n21181) );
  NOR4_X1 U24119 ( .A1(n21184), .A2(n21183), .A3(n21182), .A4(n21181), .ZN(
        n21310) );
  AOI22_X1 U24120 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(keyinput_f77), .B1(
        P1_EBX_REG_12__SCAN_IN), .B2(keyinput_f103), .ZN(n21185) );
  OAI221_X1 U24121 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(keyinput_f77), .C1(
        P1_EBX_REG_12__SCAN_IN), .C2(keyinput_f103), .A(n21185), .ZN(n21194)
         );
  AOI22_X1 U24122 ( .A1(DATAI_17_), .A2(keyinput_f15), .B1(
        P1_EBX_REG_7__SCAN_IN), .B2(keyinput_f108), .ZN(n21186) );
  OAI221_X1 U24123 ( .B1(DATAI_17_), .B2(keyinput_f15), .C1(
        P1_EBX_REG_7__SCAN_IN), .C2(keyinput_f108), .A(n21186), .ZN(n21193) );
  AOI22_X1 U24124 ( .A1(keyinput_f41), .A2(P1_M_IO_N_REG_SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(keyinput_f84), .ZN(n21187) );
  OAI221_X1 U24125 ( .B1(keyinput_f41), .B2(P1_M_IO_N_REG_SCAN_IN), .C1(
        P1_EBX_REG_31__SCAN_IN), .C2(keyinput_f84), .A(n21187), .ZN(n21192) );
  AOI22_X1 U24126 ( .A1(n21190), .A2(keyinput_f39), .B1(n21189), .B2(
        keyinput_f45), .ZN(n21188) );
  OAI221_X1 U24127 ( .B1(n21190), .B2(keyinput_f39), .C1(n21189), .C2(
        keyinput_f45), .A(n21188), .ZN(n21191) );
  NOR4_X1 U24128 ( .A1(n21194), .A2(n21193), .A3(n21192), .A4(n21191), .ZN(
        n21243) );
  INV_X1 U24129 ( .A(DATAI_2_), .ZN(n21197) );
  AOI22_X1 U24130 ( .A1(n21197), .A2(keyinput_f30), .B1(n21196), .B2(
        keyinput_f96), .ZN(n21195) );
  OAI221_X1 U24131 ( .B1(n21197), .B2(keyinput_f30), .C1(n21196), .C2(
        keyinput_f96), .A(n21195), .ZN(n21208) );
  INV_X1 U24132 ( .A(DATAI_28_), .ZN(n21199) );
  AOI22_X1 U24133 ( .A1(n13486), .A2(keyinput_f17), .B1(n21199), .B2(
        keyinput_f4), .ZN(n21198) );
  OAI221_X1 U24134 ( .B1(n13486), .B2(keyinput_f17), .C1(n21199), .C2(
        keyinput_f4), .A(n21198), .ZN(n21207) );
  AOI22_X1 U24135 ( .A1(n21202), .A2(keyinput_f99), .B1(keyinput_f24), .B2(
        n21201), .ZN(n21200) );
  OAI221_X1 U24136 ( .B1(n21202), .B2(keyinput_f99), .C1(n21201), .C2(
        keyinput_f24), .A(n21200), .ZN(n21206) );
  AOI22_X1 U24137 ( .A1(n14926), .A2(keyinput_f7), .B1(n21204), .B2(
        keyinput_f105), .ZN(n21203) );
  OAI221_X1 U24138 ( .B1(n14926), .B2(keyinput_f7), .C1(n21204), .C2(
        keyinput_f105), .A(n21203), .ZN(n21205) );
  NOR4_X1 U24139 ( .A1(n21208), .A2(n21207), .A3(n21206), .A4(n21205), .ZN(
        n21242) );
  INV_X1 U24140 ( .A(DATAI_6_), .ZN(n21211) );
  INV_X1 U24141 ( .A(DATAI_14_), .ZN(n21210) );
  AOI22_X1 U24142 ( .A1(n21211), .A2(keyinput_f26), .B1(n21210), .B2(
        keyinput_f18), .ZN(n21209) );
  OAI221_X1 U24143 ( .B1(n21211), .B2(keyinput_f26), .C1(n21210), .C2(
        keyinput_f18), .A(n21209), .ZN(n21223) );
  AOI22_X1 U24144 ( .A1(n14851), .A2(keyinput_f93), .B1(keyinput_f53), .B2(
        n21213), .ZN(n21212) );
  OAI221_X1 U24145 ( .B1(n14851), .B2(keyinput_f93), .C1(n21213), .C2(
        keyinput_f53), .A(n21212), .ZN(n21222) );
  AOI22_X1 U24146 ( .A1(n21216), .A2(keyinput_f92), .B1(keyinput_f95), .B2(
        n21215), .ZN(n21214) );
  OAI221_X1 U24147 ( .B1(n21216), .B2(keyinput_f92), .C1(n21215), .C2(
        keyinput_f95), .A(n21214), .ZN(n21221) );
  INV_X1 U24148 ( .A(keyinput_f51), .ZN(n21218) );
  AOI22_X1 U24149 ( .A1(n21219), .A2(keyinput_f64), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(n21218), .ZN(n21217) );
  OAI221_X1 U24150 ( .B1(n21219), .B2(keyinput_f64), .C1(n21218), .C2(
        P1_BYTEENABLE_REG_3__SCAN_IN), .A(n21217), .ZN(n21220) );
  NOR4_X1 U24151 ( .A1(n21223), .A2(n21222), .A3(n21221), .A4(n21220), .ZN(
        n21241) );
  AOI22_X1 U24152 ( .A1(n21226), .A2(keyinput_f73), .B1(keyinput_f68), .B2(
        n21225), .ZN(n21224) );
  OAI221_X1 U24153 ( .B1(n21226), .B2(keyinput_f73), .C1(n21225), .C2(
        keyinput_f68), .A(n21224), .ZN(n21239) );
  AOI22_X1 U24154 ( .A1(n21229), .A2(keyinput_f78), .B1(n21228), .B2(
        keyinput_f79), .ZN(n21227) );
  OAI221_X1 U24155 ( .B1(n21229), .B2(keyinput_f78), .C1(n21228), .C2(
        keyinput_f79), .A(n21227), .ZN(n21238) );
  AOI22_X1 U24156 ( .A1(n21232), .A2(keyinput_f59), .B1(keyinput_f62), .B2(
        n21231), .ZN(n21230) );
  OAI221_X1 U24157 ( .B1(n21232), .B2(keyinput_f59), .C1(n21231), .C2(
        keyinput_f62), .A(n21230), .ZN(n21237) );
  AOI22_X1 U24158 ( .A1(n21235), .A2(keyinput_f22), .B1(n21234), .B2(
        keyinput_f121), .ZN(n21233) );
  OAI221_X1 U24159 ( .B1(n21235), .B2(keyinput_f22), .C1(n21234), .C2(
        keyinput_f121), .A(n21233), .ZN(n21236) );
  NOR4_X1 U24160 ( .A1(n21239), .A2(n21238), .A3(n21237), .A4(n21236), .ZN(
        n21240) );
  NAND4_X1 U24161 ( .A1(n21243), .A2(n21242), .A3(n21241), .A4(n21240), .ZN(
        n21308) );
  AOI22_X1 U24162 ( .A1(n21246), .A2(keyinput_f75), .B1(n21245), .B2(
        keyinput_f104), .ZN(n21244) );
  OAI221_X1 U24163 ( .B1(n21246), .B2(keyinput_f75), .C1(n21245), .C2(
        keyinput_f104), .A(n21244), .ZN(n21307) );
  OAI22_X1 U24164 ( .A1(n21249), .A2(keyinput_f54), .B1(n21248), .B2(
        keyinput_f33), .ZN(n21247) );
  AOI221_X1 U24165 ( .B1(n21249), .B2(keyinput_f54), .C1(keyinput_f33), .C2(
        n21248), .A(n21247), .ZN(n21258) );
  OAI22_X1 U24166 ( .A1(n21252), .A2(keyinput_f106), .B1(n21251), .B2(
        keyinput_f13), .ZN(n21250) );
  AOI221_X1 U24167 ( .B1(n21252), .B2(keyinput_f106), .C1(keyinput_f13), .C2(
        n21251), .A(n21250), .ZN(n21257) );
  OAI22_X1 U24168 ( .A1(n21255), .A2(keyinput_f101), .B1(n21254), .B2(
        keyinput_f34), .ZN(n21253) );
  AOI221_X1 U24169 ( .B1(n21255), .B2(keyinput_f101), .C1(keyinput_f34), .C2(
        n21254), .A(n21253), .ZN(n21256) );
  NAND3_X1 U24170 ( .A1(n21258), .A2(n21257), .A3(n21256), .ZN(n21306) );
  OAI22_X1 U24171 ( .A1(n14930), .A2(keyinput_f123), .B1(n21260), .B2(
        keyinput_f86), .ZN(n21259) );
  AOI221_X1 U24172 ( .B1(n14930), .B2(keyinput_f123), .C1(keyinput_f86), .C2(
        n21260), .A(n21259), .ZN(n21304) );
  XNOR2_X1 U24173 ( .A(n21261), .B(keyinput_f47), .ZN(n21272) );
  XNOR2_X1 U24174 ( .A(keyinput_f49), .B(n21262), .ZN(n21271) );
  AOI22_X1 U24175 ( .A1(n21265), .A2(keyinput_f16), .B1(n21264), .B2(
        keyinput_f122), .ZN(n21263) );
  OAI221_X1 U24176 ( .B1(n21265), .B2(keyinput_f16), .C1(n21264), .C2(
        keyinput_f122), .A(n21263), .ZN(n21270) );
  INV_X1 U24177 ( .A(DATAI_5_), .ZN(n21268) );
  AOI22_X1 U24178 ( .A1(n21268), .A2(keyinput_f27), .B1(n21267), .B2(
        keyinput_f111), .ZN(n21266) );
  OAI221_X1 U24179 ( .B1(n21268), .B2(keyinput_f27), .C1(n21267), .C2(
        keyinput_f111), .A(n21266), .ZN(n21269) );
  NOR4_X1 U24180 ( .A1(n21272), .A2(n21271), .A3(n21270), .A4(n21269), .ZN(
        n21303) );
  INV_X1 U24181 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21274) );
  AOI22_X1 U24182 ( .A1(n15098), .A2(keyinput_f67), .B1(keyinput_f38), .B2(
        n21274), .ZN(n21273) );
  OAI221_X1 U24183 ( .B1(n15098), .B2(keyinput_f67), .C1(n21274), .C2(
        keyinput_f38), .A(n21273), .ZN(n21287) );
  AOI22_X1 U24184 ( .A1(n21277), .A2(keyinput_f29), .B1(n21276), .B2(
        keyinput_f74), .ZN(n21275) );
  OAI221_X1 U24185 ( .B1(n21277), .B2(keyinput_f29), .C1(n21276), .C2(
        keyinput_f74), .A(n21275), .ZN(n21286) );
  AOI22_X1 U24186 ( .A1(n21280), .A2(keyinput_f20), .B1(keyinput_f6), .B2(
        n21279), .ZN(n21278) );
  OAI221_X1 U24187 ( .B1(n21280), .B2(keyinput_f20), .C1(n21279), .C2(
        keyinput_f6), .A(n21278), .ZN(n21285) );
  AOI22_X1 U24188 ( .A1(n21283), .A2(keyinput_f98), .B1(keyinput_f23), .B2(
        n21282), .ZN(n21281) );
  OAI221_X1 U24189 ( .B1(n21283), .B2(keyinput_f98), .C1(n21282), .C2(
        keyinput_f23), .A(n21281), .ZN(n21284) );
  NOR4_X1 U24190 ( .A1(n21287), .A2(n21286), .A3(n21285), .A4(n21284), .ZN(
        n21302) );
  AOI22_X1 U24191 ( .A1(n21290), .A2(keyinput_f32), .B1(n21289), .B2(
        keyinput_f97), .ZN(n21288) );
  OAI221_X1 U24192 ( .B1(n21290), .B2(keyinput_f32), .C1(n21289), .C2(
        keyinput_f97), .A(n21288), .ZN(n21300) );
  AOI22_X1 U24193 ( .A1(n14996), .A2(keyinput_f55), .B1(keyinput_f76), .B2(
        n21292), .ZN(n21291) );
  OAI221_X1 U24194 ( .B1(n14996), .B2(keyinput_f55), .C1(n21292), .C2(
        keyinput_f76), .A(n21291), .ZN(n21299) );
  AOI22_X1 U24195 ( .A1(n21294), .A2(keyinput_f87), .B1(keyinput_f12), .B2(
        n14950), .ZN(n21293) );
  OAI221_X1 U24196 ( .B1(n21294), .B2(keyinput_f87), .C1(n14950), .C2(
        keyinput_f12), .A(n21293), .ZN(n21298) );
  AOI22_X1 U24197 ( .A1(n13685), .A2(keyinput_f82), .B1(n21296), .B2(
        keyinput_f109), .ZN(n21295) );
  OAI221_X1 U24198 ( .B1(n13685), .B2(keyinput_f82), .C1(n21296), .C2(
        keyinput_f109), .A(n21295), .ZN(n21297) );
  NOR4_X1 U24199 ( .A1(n21300), .A2(n21299), .A3(n21298), .A4(n21297), .ZN(
        n21301) );
  NAND4_X1 U24200 ( .A1(n21304), .A2(n21303), .A3(n21302), .A4(n21301), .ZN(
        n21305) );
  NOR4_X1 U24201 ( .A1(n21308), .A2(n21307), .A3(n21306), .A4(n21305), .ZN(
        n21309) );
  NAND4_X1 U24202 ( .A1(n21312), .A2(n21311), .A3(n21310), .A4(n21309), .ZN(
        n21314) );
  AOI21_X1 U24203 ( .B1(keyinput_f81), .B2(n21314), .A(keyinput_g81), .ZN(
        n21316) );
  INV_X1 U24204 ( .A(keyinput_f81), .ZN(n21313) );
  AOI21_X1 U24205 ( .B1(n21314), .B2(n21313), .A(P1_REIP_REG_2__SCAN_IN), .ZN(
        n21315) );
  AOI22_X1 U24206 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n21316), .B1(keyinput_g81), .B2(n21315), .ZN(n21317) );
  AOI21_X1 U24207 ( .B1(n21319), .B2(n21318), .A(n21317), .ZN(n21322) );
  AOI22_X1 U24208 ( .A1(n21320), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16710), .ZN(n21321) );
  XNOR2_X1 U24209 ( .A(n21322), .B(n21321), .ZN(U355) );
  INV_X2 U11407 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13827) );
  INV_X2 U11390 ( .A(n12959), .ZN(n12508) );
  NAND2_X2 U11337 ( .A1(n10711), .A2(n10710), .ZN(n14134) );
  NAND2_X1 U14642 ( .A1(n13634), .A2(n13633), .ZN(n13632) );
  AND2_X2 U11984 ( .A1(n13179), .A2(n20012), .ZN(n11538) );
  CLKBUF_X2 U11262 ( .A(n9943), .Z(n9815) );
  CLKBUF_X1 U11286 ( .A(n10653), .Z(n9817) );
  NAND2_X2 U11297 ( .A1(n11508), .A2(n10738), .ZN(n10751) );
  CLKBUF_X1 U11299 ( .A(n14462), .Z(n9811) );
  CLKBUF_X1 U11316 ( .A(n14462), .Z(n14236) );
  CLKBUF_X1 U11326 ( .A(n12252), .Z(n12253) );
  CLKBUF_X1 U11340 ( .A(n11517), .Z(n11690) );
  CLKBUF_X1 U11355 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n9932) );
  CLKBUF_X2 U11384 ( .A(n13993), .Z(n14630) );
  CLKBUF_X1 U11406 ( .A(n19312), .Z(n19324) );
  CLKBUF_X1 U11684 ( .A(n10840), .Z(n13472) );
  CLKBUF_X1 U11765 ( .A(n18951), .Z(n18944) );
endmodule

