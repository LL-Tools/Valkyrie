

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842;

  CLKBUF_X2 U3413 ( .A(n3243), .Z(n4583) );
  CLKBUF_X2 U3414 ( .A(n3342), .Z(n3317) );
  CLKBUF_X2 U3415 ( .A(n3396), .Z(n3917) );
  CLKBUF_X2 U3416 ( .A(n3390), .Z(n3894) );
  CLKBUF_X2 U3417 ( .A(n3318), .Z(n3919) );
  CLKBUF_X2 U3418 ( .A(n3306), .Z(n3391) );
  CLKBUF_X2 U3419 ( .A(n3325), .Z(n3889) );
  CLKBUF_X2 U3420 ( .A(n3319), .Z(n3909) );
  CLKBUF_X1 U3421 ( .A(n3284), .Z(n4508) );
  NOR2_X1 U3422 ( .A1(n4554), .A2(n2995), .ZN(n3282) );
  AND2_X2 U3423 ( .A1(n4406), .A2(n3005), .ZN(n3319) );
  AND2_X1 U3424 ( .A1(n2989), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3058)
         );
  CLKBUF_X2 U3425 ( .A(n3916), .Z(n3895) );
  AND2_X1 U3426 ( .A1(n4554), .A2(n5610), .ZN(n4077) );
  NAND2_X1 U3427 ( .A1(n3157), .A2(n3156), .ZN(n3265) );
  INV_X1 U3428 ( .A(n4036), .ZN(n3264) );
  CLKBUF_X3 U3429 ( .A(n3943), .Z(n4480) );
  OR2_X2 U3430 ( .A1(n6668), .A2(n5253), .ZN(n6151) );
  AND2_X2 U3431 ( .A1(n6151), .A2(n5301), .ZN(n6189) );
  INV_X1 U3432 ( .A(n5833), .ZN(n6336) );
  INV_X1 U3433 ( .A(n6345), .ZN(n6312) );
  NAND2_X2 U3434 ( .A1(n6151), .A2(n5255), .ZN(n6199) );
  NOR2_X2 U3435 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n3144), .ZN(n3151)
         );
  OR2_X2 U3436 ( .A1(n6581), .A2(n6587), .ZN(n4432) );
  AND2_X1 U3437 ( .A1(n5300), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5301) );
  INV_X4 U3438 ( .A(n5756), .ZN(n6025) );
  CLKBUF_X1 U3439 ( .A(n3273), .Z(n4472) );
  CLKBUF_X2 U3440 ( .A(n4212), .Z(n5267) );
  INV_X1 U3441 ( .A(n3282), .ZN(n3963) );
  CLKBUF_X2 U3442 ( .A(n3303), .Z(n3920) );
  CLKBUF_X2 U3443 ( .A(n3244), .Z(n3911) );
  OR2_X1 U3444 ( .A1(n5845), .A2(n6316), .ZN(n3002) );
  NAND2_X1 U34450 ( .A1(n5789), .A2(n3041), .ZN(n5783) );
  NAND2_X1 U34460 ( .A1(n5791), .A2(n5790), .ZN(n5789) );
  CLKBUF_X1 U34470 ( .A(n5334), .Z(n5347) );
  NAND2_X1 U34480 ( .A1(n6318), .A2(n3994), .ZN(n5138) );
  AND2_X1 U3449 ( .A1(n3045), .A2(n3115), .ZN(n3050) );
  AND2_X1 U3450 ( .A1(n3116), .A2(n5801), .ZN(n3115) );
  INV_X4 U34510 ( .A(n6189), .ZN(n6217) );
  NAND2_X1 U34520 ( .A1(n2978), .A2(n5831), .ZN(n3118) );
  AND2_X1 U34530 ( .A1(n3568), .A2(n4476), .ZN(n4709) );
  INV_X2 U3454 ( .A(n5756), .ZN(n5781) );
  OAI211_X1 U34550 ( .C1(n3001), .C2(n4425), .A(n2998), .B(n3950), .ZN(n6337)
         );
  NAND4_X1 U34560 ( .A1(n3590), .A2(n4519), .A3(n3140), .A4(n3591), .ZN(n3581)
         );
  NAND2_X1 U3457 ( .A1(n3831), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3881)
         );
  NAND2_X1 U3458 ( .A1(n3375), .A2(n3374), .ZN(n3591) );
  CLKBUF_X1 U34590 ( .A(n5612), .Z(n5649) );
  OAI21_X2 U34600 ( .B1(n3947), .B2(n4060), .A(n3946), .ZN(n4385) );
  NAND2_X1 U34610 ( .A1(n3550), .A2(n3549), .ZN(n3947) );
  CLKBUF_X1 U34620 ( .A(n4484), .Z(n5552) );
  NAND2_X1 U34630 ( .A1(n5244), .A2(n5243), .ZN(n6668) );
  XNOR2_X1 U34640 ( .A(n3405), .B(n4734), .ZN(n4484) );
  AOI21_X2 U34650 ( .B1(n3019), .B2(n4091), .A(n4090), .ZN(n6581) );
  NAND2_X1 U3466 ( .A1(n3014), .A2(n3013), .ZN(n3019) );
  OR2_X1 U3467 ( .A1(n3367), .A2(n3142), .ZN(n3377) );
  NOR2_X1 U34680 ( .A1(n4459), .A2(n4456), .ZN(n4141) );
  NAND2_X1 U34690 ( .A1(n4088), .A2(n4087), .ZN(n4091) );
  NAND2_X1 U34700 ( .A1(n3338), .A2(n3337), .ZN(n3548) );
  NOR2_X1 U34710 ( .A1(n4089), .A2(n4237), .ZN(n4090) );
  NAND2_X1 U34720 ( .A1(n3216), .A2(n3215), .ZN(n4108) );
  INV_X2 U34730 ( .A(n4110), .ZN(n4132) );
  NAND2_X1 U34740 ( .A1(n3272), .A2(n3271), .ZN(n4067) );
  OR2_X1 U3475 ( .A1(n3316), .A2(n3315), .ZN(n3999) );
  NAND2_X1 U3476 ( .A1(n3006), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3007) );
  BUF_X2 U3477 ( .A(n3265), .Z(n5610) );
  INV_X1 U3478 ( .A(n4244), .ZN(n4527) );
  AND3_X2 U3479 ( .A1(n3134), .A2(n3202), .A3(n3138), .ZN(n4244) );
  INV_X1 U3480 ( .A(n3265), .ZN(n2965) );
  AND4_X1 U3481 ( .A1(n3260), .A2(n3259), .A3(n3262), .A4(n3261), .ZN(n3302)
         );
  NAND2_X1 U3482 ( .A1(n3057), .A2(n3056), .ZN(n3284) );
  NAND4_X2 U3483 ( .A1(n3262), .A2(n3261), .A3(n3260), .A4(n3259), .ZN(n3271)
         );
  AND4_X1 U3484 ( .A1(n3179), .A2(n3178), .A3(n3177), .A4(n3176), .ZN(n3260)
         );
  AND4_X1 U3485 ( .A1(n3187), .A2(n3186), .A3(n3185), .A4(n3184), .ZN(n3262)
         );
  AND4_X1 U3486 ( .A1(n3191), .A2(n3190), .A3(n3189), .A4(n3188), .ZN(n3261)
         );
  AND4_X1 U3487 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n3259)
         );
  AND4_X1 U3488 ( .A1(n3161), .A2(n3160), .A3(n3165), .A4(n3158), .ZN(n3057)
         );
  AND4_X1 U3489 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .ZN(n3157)
         );
  AND4_X1 U3490 ( .A1(n3155), .A2(n3154), .A3(n3153), .A4(n3152), .ZN(n3156)
         );
  AND4_X1 U3491 ( .A1(n3159), .A2(n3164), .A3(n3163), .A4(n3162), .ZN(n3056)
         );
  BUF_X2 U3492 ( .A(n3237), .Z(n3910) );
  BUF_X2 U3493 ( .A(n3341), .Z(n2966) );
  AND2_X2 U3494 ( .A1(n3058), .A2(n4401), .ZN(n3318) );
  BUF_X2 U3495 ( .A(n3343), .Z(n3305) );
  AND2_X2 U3496 ( .A1(n3150), .A2(n4578), .ZN(n3348) );
  AND2_X1 U3497 ( .A1(n4033), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3150)
         );
  CLKBUF_X1 U3498 ( .A(n5251), .Z(n3934) );
  AND2_X1 U3499 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4580) );
  NOR2_X2 U3500 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4578) );
  NOR2_X1 U3501 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5251) );
  AND2_X4 U3502 ( .A1(n3283), .A2(n4554), .ZN(n4110) );
  NAND2_X1 U3503 ( .A1(n3118), .A2(n4017), .ZN(n3116) );
  NAND3_X1 U3504 ( .A1(n4519), .A2(n3590), .A3(n3591), .ZN(n3593) );
  AND2_X1 U3505 ( .A1(n4081), .A2(n4084), .ZN(n4076) );
  AND2_X2 U3506 ( .A1(n4402), .A2(n4578), .ZN(n3325) );
  OR2_X1 U3507 ( .A1(n4548), .A2(n6575), .ZN(n3139) );
  NOR2_X1 U3508 ( .A1(n4397), .A2(n4119), .ZN(n4267) );
  AND2_X1 U3509 ( .A1(n4249), .A2(n4302), .ZN(n4364) );
  AND2_X1 U3510 ( .A1(n3216), .A2(n4548), .ZN(n3194) );
  NAND2_X1 U3511 ( .A1(n3053), .A2(n3052), .ZN(n4008) );
  INV_X1 U3512 ( .A(n3580), .ZN(n3052) );
  INV_X1 U3513 ( .A(n3581), .ZN(n3053) );
  AOI21_X1 U3514 ( .B1(n3273), .B2(n3283), .A(n3263), .ZN(n3270) );
  AOI21_X1 U3515 ( .B1(n4073), .B2(n4072), .A(n4071), .ZN(n4081) );
  INV_X1 U3516 ( .A(n4070), .ZN(n4072) );
  INV_X1 U3517 ( .A(n4208), .ZN(n5257) );
  INV_X1 U3518 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n2989) );
  NOR2_X1 U3519 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3145) );
  OAI21_X1 U3520 ( .B1(n3073), .B2(n4023), .A(n4027), .ZN(n3071) );
  NOR2_X1 U3521 ( .A1(n2971), .A2(n3063), .ZN(n3061) );
  INV_X1 U3522 ( .A(n3064), .ZN(n3063) );
  AND2_X1 U3523 ( .A1(n3044), .A2(n4020), .ZN(n3043) );
  NAND2_X1 U3524 ( .A1(n3128), .A2(n3050), .ZN(n2996) );
  INV_X1 U3525 ( .A(n3128), .ZN(n3049) );
  AND3_X1 U3526 ( .A1(n2965), .A2(n4244), .A3(n3362), .ZN(n4393) );
  NAND2_X1 U3527 ( .A1(n3594), .A2(n3593), .ZN(n3966) );
  NAND2_X1 U3528 ( .A1(n6048), .A2(n4489), .ZN(n4499) );
  NAND2_X1 U3529 ( .A1(n3409), .A2(n3408), .ZN(n4734) );
  INV_X1 U3530 ( .A(n3139), .ZN(n3720) );
  NAND2_X1 U3531 ( .A1(n4363), .A2(n4362), .ZN(n4470) );
  OR2_X1 U3532 ( .A1(n5244), .A2(n4310), .ZN(n6287) );
  AOI21_X1 U3533 ( .B1(n5251), .B2(n5699), .A(n3849), .ZN(n5348) );
  OR3_X1 U3534 ( .A1(n5705), .A2(n5756), .A3(n4028), .ZN(n5666) );
  NAND2_X1 U3535 ( .A1(n3004), .A2(n3003), .ZN(n5705) );
  INV_X1 U3536 ( .A(n3071), .ZN(n3003) );
  NAND2_X1 U3537 ( .A1(n5754), .A2(n3072), .ZN(n3004) );
  OAI21_X1 U3538 ( .B1(n5754), .B2(n3071), .A(n3069), .ZN(n5703) );
  AND2_X1 U3539 ( .A1(n3070), .A2(n5704), .ZN(n3069) );
  OR2_X1 U3540 ( .A1(n3071), .A2(n3072), .ZN(n3070) );
  AND3_X1 U3541 ( .A1(n4279), .A2(n5961), .A3(n3025), .ZN(n5216) );
  NOR2_X1 U3542 ( .A1(n3026), .A2(n2973), .ZN(n3025) );
  NOR2_X1 U3543 ( .A1(n2971), .A2(n5747), .ZN(n5746) );
  NAND2_X1 U3544 ( .A1(n5986), .A2(n5982), .ZN(n6387) );
  NAND2_X1 U3545 ( .A1(n4253), .A2(n4468), .ZN(n4274) );
  INV_X1 U3546 ( .A(n6587), .ZN(n4468) );
  AND4_X1 U3547 ( .A1(n3232), .A2(n3231), .A3(n3230), .A4(n3229), .ZN(n3252)
         );
  AND4_X1 U3548 ( .A1(n3236), .A2(n3235), .A3(n3234), .A4(n3233), .ZN(n3251)
         );
  INV_X1 U3549 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6575) );
  INV_X1 U3550 ( .A(n6351), .ZN(n6438) );
  AND2_X1 U3551 ( .A1(n3548), .A2(n6579), .ZN(n3121) );
  INV_X1 U3552 ( .A(n5454), .ZN(n3707) );
  INV_X1 U3553 ( .A(n5468), .ZN(n3079) );
  NAND2_X1 U3554 ( .A1(n3123), .A2(n2974), .ZN(n3073) );
  AOI21_X1 U3555 ( .B1(n5747), .B2(n3065), .A(n4226), .ZN(n3064) );
  NAND2_X1 U3556 ( .A1(n3042), .A2(n5830), .ZN(n3045) );
  OR2_X1 U3557 ( .A1(n3339), .A2(n6579), .ZN(n4006) );
  NAND2_X1 U3558 ( .A1(n4256), .A2(n3999), .ZN(n3339) );
  NAND2_X1 U3559 ( .A1(n3255), .A2(n2965), .ZN(n3256) );
  INV_X1 U3560 ( .A(n3364), .ZN(n3255) );
  OR2_X1 U3561 ( .A1(n4472), .A2(n3963), .ZN(n3287) );
  INV_X1 U3562 ( .A(n3007), .ZN(n3403) );
  INV_X1 U3563 ( .A(n3951), .ZN(n3960) );
  CLKBUF_X1 U3564 ( .A(n3291), .Z(n3292) );
  NOR2_X1 U3565 ( .A1(n3040), .A2(n3039), .ZN(n3038) );
  INV_X1 U3566 ( .A(n5373), .ZN(n3039) );
  XNOR2_X1 U3567 ( .A(n4008), .B(n3028), .ZN(n3995) );
  INV_X1 U3568 ( .A(n3458), .ZN(n3028) );
  INV_X1 U3569 ( .A(n3459), .ZN(n3462) );
  AND3_X1 U3570 ( .A1(n4606), .A2(n4699), .A3(n4454), .ZN(n4710) );
  INV_X1 U3571 ( .A(n5251), .ZN(n3908) );
  AND2_X1 U3572 ( .A1(n3553), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3556) );
  INV_X1 U3573 ( .A(n5374), .ZN(n3096) );
  NOR2_X1 U3574 ( .A1(n5384), .A2(n3098), .ZN(n3097) );
  INV_X1 U3575 ( .A(n4262), .ZN(n3098) );
  AND2_X1 U3576 ( .A1(n5482), .A2(n5464), .ZN(n3109) );
  NAND2_X1 U3577 ( .A1(n3115), .A2(n3117), .ZN(n3112) );
  NOR2_X1 U3578 ( .A1(n3106), .A2(n3105), .ZN(n3104) );
  INV_X1 U3579 ( .A(n6028), .ZN(n3105) );
  NAND2_X1 U3580 ( .A1(n4008), .A2(n4007), .ZN(n4013) );
  NOR2_X1 U3581 ( .A1(n4006), .A2(n4060), .ZN(n4007) );
  OR2_X1 U3582 ( .A1(n4160), .A2(n3107), .ZN(n3106) );
  INV_X1 U3583 ( .A(n5191), .ZN(n3107) );
  NOR2_X1 U3584 ( .A1(n3129), .A2(n3127), .ZN(n3126) );
  INV_X1 U3585 ( .A(n5137), .ZN(n3129) );
  INV_X1 U3586 ( .A(n4136), .ZN(n4201) );
  OR2_X1 U3587 ( .A1(n3354), .A2(n3353), .ZN(n3940) );
  INV_X1 U3588 ( .A(n4077), .ZN(n4060) );
  NAND2_X1 U3589 ( .A1(n4484), .A2(n6579), .ZN(n3422) );
  AOI21_X1 U3590 ( .B1(n4075), .B2(n4076), .A(n4074), .ZN(n4080) );
  AND2_X1 U3591 ( .A1(n4067), .A2(n4066), .ZN(n4068) );
  INV_X1 U3592 ( .A(n4080), .ZN(n3018) );
  NOR2_X1 U3593 ( .A1(n4093), .A2(n4094), .ZN(n4254) );
  AND2_X1 U3594 ( .A1(n4239), .A2(n4238), .ZN(n4910) );
  CLKBUF_X1 U3595 ( .A(n4248), .Z(n4911) );
  AND2_X2 U3596 ( .A1(n6151), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5545) );
  OR2_X1 U3597 ( .A1(n5260), .A2(n5259), .ZN(n3136) );
  AND2_X1 U3598 ( .A1(n4188), .A2(n4187), .ZN(n5434) );
  NOR2_X1 U3599 ( .A1(n6002), .A2(n5606), .ZN(n5973) );
  INV_X1 U3600 ( .A(n4357), .ZN(n5269) );
  NOR2_X2 U3601 ( .A1(n3830), .A2(n5700), .ZN(n3831) );
  NAND2_X1 U3602 ( .A1(n3753), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3769)
         );
  INV_X1 U3603 ( .A(n3754), .ZN(n3753) );
  CLKBUF_X1 U3604 ( .A(n5452), .Z(n5467) );
  INV_X1 U3605 ( .A(n5604), .ZN(n3078) );
  NAND2_X1 U3606 ( .A1(n5138), .A2(n5137), .ZN(n5136) );
  NOR2_X1 U3607 ( .A1(n5267), .A2(EBX_REG_29__SCAN_IN), .ZN(n4215) );
  NAND2_X1 U3608 ( .A1(n5781), .A2(n6775), .ZN(n3133) );
  NAND2_X1 U3609 ( .A1(n5703), .A2(n3133), .ZN(n5684) );
  AND2_X1 U3610 ( .A1(n6025), .A2(n4227), .ZN(n4228) );
  NOR2_X1 U3611 ( .A1(n5417), .A2(n4192), .ZN(n5404) );
  NOR2_X1 U3612 ( .A1(n3061), .A2(n3059), .ZN(n5728) );
  NAND2_X1 U3613 ( .A1(n3062), .A2(n3060), .ZN(n3059) );
  INV_X1 U3614 ( .A(n5729), .ZN(n3060) );
  NOR2_X1 U3615 ( .A1(n3125), .A2(n4019), .ZN(n3068) );
  NAND2_X1 U3616 ( .A1(n5781), .A2(n6796), .ZN(n3041) );
  OR2_X1 U3617 ( .A1(n6000), .A2(n6001), .ZN(n6002) );
  INV_X1 U3618 ( .A(n4017), .ZN(n3117) );
  NAND2_X1 U3619 ( .A1(n5829), .A2(n5830), .ZN(n4014) );
  NAND2_X1 U3620 ( .A1(n5231), .A2(n6579), .ZN(n4102) );
  INV_X1 U3621 ( .A(n4212), .ZN(n4901) );
  NAND2_X1 U3622 ( .A1(n3012), .A2(n3011), .ZN(n5982) );
  INV_X1 U3623 ( .A(n4267), .ZN(n3011) );
  NAND2_X1 U3624 ( .A1(n3119), .A2(n3548), .ZN(n3549) );
  XNOR2_X1 U3625 ( .A(n3558), .B(n3559), .ZN(n3943) );
  NOR2_X1 U3626 ( .A1(n5033), .A2(n4480), .ZN(n5045) );
  NOR2_X1 U3627 ( .A1(n4926), .A2(n4925), .ZN(n5088) );
  AND2_X1 U3628 ( .A1(n4480), .A2(n5044), .ZN(n6054) );
  NAND2_X1 U3629 ( .A1(n4499), .A2(n6579), .ZN(n4926) );
  INV_X1 U3630 ( .A(n5043), .ZN(n5044) );
  AND2_X1 U3631 ( .A1(n4480), .A2(n5043), .ZN(n4922) );
  INV_X1 U3632 ( .A(n5038), .ZN(n6499) );
  AND2_X1 U3633 ( .A1(n4599), .A2(n4598), .ZN(n4915) );
  OR2_X1 U3634 ( .A1(n4241), .A2(n3963), .ZN(n4919) );
  OR2_X1 U3635 ( .A1(n5311), .A2(n5608), .ZN(n4224) );
  AND2_X2 U3636 ( .A1(n4124), .A2(n4468), .ZN(n6243) );
  OR2_X1 U3637 ( .A1(n4467), .A2(n5267), .ZN(n4122) );
  XNOR2_X1 U3638 ( .A(n3939), .B(n3938), .ZN(n5250) );
  OR2_X1 U3639 ( .A1(n5334), .A2(n2981), .ZN(n3939) );
  NOR2_X2 U3640 ( .A1(n5656), .A2(n5239), .ZN(n5650) );
  OAI21_X1 U3641 ( .B1(n4470), .B2(n4469), .A(n4468), .ZN(n4471) );
  INV_X2 U3642 ( .A(n6247), .ZN(n5658) );
  OR2_X1 U3643 ( .A1(n4432), .A2(n4919), .ZN(n6307) );
  XNOR2_X1 U3644 ( .A(n5314), .B(n3082), .ZN(n5663) );
  OR2_X1 U3645 ( .A1(n4432), .A2(n4914), .ZN(n6316) );
  INV_X1 U3646 ( .A(n6316), .ZN(n6340) );
  XNOR2_X1 U3647 ( .A(n4031), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5845)
         );
  NAND2_X1 U3648 ( .A1(n5844), .A2(n3024), .ZN(n3023) );
  INV_X1 U3649 ( .A(n5842), .ZN(n3024) );
  NOR2_X1 U3650 ( .A1(n5905), .A2(n5219), .ZN(n5890) );
  OR2_X1 U3651 ( .A1(n4274), .A2(n4258), .ZN(n6351) );
  INV_X1 U3652 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5152) );
  CLKBUF_X1 U3654 ( .A(n4482), .Z(n4483) );
  CLKBUF_X1 U3655 ( .A(n3955), .Z(n6043) );
  INV_X1 U3656 ( .A(n6497), .ZN(n6666) );
  NAND2_X1 U3657 ( .A1(n4497), .A2(n6054), .ZN(n6565) );
  NAND2_X1 U3658 ( .A1(n4059), .A2(n4058), .ZN(n4073) );
  CLKBUF_X2 U3659 ( .A(n3324), .Z(n3918) );
  OR2_X1 U3660 ( .A1(n3444), .A2(n3443), .ZN(n3987) );
  NOR2_X1 U3661 ( .A1(n4554), .A2(n3254), .ZN(n3364) );
  AND2_X1 U3662 ( .A1(n3122), .A2(n3120), .ZN(n3340) );
  OR2_X1 U3663 ( .A1(n3420), .A2(n3419), .ZN(n3970) );
  AND2_X1 U3664 ( .A1(n4235), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4040) );
  NAND2_X1 U3665 ( .A1(n3302), .A2(n3265), .ZN(n4036) );
  INV_X1 U3666 ( .A(n5270), .ZN(n2995) );
  NAND2_X1 U3667 ( .A1(n3085), .A2(n3084), .ZN(n3083) );
  INV_X1 U3668 ( .A(n5335), .ZN(n3084) );
  NOR2_X1 U3669 ( .A1(n3086), .A2(n5315), .ZN(n3085) );
  INV_X1 U3670 ( .A(n5325), .ZN(n3086) );
  AND2_X1 U3671 ( .A1(n3708), .A2(n2980), .ZN(n5346) );
  INV_X1 U3672 ( .A(n5362), .ZN(n3037) );
  OR2_X1 U3673 ( .A1(n3807), .A2(n3806), .ZN(n3823) );
  NAND2_X1 U3674 ( .A1(n2979), .A2(n3707), .ZN(n3040) );
  INV_X1 U3675 ( .A(n3089), .ZN(n3088) );
  INV_X1 U3676 ( .A(n5383), .ZN(n3087) );
  NAND2_X1 U3677 ( .A1(n3772), .A2(n3090), .ZN(n3089) );
  INV_X1 U3678 ( .A(n3091), .ZN(n3090) );
  AND2_X1 U3679 ( .A1(n5407), .A2(n5203), .ZN(n3772) );
  NAND2_X1 U3680 ( .A1(n5421), .A2(n3092), .ZN(n3091) );
  NAND2_X1 U3681 ( .A1(n3708), .A2(n3707), .ZN(n5436) );
  INV_X1 U3682 ( .A(n3902), .ZN(n3932) );
  AOI21_X1 U3683 ( .B1(n3623), .B2(n5805), .A(n2969), .ZN(n3029) );
  NAND2_X1 U3684 ( .A1(n3688), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3690)
         );
  INV_X1 U3685 ( .A(n3687), .ZN(n3688) );
  NOR2_X1 U3686 ( .A1(n4400), .A2(n6579), .ZN(n3902) );
  OR2_X1 U3687 ( .A1(n3674), .A2(n3081), .ZN(n3080) );
  INV_X1 U3688 ( .A(n5603), .ZN(n3081) );
  OR2_X1 U3689 ( .A1(n5487), .A2(n5654), .ZN(n3674) );
  AND2_X1 U3690 ( .A1(n4824), .A2(n3605), .ZN(n3611) );
  AND3_X1 U3691 ( .A1(n3604), .A2(n4709), .A3(n4710), .ZN(n3605) );
  NAND2_X1 U3692 ( .A1(n3611), .A2(n3610), .ZN(n3623) );
  XNOR2_X1 U3693 ( .A(n3525), .B(n3524), .ZN(n3977) );
  INV_X1 U3694 ( .A(n3593), .ZN(n3447) );
  AND2_X1 U3695 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3460), .ZN(n3572)
         );
  INV_X1 U3696 ( .A(n3284), .ZN(n3551) );
  INV_X1 U3697 ( .A(n3073), .ZN(n3072) );
  INV_X1 U3698 ( .A(n5917), .ZN(n3026) );
  AND2_X1 U3699 ( .A1(n3055), .A2(n2970), .ZN(n3062) );
  NAND2_X1 U3700 ( .A1(n3064), .A2(n3066), .ZN(n3055) );
  AND2_X1 U3701 ( .A1(n4189), .A2(n5432), .ZN(n5416) );
  AOI21_X1 U3702 ( .B1(n4023), .B2(n3124), .A(n2976), .ZN(n3123) );
  INV_X1 U3703 ( .A(n4021), .ZN(n3124) );
  AOI21_X1 U3704 ( .B1(n5195), .B2(n3131), .A(n2977), .ZN(n3130) );
  INV_X1 U3705 ( .A(n4005), .ZN(n3131) );
  OR2_X1 U3706 ( .A1(n3402), .A2(n3401), .ZN(n3951) );
  OR2_X1 U3707 ( .A1(n3331), .A2(n3330), .ZN(n3944) );
  NAND2_X1 U3708 ( .A1(n3277), .A2(n3276), .ZN(n3380) );
  OAI21_X1 U3709 ( .B1(n6039), .B2(STATE2_REG_0__SCAN_IN), .A(n3371), .ZN(
        n3557) );
  OR2_X1 U3710 ( .A1(n4472), .A2(n3640), .ZN(n4400) );
  AND4_X1 U3711 ( .A1(n4116), .A2(n4115), .A3(n4114), .A4(n4113), .ZN(n4118)
         );
  OAI21_X1 U3712 ( .B1(n3379), .B2(n3378), .A(n3377), .ZN(n3388) );
  AND2_X1 U3713 ( .A1(n3222), .A2(n3221), .ZN(n3225) );
  AOI22_X1 U3714 ( .A1(n3342), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3319), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3209) );
  AND2_X1 U3715 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3381) );
  NAND2_X1 U3716 ( .A1(n3396), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U3717 ( .A1(n3348), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3232) );
  OR2_X1 U3718 ( .A1(n3271), .A2(n6579), .ZN(n3410) );
  INV_X1 U3719 ( .A(n3005), .ZN(n4571) );
  INV_X1 U3720 ( .A(n4554), .ZN(n4120) );
  OR2_X1 U3721 ( .A1(n6150), .A2(n5281), .ZN(n5492) );
  INV_X1 U3722 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6170) );
  INV_X1 U3723 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5519) );
  INV_X1 U3724 ( .A(n5242), .ZN(n5530) );
  INV_X1 U3725 ( .A(n6143), .ZN(n6214) );
  AND2_X1 U3726 ( .A1(n4166), .A2(n4165), .ZN(n6028) );
  AND2_X2 U3727 ( .A1(n4401), .A2(n3005), .ZN(n3324) );
  NAND2_X1 U3728 ( .A1(n3884), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4100)
         );
  INV_X1 U3729 ( .A(n3796), .ZN(n3797) );
  OR2_X2 U3730 ( .A1(n3738), .A2(n3737), .ZN(n3754) );
  NOR2_X2 U3731 ( .A1(n3690), .A2(n5472), .ZN(n3691) );
  NAND2_X1 U3732 ( .A1(n5802), .A2(n3623), .ZN(n5604) );
  AND2_X1 U3733 ( .A1(n3606), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3607)
         );
  NAND2_X1 U3734 ( .A1(n3607), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3634)
         );
  OR2_X1 U3735 ( .A1(n5804), .A2(n5805), .ZN(n5802) );
  NOR2_X1 U3736 ( .A1(n3508), .A2(n6181), .ZN(n3477) );
  NAND2_X1 U3737 ( .A1(n3503), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3508)
         );
  NOR2_X2 U3738 ( .A1(n3586), .A2(n5519), .ZN(n3503) );
  NAND2_X1 U3739 ( .A1(n3995), .A2(n3664), .ZN(n3027) );
  NOR2_X1 U3740 ( .A1(n5517), .A2(n3908), .ZN(n3461) );
  OR2_X1 U3741 ( .A1(n4726), .A2(n3639), .ZN(n3603) );
  NAND2_X1 U3742 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3595) );
  OAI211_X1 U3743 ( .C1(n3600), .C2(n4412), .A(n3561), .B(n3560), .ZN(n4376)
         );
  OR3_X1 U3744 ( .A1(n5863), .A2(n5223), .A3(n5847), .ZN(n5840) );
  AND2_X1 U3745 ( .A1(n2982), .A2(n3095), .ZN(n3094) );
  INV_X1 U3746 ( .A(n5365), .ZN(n3095) );
  AND2_X1 U3747 ( .A1(n4203), .A2(n4202), .ZN(n5374) );
  NAND2_X1 U3748 ( .A1(n5406), .A2(n3097), .ZN(n5386) );
  OR2_X1 U3749 ( .A1(n3061), .A2(n3054), .ZN(n5730) );
  INV_X1 U3750 ( .A(n3062), .ZN(n3054) );
  INV_X1 U3751 ( .A(n5434), .ZN(n3108) );
  NAND2_X1 U3752 ( .A1(n5769), .A2(n2984), .ZN(n5766) );
  AND2_X1 U3753 ( .A1(n5481), .A2(n5482), .ZN(n5484) );
  INV_X1 U3754 ( .A(n5754), .ZN(n5755) );
  NAND2_X1 U3755 ( .A1(n3048), .A2(n3046), .ZN(n3111) );
  NAND2_X1 U3756 ( .A1(n2967), .A2(n3047), .ZN(n3046) );
  INV_X1 U3757 ( .A(n3050), .ZN(n3047) );
  NAND2_X1 U3758 ( .A1(n3103), .A2(n2968), .ZN(n6000) );
  INV_X1 U3759 ( .A(n5081), .ZN(n3102) );
  NAND2_X1 U3760 ( .A1(n3103), .A2(n3104), .ZN(n6031) );
  NOR2_X1 U3761 ( .A1(n4828), .A2(n3106), .ZN(n6029) );
  NOR2_X1 U3762 ( .A1(n4828), .A2(n4160), .ZN(n5192) );
  AND2_X1 U3763 ( .A1(n6355), .A2(n6413), .ZN(n6349) );
  NAND2_X1 U3764 ( .A1(n4878), .A2(n3984), .ZN(n6320) );
  NAND2_X1 U3765 ( .A1(n6320), .A2(n6319), .ZN(n6318) );
  NAND2_X1 U3766 ( .A1(n4880), .A2(n4879), .ZN(n4878) );
  NAND2_X1 U3767 ( .A1(n4653), .A2(n4652), .ZN(n2994) );
  NOR2_X1 U3768 ( .A1(n6429), .A2(n6432), .ZN(n6413) );
  NAND2_X1 U3769 ( .A1(n2999), .A2(n3942), .ZN(n2998) );
  INV_X1 U3770 ( .A(n4274), .ZN(n3012) );
  NAND2_X1 U3771 ( .A1(n3943), .A2(n4077), .ZN(n3001) );
  NAND2_X1 U3772 ( .A1(n3012), .A2(n4577), .ZN(n6432) );
  CLKBUF_X1 U3773 ( .A(n3302), .Z(n4256) );
  INV_X1 U3774 ( .A(n3591), .ZN(n3076) );
  INV_X1 U3775 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4581) );
  OR3_X1 U3776 ( .A1(n4369), .A2(n4470), .A3(n4368), .ZN(n4891) );
  OR2_X1 U3777 ( .A1(n5552), .A2(n6056), .ZN(n4841) );
  AND2_X1 U3778 ( .A1(n4616), .A2(n4727), .ZN(n4619) );
  OR2_X1 U3779 ( .A1(n5552), .A2(n4719), .ZN(n4996) );
  BUF_X1 U3780 ( .A(n3966), .Z(n4726) );
  INV_X1 U3781 ( .A(n4480), .ZN(n4738) );
  AND3_X1 U3782 ( .A1(n6811), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6500) );
  INV_X1 U3783 ( .A(n6572), .ZN(n5128) );
  AND2_X1 U3784 ( .A1(n5045), .A2(n5044), .ZN(n5095) );
  AND2_X1 U3785 ( .A1(n4499), .A2(n4498), .ZN(n4555) );
  NAND2_X1 U3786 ( .A1(n4069), .A2(n3015), .ZN(n3014) );
  OR2_X1 U3787 ( .A1(n4080), .A2(n4079), .ZN(n3015) );
  AOI21_X1 U3788 ( .B1(n4079), .B2(n3016), .A(n2975), .ZN(n3013) );
  NAND2_X1 U3789 ( .A1(n3018), .A2(n3017), .ZN(n3016) );
  INV_X1 U3790 ( .A(n4068), .ZN(n3017) );
  NAND2_X1 U3791 ( .A1(n4075), .A2(n4077), .ZN(n4089) );
  NAND2_X1 U3792 ( .A1(n4086), .A2(n4085), .ZN(n4237) );
  OR2_X1 U3793 ( .A1(n4083), .A2(n4082), .ZN(n4086) );
  AND2_X1 U3794 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6444), .ZN(n4082)
         );
  NAND2_X2 U3795 ( .A1(n3410), .A2(n3007), .ZN(n4088) );
  INV_X1 U3796 ( .A(n4237), .ZN(n4087) );
  AND2_X1 U3797 ( .A1(n5254), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4092) );
  NAND2_X1 U3798 ( .A1(n4120), .A2(n3006), .ZN(n5242) );
  INV_X1 U3799 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6812) );
  NAND2_X1 U3800 ( .A1(n6151), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6143) );
  AND2_X1 U3801 ( .A1(n5545), .A2(n5299), .ZN(n6222) );
  AND2_X1 U3802 ( .A1(n5545), .A2(n5268), .ZN(n6211) );
  INV_X1 U3803 ( .A(n6222), .ZN(n6171) );
  INV_X1 U3804 ( .A(n6150), .ZN(n6207) );
  XNOR2_X1 U3805 ( .A(n5265), .B(n5264), .ZN(n5843) );
  OR2_X1 U3806 ( .A1(n5323), .A2(n5322), .ZN(n5857) );
  AND2_X1 U3807 ( .A1(n6249), .A2(n4474), .ZN(n6246) );
  INV_X1 U3808 ( .A(n6246), .ZN(n4711) );
  AND2_X1 U3809 ( .A1(n4434), .A2(n5269), .ZN(n6261) );
  NAND2_X1 U3810 ( .A1(n6307), .A2(n4433), .ZN(n4434) );
  AND2_X1 U3811 ( .A1(n4309), .A2(n6307), .ZN(n6305) );
  INV_X1 U3812 ( .A(n6287), .ZN(n6304) );
  AOI21_X1 U3813 ( .B1(n5315), .B2(n5313), .A(n5314), .ZN(n5672) );
  OAI21_X1 U3814 ( .B1(n5324), .B2(n5325), .A(n5313), .ZN(n5682) );
  AND2_X1 U3815 ( .A1(n3881), .A2(n3833), .ZN(n5699) );
  NAND2_X1 U3816 ( .A1(n5347), .A2(n3034), .ZN(n5697) );
  NAND2_X1 U3817 ( .A1(n3036), .A2(n3035), .ZN(n3034) );
  INV_X1 U3818 ( .A(n5348), .ZN(n3035) );
  INV_X1 U3819 ( .A(n5361), .ZN(n3036) );
  INV_X1 U3820 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U3821 ( .A1(n5196), .A2(n5195), .ZN(n5194) );
  NAND2_X1 U3822 ( .A1(n5136), .A2(n4005), .ZN(n5196) );
  NAND2_X1 U3823 ( .A1(n6316), .A2(n4096), .ZN(n5833) );
  OR2_X1 U3824 ( .A1(n5838), .A2(n5839), .ZN(n3101) );
  INV_X1 U3825 ( .A(n5837), .ZN(n5838) );
  XNOR2_X1 U3826 ( .A(n5212), .B(n5839), .ZN(n5665) );
  NAND2_X1 U3827 ( .A1(n5703), .A2(n3132), .ZN(n5677) );
  AND2_X1 U3828 ( .A1(n2985), .A2(n3133), .ZN(n3132) );
  INV_X1 U3829 ( .A(n5684), .ZN(n5695) );
  NAND2_X1 U3830 ( .A1(n5954), .A2(n4272), .ZN(n5902) );
  NAND2_X1 U3831 ( .A1(n5216), .A2(n5215), .ZN(n5905) );
  XNOR2_X1 U3832 ( .A(n4231), .B(n4230), .ZN(n5210) );
  NOR2_X1 U3833 ( .A1(n5728), .A2(n4228), .ZN(n4231) );
  NOR2_X1 U3834 ( .A1(n5746), .A2(n3066), .ZN(n5738) );
  INV_X1 U3835 ( .A(n5902), .ZN(n5935) );
  AOI21_X1 U3836 ( .B1(n4014), .B2(n3114), .A(n3117), .ZN(n3113) );
  INV_X1 U3837 ( .A(n3118), .ZN(n3114) );
  AND2_X1 U3838 ( .A1(n5961), .A2(n5960), .ZN(n6033) );
  AND2_X1 U3839 ( .A1(n6387), .A2(n4426), .ZN(n6428) );
  NAND2_X1 U3840 ( .A1(n4377), .A2(n4901), .ZN(n4379) );
  OR2_X1 U3841 ( .A1(n4274), .A2(n4261), .ZN(n6434) );
  AOI21_X1 U3842 ( .B1(n3010), .B2(n4416), .A(n3008), .ZN(n6391) );
  NOR2_X1 U3843 ( .A1(n3012), .A2(n3009), .ZN(n3008) );
  OR2_X1 U3844 ( .A1(n4274), .A2(n4592), .ZN(n5986) );
  INV_X1 U3845 ( .A(n3552), .ZN(n6490) );
  AND2_X1 U3846 ( .A1(n4480), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6042) );
  INV_X1 U3847 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5254) );
  INV_X1 U3848 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4412) );
  AND2_X2 U3849 ( .A1(n2997), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4406)
         );
  INV_X1 U3850 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n2997) );
  INV_X1 U3851 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5234) );
  OR2_X1 U3852 ( .A1(n6581), .A2(n4986), .ZN(n6048) );
  NOR2_X1 U3853 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5231) );
  NAND2_X1 U3854 ( .A1(n4619), .A2(n5044), .ZN(n4993) );
  INV_X1 U3855 ( .A(n4872), .ZN(n4647) );
  OAI21_X1 U3856 ( .B1(n4724), .B2(n4722), .A(n4721), .ZN(n6464) );
  NAND2_X1 U3857 ( .A1(n5157), .A2(n5156), .ZN(n5183) );
  AND2_X1 U3858 ( .A1(n4555), .A2(n4527), .ZN(n6476) );
  AND2_X1 U3859 ( .A1(n6055), .A2(n4737), .ZN(n6484) );
  NAND2_X1 U3860 ( .A1(n6055), .A2(n4922), .ZN(n6679) );
  OAI21_X1 U3861 ( .B1(n6063), .B2(n6062), .A(n6061), .ZN(n6092) );
  NOR2_X1 U3862 ( .A1(n4503), .A2(n4926), .ZN(n6480) );
  NOR2_X1 U3863 ( .A1(n4512), .A2(n4926), .ZN(n6452) );
  NOR2_X1 U3864 ( .A1(n4553), .A2(n4926), .ZN(n6547) );
  NOR2_X1 U3865 ( .A1(n4615), .A2(n4926), .ZN(n6558) );
  NOR2_X1 U3866 ( .A1(n6750), .A2(n4926), .ZN(n6568) );
  NOR2_X1 U3867 ( .A1(n4490), .A2(n4926), .ZN(n6468) );
  AND2_X1 U3868 ( .A1(n4765), .A2(n4764), .ZN(n4817) );
  OAI21_X1 U3869 ( .B1(n4761), .B2(n4760), .A(n4759), .ZN(n4816) );
  INV_X1 U3870 ( .A(n4823), .ZN(n4695) );
  OAI21_X1 U3871 ( .B1(n4669), .B2(n4758), .A(n6499), .ZN(n4692) );
  OR4_X1 U3872 ( .A1(n4952), .A2(n5155), .A3(n4990), .A4(n4951), .ZN(n4978) );
  INV_X1 U3873 ( .A(n6469), .ZN(n6494) );
  INV_X1 U3874 ( .A(n6468), .ZN(n6505) );
  INV_X1 U3875 ( .A(n6547), .ZN(n6510) );
  INV_X1 U3876 ( .A(n6472), .ZN(n6544) );
  INV_X1 U3877 ( .A(n6552), .ZN(n6682) );
  INV_X1 U3878 ( .A(n6476), .ZN(n6676) );
  INV_X1 U3879 ( .A(n6483), .ZN(n6511) );
  INV_X1 U3880 ( .A(n6450), .ZN(n6518) );
  INV_X1 U3881 ( .A(n6452), .ZN(n6525) );
  INV_X1 U3882 ( .A(n6558), .ZN(n6530) );
  INV_X1 U3883 ( .A(n6459), .ZN(n6531) );
  INV_X1 U3884 ( .A(n6463), .ZN(n6537) );
  INV_X1 U3885 ( .A(n6568), .ZN(n6543) );
  INV_X1 U3886 ( .A(n5112), .ZN(n6563) );
  OAI211_X1 U3887 ( .C1(n6666), .C2(n4524), .A(n4522), .B(n6499), .ZN(n4552)
         );
  OR2_X1 U3888 ( .A1(n4917), .A2(n4916), .ZN(n6574) );
  NAND2_X1 U3889 ( .A1(n4092), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U3890 ( .A1(n5663), .A2(n6240), .ZN(n4225) );
  NOR2_X1 U3891 ( .A1(n5656), .A2(n4548), .ZN(n5238) );
  INV_X1 U3892 ( .A(n5663), .ZN(n5615) );
  NAND2_X1 U3893 ( .A1(n3002), .A2(n2972), .ZN(U2955) );
  OAI21_X1 U3894 ( .B1(n5697), .B2(n5779), .A(n3031), .ZN(U2960) );
  INV_X1 U3895 ( .A(n3032), .ZN(n3031) );
  OAI21_X1 U3896 ( .B1(n5880), .B2(n6316), .A(n3033), .ZN(n3032) );
  AOI21_X1 U3897 ( .B1(n6312), .B2(n5699), .A(n5698), .ZN(n3033) );
  INV_X1 U3898 ( .A(n2991), .ZN(n2990) );
  OAI21_X1 U3899 ( .B1(n5778), .B2(n5779), .A(n5776), .ZN(n2991) );
  OAI211_X1 U3900 ( .C1(n5845), .C2(n6351), .A(n3022), .B(n3020), .ZN(U2987)
         );
  OAI21_X1 U3901 ( .B1(n5837), .B2(n3021), .A(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n3020) );
  NOR2_X1 U3902 ( .A1(n5841), .A2(n3023), .ZN(n3022) );
  NOR2_X1 U3903 ( .A1(n5962), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3021)
         );
  OAI21_X1 U3904 ( .B1(n5665), .B2(n6351), .A(n3074), .ZN(U2988) );
  AND2_X1 U3905 ( .A1(n3100), .A2(n3075), .ZN(n3074) );
  AND2_X1 U3906 ( .A1(n3101), .A2(n5225), .ZN(n3100) );
  OR2_X1 U3907 ( .A1(n5311), .A2(n6434), .ZN(n3075) );
  AND2_X1 U3908 ( .A1(n5955), .A2(n2993), .ZN(n2992) );
  OR2_X1 U3909 ( .A1(n5958), .A2(n5957), .ZN(n2993) );
  AND2_X1 U3910 ( .A1(n3301), .A2(n3379), .ZN(n3552) );
  NAND2_X1 U3911 ( .A1(n5324), .A2(n5325), .ZN(n5313) );
  INV_X1 U3912 ( .A(n3963), .ZN(n5279) );
  NOR2_X1 U3913 ( .A1(n5452), .A2(n3040), .ZN(n5372) );
  AND2_X1 U3914 ( .A1(n3112), .A2(n4018), .ZN(n2967) );
  INV_X1 U3915 ( .A(n5270), .ZN(n3006) );
  AND2_X1 U3916 ( .A1(n3104), .A2(n3102), .ZN(n2968) );
  OR2_X1 U3917 ( .A1(n3080), .A2(n3079), .ZN(n2969) );
  INV_X1 U3918 ( .A(n3546), .ZN(n3119) );
  NAND2_X1 U3919 ( .A1(n5756), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n2970) );
  AND2_X1 U3920 ( .A1(n3067), .A2(n3123), .ZN(n2971) );
  NAND2_X1 U3921 ( .A1(n3027), .A2(n3463), .ZN(n4707) );
  INV_X1 U3922 ( .A(n4133), .ZN(n4173) );
  NOR2_X1 U3923 ( .A1(n3078), .A2(n3080), .ZN(n5466) );
  NAND2_X1 U3924 ( .A1(n5406), .A2(n4262), .ZN(n4263) );
  NAND2_X1 U3925 ( .A1(n3128), .A2(n3130), .ZN(n5829) );
  INV_X1 U3926 ( .A(n3113), .ZN(n5800) );
  NOR2_X1 U3927 ( .A1(n5436), .A2(n3091), .ZN(n5202) );
  NAND2_X1 U3928 ( .A1(n5604), .A2(n5603), .ZN(n5485) );
  NOR2_X1 U3929 ( .A1(n5334), .A2(n5335), .ZN(n5324) );
  INV_X1 U3930 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4033) );
  INV_X1 U3931 ( .A(n4107), .ZN(n3082) );
  AND2_X1 U3932 ( .A1(n3253), .A2(n4394), .ZN(n3281) );
  AND2_X1 U3933 ( .A1(n4106), .A2(n4105), .ZN(n2972) );
  AND2_X1 U3934 ( .A1(n6387), .A2(n4276), .ZN(n2973) );
  OR2_X1 U3935 ( .A1(n5781), .A2(n4026), .ZN(n2974) );
  AND2_X1 U3936 ( .A1(n4080), .A2(n4068), .ZN(n2975) );
  OR2_X1 U3937 ( .A1(n5436), .A2(n5435), .ZN(n3093) );
  NAND2_X1 U3938 ( .A1(n5406), .A2(n2982), .ZN(n3099) );
  INV_X1 U3939 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6579) );
  AND2_X1 U3940 ( .A1(n5756), .A2(n4024), .ZN(n2976) );
  INV_X1 U3941 ( .A(n4023), .ZN(n3125) );
  AND2_X1 U3942 ( .A1(n4012), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n2977)
         );
  OR2_X1 U3943 ( .A1(n5436), .A2(n3089), .ZN(n5201) );
  OR2_X1 U3944 ( .A1(n5781), .A2(n4015), .ZN(n2978) );
  AND2_X1 U3945 ( .A1(n3088), .A2(n3087), .ZN(n2979) );
  INV_X1 U3946 ( .A(n5830), .ZN(n3051) );
  AND2_X1 U3947 ( .A1(n3038), .A2(n3037), .ZN(n2980) );
  OR2_X1 U3948 ( .A1(n3083), .A2(n3082), .ZN(n2981) );
  NAND2_X1 U3949 ( .A1(n5481), .A2(n3109), .ZN(n5431) );
  AND2_X1 U3950 ( .A1(n5973), .A2(n5972), .ZN(n5481) );
  AND2_X1 U3951 ( .A1(n3097), .A2(n3096), .ZN(n2982) );
  INV_X1 U3952 ( .A(n5435), .ZN(n3092) );
  OR2_X1 U3953 ( .A1(n4701), .A2(n4795), .ZN(n4828) );
  INV_X1 U3954 ( .A(n4828), .ZN(n3103) );
  AND2_X1 U3955 ( .A1(n3959), .A2(n3958), .ZN(n4652) );
  AND2_X1 U3956 ( .A1(n5719), .A2(n5720), .ZN(n2983) );
  INV_X1 U3957 ( .A(n3010), .ZN(n5988) );
  NAND2_X1 U3958 ( .A1(n6432), .A2(n5982), .ZN(n3010) );
  AND2_X1 U3959 ( .A1(n5781), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n2984)
         );
  AND2_X1 U3960 ( .A1(n5781), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n2985)
         );
  AND2_X1 U3961 ( .A1(n5781), .A2(n5757), .ZN(n2986) );
  AND2_X1 U3962 ( .A1(n3109), .A2(n3108), .ZN(n2987) );
  AND2_X2 U3963 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3005) );
  XNOR2_X1 U3964 ( .A(n4414), .B(n4131), .ZN(n4377) );
  AND2_X1 U3965 ( .A1(n3001), .A2(n3000), .ZN(n2988) );
  OR2_X1 U3966 ( .A1(n4102), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6435) );
  INV_X1 U3967 ( .A(n6435), .ZN(n3009) );
  INV_X1 U3968 ( .A(n6654), .ZN(n6652) );
  NAND2_X1 U3969 ( .A1(n5777), .A2(n2990), .ZN(U2969) );
  NAND2_X1 U3970 ( .A1(n5956), .A2(n2992), .ZN(U3001) );
  OAI21_X2 U3971 ( .B1(n3966), .B2(n4060), .A(n3965), .ZN(n3967) );
  XNOR2_X2 U3972 ( .A(n3077), .B(n3404), .ZN(n3590) );
  NAND2_X1 U3973 ( .A1(n3422), .A2(n3421), .ZN(n4519) );
  NAND2_X1 U3974 ( .A1(n2994), .A2(n3968), .ZN(n6329) );
  OAI21_X1 U3975 ( .B1(n4652), .B2(n4653), .A(n2994), .ZN(n4654) );
  INV_X1 U3976 ( .A(n5766), .ZN(n5772) );
  NOR2_X1 U3977 ( .A1(n5783), .A2(n2986), .ZN(n5769) );
  NAND3_X1 U3978 ( .A1(n2996), .A2(n3043), .A3(n2967), .ZN(n5754) );
  INV_X1 U3979 ( .A(n4425), .ZN(n2999) );
  NAND2_X1 U3980 ( .A1(n6337), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3956)
         );
  INV_X1 U3981 ( .A(n3942), .ZN(n3000) );
  AND2_X2 U3982 ( .A1(n3005), .A2(n4402), .ZN(n3306) );
  AND2_X2 U3983 ( .A1(n3150), .A2(n3005), .ZN(n3341) );
  NOR2_X1 U3984 ( .A1(n4579), .A2(n3005), .ZN(n4586) );
  NOR2_X4 U3985 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4401) );
  NAND2_X1 U3986 ( .A1(n5804), .A2(n3623), .ZN(n3030) );
  NAND2_X1 U3987 ( .A1(n3030), .A2(n3029), .ZN(n5452) );
  NAND2_X1 U3988 ( .A1(n3708), .A2(n3038), .ZN(n5360) );
  NAND2_X1 U3989 ( .A1(n3303), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U3990 ( .A1(n3303), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U3991 ( .A1(n3303), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U3992 ( .A1(n3341), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3198) );
  AOI22_X1 U3993 ( .A1(n3341), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U3994 ( .A1(n3341), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U3995 ( .A1(n3390), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3168) );
  AND2_X2 U3996 ( .A1(n4406), .A2(n4578), .ZN(n3303) );
  INV_X1 U3997 ( .A(n3130), .ZN(n3042) );
  NAND3_X1 U3998 ( .A1(n3045), .A2(n3115), .A3(n3051), .ZN(n3044) );
  NAND3_X1 U3999 ( .A1(n2967), .A2(n5830), .A3(n3049), .ZN(n3048) );
  INV_X2 U4000 ( .A(n4013), .ZN(n5756) );
  NAND2_X1 U4001 ( .A1(n3265), .A2(n3551), .ZN(n3273) );
  AND2_X2 U4002 ( .A1(n3058), .A2(n4402), .ZN(n3390) );
  AND2_X2 U4003 ( .A1(n4406), .A2(n3058), .ZN(n3396) );
  AND2_X2 U4004 ( .A1(n3150), .A2(n3058), .ZN(n3342) );
  INV_X1 U4005 ( .A(n3065), .ZN(n3066) );
  NAND2_X1 U4006 ( .A1(n5756), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3065) );
  NAND2_X1 U4007 ( .A1(n3111), .A2(n3068), .ZN(n3067) );
  INV_X1 U4008 ( .A(n3111), .ZN(n5795) );
  AND2_X2 U4009 ( .A1(n4578), .A2(n4401), .ZN(n3244) );
  NOR2_X1 U4010 ( .A1(n3280), .A2(n3141), .ZN(n4248) );
  OAI21_X1 U4011 ( .B1(n3280), .B2(n4554), .A(n3403), .ZN(n3275) );
  NAND2_X1 U4012 ( .A1(n3269), .A2(n3270), .ZN(n3280) );
  XNOR2_X1 U4013 ( .A(n3590), .B(n3076), .ZN(n3955) );
  OAI22_X2 U4014 ( .A1(n4482), .A2(STATE2_REG_0__SCAN_IN), .B1(n3960), .B2(
        n3410), .ZN(n3077) );
  INV_X1 U4015 ( .A(n5452), .ZN(n3708) );
  NOR2_X1 U4016 ( .A1(n5334), .A2(n3083), .ZN(n5314) );
  INV_X1 U4017 ( .A(n3093), .ZN(n5437) );
  AND2_X2 U4018 ( .A1(n5406), .A2(n3094), .ZN(n5364) );
  INV_X1 U4019 ( .A(n3099), .ZN(n5376) );
  NAND2_X1 U4020 ( .A1(n5481), .A2(n2987), .ZN(n5417) );
  INV_X1 U4021 ( .A(n4455), .ZN(n4142) );
  NAND2_X1 U4022 ( .A1(n3110), .A2(n4131), .ZN(n4455) );
  NAND2_X1 U4023 ( .A1(n4414), .A2(n4901), .ZN(n3110) );
  NAND2_X1 U4024 ( .A1(n4014), .A2(n5831), .ZN(n5811) );
  NAND2_X1 U4025 ( .A1(n3119), .A2(n3548), .ZN(n3122) );
  NAND3_X1 U4026 ( .A1(n3301), .A2(n3379), .A3(n6579), .ZN(n3545) );
  NAND3_X1 U4027 ( .A1(n3301), .A2(n3379), .A3(n3121), .ZN(n3120) );
  NAND2_X1 U4028 ( .A1(n5138), .A2(n3126), .ZN(n3128) );
  INV_X1 U4029 ( .A(n5195), .ZN(n3127) );
  NAND2_X1 U4030 ( .A1(n5261), .A2(n3136), .ZN(n5265) );
  AND3_X1 U4031 ( .A1(n4710), .A2(n4709), .A3(n4708), .ZN(n4825) );
  NAND2_X1 U4032 ( .A1(n4142), .A2(n4141), .ZN(n4457) );
  NAND2_X1 U4033 ( .A1(n5250), .A2(n6332), .ZN(n4106) );
  NAND2_X1 U4034 ( .A1(n5364), .A2(n5349), .ZN(n5351) );
  CLKBUF_X1 U4035 ( .A(n5346), .Z(n5361) );
  NAND2_X1 U4036 ( .A1(n3377), .A2(n3376), .ZN(n3369) );
  OAI22_X1 U4037 ( .A1(n5666), .A2(n4030), .B1(n5703), .B2(n4029), .ZN(n4031)
         );
  MUX2_X1 U4038 ( .A(n5666), .B(n5667), .S(n5223), .Z(n5212) );
  OAI21_X1 U4039 ( .B1(n3611), .B2(n3610), .A(n3623), .ZN(n5804) );
  AND2_X2 U4040 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4402) );
  NAND2_X1 U4041 ( .A1(n5322), .A2(n4216), .ZN(n4219) );
  AND2_X1 U4042 ( .A1(n6043), .A2(n4519), .ZN(n4659) );
  OR2_X1 U4043 ( .A1(n6043), .A2(n4726), .ZN(n5033) );
  AND2_X1 U4044 ( .A1(n6243), .A2(n4548), .ZN(n6240) );
  INV_X2 U4045 ( .A(n6240), .ZN(n5609) );
  NAND2_X1 U4046 ( .A1(n4248), .A2(n4120), .ZN(n4255) );
  AND4_X1 U4047 ( .A1(n3198), .A2(n3197), .A3(n3196), .A4(n3195), .ZN(n3134)
         );
  AND2_X1 U4048 ( .A1(n4224), .A2(n4223), .ZN(n3135) );
  AND2_X1 U4049 ( .A1(n4417), .A2(n5223), .ZN(n3137) );
  AND3_X1 U4050 ( .A1(n3201), .A2(n3200), .A3(n3199), .ZN(n3138) );
  INV_X1 U4051 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4370) );
  AND2_X1 U4052 ( .A1(n3569), .A2(n3524), .ZN(n3140) );
  OR2_X1 U4053 ( .A1(n4036), .A2(n5270), .ZN(n3141) );
  NOR2_X1 U4054 ( .A1(n3366), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3142)
         );
  OR2_X1 U4055 ( .A1(n6598), .A2(n6497), .ZN(n5779) );
  AND3_X1 U4056 ( .A1(n3543), .A2(n3542), .A3(n3541), .ZN(n3143) );
  NOR2_X1 U4057 ( .A1(n2965), .A2(n3284), .ZN(n3192) );
  XNOR2_X1 U4058 ( .A(n4581), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4070)
         );
  AND2_X1 U4059 ( .A1(n5781), .A2(n5984), .ZN(n4019) );
  NAND2_X1 U4060 ( .A1(n5270), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4035) );
  NAND2_X1 U4061 ( .A1(n3266), .A2(n4244), .ZN(n3267) );
  OR2_X1 U4062 ( .A1(n3432), .A2(n3431), .ZN(n3986) );
  INV_X1 U4063 ( .A(n4019), .ZN(n4020) );
  INV_X1 U4064 ( .A(n4035), .ZN(n3272) );
  AND2_X1 U4065 ( .A1(n4708), .A2(n4826), .ZN(n3604) );
  OR2_X1 U4066 ( .A1(n3457), .A2(n3456), .ZN(n3997) );
  AOI22_X1 U4067 ( .A1(n4075), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4088), 
        .B2(n3997), .ZN(n3580) );
  NAND2_X1 U4068 ( .A1(n3324), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3178)
         );
  AND2_X1 U4069 ( .A1(n4370), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4084)
         );
  OR2_X1 U4070 ( .A1(n3843), .A2(n3842), .ZN(n3850) );
  INV_X1 U4071 ( .A(n3885), .ZN(n3884) );
  NOR2_X1 U4072 ( .A1(n3462), .A2(n3461), .ZN(n3463) );
  NAND2_X1 U4073 ( .A1(n3318), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3230) );
  INV_X1 U4074 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6791) );
  INV_X1 U4075 ( .A(n4084), .ZN(n4085) );
  NOR2_X1 U4076 ( .A1(n3137), .A2(n4215), .ZN(n4216) );
  AND2_X1 U4077 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5282), .ZN(n5456) );
  INV_X1 U4078 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6181) );
  AND2_X1 U4079 ( .A1(n4180), .A2(n4179), .ZN(n5972) );
  INV_X1 U4080 ( .A(n4173), .ZN(n4210) );
  INV_X1 U4081 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5472) );
  NOR2_X1 U4082 ( .A1(n6812), .A2(n3634), .ZN(n3651) );
  AND2_X1 U4083 ( .A1(n4707), .A2(n3523), .ZN(n4824) );
  INV_X1 U4084 ( .A(n3595), .ZN(n3460) );
  AND2_X1 U4085 ( .A1(n6575), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3936) );
  AND2_X1 U4086 ( .A1(n4267), .A2(n4250), .ZN(n4577) );
  AND2_X1 U4087 ( .A1(n3406), .A2(n4556), .ZN(n6065) );
  INV_X1 U4088 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4895) );
  NAND2_X1 U4089 ( .A1(n3547), .A2(n3546), .ZN(n3550) );
  AND2_X1 U4090 ( .A1(n4185), .A2(n4184), .ZN(n5464) );
  NOR2_X1 U4091 ( .A1(n3529), .A2(n6170), .ZN(n3606) );
  XNOR2_X1 U4092 ( .A(n4101), .B(n5290), .ZN(n5300) );
  INV_X1 U4093 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5535) );
  INV_X1 U4094 ( .A(n3556), .ZN(n3600) );
  INV_X1 U4095 ( .A(n4104), .ZN(n4105) );
  NAND2_X1 U4096 ( .A1(n3797), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3828)
         );
  NAND2_X1 U4097 ( .A1(n3691), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3738)
         );
  NAND2_X1 U4098 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n3651), .ZN(n3687)
         );
  NAND2_X1 U4099 ( .A1(n3477), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3529)
         );
  NOR2_X1 U4100 ( .A1(n4713), .A2(n4714), .ZN(n4792) );
  NOR2_X1 U4101 ( .A1(n3575), .A2(n5535), .ZN(n3582) );
  INV_X1 U4102 ( .A(n6395), .ZN(n5962) );
  NAND2_X1 U4103 ( .A1(n6349), .A2(n4268), .ZN(n5983) );
  INV_X1 U4104 ( .A(n4841), .ZN(n4834) );
  NAND2_X1 U4105 ( .A1(n4619), .A2(n5043), .ZN(n4872) );
  INV_X1 U4106 ( .A(n4996), .ZN(n4987) );
  INV_X1 U4107 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6811) );
  AND2_X1 U4108 ( .A1(n5552), .A2(n3552), .ZN(n5036) );
  INV_X1 U4109 ( .A(n5095), .ZN(n5130) );
  AND2_X1 U4110 ( .A1(n4487), .A2(n6562), .ZN(n4491) );
  INV_X1 U4111 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4889) );
  INV_X1 U4112 ( .A(n6456), .ZN(n6555) );
  INV_X1 U4113 ( .A(n6199), .ZN(n6190) );
  NOR2_X1 U4114 ( .A1(n5300), .A2(n5254), .ZN(n5255) );
  INV_X1 U4115 ( .A(n5608), .ZN(n6239) );
  INV_X2 U4116 ( .A(n6249), .ZN(n5656) );
  AND2_X1 U4117 ( .A1(n6249), .A2(n4473), .ZN(n6247) );
  INV_X1 U4118 ( .A(n6307), .ZN(n6301) );
  AND3_X1 U4119 ( .A1(n3673), .A2(n3672), .A3(n3671), .ZN(n5654) );
  NAND2_X1 U4120 ( .A1(n3582), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3586)
         );
  NAND2_X1 U4121 ( .A1(n3572), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3575)
         );
  INV_X1 U4122 ( .A(n4229), .ZN(n4230) );
  AND2_X1 U4123 ( .A1(n6036), .A2(n5941), .ZN(n5954) );
  NAND2_X1 U4124 ( .A1(n5983), .A2(n6014), .ZN(n6036) );
  NAND2_X1 U4125 ( .A1(n6354), .A2(n6392), .ZN(n6419) );
  INV_X1 U4126 ( .A(n6434), .ZN(n6422) );
  NAND2_X1 U4127 ( .A1(n6575), .A2(n4986), .ZN(n6497) );
  OAI211_X1 U4128 ( .C1(n6666), .C2(n4837), .A(n4624), .B(n6499), .ZN(n4648)
         );
  INV_X1 U4129 ( .A(n4993), .ZN(n5029) );
  AND2_X1 U4130 ( .A1(n4728), .A2(n4727), .ZN(n6461) );
  OAI21_X1 U4131 ( .B1(n4743), .B2(n4742), .A(n4741), .ZN(n4780) );
  AND2_X1 U4132 ( .A1(n6043), .A2(n4660), .ZN(n6055) );
  OAI21_X1 U4133 ( .B1(n6501), .B2(n6500), .A(n6499), .ZN(n6686) );
  INV_X1 U4134 ( .A(n6680), .ZN(n6539) );
  OR2_X1 U4135 ( .A1(n4926), .A2(n4492), .ZN(n5038) );
  OAI22_X1 U4136 ( .A1(n5094), .A2(n5093), .B1(n5092), .B2(n5091), .ZN(n5132)
         );
  INV_X1 U4137 ( .A(n5033), .ZN(n4497) );
  INV_X1 U4138 ( .A(n6565), .ZN(n4820) );
  NOR2_X1 U4139 ( .A1(n4526), .A2(n4926), .ZN(n6552) );
  NOR2_X1 U4140 ( .A1(n4706), .A2(n4926), .ZN(n6463) );
  INV_X1 U4141 ( .A(n4953), .ZN(n4982) );
  AND2_X1 U4142 ( .A1(n4659), .A2(n4738), .ZN(n4670) );
  INV_X1 U4143 ( .A(n4833), .ZN(n4874) );
  AND2_X1 U4144 ( .A1(n6579), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5252) );
  INV_X1 U4145 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6104) );
  INV_X1 U4146 ( .A(n6211), .ZN(n6184) );
  INV_X1 U4147 ( .A(n5558), .ZN(n6218) );
  NAND2_X1 U4148 ( .A1(n6243), .A2(n5611), .ZN(n5608) );
  NAND2_X1 U4149 ( .A1(n6287), .A2(n4471), .ZN(n6249) );
  OR2_X1 U4150 ( .A1(n4602), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6263) );
  INV_X1 U4151 ( .A(n6261), .ZN(n6278) );
  INV_X1 U4152 ( .A(n6305), .ZN(n6298) );
  OAI21_X1 U4153 ( .B1(n3092), .B2(n5453), .A(n3093), .ZN(n5753) );
  NAND2_X1 U4154 ( .A1(n5833), .A2(n4387), .ZN(n6345) );
  AND2_X1 U4155 ( .A1(n4281), .A2(n4280), .ZN(n4282) );
  INV_X1 U4156 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6444) );
  AOI22_X1 U4157 ( .A1(n4623), .A2(n4618), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4837), .ZN(n4651) );
  AOI211_X2 U4158 ( .C1(n4992), .C2(n4991), .A(n6060), .B(n4990), .ZN(n5032)
         );
  OR2_X1 U4159 ( .A1(n6043), .A2(n4725), .ZN(n6467) );
  NAND3_X1 U4160 ( .A1(n6055), .A2(n5043), .A3(n4738), .ZN(n5189) );
  AOI22_X1 U4161 ( .A1(n4736), .A2(n4742), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5153), .ZN(n4783) );
  AOI21_X1 U4162 ( .B1(n6500), .B2(STATE2_REG_2__SCAN_IN), .A(n6493), .ZN(
        n6683) );
  NAND2_X1 U4163 ( .A1(n5045), .A2(n5043), .ZN(n6099) );
  AOI211_X2 U4164 ( .C1(n5040), .C2(n5041), .A(n5039), .B(n5038), .ZN(n5080)
         );
  AOI21_X1 U4165 ( .B1(n5090), .B2(n5093), .A(n5089), .ZN(n5135) );
  NAND2_X1 U4166 ( .A1(n4497), .A2(n4922), .ZN(n6572) );
  NAND2_X1 U4167 ( .A1(n4670), .A2(n5043), .ZN(n4823) );
  INV_X1 U4168 ( .A(n6480), .ZN(n6517) );
  NAND2_X1 U4169 ( .A1(n4670), .A2(n5044), .ZN(n4985) );
  NAND2_X1 U4170 ( .A1(n4659), .A2(n4922), .ZN(n4953) );
  INV_X1 U4171 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n4986) );
  INV_X1 U4172 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6100) );
  INV_X1 U4173 ( .A(n6647), .ZN(n6645) );
  NAND2_X1 U4174 ( .A1(n4225), .A2(n3135), .ZN(U2829) );
  AOI22_X1 U4175 ( .A1(n3342), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3319), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3148) );
  INV_X1 U4176 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3144) );
  AND2_X2 U4177 ( .A1(n3151), .A2(n4401), .ZN(n3237) );
  AND2_X2 U4178 ( .A1(n4580), .A2(n3145), .ZN(n3343) );
  AOI22_X1 U4179 ( .A1(n3237), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U4180 ( .A1(n3390), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3146) );
  AND2_X2 U4181 ( .A1(n4406), .A2(n3151), .ZN(n3242) );
  AOI22_X1 U4182 ( .A1(n3348), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3155) );
  AND2_X2 U4183 ( .A1(n3151), .A2(n4402), .ZN(n3243) );
  AOI22_X1 U4184 ( .A1(n3396), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3243), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4185 ( .A1(n3244), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4186 ( .A1(n3318), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3325), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4187 ( .A1(n3348), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4188 ( .A1(n3342), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4189 ( .A1(n3396), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4190 ( .A1(n3341), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4191 ( .A1(n3319), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3243), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4192 ( .A1(n3242), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3325), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4193 ( .A1(n3390), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3162) );
  NAND2_X1 U4194 ( .A1(n2965), .A2(n3284), .ZN(n3216) );
  AOI22_X1 U4195 ( .A1(n3348), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3396), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U4196 ( .A1(n3319), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U4197 ( .A1(n3318), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3166) );
  NAND4_X1 U4198 ( .A1(n3169), .A2(n3168), .A3(n3167), .A4(n3166), .ZN(n3175)
         );
  AOI22_X1 U4199 ( .A1(n3242), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3243), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4200 ( .A1(n3342), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3325), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4201 ( .A1(n3237), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4202 ( .A1(n3341), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3170) );
  NAND4_X1 U4203 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3174)
         );
  OR2_X2 U4204 ( .A1(n3175), .A2(n3174), .ZN(n4548) );
  NAND2_X1 U4205 ( .A1(n3318), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3179) );
  NAND2_X1 U4206 ( .A1(n3244), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3177) );
  NAND2_X1 U4207 ( .A1(n3325), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U4208 ( .A1(n3237), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U4209 ( .A1(n3390), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3182)
         );
  NAND2_X1 U4210 ( .A1(n3343), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3181) );
  NAND2_X1 U4211 ( .A1(n3306), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3180)
         );
  NAND2_X1 U4212 ( .A1(n3342), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3187)
         );
  NAND2_X1 U4213 ( .A1(n3341), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3185)
         );
  NAND2_X1 U4214 ( .A1(n3319), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3184)
         );
  NAND2_X1 U4215 ( .A1(n3396), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3191) );
  NAND2_X1 U4216 ( .A1(n3348), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3190) );
  NAND2_X1 U4217 ( .A1(n3242), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U4218 ( .A1(n3243), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3188) );
  NAND2_X1 U4219 ( .A1(n3302), .A2(n3192), .ZN(n3193) );
  NAND2_X1 U4220 ( .A1(n3194), .A2(n3193), .ZN(n3291) );
  INV_X1 U4221 ( .A(n3291), .ZN(n3214) );
  AOI22_X1 U4222 ( .A1(n3348), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4223 ( .A1(n3390), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3196) );
  AOI22_X1 U4224 ( .A1(n3342), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3195) );
  BUF_X4 U4225 ( .A(n3242), .Z(n3916) );
  AOI22_X1 U4226 ( .A1(n3916), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3243), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3202) );
  AOI22_X1 U4227 ( .A1(n3319), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4228 ( .A1(n3306), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4229 ( .A1(n3396), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3325), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4230 ( .A1(n3348), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4231 ( .A1(n3396), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3243), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4232 ( .A1(n3244), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3204) );
  AOI22_X1 U4233 ( .A1(n3318), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3325), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3203) );
  NAND4_X1 U4234 ( .A1(n3206), .A2(n3205), .A3(n3204), .A4(n3203), .ZN(n3212)
         );
  AOI22_X1 U4235 ( .A1(n3341), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4236 ( .A1(n3237), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3208) );
  AOI22_X1 U4237 ( .A1(n3390), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3207) );
  NAND4_X1 U4238 ( .A1(n3210), .A2(n3209), .A3(n3208), .A4(n3207), .ZN(n3211)
         );
  OR2_X2 U4239 ( .A1(n3212), .A2(n3211), .ZN(n3283) );
  NAND2_X1 U4240 ( .A1(n4244), .A2(n3283), .ZN(n4111) );
  INV_X1 U4241 ( .A(n4111), .ZN(n3213) );
  NAND2_X1 U4242 ( .A1(n3214), .A2(n3213), .ZN(n4093) );
  INV_X1 U4243 ( .A(n4093), .ZN(n3257) );
  AND2_X1 U4244 ( .A1(n3302), .A2(n4548), .ZN(n3215) );
  AOI22_X1 U4245 ( .A1(n3342), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3319), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3219) );
  AOI22_X1 U4246 ( .A1(n3237), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4247 ( .A1(n3390), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3217) );
  NAND4_X1 U4248 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n3228)
         );
  AOI22_X1 U4249 ( .A1(n3348), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3242), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U4250 ( .A1(n3396), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4251 ( .A1(n3243), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U4252 ( .A1(n3244), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3224) );
  AOI22_X1 U4253 ( .A1(n3318), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3325), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3223) );
  NAND4_X1 U4254 ( .A1(n3226), .A2(n3225), .A3(n3224), .A4(n3223), .ZN(n3227)
         );
  OR2_X4 U4255 ( .A1(n3228), .A2(n3227), .ZN(n4554) );
  NAND2_X1 U4256 ( .A1(n3325), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4257 ( .A1(n3341), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3236)
         );
  NAND2_X1 U4258 ( .A1(n3342), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3235)
         );
  NAND2_X1 U4259 ( .A1(n3319), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3234)
         );
  NAND2_X1 U4260 ( .A1(n3306), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3233)
         );
  NAND2_X1 U4261 ( .A1(n3390), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3240)
         );
  NAND2_X1 U4262 ( .A1(n3237), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U4263 ( .A1(n3343), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3238) );
  AND4_X1 U4264 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(n3250)
         );
  NAND2_X1 U4265 ( .A1(n3242), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3248) );
  NAND2_X1 U4266 ( .A1(n3243), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3247) );
  NAND2_X1 U4267 ( .A1(n3244), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U4268 ( .A1(n3324), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3245)
         );
  AND4_X1 U4269 ( .A1(n3248), .A2(n3247), .A3(n3246), .A4(n3245), .ZN(n3249)
         );
  NAND4_X4 U4270 ( .A1(n3252), .A2(n3251), .A3(n3250), .A4(n3249), .ZN(n5270)
         );
  NAND2_X1 U4271 ( .A1(n4108), .A2(n3282), .ZN(n3253) );
  NAND2_X1 U4272 ( .A1(n3264), .A2(n4110), .ZN(n4394) );
  NAND2_X1 U4273 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n4286) );
  OAI21_X1 U4274 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_1__SCAN_IN), .A(
        n4286), .ZN(n4232) );
  INV_X1 U4275 ( .A(n4232), .ZN(n3254) );
  NAND3_X1 U4276 ( .A1(n3257), .A2(n3281), .A3(n3256), .ZN(n3258) );
  NAND2_X1 U4277 ( .A1(n3258), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3277) );
  OAI21_X1 U4278 ( .B1(n3284), .B2(n3271), .A(n4548), .ZN(n3263) );
  NAND2_X1 U4279 ( .A1(n3264), .A2(n4527), .ZN(n3268) );
  NAND2_X1 U4280 ( .A1(n3265), .A2(n3284), .ZN(n3266) );
  NAND2_X1 U4281 ( .A1(n3268), .A2(n3267), .ZN(n3269) );
  NAND2_X1 U4282 ( .A1(n4075), .A2(n4472), .ZN(n3274) );
  AND2_X1 U4283 ( .A1(n3275), .A2(n3274), .ZN(n3276) );
  NAND2_X1 U4284 ( .A1(n3380), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3279) );
  MUX2_X1 U4285 ( .A(n4092), .B(n4102), .S(n5152), .Z(n3278) );
  NAND2_X1 U4286 ( .A1(n3279), .A2(n3278), .ZN(n3300) );
  INV_X1 U4287 ( .A(n3300), .ZN(n3298) );
  NAND2_X1 U4288 ( .A1(n3280), .A2(n5530), .ZN(n4117) );
  NAND2_X1 U4289 ( .A1(n3271), .A2(n4548), .ZN(n3640) );
  INV_X1 U4290 ( .A(n3640), .ZN(n3286) );
  NOR2_X1 U4291 ( .A1(n3283), .A2(n4508), .ZN(n3285) );
  NAND3_X1 U4292 ( .A1(n3286), .A2(n4244), .A3(n3285), .ZN(n4590) );
  AND2_X1 U4293 ( .A1(n5231), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4300) );
  INV_X1 U4294 ( .A(n3283), .ZN(n3362) );
  NAND2_X1 U4295 ( .A1(n3362), .A2(n5270), .ZN(n4133) );
  NAND4_X1 U4296 ( .A1(n3287), .A2(n4590), .A3(n4300), .A4(n4133), .ZN(n3290)
         );
  AND2_X1 U4297 ( .A1(n3006), .A2(n4554), .ZN(n5544) );
  NAND2_X1 U4298 ( .A1(n5544), .A2(n4036), .ZN(n3289) );
  NAND2_X1 U4299 ( .A1(n4527), .A2(n5270), .ZN(n3288) );
  NAND2_X1 U4300 ( .A1(n3289), .A2(n3288), .ZN(n4112) );
  NOR2_X1 U4301 ( .A1(n3290), .A2(n4112), .ZN(n3296) );
  NAND2_X1 U4302 ( .A1(n4472), .A2(n3271), .ZN(n3293) );
  NAND2_X1 U4303 ( .A1(n3293), .A2(n3283), .ZN(n3294) );
  OAI21_X1 U4304 ( .B1(n3292), .B2(n3294), .A(n4554), .ZN(n3295) );
  NAND4_X1 U4305 ( .A1(n4117), .A2(n3281), .A3(n3296), .A4(n3295), .ZN(n3299)
         );
  INV_X1 U4306 ( .A(n3299), .ZN(n3297) );
  NAND2_X1 U4307 ( .A1(n3298), .A2(n3297), .ZN(n3301) );
  NAND2_X2 U4308 ( .A1(n3300), .A2(n3299), .ZN(n3379) );
  AOI22_X1 U4309 ( .A1(n3303), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4311 ( .A1(n3304), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4312 ( .A1(n3237), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4313 ( .A1(n3894), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3307) );
  NAND4_X1 U4314 ( .A1(n3310), .A2(n3309), .A3(n3308), .A4(n3307), .ZN(n3316)
         );
  AOI22_X1 U4315 ( .A1(n2966), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3317), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4316 ( .A1(n3895), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3243), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4317 ( .A1(n3244), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4318 ( .A1(n3917), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3311) );
  NAND4_X1 U4319 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3315)
         );
  INV_X1 U4320 ( .A(n3999), .ZN(n4009) );
  NAND2_X1 U4321 ( .A1(n4009), .A2(n4256), .ZN(n3332) );
  AOI22_X1 U4322 ( .A1(n3317), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3894), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4323 ( .A1(n3303), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4324 ( .A1(n3916), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3319), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4325 ( .A1(n3391), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3320) );
  NAND4_X1 U4326 ( .A1(n3323), .A2(n3322), .A3(n3321), .A4(n3320), .ZN(n3331)
         );
  BUF_X1 U4327 ( .A(n3348), .Z(n3872) );
  AOI22_X1 U4328 ( .A1(n3872), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3237), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4329 ( .A1(n3917), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3243), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4330 ( .A1(n2966), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3244), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3327) );
  AOI22_X1 U4331 ( .A1(n3918), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3326) );
  NAND4_X1 U4332 ( .A1(n3329), .A2(n3328), .A3(n3327), .A4(n3326), .ZN(n3330)
         );
  MUX2_X1 U4333 ( .A(n3339), .B(n3332), .S(n3944), .Z(n3333) );
  INV_X1 U4334 ( .A(n3333), .ZN(n3334) );
  NAND2_X1 U4335 ( .A1(n3334), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3546) );
  INV_X2 U4336 ( .A(n4067), .ZN(n4075) );
  NAND2_X1 U4337 ( .A1(n4075), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3338) );
  INV_X1 U4338 ( .A(n3944), .ZN(n3335) );
  OAI211_X1 U4339 ( .C1(n3335), .C2(n5270), .A(n3339), .B(
        STATE2_REG_0__SCAN_IN), .ZN(n3336) );
  INV_X1 U4340 ( .A(n3336), .ZN(n3337) );
  NAND2_X1 U4341 ( .A1(n3340), .A2(n4006), .ZN(n3372) );
  INV_X1 U4342 ( .A(n3372), .ZN(n3358) );
  NAND2_X1 U4343 ( .A1(n4075), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4344 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n2966), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4345 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3317), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4346 ( .A1(n3894), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4347 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n3911), .B1(n3918), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3344) );
  NAND4_X1 U4348 ( .A1(n3347), .A2(n3346), .A3(n3345), .A4(n3344), .ZN(n3354)
         );
  AOI22_X1 U4349 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n3304), .B1(n3895), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4350 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n3917), .B1(n4583), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4351 ( .A1(n3919), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4352 ( .A1(n3237), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3349) );
  NAND4_X1 U4353 ( .A1(n3352), .A2(n3351), .A3(n3350), .A4(n3349), .ZN(n3353)
         );
  NAND2_X1 U4354 ( .A1(n3403), .A2(n3940), .ZN(n3355) );
  OAI211_X1 U4355 ( .C1(n3999), .C2(n3410), .A(n3356), .B(n3355), .ZN(n3373)
         );
  INV_X1 U4356 ( .A(n3373), .ZN(n3357) );
  NAND2_X1 U4357 ( .A1(n3358), .A2(n3357), .ZN(n3559) );
  NOR2_X1 U4358 ( .A1(n4111), .A2(n5610), .ZN(n3360) );
  INV_X1 U4359 ( .A(n4108), .ZN(n3359) );
  NAND2_X1 U4360 ( .A1(n3360), .A2(n3359), .ZN(n4241) );
  INV_X1 U4361 ( .A(n4241), .ZN(n3361) );
  NAND2_X1 U4362 ( .A1(n3361), .A2(n5270), .ZN(n4301) );
  NAND2_X1 U4363 ( .A1(n4548), .A2(n4508), .ZN(n5239) );
  NOR2_X1 U4364 ( .A1(n5242), .A2(n5239), .ZN(n3363) );
  NAND2_X1 U4365 ( .A1(n3363), .A2(n4393), .ZN(n4259) );
  OAI211_X1 U4366 ( .C1(n3364), .C2(n4301), .A(n4255), .B(n4259), .ZN(n3365)
         );
  NAND2_X1 U4367 ( .A1(n3365), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3367) );
  XNOR2_X1 U4368 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5092) );
  OAI22_X1 U4369 ( .A1(n4102), .A2(n5092), .B1(n4092), .B2(n4889), .ZN(n3366)
         );
  AOI21_X1 U4370 ( .B1(n3380), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3366), 
        .ZN(n3368) );
  NAND2_X1 U4371 ( .A1(n3368), .A2(n3367), .ZN(n3376) );
  XNOR2_X2 U4372 ( .A(n3369), .B(n3379), .ZN(n6039) );
  INV_X1 U4373 ( .A(n3410), .ZN(n3370) );
  NAND2_X1 U4374 ( .A1(n3370), .A2(n3940), .ZN(n3371) );
  NAND2_X1 U4375 ( .A1(n3559), .A2(n3557), .ZN(n3375) );
  NAND2_X1 U4376 ( .A1(n3372), .A2(n3373), .ZN(n3374) );
  INV_X1 U4377 ( .A(n3376), .ZN(n3378) );
  INV_X1 U4378 ( .A(n4102), .ZN(n6667) );
  NAND2_X1 U4379 ( .A1(n3381), .A2(n4895), .ZN(n4720) );
  INV_X1 U4380 ( .A(n3381), .ZN(n3382) );
  NAND2_X1 U4381 ( .A1(n3382), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4382 ( .A1(n4720), .A2(n3383), .ZN(n4763) );
  NAND2_X1 U4383 ( .A1(n6667), .A2(n4763), .ZN(n3384) );
  OAI21_X1 U4384 ( .B1(n4092), .B2(n4895), .A(n3384), .ZN(n3385) );
  AOI21_X1 U4385 ( .B1(n3380), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3385), 
        .ZN(n3387) );
  INV_X1 U4386 ( .A(n3387), .ZN(n3386) );
  OR2_X1 U4387 ( .A1(n3388), .A2(n3386), .ZN(n3389) );
  NAND2_X1 U4388 ( .A1(n3388), .A2(n3386), .ZN(n3405) );
  NAND2_X1 U4389 ( .A1(n3389), .A2(n3405), .ZN(n4482) );
  AOI22_X1 U4390 ( .A1(n2966), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4391 ( .A1(n3317), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4392 ( .A1(n3910), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4393 ( .A1(n3894), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3392) );
  NAND4_X1 U4394 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3402)
         );
  AOI22_X1 U4395 ( .A1(n3304), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4396 ( .A1(n3917), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4397 ( .A1(n3911), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4398 ( .A1(n3919), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3397) );
  NAND4_X1 U4399 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3401)
         );
  AOI22_X1 U4400 ( .A1(n4075), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3403), 
        .B2(n3951), .ZN(n3404) );
  NAND2_X1 U4401 ( .A1(n3380), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3409) );
  NAND2_X1 U4402 ( .A1(n6500), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U4403 ( .A1(n6677), .A2(n6811), .ZN(n3406) );
  NAND3_X1 U4404 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4950) );
  INV_X1 U4405 ( .A(n4950), .ZN(n4524) );
  NAND2_X1 U4406 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4524), .ZN(n4556) );
  NOR2_X1 U4407 ( .A1(n4092), .A2(n6811), .ZN(n3407) );
  AOI21_X1 U4408 ( .B1(n6065), .B2(n6667), .A(n3407), .ZN(n3408) );
  AOI22_X1 U4409 ( .A1(n2966), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3317), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4410 ( .A1(n3894), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3413) );
  AOI22_X1 U4411 ( .A1(n3895), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4412 ( .A1(n3911), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3411) );
  NAND4_X1 U4413 ( .A1(n3414), .A2(n3413), .A3(n3412), .A4(n3411), .ZN(n3420)
         );
  AOI22_X1 U4414 ( .A1(n3917), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4415 ( .A1(n3909), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4416 ( .A1(n4583), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4417 ( .A1(n3304), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3415) );
  NAND4_X1 U4418 ( .A1(n3418), .A2(n3417), .A3(n3416), .A4(n3415), .ZN(n3419)
         );
  AOI22_X1 U4419 ( .A1(n4075), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4088), 
        .B2(n3970), .ZN(n3421) );
  NAND2_X1 U4420 ( .A1(n4075), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4421 ( .A1(n3304), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4422 ( .A1(n3917), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4423 ( .A1(n2966), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4424 ( .A1(n3920), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3423) );
  NAND4_X1 U4425 ( .A1(n3426), .A2(n3425), .A3(n3424), .A4(n3423), .ZN(n3432)
         );
  AOI22_X1 U4426 ( .A1(n3909), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4427 ( .A1(n3894), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4428 ( .A1(n4583), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4429 ( .A1(n3317), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3427) );
  NAND4_X1 U4430 ( .A1(n3430), .A2(n3429), .A3(n3428), .A4(n3427), .ZN(n3431)
         );
  NAND2_X1 U4431 ( .A1(n4088), .A2(n3986), .ZN(n3433) );
  NAND2_X1 U4432 ( .A1(n3434), .A2(n3433), .ZN(n3569) );
  NAND2_X1 U4433 ( .A1(n4075), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4434 ( .A1(n2966), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4435 ( .A1(n3317), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3437) );
  AOI22_X1 U4436 ( .A1(n3910), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3436) );
  AOI22_X1 U4437 ( .A1(n3894), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3435) );
  NAND4_X1 U4438 ( .A1(n3438), .A2(n3437), .A3(n3436), .A4(n3435), .ZN(n3444)
         );
  AOI22_X1 U4439 ( .A1(n3304), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4440 ( .A1(n3917), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3441) );
  INV_X1 U4441 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6825) );
  AOI22_X1 U4442 ( .A1(n3911), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4443 ( .A1(n3919), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3439) );
  NAND4_X1 U4444 ( .A1(n3442), .A2(n3441), .A3(n3440), .A4(n3439), .ZN(n3443)
         );
  NAND2_X1 U4445 ( .A1(n4088), .A2(n3987), .ZN(n3445) );
  NAND2_X1 U4446 ( .A1(n3446), .A2(n3445), .ZN(n3524) );
  AOI22_X1 U4447 ( .A1(n2966), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4448 ( .A1(n3317), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4449 ( .A1(n3910), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4450 ( .A1(n3894), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4451 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3457)
         );
  AOI22_X1 U4452 ( .A1(n3304), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4453 ( .A1(n3917), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4454 ( .A1(n3911), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4455 ( .A1(n3919), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3452) );
  NAND4_X1 U4456 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(n3456)
         );
  AOI22_X1 U4457 ( .A1(n4075), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4088), 
        .B2(n3999), .ZN(n3458) );
  NOR2_X2 U4458 ( .A1(n4508), .A2(n6575), .ZN(n3664) );
  AOI22_X1 U4459 ( .A1(n3720), .A2(EAX_REG_7__SCAN_IN), .B1(n3936), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3459) );
  XNOR2_X1 U4460 ( .A(n3586), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5517) );
  XNOR2_X1 U4461 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3529), .ZN(n6311)
         );
  AOI22_X1 U4462 ( .A1(n3920), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4463 ( .A1(n3304), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4464 ( .A1(n2966), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4465 ( .A1(n3919), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3464) );
  NAND4_X1 U4466 ( .A1(n3467), .A2(n3466), .A3(n3465), .A4(n3464), .ZN(n3473)
         );
  AOI22_X1 U4467 ( .A1(n3917), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4468 ( .A1(n3909), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4469 ( .A1(n3894), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4470 ( .A1(n3317), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3468) );
  NAND4_X1 U4471 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3472)
         );
  OR2_X1 U4472 ( .A1(n3473), .A2(n3472), .ZN(n3474) );
  AOI22_X1 U4473 ( .A1(n3664), .A2(n3474), .B1(n3936), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3476) );
  NAND2_X1 U4474 ( .A1(n3720), .A2(EAX_REG_11__SCAN_IN), .ZN(n3475) );
  OAI211_X1 U4475 ( .C1(n6311), .C2(n3908), .A(n3476), .B(n3475), .ZN(n6175)
         );
  XNOR2_X1 U4476 ( .A(n3477), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5825)
         );
  NAND2_X1 U4477 ( .A1(n5825), .A2(n5251), .ZN(n3492) );
  AOI22_X1 U4478 ( .A1(n3304), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4479 ( .A1(n3920), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4480 ( .A1(n3918), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4481 ( .A1(n3894), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3478) );
  NAND4_X1 U4482 ( .A1(n3481), .A2(n3480), .A3(n3479), .A4(n3478), .ZN(n3487)
         );
  AOI22_X1 U4483 ( .A1(n2966), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3317), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4484 ( .A1(n3917), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4485 ( .A1(n3895), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4486 ( .A1(n3910), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3482) );
  NAND4_X1 U4487 ( .A1(n3485), .A2(n3484), .A3(n3483), .A4(n3482), .ZN(n3486)
         );
  OAI21_X1 U4488 ( .B1(n3487), .B2(n3486), .A(n3664), .ZN(n3490) );
  NAND2_X1 U4489 ( .A1(n3720), .A2(EAX_REG_10__SCAN_IN), .ZN(n3489) );
  NAND2_X1 U4490 ( .A1(n3936), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3488)
         );
  AND3_X1 U4491 ( .A1(n3490), .A2(n3489), .A3(n3488), .ZN(n3491) );
  NAND2_X1 U4492 ( .A1(n3492), .A2(n3491), .ZN(n5144) );
  AOI22_X1 U4493 ( .A1(n3894), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4494 ( .A1(n3872), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4495 ( .A1(n3909), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4496 ( .A1(n3910), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3493) );
  NAND4_X1 U4497 ( .A1(n3496), .A2(n3495), .A3(n3494), .A4(n3493), .ZN(n3502)
         );
  AOI22_X1 U4498 ( .A1(n3917), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4499 ( .A1(n3317), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4500 ( .A1(n3919), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4501 ( .A1(n2966), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3497) );
  NAND4_X1 U4502 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3501)
         );
  OAI21_X1 U4503 ( .B1(n3502), .B2(n3501), .A(n3664), .ZN(n3507) );
  NAND2_X1 U4504 ( .A1(n3720), .A2(EAX_REG_8__SCAN_IN), .ZN(n3506) );
  XNOR2_X1 U4505 ( .A(n3503), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U4506 ( .A1(n5507), .A2(n5251), .ZN(n3505) );
  NAND2_X1 U4507 ( .A1(n3936), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3504)
         );
  NAND4_X1 U4508 ( .A1(n3507), .A2(n3506), .A3(n3505), .A4(n3504), .ZN(n4712)
         );
  XNOR2_X1 U4509 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3508), .ZN(n6188) );
  AOI22_X1 U4510 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3917), .B1(n3919), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4511 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n3895), .B1(n4583), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4512 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n3909), .B1(n3918), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4513 ( .A1(n3391), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3509) );
  NAND4_X1 U4514 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), .ZN(n3518)
         );
  AOI22_X1 U4515 ( .A1(n2966), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4516 ( .A1(n3894), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4517 ( .A1(n3317), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4518 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(n3304), .B1(n3889), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3513) );
  NAND4_X1 U4519 ( .A1(n3516), .A2(n3515), .A3(n3514), .A4(n3513), .ZN(n3517)
         );
  OAI21_X1 U4520 ( .B1(n3518), .B2(n3517), .A(n3664), .ZN(n3521) );
  NAND2_X1 U4521 ( .A1(n3720), .A2(EAX_REG_9__SCAN_IN), .ZN(n3520) );
  NAND2_X1 U4522 ( .A1(n3936), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3519)
         );
  AND3_X1 U4523 ( .A1(n3521), .A2(n3520), .A3(n3519), .ZN(n3522) );
  OAI21_X1 U4524 ( .B1(n6188), .B2(n3908), .A(n3522), .ZN(n4791) );
  AND4_X1 U4525 ( .A1(n6175), .A2(n5144), .A3(n4712), .A4(n4791), .ZN(n3523)
         );
  NAND2_X1 U4526 ( .A1(n3447), .A2(n3569), .ZN(n3525) );
  NAND2_X1 U4527 ( .A1(n3977), .A2(n3664), .ZN(n3528) );
  XNOR2_X1 U4528 ( .A(n3575), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5533) );
  INV_X1 U4529 ( .A(n3936), .ZN(n3669) );
  OAI22_X1 U4530 ( .A1(n5533), .A2(n3908), .B1(n3669), .B2(n5535), .ZN(n3526)
         );
  AOI21_X1 U4531 ( .B1(n3720), .B2(EAX_REG_5__SCAN_IN), .A(n3526), .ZN(n3527)
         );
  NAND2_X1 U4532 ( .A1(n3528), .A2(n3527), .ZN(n4708) );
  INV_X1 U4533 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3530) );
  XNOR2_X1 U4534 ( .A(n3606), .B(n3530), .ZN(n6162) );
  OR2_X1 U4535 ( .A1(n6162), .A2(n3908), .ZN(n3544) );
  AOI22_X1 U4536 ( .A1(n3317), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3917), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4537 ( .A1(n3895), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4538 ( .A1(n3894), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4539 ( .A1(n3910), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3531) );
  NAND4_X1 U4540 ( .A1(n3534), .A2(n3533), .A3(n3532), .A4(n3531), .ZN(n3540)
         );
  AOI22_X1 U4541 ( .A1(n2966), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4542 ( .A1(n3909), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4543 ( .A1(n4583), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4544 ( .A1(n3872), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3535) );
  NAND4_X1 U4545 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .ZN(n3539)
         );
  OAI21_X1 U4546 ( .B1(n3540), .B2(n3539), .A(n3664), .ZN(n3543) );
  NAND2_X1 U4547 ( .A1(n3720), .A2(EAX_REG_12__SCAN_IN), .ZN(n3542) );
  NAND2_X1 U4548 ( .A1(n3936), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3541)
         );
  NAND2_X1 U4549 ( .A1(n3544), .A2(n3143), .ZN(n4826) );
  NAND2_X1 U4550 ( .A1(n3545), .A2(n3548), .ZN(n3547) );
  AOI21_X1 U4551 ( .B1(n5043), .B2(n3551), .A(n6575), .ZN(n4384) );
  INV_X1 U4552 ( .A(n3664), .ZN(n3639) );
  AOI22_X1 U4553 ( .A1(n3720), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6575), .ZN(n3555) );
  INV_X1 U4554 ( .A(n5239), .ZN(n3553) );
  NAND2_X1 U4555 ( .A1(n3556), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3554) );
  OAI211_X1 U4556 ( .C1(n6490), .C2(n3639), .A(n3555), .B(n3554), .ZN(n4383)
         );
  MUX2_X1 U4557 ( .A(n3934), .B(n4384), .S(n4383), .Z(n4375) );
  INV_X1 U4558 ( .A(n3557), .ZN(n3558) );
  NAND2_X1 U4559 ( .A1(n4480), .A2(n3664), .ZN(n3561) );
  AOI22_X1 U4560 ( .A1(n3720), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6575), .ZN(n3560) );
  NAND2_X1 U4561 ( .A1(n4375), .A2(n4376), .ZN(n4374) );
  INV_X1 U4562 ( .A(n4374), .ZN(n3564) );
  OAI21_X1 U4563 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3595), .ZN(n6344) );
  AOI22_X1 U4564 ( .A1(n3936), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n3934), 
        .B2(n6344), .ZN(n3563) );
  NAND2_X1 U4565 ( .A1(n3720), .A2(EAX_REG_2__SCAN_IN), .ZN(n3562) );
  OAI211_X1 U4566 ( .C1(n3600), .C2(n5234), .A(n3563), .B(n3562), .ZN(n3566)
         );
  NAND2_X1 U4567 ( .A1(n3564), .A2(n3566), .ZN(n3565) );
  AOI21_X1 U4568 ( .B1(n6043), .B2(n3664), .A(n3936), .ZN(n4477) );
  NAND2_X1 U4569 ( .A1(n3565), .A2(n4477), .ZN(n3568) );
  INV_X1 U4570 ( .A(n3566), .ZN(n3567) );
  NAND2_X1 U4571 ( .A1(n4374), .A2(n3567), .ZN(n4476) );
  XNOR2_X1 U4572 ( .A(n3593), .B(n3569), .ZN(n3969) );
  NAND2_X1 U4573 ( .A1(n3969), .A2(n3664), .ZN(n3579) );
  NAND2_X1 U4574 ( .A1(n6575), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3571)
         );
  NAND2_X1 U4575 ( .A1(n3720), .A2(EAX_REG_4__SCAN_IN), .ZN(n3570) );
  OAI211_X1 U4576 ( .C1(n3600), .C2(n4370), .A(n3571), .B(n3570), .ZN(n3576)
         );
  INV_X1 U4577 ( .A(n3572), .ZN(n3597) );
  INV_X1 U4578 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3573) );
  NAND2_X1 U4579 ( .A1(n3597), .A2(n3573), .ZN(n3574) );
  NAND2_X1 U4580 ( .A1(n3575), .A2(n3574), .ZN(n6335) );
  MUX2_X1 U4581 ( .A(n3576), .B(n6335), .S(n3934), .Z(n3577) );
  INV_X1 U4582 ( .A(n3577), .ZN(n3578) );
  NAND2_X1 U4583 ( .A1(n3579), .A2(n3578), .ZN(n4606) );
  INV_X1 U4584 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3589) );
  NAND2_X1 U4585 ( .A1(n3581), .A2(n3580), .ZN(n3985) );
  NAND2_X1 U4586 ( .A1(n3985), .A2(n3664), .ZN(n3588) );
  INV_X1 U4587 ( .A(n3582), .ZN(n3584) );
  INV_X1 U4588 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3583) );
  NAND2_X1 U4589 ( .A1(n3584), .A2(n3583), .ZN(n3585) );
  NAND2_X1 U4590 ( .A1(n3586), .A2(n3585), .ZN(n6325) );
  AOI22_X1 U4591 ( .A1(n6325), .A2(n5251), .B1(n3936), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3587) );
  OAI211_X1 U4592 ( .C1(n3139), .C2(n3589), .A(n3588), .B(n3587), .ZN(n4699)
         );
  NAND2_X1 U4593 ( .A1(n3591), .A2(n3590), .ZN(n3592) );
  INV_X1 U4594 ( .A(n4519), .ZN(n4660) );
  NAND2_X1 U4595 ( .A1(n3592), .A2(n4660), .ZN(n3594) );
  INV_X1 U4596 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U4597 ( .A1(n5546), .A2(n3595), .ZN(n3596) );
  NAND2_X1 U4598 ( .A1(n3597), .A2(n3596), .ZN(n5547) );
  AOI22_X1 U4599 ( .A1(n5547), .A2(n3934), .B1(n3936), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3599) );
  NAND2_X1 U4600 ( .A1(n3720), .A2(EAX_REG_3__SCAN_IN), .ZN(n3598) );
  OAI211_X1 U4601 ( .C1(n3600), .C2(n4581), .A(n3599), .B(n3598), .ZN(n3601)
         );
  INV_X1 U4602 ( .A(n3601), .ZN(n3602) );
  NAND2_X1 U4603 ( .A1(n3603), .A2(n3602), .ZN(n4454) );
  NAND2_X1 U4604 ( .A1(n3720), .A2(EAX_REG_13__SCAN_IN), .ZN(n3609) );
  OAI21_X1 U4605 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3607), .A(n3634), 
        .ZN(n6155) );
  AOI22_X1 U4606 ( .A1(n5251), .A2(n6155), .B1(n3936), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3608) );
  NAND2_X1 U4607 ( .A1(n3609), .A2(n3608), .ZN(n3610) );
  AOI22_X1 U4608 ( .A1(n3317), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4609 ( .A1(n3917), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4610 ( .A1(n3304), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4611 ( .A1(n3911), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3612) );
  NAND4_X1 U4612 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3621)
         );
  AOI22_X1 U4613 ( .A1(n3894), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4614 ( .A1(n2966), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4615 ( .A1(n3895), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4616 ( .A1(n3391), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3616) );
  NAND4_X1 U4617 ( .A1(n3619), .A2(n3618), .A3(n3617), .A4(n3616), .ZN(n3620)
         );
  OR2_X1 U4618 ( .A1(n3621), .A2(n3620), .ZN(n3622) );
  NAND2_X1 U4619 ( .A1(n3664), .A2(n3622), .ZN(n5805) );
  AOI22_X1 U4620 ( .A1(n2966), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4621 ( .A1(n3872), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4622 ( .A1(n3919), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4623 ( .A1(n4583), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3624) );
  NAND4_X1 U4624 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3624), .ZN(n3633)
         );
  AOI22_X1 U4625 ( .A1(n3317), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3894), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4626 ( .A1(n3920), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4627 ( .A1(n3917), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4628 ( .A1(n3391), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3628) );
  NAND4_X1 U4629 ( .A1(n3631), .A2(n3630), .A3(n3629), .A4(n3628), .ZN(n3632)
         );
  NOR2_X1 U4630 ( .A1(n3633), .A2(n3632), .ZN(n3638) );
  INV_X1 U4631 ( .A(n3634), .ZN(n3635) );
  INV_X1 U4632 ( .A(n3651), .ZN(n3667) );
  OAI21_X1 U4633 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n3635), .A(n3667), 
        .ZN(n6136) );
  AOI22_X1 U4634 ( .A1(n5251), .A2(n6136), .B1(n3936), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4635 ( .A1(n3720), .A2(EAX_REG_14__SCAN_IN), .ZN(n3636) );
  OAI211_X1 U4636 ( .C1(n3639), .C2(n3638), .A(n3637), .B(n3636), .ZN(n5603)
         );
  AOI22_X1 U4637 ( .A1(n3920), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4638 ( .A1(n3872), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4639 ( .A1(n2966), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4640 ( .A1(n4583), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3641) );
  NAND4_X1 U4641 ( .A1(n3644), .A2(n3643), .A3(n3642), .A4(n3641), .ZN(n3650)
         );
  AOI22_X1 U4642 ( .A1(n3317), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4643 ( .A1(n3917), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4644 ( .A1(n3894), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4645 ( .A1(n3889), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3645) );
  NAND4_X1 U4646 ( .A1(n3648), .A2(n3647), .A3(n3646), .A4(n3645), .ZN(n3649)
         );
  OR2_X1 U4647 ( .A1(n3650), .A2(n3649), .ZN(n3655) );
  INV_X1 U4648 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4317) );
  INV_X1 U4649 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3652) );
  XNOR2_X1 U4650 ( .A(n3687), .B(n3652), .ZN(n5785) );
  AOI22_X1 U4651 ( .A1(n5785), .A2(n3934), .B1(PHYADDRPOINTER_REG_16__SCAN_IN), 
        .B2(n3936), .ZN(n3653) );
  OAI21_X1 U4652 ( .B1(n3139), .B2(n4317), .A(n3653), .ZN(n3654) );
  AOI21_X1 U4653 ( .B1(n3902), .B2(n3655), .A(n3654), .ZN(n5487) );
  AOI22_X1 U4654 ( .A1(n3895), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4655 ( .A1(n2966), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4656 ( .A1(n3920), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4657 ( .A1(n3894), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3656) );
  NAND4_X1 U4658 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(n3666)
         );
  AOI22_X1 U4659 ( .A1(n3872), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4660 ( .A1(n3317), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4661 ( .A1(n3919), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4662 ( .A1(n3917), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3660) );
  NAND4_X1 U4663 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3660), .ZN(n3665)
         );
  OAI21_X1 U4664 ( .B1(n3666), .B2(n3665), .A(n3664), .ZN(n3673) );
  NAND2_X1 U4665 ( .A1(n3720), .A2(EAX_REG_15__SCAN_IN), .ZN(n3672) );
  INV_X1 U4666 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U4667 ( .A1(n6757), .A2(n3667), .ZN(n3668) );
  AND2_X1 U4668 ( .A1(n3668), .A2(n3687), .ZN(n6127) );
  OAI22_X1 U4669 ( .A1(n6127), .A2(n3908), .B1(n6757), .B2(n3669), .ZN(n3670)
         );
  INV_X1 U4670 ( .A(n3670), .ZN(n3671) );
  AOI22_X1 U4671 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n3917), .B1(n3910), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4672 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n3872), .B1(n4583), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4673 ( .A1(n3909), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4674 ( .A1(n3317), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3675) );
  NAND4_X1 U4675 ( .A1(n3678), .A2(n3677), .A3(n3676), .A4(n3675), .ZN(n3684)
         );
  AOI22_X1 U4676 ( .A1(n2966), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4677 ( .A1(n3894), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4678 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n3895), .B1(n3918), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4679 ( .A1(n3920), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3679) );
  NAND4_X1 U4680 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(n3683)
         );
  NOR2_X1 U4681 ( .A1(n3684), .A2(n3683), .ZN(n3686) );
  AOI22_X1 U4682 ( .A1(n3720), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6575), .ZN(n3685) );
  OAI21_X1 U4683 ( .B1(n3932), .B2(n3686), .A(n3685), .ZN(n3689) );
  XNOR2_X1 U4684 ( .A(n3690), .B(n5472), .ZN(n5774) );
  MUX2_X1 U4685 ( .A(n3689), .B(n5774), .S(n3934), .Z(n5468) );
  INV_X1 U4686 ( .A(n3691), .ZN(n3692) );
  INV_X1 U4687 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U4688 ( .A1(n3692), .A2(n5762), .ZN(n3693) );
  AND2_X1 U4689 ( .A1(n3738), .A2(n3693), .ZN(n5760) );
  AOI22_X1 U4690 ( .A1(n3894), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4691 ( .A1(n3909), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4692 ( .A1(n3872), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4693 ( .A1(n3917), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3694) );
  NAND4_X1 U4694 ( .A1(n3697), .A2(n3696), .A3(n3695), .A4(n3694), .ZN(n3703)
         );
  AOI22_X1 U4695 ( .A1(n3317), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4696 ( .A1(n4583), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4697 ( .A1(n2966), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4698 ( .A1(n3911), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3698) );
  NAND4_X1 U4699 ( .A1(n3701), .A2(n3700), .A3(n3699), .A4(n3698), .ZN(n3702)
         );
  OR2_X1 U4700 ( .A1(n3703), .A2(n3702), .ZN(n3705) );
  INV_X1 U4701 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4321) );
  OAI22_X1 U4702 ( .A1(n3139), .A2(n4321), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5762), .ZN(n3704) );
  AOI21_X1 U4703 ( .B1(n3902), .B2(n3705), .A(n3704), .ZN(n3706) );
  MUX2_X1 U4704 ( .A(n5760), .B(n3706), .S(n3908), .Z(n5454) );
  AOI22_X1 U4705 ( .A1(n2966), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4706 ( .A1(n3317), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4707 ( .A1(n3910), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4708 ( .A1(n3894), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3709) );
  NAND4_X1 U4709 ( .A1(n3712), .A2(n3711), .A3(n3710), .A4(n3709), .ZN(n3718)
         );
  AOI22_X1 U4710 ( .A1(n3872), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4711 ( .A1(n3917), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4712 ( .A1(n3911), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4713 ( .A1(n3919), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3713) );
  NAND4_X1 U4714 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(n3717)
         );
  NOR2_X1 U4715 ( .A1(n3718), .A2(n3717), .ZN(n3722) );
  INV_X1 U4716 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5748) );
  AOI21_X1 U4717 ( .B1(n5748), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3719) );
  AOI21_X1 U4718 ( .B1(n3720), .B2(EAX_REG_19__SCAN_IN), .A(n3719), .ZN(n3721)
         );
  OAI21_X1 U4719 ( .B1(n3932), .B2(n3722), .A(n3721), .ZN(n3724) );
  XNOR2_X1 U4720 ( .A(n3738), .B(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5750)
         );
  NAND2_X1 U4721 ( .A1(n5750), .A2(n3934), .ZN(n3723) );
  NAND2_X1 U4722 ( .A1(n3724), .A2(n3723), .ZN(n5435) );
  AOI22_X1 U4723 ( .A1(n3317), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3728) );
  AOI22_X1 U4724 ( .A1(n3872), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4725 ( .A1(n3917), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4726 ( .A1(n3920), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3725) );
  NAND4_X1 U4727 ( .A1(n3728), .A2(n3727), .A3(n3726), .A4(n3725), .ZN(n3734)
         );
  AOI22_X1 U4728 ( .A1(n3894), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4729 ( .A1(n3909), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4730 ( .A1(n4583), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4731 ( .A1(n2966), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3729) );
  NAND4_X1 U4732 ( .A1(n3732), .A2(n3731), .A3(n3730), .A4(n3729), .ZN(n3733)
         );
  NOR2_X1 U4733 ( .A1(n3734), .A2(n3733), .ZN(n3736) );
  AOI22_X1 U4734 ( .A1(n3720), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6575), .ZN(n3735) );
  OAI21_X1 U4735 ( .B1(n3932), .B2(n3736), .A(n3735), .ZN(n3740) );
  INV_X1 U4736 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5740) );
  OAI21_X1 U4737 ( .B1(n3738), .B2(n5748), .A(n5740), .ZN(n3739) );
  NAND2_X1 U4738 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3737) );
  NAND2_X1 U4739 ( .A1(n3739), .A2(n3754), .ZN(n5739) );
  MUX2_X1 U4740 ( .A(n3740), .B(n5739), .S(n3934), .Z(n5421) );
  AOI22_X1 U4741 ( .A1(n2966), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4742 ( .A1(n3909), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4743 ( .A1(n3872), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3742) );
  AOI22_X1 U4744 ( .A1(n3910), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3741) );
  NAND4_X1 U4745 ( .A1(n3744), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(n3750)
         );
  AOI22_X1 U4746 ( .A1(n3917), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4747 ( .A1(n3317), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4748 ( .A1(n3918), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4749 ( .A1(n3894), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3745) );
  NAND4_X1 U4750 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3749)
         );
  NOR2_X1 U4751 ( .A1(n3750), .A2(n3749), .ZN(n3752) );
  AOI22_X1 U4752 ( .A1(n3720), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6575), .ZN(n3751) );
  OAI21_X1 U4753 ( .B1(n3932), .B2(n3752), .A(n3751), .ZN(n3756) );
  INV_X1 U4754 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6745) );
  NAND2_X1 U4755 ( .A1(n3754), .A2(n6745), .ZN(n3755) );
  NAND2_X1 U4756 ( .A1(n3769), .A2(n3755), .ZN(n5732) );
  MUX2_X1 U4757 ( .A(n3756), .B(n5732), .S(n3934), .Z(n5407) );
  AOI22_X1 U4758 ( .A1(n3872), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3894), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4759 ( .A1(n2966), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4760 ( .A1(n3917), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4761 ( .A1(n3918), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3757) );
  NAND4_X1 U4762 ( .A1(n3760), .A2(n3759), .A3(n3758), .A4(n3757), .ZN(n3766)
         );
  AOI22_X1 U4763 ( .A1(n3909), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4764 ( .A1(n3317), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4765 ( .A1(n3916), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4766 ( .A1(n3391), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3761) );
  NAND4_X1 U4767 ( .A1(n3764), .A2(n3763), .A3(n3762), .A4(n3761), .ZN(n3765)
         );
  NOR2_X1 U4768 ( .A1(n3766), .A2(n3765), .ZN(n3768) );
  AOI22_X1 U4769 ( .A1(n3720), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6575), .ZN(n3767) );
  OAI21_X1 U4770 ( .B1(n3932), .B2(n3768), .A(n3767), .ZN(n3771) );
  OR2_X2 U4771 ( .A1(n3769), .A2(n6791), .ZN(n3796) );
  NAND2_X1 U4772 ( .A1(n3769), .A2(n6791), .ZN(n3770) );
  NAND2_X1 U4773 ( .A1(n3796), .A2(n3770), .ZN(n5399) );
  MUX2_X1 U4774 ( .A(n3771), .B(n5399), .S(n3934), .Z(n5203) );
  AOI22_X1 U4775 ( .A1(n3304), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4776 ( .A1(n2966), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4777 ( .A1(n3894), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4778 ( .A1(n4583), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3773) );
  NAND4_X1 U4779 ( .A1(n3776), .A2(n3775), .A3(n3774), .A4(n3773), .ZN(n3782)
         );
  AOI22_X1 U4780 ( .A1(n3317), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4781 ( .A1(n3917), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4782 ( .A1(n3910), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4783 ( .A1(n3911), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3777) );
  NAND4_X1 U4784 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3781)
         );
  NOR2_X1 U4785 ( .A1(n3782), .A2(n3781), .ZN(n3809) );
  AOI22_X1 U4786 ( .A1(n3317), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3917), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4787 ( .A1(n3304), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4788 ( .A1(n2966), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4789 ( .A1(n3894), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3783) );
  NAND4_X1 U4790 ( .A1(n3786), .A2(n3785), .A3(n3784), .A4(n3783), .ZN(n3792)
         );
  AOI22_X1 U4791 ( .A1(n3919), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4792 ( .A1(n3909), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4793 ( .A1(n3918), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4794 ( .A1(n3910), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3787) );
  NAND4_X1 U4795 ( .A1(n3790), .A2(n3789), .A3(n3788), .A4(n3787), .ZN(n3791)
         );
  NOR2_X1 U4796 ( .A1(n3792), .A2(n3791), .ZN(n3808) );
  XOR2_X1 U4797 ( .A(n3809), .B(n3808), .Z(n3794) );
  INV_X1 U4798 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4324) );
  INV_X1 U4799 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5724) );
  OAI22_X1 U4800 ( .A1(n3139), .A2(n4324), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5724), .ZN(n3793) );
  AOI21_X1 U4801 ( .B1(n3902), .B2(n3794), .A(n3793), .ZN(n3795) );
  XNOR2_X1 U4802 ( .A(n3796), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5722)
         );
  MUX2_X1 U4803 ( .A(n3795), .B(n5722), .S(n3934), .Z(n5383) );
  XNOR2_X1 U4804 ( .A(n3828), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5717)
         );
  AOI22_X1 U4805 ( .A1(n2966), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4806 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n3317), .B1(n3909), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4807 ( .A1(n3910), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4808 ( .A1(n3894), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3798) );
  NAND4_X1 U4809 ( .A1(n3801), .A2(n3800), .A3(n3799), .A4(n3798), .ZN(n3807)
         );
  AOI22_X1 U4810 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n3872), .B1(n3895), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4811 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n3917), .B1(n4583), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4812 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(n3911), .B1(n3918), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4813 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n3919), .B1(n3889), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3802) );
  NAND4_X1 U4814 ( .A1(n3805), .A2(n3804), .A3(n3803), .A4(n3802), .ZN(n3806)
         );
  NOR2_X1 U4815 ( .A1(n3809), .A2(n3808), .ZN(n3824) );
  XOR2_X1 U4816 ( .A(n3823), .B(n3824), .Z(n3810) );
  NAND2_X1 U4817 ( .A1(n3810), .A2(n3902), .ZN(n3812) );
  AOI22_X1 U4818 ( .A1(n3720), .A2(EAX_REG_24__SCAN_IN), .B1(n3936), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3811) );
  OAI211_X1 U4819 ( .C1(n5717), .C2(n3908), .A(n3812), .B(n3811), .ZN(n5373)
         );
  AOI22_X1 U4820 ( .A1(n2966), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4821 ( .A1(n3317), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4822 ( .A1(n3910), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4823 ( .A1(n3894), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3813) );
  NAND4_X1 U4824 ( .A1(n3816), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(n3822)
         );
  AOI22_X1 U4825 ( .A1(n3304), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4826 ( .A1(n3917), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4827 ( .A1(n3911), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4828 ( .A1(n3919), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3817) );
  NAND4_X1 U4829 ( .A1(n3820), .A2(n3819), .A3(n3818), .A4(n3817), .ZN(n3821)
         );
  NOR2_X1 U4830 ( .A1(n3822), .A2(n3821), .ZN(n3845) );
  NAND2_X1 U4831 ( .A1(n3824), .A2(n3823), .ZN(n3844) );
  XOR2_X1 U4832 ( .A(n3845), .B(n3844), .Z(n3827) );
  INV_X1 U4833 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3825) );
  OAI22_X1 U4834 ( .A1(n3139), .A2(n3825), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5700), .ZN(n3826) );
  AOI21_X1 U4835 ( .B1(n3827), .B2(n3902), .A(n3826), .ZN(n3829) );
  INV_X1 U4836 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5713) );
  OR2_X2 U4837 ( .A1(n3828), .A2(n5713), .ZN(n3830) );
  XNOR2_X1 U4838 ( .A(n3830), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5702)
         );
  MUX2_X1 U4839 ( .A(n3829), .B(n5702), .S(n3934), .Z(n5362) );
  INV_X1 U4840 ( .A(n3831), .ZN(n3832) );
  INV_X1 U4841 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U4842 ( .A1(n3832), .A2(n5696), .ZN(n3833) );
  AOI22_X1 U4843 ( .A1(n2966), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4844 ( .A1(n3317), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4845 ( .A1(n3910), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4846 ( .A1(n3894), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3834) );
  NAND4_X1 U4847 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3843)
         );
  AOI22_X1 U4848 ( .A1(n3872), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4849 ( .A1(n3917), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4850 ( .A1(n3911), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4851 ( .A1(n3919), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3838) );
  NAND4_X1 U4852 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(n3842)
         );
  NOR2_X1 U4853 ( .A1(n3845), .A2(n3844), .ZN(n3851) );
  XOR2_X1 U4854 ( .A(n3850), .B(n3851), .Z(n3848) );
  INV_X1 U4855 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6282) );
  NOR2_X1 U4856 ( .A1(n6104), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3846)
         );
  OAI22_X1 U4857 ( .A1(n3139), .A2(n6282), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3846), .ZN(n3847) );
  AOI21_X1 U4858 ( .B1(n3848), .B2(n3902), .A(n3847), .ZN(n3849) );
  NAND2_X1 U4859 ( .A1(n5346), .A2(n5348), .ZN(n5334) );
  NAND2_X1 U4860 ( .A1(n3851), .A2(n3850), .ZN(n3866) );
  AOI22_X1 U4861 ( .A1(n2966), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3317), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4862 ( .A1(n3917), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3919), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4863 ( .A1(n3916), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4864 ( .A1(n3910), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3852) );
  NAND4_X1 U4865 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3861)
         );
  AOI22_X1 U4866 ( .A1(n3920), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4867 ( .A1(n3911), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4868 ( .A1(n3304), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4869 ( .A1(n3894), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3856) );
  NAND4_X1 U4870 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3860)
         );
  NOR2_X1 U4871 ( .A1(n3861), .A2(n3860), .ZN(n3867) );
  XOR2_X1 U4872 ( .A(n3866), .B(n3867), .Z(n3864) );
  INV_X1 U4873 ( .A(EAX_REG_27__SCAN_IN), .ZN(n3862) );
  INV_X1 U4874 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5688) );
  OAI22_X1 U4875 ( .A1(n3139), .A2(n3862), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5688), .ZN(n3863) );
  AOI21_X1 U4876 ( .B1(n3864), .B2(n3902), .A(n3863), .ZN(n3865) );
  XNOR2_X1 U4877 ( .A(n3881), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5686)
         );
  MUX2_X1 U4878 ( .A(n3865), .B(n5686), .S(n5251), .Z(n5335) );
  NOR2_X1 U4879 ( .A1(n3867), .A2(n3866), .ZN(n3888) );
  AOI22_X1 U4880 ( .A1(n2966), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4881 ( .A1(n3317), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4882 ( .A1(n3910), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4883 ( .A1(n3894), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3868) );
  NAND4_X1 U4884 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3878)
         );
  AOI22_X1 U4885 ( .A1(n3872), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4886 ( .A1(n3917), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4887 ( .A1(n3911), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4888 ( .A1(n3919), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3873) );
  NAND4_X1 U4889 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3877)
         );
  OR2_X1 U4890 ( .A1(n3878), .A2(n3877), .ZN(n3887) );
  XNOR2_X1 U4891 ( .A(n3888), .B(n3887), .ZN(n3880) );
  AOI22_X1 U4892 ( .A1(n3720), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6575), .ZN(n3879) );
  OAI21_X1 U4893 ( .B1(n3880), .B2(n3932), .A(n3879), .ZN(n3883) );
  NOR2_X1 U4894 ( .A1(n3881), .A2(n5688), .ZN(n3882) );
  INV_X1 U4895 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5327) );
  OR3_X2 U4896 ( .A1(n3881), .A2(n5688), .A3(n5327), .ZN(n3885) );
  OAI21_X1 U4897 ( .B1(n3882), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n3885), 
        .ZN(n5674) );
  MUX2_X1 U4898 ( .A(n3883), .B(n5674), .S(n5251), .Z(n5325) );
  INV_X1 U4899 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U4900 ( .A1(n3885), .A2(n6827), .ZN(n3886) );
  NAND2_X1 U4901 ( .A1(n4100), .A2(n3886), .ZN(n5670) );
  INV_X1 U4902 ( .A(EAX_REG_29__SCAN_IN), .ZN(n3906) );
  NAND2_X1 U4903 ( .A1(n3888), .A2(n3887), .ZN(n3927) );
  AOI22_X1 U4904 ( .A1(n2966), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4905 ( .A1(n3918), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4906 ( .A1(n3910), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4907 ( .A1(n3920), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4908 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3901)
         );
  AOI22_X1 U4909 ( .A1(n3317), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3894), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4910 ( .A1(n3304), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4911 ( .A1(n3917), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4912 ( .A1(n3919), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3911), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3896) );
  NAND4_X1 U4913 ( .A1(n3899), .A2(n3898), .A3(n3897), .A4(n3896), .ZN(n3900)
         );
  NOR2_X1 U4914 ( .A1(n3901), .A2(n3900), .ZN(n3928) );
  XOR2_X1 U4915 ( .A(n3927), .B(n3928), .Z(n3903) );
  NAND2_X1 U4916 ( .A1(n3903), .A2(n3902), .ZN(n3905) );
  OAI21_X1 U4917 ( .B1(n6104), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6575), 
        .ZN(n3904) );
  OAI211_X1 U4918 ( .C1(n3139), .C2(n3906), .A(n3905), .B(n3904), .ZN(n3907)
         );
  OAI21_X1 U4919 ( .B1(n3908), .B2(n5670), .A(n3907), .ZN(n5315) );
  AOI22_X1 U4920 ( .A1(n3317), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3909), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4921 ( .A1(n3894), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3910), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4922 ( .A1(n3911), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4923 ( .A1(n2966), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3912) );
  NAND4_X1 U4924 ( .A1(n3915), .A2(n3914), .A3(n3913), .A4(n3912), .ZN(n3926)
         );
  AOI22_X1 U4925 ( .A1(n3872), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3916), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4926 ( .A1(n3917), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4927 ( .A1(n3919), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3918), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4928 ( .A1(n3920), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3343), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3921) );
  NAND4_X1 U4929 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3925)
         );
  NOR2_X1 U4930 ( .A1(n3926), .A2(n3925), .ZN(n3930) );
  NOR2_X1 U4931 ( .A1(n3928), .A2(n3927), .ZN(n3929) );
  XOR2_X1 U4932 ( .A(n3930), .B(n3929), .Z(n3933) );
  AOI22_X1 U4933 ( .A1(n3720), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6575), .ZN(n3931) );
  OAI21_X1 U4934 ( .B1(n3933), .B2(n3932), .A(n3931), .ZN(n3935) );
  INV_X1 U4935 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4099) );
  XNOR2_X1 U4936 ( .A(n4100), .B(n4099), .ZN(n5661) );
  MUX2_X1 U4937 ( .A(n3935), .B(n5661), .S(n3934), .Z(n4107) );
  AOI22_X1 U4938 ( .A1(n3720), .A2(EAX_REG_31__SCAN_IN), .B1(n3936), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3937) );
  INV_X1 U4939 ( .A(n3937), .ZN(n3938) );
  NAND2_X1 U4940 ( .A1(n5252), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6598) );
  INV_X2 U4941 ( .A(n5779), .ZN(n6332) );
  NAND2_X1 U4942 ( .A1(n3944), .A2(n3940), .ZN(n3961) );
  OAI21_X1 U4943 ( .B1(n3940), .B2(n3944), .A(n3961), .ZN(n3941) );
  OAI211_X1 U4944 ( .C1(n3941), .C2(n3963), .A(n3213), .B(n5610), .ZN(n3942)
         );
  NAND2_X1 U4945 ( .A1(n3006), .A2(n3283), .ZN(n3952) );
  OAI21_X1 U4946 ( .B1(n3963), .B2(n3944), .A(n3952), .ZN(n3945) );
  INV_X1 U4947 ( .A(n3945), .ZN(n3946) );
  NAND2_X1 U4948 ( .A1(n4385), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3948)
         );
  INV_X1 U4949 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U4950 ( .A1(n3948), .A2(n6389), .ZN(n3949) );
  AND2_X1 U4951 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U4952 ( .A1(n4385), .A2(n6430), .ZN(n3950) );
  NAND2_X1 U4953 ( .A1(n3949), .A2(n3950), .ZN(n4425) );
  XNOR2_X1 U4954 ( .A(n3961), .B(n3951), .ZN(n3953) );
  OAI21_X1 U4955 ( .B1(n3953), .B2(n3963), .A(n3952), .ZN(n3954) );
  AOI21_X1 U4956 ( .B1(n3955), .B2(n4077), .A(n3954), .ZN(n6339) );
  NAND2_X1 U4957 ( .A1(n3956), .A2(n6339), .ZN(n3959) );
  INV_X1 U4958 ( .A(n6337), .ZN(n3957) );
  INV_X1 U4959 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U4960 ( .A1(n3957), .A2(n6388), .ZN(n3958) );
  NAND2_X1 U4961 ( .A1(n3961), .A2(n3960), .ZN(n3971) );
  INV_X1 U4962 ( .A(n3970), .ZN(n3962) );
  XNOR2_X1 U4963 ( .A(n3971), .B(n3962), .ZN(n3964) );
  NAND2_X1 U4964 ( .A1(n3964), .A2(n5279), .ZN(n3965) );
  INV_X1 U4965 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4266) );
  XNOR2_X1 U4966 ( .A(n3967), .B(n4266), .ZN(n4653) );
  NAND2_X1 U4967 ( .A1(n3967), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3968)
         );
  NAND2_X1 U4968 ( .A1(n3969), .A2(n4077), .ZN(n3974) );
  NAND2_X1 U4969 ( .A1(n3971), .A2(n3970), .ZN(n3989) );
  XNOR2_X1 U4970 ( .A(n3989), .B(n3986), .ZN(n3972) );
  NAND2_X1 U4971 ( .A1(n3972), .A2(n5279), .ZN(n3973) );
  NAND2_X1 U4972 ( .A1(n3974), .A2(n3973), .ZN(n3975) );
  INV_X1 U4973 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4265) );
  XNOR2_X1 U4974 ( .A(n3975), .B(n4265), .ZN(n6328) );
  NAND2_X1 U4975 ( .A1(n6329), .A2(n6328), .ZN(n6327) );
  NAND2_X1 U4976 ( .A1(n3975), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3976)
         );
  NAND2_X1 U4977 ( .A1(n6327), .A2(n3976), .ZN(n4880) );
  NAND2_X1 U4978 ( .A1(n3977), .A2(n4077), .ZN(n3982) );
  INV_X1 U4979 ( .A(n3986), .ZN(n3978) );
  OR2_X1 U4980 ( .A1(n3989), .A2(n3978), .ZN(n3979) );
  XNOR2_X1 U4981 ( .A(n3979), .B(n3987), .ZN(n3980) );
  NAND2_X1 U4982 ( .A1(n3980), .A2(n5279), .ZN(n3981) );
  NAND2_X1 U4983 ( .A1(n3982), .A2(n3981), .ZN(n3983) );
  INV_X1 U4984 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6742) );
  XNOR2_X1 U4985 ( .A(n3983), .B(n6742), .ZN(n4879) );
  NAND2_X1 U4986 ( .A1(n3983), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3984)
         );
  NAND3_X1 U4987 ( .A1(n4008), .A2(n4077), .A3(n3985), .ZN(n3992) );
  NAND2_X1 U4988 ( .A1(n3987), .A2(n3986), .ZN(n3988) );
  OR2_X1 U4989 ( .A1(n3989), .A2(n3988), .ZN(n3996) );
  XNOR2_X1 U4990 ( .A(n3996), .B(n3997), .ZN(n3990) );
  NAND2_X1 U4991 ( .A1(n3990), .A2(n5279), .ZN(n3991) );
  NAND2_X1 U4992 ( .A1(n3992), .A2(n3991), .ZN(n3993) );
  INV_X1 U4993 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6399) );
  XNOR2_X1 U4994 ( .A(n3993), .B(n6399), .ZN(n6319) );
  NAND2_X1 U4995 ( .A1(n3993), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3994)
         );
  NAND2_X1 U4996 ( .A1(n3995), .A2(n4077), .ZN(n4002) );
  INV_X1 U4997 ( .A(n3996), .ZN(n3998) );
  NAND2_X1 U4998 ( .A1(n3998), .A2(n3997), .ZN(n4010) );
  XNOR2_X1 U4999 ( .A(n4010), .B(n3999), .ZN(n4000) );
  NAND2_X1 U5000 ( .A1(n4000), .A2(n5279), .ZN(n4001) );
  NAND2_X1 U5001 ( .A1(n4002), .A2(n4001), .ZN(n4004) );
  INV_X1 U5002 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4003) );
  XNOR2_X1 U5003 ( .A(n4004), .B(n4003), .ZN(n5137) );
  NAND2_X1 U5004 ( .A1(n4004), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4005)
         );
  OR3_X1 U5005 ( .A1(n4010), .A2(n4009), .A3(n3963), .ZN(n4011) );
  NAND2_X1 U5006 ( .A1(n4013), .A2(n4011), .ZN(n4012) );
  INV_X1 U5007 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4155) );
  XNOR2_X1 U5008 ( .A(n4012), .B(n4155), .ZN(n5195) );
  INV_X1 U5009 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6367) );
  NAND2_X1 U5010 ( .A1(n5781), .A2(n6367), .ZN(n5830) );
  NAND2_X1 U5011 ( .A1(n5756), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5831)
         );
  INV_X1 U5012 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5812) );
  INV_X1 U5013 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6037) );
  INV_X1 U5014 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5810) );
  AND3_X1 U5015 ( .A1(n5812), .A2(n6037), .A3(n5810), .ZN(n4015) );
  NAND2_X1 U5016 ( .A1(n6025), .A2(n5810), .ZN(n5809) );
  NAND2_X1 U5017 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U5018 ( .A1(n6025), .A2(n5814), .ZN(n4016) );
  AND2_X1 U5019 ( .A1(n5809), .A2(n4016), .ZN(n4017) );
  XNOR2_X1 U5020 ( .A(n6025), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5801)
         );
  INV_X1 U5021 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U5022 ( .A1(n6025), .A2(n6005), .ZN(n4018) );
  INV_X1 U5023 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5984) );
  OAI21_X1 U5024 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5756), .ZN(n4021) );
  NAND4_X1 U5025 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(INSTADDRPOINTER_REG_15__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4022) );
  NAND2_X1 U5026 ( .A1(n6025), .A2(n4022), .ZN(n4023) );
  INV_X1 U5027 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5957) );
  INV_X1 U5028 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5940) );
  INV_X1 U5029 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5757) );
  NAND3_X1 U5030 ( .A1(n5957), .A2(n5940), .A3(n5757), .ZN(n4024) );
  INV_X1 U5031 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5720) );
  INV_X1 U5032 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4227) );
  INV_X1 U5033 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6734) );
  INV_X1 U5034 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5892) );
  NAND4_X1 U5035 ( .A1(n5720), .A2(n4227), .A3(n6734), .A4(n5892), .ZN(n4025)
         );
  INV_X1 U5036 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5938) );
  INV_X1 U5037 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U5038 ( .A1(n5938), .A2(n5736), .ZN(n5921) );
  NOR2_X1 U5039 ( .A1(n4025), .A2(n5921), .ZN(n4026) );
  AND2_X1 U5040 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4275) );
  AND2_X1 U5041 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5709) );
  AND2_X1 U5042 ( .A1(n4275), .A2(n5709), .ZN(n5900) );
  AND2_X1 U5043 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U5044 ( .A1(n5900), .A2(n5217), .ZN(n5221) );
  NAND2_X1 U5045 ( .A1(n6025), .A2(n5221), .ZN(n4027) );
  AND2_X1 U5046 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5213) );
  AND2_X1 U5047 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U5048 ( .A1(n5213), .A2(n5220), .ZN(n4028) );
  NAND2_X1 U5049 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4030) );
  XNOR2_X1 U5050 ( .A(n5781), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5704)
         );
  INV_X1 U5051 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U5052 ( .A1(n5756), .A2(n5877), .ZN(n5693) );
  NOR3_X1 U5053 ( .A1(n5693), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5211) );
  INV_X1 U5054 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5839) );
  INV_X1 U5055 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5223) );
  NAND3_X1 U5056 ( .A1(n5211), .A2(n5839), .A3(n5223), .ZN(n4029) );
  NAND2_X1 U5057 ( .A1(n4088), .A2(n4554), .ZN(n4032) );
  NAND2_X1 U5058 ( .A1(n4032), .A2(n5610), .ZN(n4039) );
  INV_X1 U5059 ( .A(n4039), .ZN(n4048) );
  XNOR2_X1 U5060 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4050) );
  NAND2_X1 U5061 ( .A1(n5152), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4049) );
  XNOR2_X1 U5062 ( .A(n4050), .B(n4049), .ZN(n4235) );
  INV_X1 U5063 ( .A(n4040), .ZN(n4047) );
  NAND2_X1 U5064 ( .A1(n4033), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4034) );
  AND2_X1 U5065 ( .A1(n4049), .A2(n4034), .ZN(n4042) );
  AOI21_X1 U5066 ( .B1(n4036), .B2(n4042), .A(n4035), .ZN(n4038) );
  NAND2_X1 U5067 ( .A1(n4120), .A2(n5610), .ZN(n4037) );
  NAND2_X1 U5068 ( .A1(n5242), .A2(n4037), .ZN(n4054) );
  OAI22_X1 U5069 ( .A1(n4040), .A2(n4039), .B1(n4038), .B2(n4054), .ZN(n4041)
         );
  OAI21_X1 U5070 ( .B1(n4089), .B2(n4235), .A(n4041), .ZN(n4045) );
  INV_X1 U5071 ( .A(n4088), .ZN(n4078) );
  INV_X1 U5072 ( .A(n4042), .ZN(n4043) );
  OAI21_X1 U5073 ( .B1(n4078), .B2(n4043), .A(n4089), .ZN(n4044) );
  NAND2_X1 U5074 ( .A1(n4045), .A2(n4044), .ZN(n4046) );
  OAI21_X1 U5075 ( .B1(n4048), .B2(n4047), .A(n4046), .ZN(n4065) );
  INV_X1 U5076 ( .A(n4049), .ZN(n4051) );
  NAND2_X1 U5077 ( .A1(n4051), .A2(n4050), .ZN(n4053) );
  NAND2_X1 U5078 ( .A1(n4889), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4052) );
  NAND2_X1 U5079 ( .A1(n4053), .A2(n4052), .ZN(n4057) );
  XNOR2_X1 U5080 ( .A(n5234), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4055)
         );
  XNOR2_X1 U5081 ( .A(n4057), .B(n4055), .ZN(n4234) );
  INV_X1 U5082 ( .A(n4054), .ZN(n4062) );
  NAND2_X1 U5083 ( .A1(n4088), .A2(n4234), .ZN(n4061) );
  OAI211_X1 U5084 ( .C1(n4234), .C2(n4067), .A(n4062), .B(n4061), .ZN(n4064)
         );
  INV_X1 U5085 ( .A(n4055), .ZN(n4056) );
  NAND2_X1 U5086 ( .A1(n4057), .A2(n4056), .ZN(n4059) );
  NAND2_X1 U5087 ( .A1(n4895), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4058) );
  XNOR2_X1 U5088 ( .A(n4073), .B(n4070), .ZN(n4233) );
  OAI22_X1 U5089 ( .A1(n4062), .A2(n4061), .B1(n4233), .B2(n4060), .ZN(n4063)
         );
  AOI21_X1 U5090 ( .B1(n4065), .B2(n4064), .A(n4063), .ZN(n4069) );
  INV_X1 U5091 ( .A(n4233), .ZN(n4066) );
  NOR2_X1 U5092 ( .A1(n4581), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4071)
         );
  NOR2_X1 U5093 ( .A1(n4370), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4074) );
  INV_X1 U5094 ( .A(n4076), .ZN(n4239) );
  AOI21_X1 U5095 ( .B1(n4078), .B2(n4077), .A(n4239), .ZN(n4079) );
  INV_X1 U5096 ( .A(n4081), .ZN(n4083) );
  AND2_X1 U5097 ( .A1(n4400), .A2(n3006), .ZN(n4094) );
  NAND2_X1 U5098 ( .A1(n4254), .A2(n3264), .ZN(n4914) );
  NAND2_X1 U5099 ( .A1(n4102), .A2(n6497), .ZN(n4095) );
  NAND2_X1 U5100 ( .A1(n4095), .A2(n6579), .ZN(n4096) );
  NAND2_X1 U5101 ( .A1(n6579), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4098) );
  NAND2_X1 U5102 ( .A1(n6104), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4097) );
  NAND2_X1 U5103 ( .A1(n4098), .A2(n4097), .ZN(n4387) );
  OR2_X2 U5104 ( .A1(n4100), .A2(n4099), .ZN(n4101) );
  INV_X1 U5105 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5290) );
  INV_X1 U5106 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6650) );
  NOR2_X1 U5107 ( .A1(n6435), .A2(n6650), .ZN(n5842) );
  AOI21_X1 U5108 ( .B1(n6336), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5842), 
        .ZN(n4103) );
  OAI21_X1 U5109 ( .B1(n6345), .B2(n5300), .A(n4103), .ZN(n4104) );
  NAND2_X1 U5110 ( .A1(n4108), .A2(n5270), .ZN(n4109) );
  MUX2_X1 U5111 ( .A(n3963), .B(n4109), .S(n4472), .Z(n4247) );
  AND2_X1 U5112 ( .A1(n5544), .A2(n4244), .ZN(n4365) );
  CLKBUF_X3 U5113 ( .A(n4132), .Z(n5418) );
  NAND2_X2 U5114 ( .A1(n4210), .A2(n5418), .ZN(n5262) );
  OAI21_X1 U5115 ( .B1(n4365), .B2(n5262), .A(n4111), .ZN(n4116) );
  INV_X1 U5116 ( .A(n4112), .ZN(n4115) );
  NAND2_X1 U5117 ( .A1(n3292), .A2(n4110), .ZN(n4114) );
  NAND2_X1 U5118 ( .A1(n5239), .A2(n4527), .ZN(n4113) );
  NAND3_X1 U5119 ( .A1(n4247), .A2(n4118), .A3(n4117), .ZN(n4397) );
  OAI21_X1 U5120 ( .B1(n5418), .B2(n5270), .A(n4590), .ZN(n4119) );
  NOR2_X1 U5121 ( .A1(n4400), .A2(n4120), .ZN(n4250) );
  NAND2_X1 U5122 ( .A1(n6581), .A2(n4577), .ZN(n4123) );
  INV_X1 U5123 ( .A(n4548), .ZN(n5611) );
  AND3_X1 U5124 ( .A1(n5611), .A2(n4256), .A3(n4508), .ZN(n4121) );
  NAND2_X1 U5125 ( .A1(n4393), .A2(n4121), .ZN(n4467) );
  NAND2_X2 U5126 ( .A1(n5270), .A2(n4554), .ZN(n4212) );
  NAND2_X1 U5127 ( .A1(n4123), .A2(n4122), .ZN(n4124) );
  NOR2_X4 U5128 ( .A1(n4132), .A2(n4212), .ZN(n4136) );
  INV_X1 U5129 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U5130 ( .A1(n4136), .A2(n4380), .ZN(n4128) );
  NAND2_X1 U5131 ( .A1(n4210), .A2(n6389), .ZN(n4126) );
  NAND2_X1 U5132 ( .A1(n4901), .A2(n4380), .ZN(n4125) );
  NAND3_X1 U5133 ( .A1(n4126), .A2(n5418), .A3(n4125), .ZN(n4127) );
  NAND2_X1 U5134 ( .A1(n4128), .A2(n4127), .ZN(n4131) );
  NAND2_X1 U5135 ( .A1(n4210), .A2(EBX_REG_0__SCAN_IN), .ZN(n4130) );
  INV_X1 U5136 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U5137 ( .A1(n5418), .A2(n6758), .ZN(n4129) );
  NAND2_X1 U5138 ( .A1(n4130), .A2(n4129), .ZN(n4414) );
  NAND2_X2 U5139 ( .A1(n4901), .A2(n5418), .ZN(n4208) );
  NAND2_X1 U5140 ( .A1(n5418), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4134)
         );
  OAI211_X1 U5141 ( .C1(n4212), .C2(EBX_REG_3__SCAN_IN), .A(n4210), .B(n4134), 
        .ZN(n4135) );
  OAI21_X1 U5142 ( .B1(n4208), .B2(EBX_REG_3__SCAN_IN), .A(n4135), .ZN(n4459)
         );
  INV_X1 U5143 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U5144 ( .A1(n4136), .A2(n6242), .ZN(n4140) );
  NAND2_X1 U5145 ( .A1(n4210), .A2(n6388), .ZN(n4138) );
  NAND2_X1 U5146 ( .A1(n4901), .A2(n6242), .ZN(n4137) );
  NAND3_X1 U5147 ( .A1(n4138), .A2(n4132), .A3(n4137), .ZN(n4139) );
  AND2_X1 U5148 ( .A1(n4140), .A2(n4139), .ZN(n4456) );
  MUX2_X1 U5149 ( .A(n4208), .B(n5418), .S(EBX_REG_5__SCAN_IN), .Z(n4143) );
  OAI21_X1 U5150 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5262), .A(n4143), 
        .ZN(n4144) );
  INV_X1 U5151 ( .A(n4144), .ZN(n4610) );
  MUX2_X1 U5152 ( .A(n4201), .B(n4210), .S(EBX_REG_4__SCAN_IN), .Z(n4147) );
  NAND2_X1 U5153 ( .A1(n4173), .A2(n5267), .ZN(n4175) );
  NAND2_X1 U5154 ( .A1(n5267), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4145)
         );
  AND2_X1 U5155 ( .A1(n4175), .A2(n4145), .ZN(n4146) );
  NAND2_X1 U5156 ( .A1(n4147), .A2(n4146), .ZN(n4611) );
  NAND2_X1 U5157 ( .A1(n4610), .A2(n4611), .ZN(n4148) );
  NOR2_X2 U5158 ( .A1(n4457), .A2(n4148), .ZN(n4703) );
  MUX2_X1 U5159 ( .A(n4201), .B(n4210), .S(EBX_REG_6__SCAN_IN), .Z(n4151) );
  NAND2_X1 U5160 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5267), .ZN(n4149)
         );
  AND2_X1 U5161 ( .A1(n4175), .A2(n4149), .ZN(n4150) );
  NAND2_X1 U5162 ( .A1(n4151), .A2(n4150), .ZN(n4702) );
  NAND2_X1 U5163 ( .A1(n4703), .A2(n4702), .ZN(n4701) );
  MUX2_X1 U5164 ( .A(n4208), .B(n5418), .S(EBX_REG_7__SCAN_IN), .Z(n4152) );
  OAI21_X1 U5165 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5262), .A(n4152), 
        .ZN(n4795) );
  MUX2_X1 U5166 ( .A(n4208), .B(n5418), .S(EBX_REG_9__SCAN_IN), .Z(n4153) );
  OAI21_X1 U5167 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5262), .A(n4153), 
        .ZN(n4154) );
  INV_X1 U5168 ( .A(n4154), .ZN(n4829) );
  INV_X1 U5169 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U5170 ( .A1(n4136), .A2(n5506), .ZN(n4159) );
  NAND2_X1 U5171 ( .A1(n4210), .A2(n4155), .ZN(n4157) );
  NAND2_X1 U5172 ( .A1(n4901), .A2(n5506), .ZN(n4156) );
  NAND3_X1 U5173 ( .A1(n4157), .A2(n5418), .A3(n4156), .ZN(n4158) );
  NAND2_X1 U5174 ( .A1(n4159), .A2(n4158), .ZN(n4830) );
  NAND2_X1 U5175 ( .A1(n4829), .A2(n4830), .ZN(n4160) );
  MUX2_X1 U5176 ( .A(n4201), .B(n4210), .S(EBX_REG_10__SCAN_IN), .Z(n4163) );
  NAND2_X1 U5177 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4212), .ZN(n4161) );
  AND2_X1 U5178 ( .A1(n4175), .A2(n4161), .ZN(n4162) );
  NAND2_X1 U5179 ( .A1(n4163), .A2(n4162), .ZN(n5191) );
  INV_X1 U5180 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U5181 ( .A1(n5257), .A2(n6237), .ZN(n4166) );
  NAND2_X1 U5182 ( .A1(n5418), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4164) );
  OAI211_X1 U5183 ( .C1(n5267), .C2(EBX_REG_11__SCAN_IN), .A(n4210), .B(n4164), 
        .ZN(n4165) );
  INV_X1 U5184 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6157) );
  MUX2_X1 U5185 ( .A(n4173), .B(n4136), .S(n6157), .Z(n4169) );
  NAND2_X1 U5186 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5267), .ZN(n4167) );
  NAND2_X1 U5187 ( .A1(n4175), .A2(n4167), .ZN(n4168) );
  NOR2_X1 U5188 ( .A1(n4169), .A2(n4168), .ZN(n5081) );
  NAND2_X1 U5189 ( .A1(n5418), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4170) );
  OAI211_X1 U5190 ( .C1(n5267), .C2(EBX_REG_13__SCAN_IN), .A(n4210), .B(n4170), 
        .ZN(n4171) );
  OAI21_X1 U5191 ( .B1(n4208), .B2(EBX_REG_13__SCAN_IN), .A(n4171), .ZN(n6001)
         );
  INV_X1 U5192 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4172) );
  MUX2_X1 U5193 ( .A(n4173), .B(n4136), .S(n4172), .Z(n4177) );
  NAND2_X1 U5194 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5267), .ZN(n4174) );
  NAND2_X1 U5195 ( .A1(n4175), .A2(n4174), .ZN(n4176) );
  NOR2_X1 U5196 ( .A1(n4177), .A2(n4176), .ZN(n5606) );
  INV_X1 U5197 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U5198 ( .A1(n5257), .A2(n6230), .ZN(n4180) );
  NAND2_X1 U5199 ( .A1(n5418), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4178) );
  OAI211_X1 U5200 ( .C1(n4212), .C2(EBX_REG_15__SCAN_IN), .A(n4210), .B(n4178), 
        .ZN(n4179) );
  MUX2_X1 U5201 ( .A(n4201), .B(n4210), .S(EBX_REG_16__SCAN_IN), .Z(n4182) );
  NAND2_X1 U5202 ( .A1(n5267), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4181) );
  NAND2_X1 U5203 ( .A1(n4182), .A2(n4181), .ZN(n5482) );
  INV_X1 U5204 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U5205 ( .A1(n5257), .A2(n5599), .ZN(n4185) );
  NAND2_X1 U5206 ( .A1(n5418), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4183) );
  OAI211_X1 U5207 ( .C1(n5267), .C2(EBX_REG_17__SCAN_IN), .A(n4210), .B(n4183), 
        .ZN(n4184) );
  INV_X1 U5208 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U5209 ( .A1(n4136), .A2(n5597), .ZN(n4188) );
  NAND2_X1 U5210 ( .A1(n4210), .A2(n5938), .ZN(n4186) );
  OAI211_X1 U5211 ( .C1(EBX_REG_19__SCAN_IN), .C2(n5267), .A(n4186), .B(n5418), 
        .ZN(n4187) );
  OR2_X1 U5212 ( .A1(n5262), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4189)
         );
  INV_X1 U5213 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U5214 ( .A1(n4901), .A2(n5598), .ZN(n5432) );
  OAI22_X1 U5215 ( .A1(n5262), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n5267), .ZN(n5419) );
  NAND2_X1 U5216 ( .A1(n5416), .A2(n5419), .ZN(n4191) );
  NAND2_X1 U5217 ( .A1(n4110), .A2(EBX_REG_20__SCAN_IN), .ZN(n4190) );
  OAI211_X1 U5218 ( .C1(n5416), .C2(n4110), .A(n4191), .B(n4190), .ZN(n4192)
         );
  MUX2_X1 U5219 ( .A(n4208), .B(n5418), .S(EBX_REG_21__SCAN_IN), .Z(n4193) );
  OAI21_X1 U5220 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5262), .A(n4193), 
        .ZN(n4194) );
  INV_X1 U5221 ( .A(n4194), .ZN(n5403) );
  AND2_X2 U5222 ( .A1(n5404), .A2(n5403), .ZN(n5406) );
  INV_X1 U5223 ( .A(EBX_REG_22__SCAN_IN), .ZN(n4195) );
  NAND2_X1 U5224 ( .A1(n4136), .A2(n4195), .ZN(n4198) );
  NAND2_X1 U5225 ( .A1(n4210), .A2(n6734), .ZN(n4196) );
  OAI211_X1 U5226 ( .C1(EBX_REG_22__SCAN_IN), .C2(n5267), .A(n4196), .B(n5418), 
        .ZN(n4197) );
  NAND2_X1 U5227 ( .A1(n4198), .A2(n4197), .ZN(n4262) );
  NAND2_X1 U5228 ( .A1(n4132), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4199) );
  OAI211_X1 U5229 ( .C1(n5267), .C2(EBX_REG_23__SCAN_IN), .A(n4133), .B(n4199), 
        .ZN(n4200) );
  OAI21_X1 U5230 ( .B1(n4208), .B2(EBX_REG_23__SCAN_IN), .A(n4200), .ZN(n5384)
         );
  MUX2_X1 U5231 ( .A(n4201), .B(n4210), .S(EBX_REG_24__SCAN_IN), .Z(n4203) );
  NAND2_X1 U5232 ( .A1(n5267), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4202) );
  MUX2_X1 U5233 ( .A(n4208), .B(n5418), .S(EBX_REG_25__SCAN_IN), .Z(n4204) );
  OAI21_X1 U5234 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5262), .A(n4204), 
        .ZN(n5365) );
  INV_X1 U5235 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6714) );
  NAND2_X1 U5236 ( .A1(n4136), .A2(n6714), .ZN(n4207) );
  NAND2_X1 U5237 ( .A1(n4210), .A2(n5877), .ZN(n4205) );
  OAI211_X1 U5238 ( .C1(EBX_REG_26__SCAN_IN), .C2(n5267), .A(n4205), .B(n4132), 
        .ZN(n4206) );
  NAND2_X1 U5239 ( .A1(n4207), .A2(n4206), .ZN(n5349) );
  MUX2_X1 U5240 ( .A(n4208), .B(n5418), .S(EBX_REG_27__SCAN_IN), .Z(n4209) );
  OAI21_X1 U5241 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5262), .A(n4209), 
        .ZN(n5336) );
  OR2_X2 U5242 ( .A1(n5351), .A2(n5336), .ZN(n5338) );
  INV_X1 U5243 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U5244 ( .A1(n4136), .A2(n5588), .ZN(n4214) );
  INV_X1 U5245 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U5246 ( .A1(n4210), .A2(n5678), .ZN(n4211) );
  OAI211_X1 U5247 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4212), .A(n4211), .B(n5418), 
        .ZN(n4213) );
  AND2_X1 U5248 ( .A1(n4214), .A2(n4213), .ZN(n5321) );
  NOR2_X4 U5249 ( .A1(n5338), .A2(n5321), .ZN(n5322) );
  INV_X1 U5250 ( .A(n5262), .ZN(n4417) );
  INV_X1 U5251 ( .A(n4219), .ZN(n4218) );
  INV_X1 U5252 ( .A(n5322), .ZN(n5260) );
  NAND2_X1 U5253 ( .A1(n4219), .A2(n4132), .ZN(n5261) );
  AOI22_X1 U5254 ( .A1(n5262), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5267), .ZN(n5258) );
  INV_X1 U5255 ( .A(n5258), .ZN(n4217) );
  OAI211_X1 U5256 ( .C1(n4218), .C2(n5260), .A(n5261), .B(n4217), .ZN(n4221)
         );
  OAI211_X1 U5257 ( .C1(n5322), .C2(n5418), .A(n4219), .B(n5258), .ZN(n4220)
         );
  NAND2_X1 U5258 ( .A1(n4221), .A2(n4220), .ZN(n5311) );
  INV_X1 U5259 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4222) );
  OR2_X1 U5260 ( .A1(n6243), .A2(n4222), .ZN(n4223) );
  XNOR2_X1 U5261 ( .A(n5781), .B(n5938), .ZN(n5747) );
  NOR2_X1 U5262 ( .A1(n5756), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4226)
         );
  XNOR2_X1 U5263 ( .A(n6025), .B(n4227), .ZN(n5729) );
  NOR2_X1 U5264 ( .A1(n5781), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5719)
         );
  AOI21_X1 U5265 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5781), .A(n5719), 
        .ZN(n4229) );
  OR2_X1 U5266 ( .A1(n4232), .A2(STATE_REG_0__SCAN_IN), .ZN(n4357) );
  NAND2_X1 U5267 ( .A1(n4554), .A2(n4357), .ZN(n4240) );
  NAND3_X1 U5268 ( .A1(n4235), .A2(n4234), .A3(n4233), .ZN(n4236) );
  NAND2_X1 U5269 ( .A1(n4237), .A2(n4236), .ZN(n4238) );
  NOR2_X1 U5270 ( .A1(n4910), .A2(READY_N), .ZN(n4361) );
  NAND2_X1 U5271 ( .A1(n4240), .A2(n4361), .ZN(n4246) );
  INV_X1 U5272 ( .A(READY_N), .ZN(n4884) );
  OAI21_X1 U5273 ( .B1(n4554), .B2(n5269), .A(n4884), .ZN(n4356) );
  OAI211_X1 U5274 ( .C1(n4241), .C2(n4356), .A(n5270), .B(n5239), .ZN(n4242)
         );
  INV_X1 U5275 ( .A(n4242), .ZN(n4243) );
  OR2_X1 U5276 ( .A1(n6581), .A2(n4243), .ZN(n4245) );
  MUX2_X1 U5277 ( .A(n4246), .B(n4245), .S(n4244), .Z(n4252) );
  NAND2_X1 U5278 ( .A1(n4254), .A2(n4247), .ZN(n4249) );
  INV_X1 U5279 ( .A(n4911), .ZN(n4302) );
  AOI21_X1 U5280 ( .B1(n6581), .B2(n4250), .A(n4364), .ZN(n4251) );
  NAND2_X1 U5281 ( .A1(n4252), .A2(n4251), .ZN(n4253) );
  NAND2_X1 U5282 ( .A1(n4254), .A2(n5530), .ZN(n4575) );
  NAND2_X1 U5283 ( .A1(n4914), .A2(n4575), .ZN(n4907) );
  INV_X1 U5284 ( .A(n4255), .ZN(n4565) );
  OAI22_X1 U5285 ( .A1(n4241), .A2(n4212), .B1(n4256), .B2(n4259), .ZN(n4257)
         );
  NOR3_X1 U5286 ( .A1(n4907), .A2(n4565), .A3(n4257), .ZN(n4258) );
  OAI21_X1 U5287 ( .B1(n4259), .B2(n3271), .A(n4919), .ZN(n4260) );
  INV_X1 U5288 ( .A(n4260), .ZN(n4261) );
  OR2_X1 U5289 ( .A1(n5406), .A2(n4262), .ZN(n4264) );
  AND2_X1 U5290 ( .A1(n4264), .A2(n4263), .ZN(n5593) );
  INV_X1 U5291 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6635) );
  NOR2_X1 U5292 ( .A1(n6435), .A2(n6635), .ZN(n5206) );
  NOR2_X1 U5293 ( .A1(n4266), .A2(n4265), .ZN(n6401) );
  INV_X1 U5294 ( .A(n6401), .ZN(n6415) );
  NOR3_X1 U5295 ( .A1(n6742), .A2(n6399), .A3(n6415), .ZN(n6355) );
  AOI21_X1 U5296 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6429) );
  INV_X1 U5297 ( .A(n4577), .ZN(n4909) );
  NAND2_X1 U5298 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U5299 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6356) );
  NOR2_X1 U5300 ( .A1(n6369), .A2(n6356), .ZN(n4268) );
  NAND2_X1 U5301 ( .A1(n4911), .A2(n4554), .ZN(n4592) );
  INV_X1 U5302 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U5303 ( .A1(n5986), .A2(n4416), .ZN(n4426) );
  AND3_X1 U5304 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6355), .ZN(n6347) );
  NAND2_X1 U5305 ( .A1(n6347), .A2(n4268), .ZN(n5959) );
  INV_X1 U5306 ( .A(n5959), .ZN(n4269) );
  NAND2_X1 U5307 ( .A1(n6428), .A2(n4269), .ZN(n6014) );
  NAND2_X1 U5308 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U5309 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4270) );
  NOR2_X1 U5310 ( .A1(n6015), .A2(n4270), .ZN(n5965) );
  AND2_X1 U5311 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4271) );
  AND2_X1 U5312 ( .A1(n5965), .A2(n4271), .ZN(n5941) );
  AND2_X1 U5313 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4272) );
  AND4_X1 U5314 ( .A1(n5935), .A2(n4275), .A3(INSTADDRPOINTER_REG_21__SCAN_IN), 
        .A4(n6734), .ZN(n4273) );
  AOI211_X1 U5315 ( .C1(n6422), .C2(n5593), .A(n5206), .B(n4273), .ZN(n4281)
         );
  INV_X1 U5316 ( .A(n4275), .ZN(n5922) );
  NOR3_X1 U5317 ( .A1(n5902), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n5922), 
        .ZN(n5911) );
  NAND2_X1 U5318 ( .A1(n6391), .A2(n6432), .ZN(n6346) );
  NAND2_X1 U5319 ( .A1(n5983), .A2(n6346), .ZN(n5961) );
  NAND3_X1 U5320 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n4275), .ZN(n4276) );
  INV_X1 U5321 ( .A(n5941), .ZN(n4277) );
  OAI21_X1 U5322 ( .B1(n4276), .B2(n4277), .A(n6346), .ZN(n4279) );
  OR2_X1 U5323 ( .A1(n4277), .A2(n5959), .ZN(n4278) );
  NAND2_X1 U5324 ( .A1(n6387), .A2(n4278), .ZN(n5917) );
  INV_X1 U5325 ( .A(n5216), .ZN(n5913) );
  OAI21_X1 U5326 ( .B1(n5911), .B2(n5913), .A(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n4280) );
  OAI21_X1 U5327 ( .B1(n5210), .B2(n6351), .A(n4282), .ZN(U2996) );
  NAND2_X1 U5328 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n4285) );
  INV_X1 U5329 ( .A(n4285), .ZN(n4283) );
  AND2_X1 U5330 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n4295) );
  NAND2_X1 U5331 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4288) );
  OAI21_X1 U5332 ( .B1(n4283), .B2(n4295), .A(n4288), .ZN(n4284) );
  OAI211_X1 U5333 ( .C1(n4884), .C2(n6100), .A(n4284), .B(n4357), .ZN(U3182)
         );
  AOI22_X1 U5334 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n4298) );
  INV_X1 U5335 ( .A(n4298), .ZN(n4292) );
  INV_X1 U5336 ( .A(n4286), .ZN(n4299) );
  NOR3_X1 U5337 ( .A1(NA_N), .A2(n4884), .A3(n4285), .ZN(n4291) );
  INV_X1 U5338 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6601) );
  INV_X1 U5339 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6101) );
  OAI211_X1 U5340 ( .C1(NA_N), .C2(n6601), .A(n4286), .B(n6101), .ZN(n4296) );
  NOR2_X1 U5341 ( .A1(NA_N), .A2(n4884), .ZN(n4287) );
  OAI21_X1 U5342 ( .B1(n4287), .B2(n6100), .A(HOLD), .ZN(n4289) );
  OAI211_X1 U5343 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n4289), .A(
        STATE_REG_0__SCAN_IN), .B(n4288), .ZN(n4290) );
  AOI222_X1 U5344 ( .A1(n4292), .A2(n4299), .B1(STATE_REG_1__SCAN_IN), .B2(
        n4291), .C1(n4296), .C2(n4290), .ZN(n4293) );
  INV_X1 U5345 ( .A(n4293), .ZN(U3183) );
  INV_X1 U5346 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4294) );
  NOR2_X2 U5347 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6100), .ZN(n6675) );
  INV_X2 U5348 ( .A(n6675), .ZN(n6663) );
  OAI21_X1 U5349 ( .B1(n4295), .B2(n4294), .A(n6663), .ZN(n4297) );
  OAI211_X1 U5350 ( .C1(n4299), .C2(n4298), .A(n4297), .B(n4296), .ZN(U3181)
         );
  INV_X1 U5351 ( .A(n4300), .ZN(n6588) );
  INV_X1 U5352 ( .A(n6581), .ZN(n4304) );
  OAI21_X1 U5353 ( .B1(n4302), .B2(n4910), .A(n4301), .ZN(n4303) );
  OAI21_X1 U5354 ( .B1(n4304), .B2(n5530), .A(n4303), .ZN(n4903) );
  OAI21_X1 U5355 ( .B1(n4903), .B2(n6587), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4305) );
  OAI21_X1 U5356 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6588), .A(n4305), .ZN(
        U2790) );
  INV_X1 U5357 ( .A(n4910), .ZN(n4306) );
  NAND3_X1 U5358 ( .A1(n4911), .A2(n4468), .A3(n4306), .ZN(n5243) );
  INV_X1 U5359 ( .A(n5243), .ZN(n4308) );
  INV_X1 U5360 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6751) );
  OR2_X2 U5361 ( .A1(n4432), .A2(n4301), .ZN(n5244) );
  NOR2_X1 U5362 ( .A1(n6497), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5441) );
  INV_X1 U5363 ( .A(n5441), .ZN(n4307) );
  OAI211_X1 U5364 ( .C1(n4308), .C2(n6751), .A(n5244), .B(n4307), .ZN(U2788)
         );
  INV_X1 U5365 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4312) );
  OR2_X1 U5366 ( .A1(n5244), .A2(READY_N), .ZN(n4309) );
  NAND2_X1 U5367 ( .A1(n6305), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4311) );
  NAND2_X1 U5368 ( .A1(n4554), .A2(n4884), .ZN(n4310) );
  NAND2_X1 U5369 ( .A1(n6304), .A2(DATAI_0_), .ZN(n4315) );
  OAI211_X1 U5370 ( .C1(n6307), .C2(n4312), .A(n4311), .B(n4315), .ZN(U2939)
         );
  INV_X1 U5371 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4314) );
  NAND2_X1 U5372 ( .A1(n6305), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4313) );
  NAND2_X1 U5373 ( .A1(n6304), .A2(DATAI_5_), .ZN(n4354) );
  OAI211_X1 U5374 ( .C1(n6307), .C2(n4314), .A(n4313), .B(n4354), .ZN(U2929)
         );
  NAND2_X1 U5375 ( .A1(n6305), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4316) );
  OAI211_X1 U5376 ( .C1(n6307), .C2(n4317), .A(n4316), .B(n4315), .ZN(U2924)
         );
  INV_X1 U5377 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4319) );
  NAND2_X1 U5378 ( .A1(n6305), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U5379 ( .A1(n6304), .A2(DATAI_7_), .ZN(n4322) );
  OAI211_X1 U5380 ( .C1(n6307), .C2(n4319), .A(n4318), .B(n4322), .ZN(U2946)
         );
  NAND2_X1 U5381 ( .A1(n6305), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4320) );
  NAND2_X1 U5382 ( .A1(n6304), .A2(DATAI_2_), .ZN(n4325) );
  OAI211_X1 U5383 ( .C1(n6307), .C2(n4321), .A(n4320), .B(n4325), .ZN(U2926)
         );
  NAND2_X1 U5384 ( .A1(n6305), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4323) );
  OAI211_X1 U5385 ( .C1(n6307), .C2(n4324), .A(n4323), .B(n4322), .ZN(U2931)
         );
  INV_X1 U5386 ( .A(EAX_REG_2__SCAN_IN), .ZN(n4327) );
  NAND2_X1 U5387 ( .A1(n6305), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4326) );
  OAI211_X1 U5388 ( .C1(n6307), .C2(n4327), .A(n4326), .B(n4325), .ZN(U2941)
         );
  INV_X1 U5389 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n4329) );
  INV_X1 U5390 ( .A(DATAI_1_), .ZN(n4553) );
  NOR2_X1 U5391 ( .A1(n6287), .A2(n4553), .ZN(n4330) );
  AOI21_X1 U5392 ( .B1(n6301), .B2(EAX_REG_1__SCAN_IN), .A(n4330), .ZN(n4328)
         );
  OAI21_X1 U5393 ( .B1(n6298), .B2(n4329), .A(n4328), .ZN(U2940) );
  INV_X1 U5394 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4332) );
  AOI21_X1 U5395 ( .B1(n6301), .B2(EAX_REG_17__SCAN_IN), .A(n4330), .ZN(n4331)
         );
  OAI21_X1 U5396 ( .B1(n6298), .B2(n4332), .A(n4331), .ZN(U2925) );
  INV_X1 U5397 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n4334) );
  INV_X1 U5398 ( .A(DATAI_4_), .ZN(n4512) );
  NOR2_X1 U5399 ( .A1(n6287), .A2(n4512), .ZN(n4341) );
  AOI21_X1 U5400 ( .B1(n6301), .B2(EAX_REG_4__SCAN_IN), .A(n4341), .ZN(n4333)
         );
  OAI21_X1 U5401 ( .B1(n6298), .B2(n4334), .A(n4333), .ZN(U2943) );
  INV_X1 U5402 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4336) );
  INV_X1 U5403 ( .A(DATAI_3_), .ZN(n4503) );
  NOR2_X1 U5404 ( .A1(n6287), .A2(n4503), .ZN(n4347) );
  AOI21_X1 U5405 ( .B1(n6301), .B2(EAX_REG_19__SCAN_IN), .A(n4347), .ZN(n4335)
         );
  OAI21_X1 U5406 ( .B1(n6298), .B2(n4336), .A(n4335), .ZN(U2927) );
  INV_X1 U5407 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n4338) );
  INV_X1 U5408 ( .A(DATAI_8_), .ZN(n6794) );
  NOR2_X1 U5409 ( .A1(n6287), .A2(n6794), .ZN(n4350) );
  AOI21_X1 U5410 ( .B1(n6301), .B2(EAX_REG_24__SCAN_IN), .A(n4350), .ZN(n4337)
         );
  OAI21_X1 U5411 ( .B1(n6298), .B2(n4338), .A(n4337), .ZN(U2932) );
  INV_X1 U5412 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n4340) );
  INV_X1 U5413 ( .A(DATAI_6_), .ZN(n4706) );
  NOR2_X1 U5414 ( .A1(n6287), .A2(n4706), .ZN(n4344) );
  AOI21_X1 U5415 ( .B1(n6301), .B2(EAX_REG_22__SCAN_IN), .A(n4344), .ZN(n4339)
         );
  OAI21_X1 U5416 ( .B1(n6298), .B2(n4340), .A(n4339), .ZN(U2930) );
  INV_X1 U5417 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n4343) );
  AOI21_X1 U5418 ( .B1(n6301), .B2(EAX_REG_20__SCAN_IN), .A(n4341), .ZN(n4342)
         );
  OAI21_X1 U5419 ( .B1(n6298), .B2(n4343), .A(n4342), .ZN(U2928) );
  INV_X1 U5420 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n4346) );
  AOI21_X1 U5421 ( .B1(n6301), .B2(EAX_REG_6__SCAN_IN), .A(n4344), .ZN(n4345)
         );
  OAI21_X1 U5422 ( .B1(n6298), .B2(n4346), .A(n4345), .ZN(U2945) );
  INV_X1 U5423 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n4349) );
  AOI21_X1 U5424 ( .B1(n6301), .B2(EAX_REG_3__SCAN_IN), .A(n4347), .ZN(n4348)
         );
  OAI21_X1 U5425 ( .B1(n6298), .B2(n4349), .A(n4348), .ZN(U2942) );
  INV_X1 U5426 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n4352) );
  AOI21_X1 U5427 ( .B1(n6301), .B2(EAX_REG_8__SCAN_IN), .A(n4350), .ZN(n4351)
         );
  OAI21_X1 U5428 ( .B1(n6298), .B2(n4352), .A(n4351), .ZN(U2947) );
  INV_X1 U5429 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n4355) );
  NAND2_X1 U5430 ( .A1(n6301), .A2(EAX_REG_5__SCAN_IN), .ZN(n4353) );
  OAI211_X1 U5431 ( .C1(n6298), .C2(n4355), .A(n4354), .B(n4353), .ZN(U2944)
         );
  NAND2_X1 U5432 ( .A1(n4592), .A2(n4241), .ZN(n4359) );
  AOI21_X1 U5433 ( .B1(n4301), .B2(n4357), .A(n4356), .ZN(n4358) );
  AND2_X1 U5434 ( .A1(n4359), .A2(n4358), .ZN(n4360) );
  MUX2_X1 U5435 ( .A(n4360), .B(n4577), .S(n6581), .Z(n4369) );
  OR2_X1 U5436 ( .A1(n6581), .A2(n4575), .ZN(n4363) );
  NAND2_X1 U5437 ( .A1(n4565), .A2(n4361), .ZN(n4362) );
  INV_X1 U5438 ( .A(n4364), .ZN(n4367) );
  INV_X1 U5439 ( .A(n4365), .ZN(n4366) );
  NAND2_X1 U5440 ( .A1(n4367), .A2(n4366), .ZN(n4368) );
  NAND2_X1 U5441 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4602) );
  NOR2_X1 U5442 ( .A1(n6579), .A2(n4602), .ZN(n4920) );
  AOI22_X1 U5443 ( .A1(n4891), .A2(n4468), .B1(FLUSH_REG_SCAN_IN), .B2(n4920), 
        .ZN(n4373) );
  INV_X1 U5444 ( .A(n4734), .ZN(n4923) );
  NOR2_X1 U5445 ( .A1(n3405), .A2(n4923), .ZN(n4371) );
  XNOR2_X1 U5446 ( .A(n4371), .B(n4370), .ZN(n6209) );
  NAND3_X1 U5447 ( .A1(n6209), .A2(n4565), .A3(n5231), .ZN(n4372) );
  NAND2_X1 U5448 ( .A1(n6579), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4921) );
  NAND2_X1 U5449 ( .A1(n4373), .A2(n4921), .ZN(n6052) );
  OAI22_X1 U5450 ( .A1(n4373), .A2(n4372), .B1(n4370), .B2(n6052), .ZN(U3455)
         );
  OAI21_X1 U5451 ( .B1(n4376), .B2(n4375), .A(n4374), .ZN(n5576) );
  OR2_X1 U5452 ( .A1(n4377), .A2(n4901), .ZN(n4378) );
  AND2_X1 U5453 ( .A1(n4379), .A2(n4378), .ZN(n4428) );
  OAI22_X1 U5454 ( .A1(n5608), .A2(n4428), .B1(n4380), .B2(n6243), .ZN(n4381)
         );
  INV_X1 U5455 ( .A(n4381), .ZN(n4382) );
  OAI21_X1 U5456 ( .B1(n5576), .B2(n5609), .A(n4382), .ZN(U2858) );
  XNOR2_X1 U5457 ( .A(n4384), .B(n4383), .ZN(n5584) );
  XNOR2_X1 U5458 ( .A(n4385), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4466)
         );
  INV_X1 U5459 ( .A(n4466), .ZN(n4391) );
  INV_X1 U5460 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4386) );
  NOR2_X1 U5461 ( .A1(n6435), .A2(n4386), .ZN(n4463) );
  INV_X1 U5462 ( .A(n4387), .ZN(n4389) );
  INV_X1 U5463 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4388) );
  AOI21_X1 U5464 ( .B1(n5833), .B2(n4389), .A(n4388), .ZN(n4390) );
  AOI211_X1 U5465 ( .C1(n4391), .C2(n6340), .A(n4463), .B(n4390), .ZN(n4392)
         );
  OAI21_X1 U5466 ( .B1(n5584), .B2(n5779), .A(n4392), .ZN(U2986) );
  INV_X1 U5467 ( .A(n6039), .ZN(n5568) );
  INV_X1 U5468 ( .A(n4393), .ZN(n4395) );
  AND3_X1 U5469 ( .A1(n4241), .A2(n4395), .A3(n4394), .ZN(n4396) );
  AND2_X1 U5470 ( .A1(n4255), .A2(n4396), .ZN(n4399) );
  INV_X1 U5471 ( .A(n4397), .ZN(n4398) );
  NAND2_X1 U5472 ( .A1(n4399), .A2(n4398), .ZN(n4589) );
  NAND2_X1 U5473 ( .A1(n5568), .A2(n4589), .ZN(n4405) );
  INV_X1 U5474 ( .A(n4400), .ZN(n4420) );
  INV_X1 U5475 ( .A(n4401), .ZN(n4403) );
  INV_X1 U5476 ( .A(n4402), .ZN(n5232) );
  NAND3_X1 U5477 ( .A1(n4420), .A2(n4403), .A3(n5232), .ZN(n4404) );
  OAI211_X1 U5478 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n4592), .A(n4405), .B(n4404), .ZN(n4890) );
  INV_X1 U5479 ( .A(n4406), .ZN(n4409) );
  NAND2_X1 U5480 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5227) );
  INV_X1 U5481 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U5482 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4407), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6389), .ZN(n5226) );
  INV_X1 U5483 ( .A(n5226), .ZN(n4408) );
  OAI22_X1 U5484 ( .A1(n6048), .A2(n4409), .B1(n5227), .B2(n4408), .ZN(n4410)
         );
  AOI21_X1 U5485 ( .B1(n5231), .B2(n4890), .A(n4410), .ZN(n4413) );
  INV_X1 U5486 ( .A(n6052), .ZN(n5236) );
  OAI21_X1 U5487 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6048), .A(n6052), 
        .ZN(n4411) );
  INV_X1 U5488 ( .A(n4411), .ZN(n4421) );
  OAI22_X1 U5489 ( .A1(n4413), .A2(n5236), .B1(n4412), .B2(n4421), .ZN(U3460)
         );
  INV_X1 U5490 ( .A(n4414), .ZN(n4415) );
  AOI21_X1 U5491 ( .B1(n4417), .B2(n4416), .A(n4415), .ZN(n5577) );
  INV_X1 U5492 ( .A(n5577), .ZN(n4418) );
  OAI222_X1 U5493 ( .A1(n4418), .A2(n5608), .B1(n6758), .B2(n6243), .C1(n5609), 
        .C2(n5584), .ZN(U2859) );
  INV_X1 U5494 ( .A(n4592), .ZN(n4419) );
  NAND2_X1 U5495 ( .A1(n4419), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4886) );
  INV_X1 U5496 ( .A(n5231), .ZN(n6050) );
  AOI22_X1 U5497 ( .A1(n3552), .A2(n4589), .B1(n4420), .B2(n4033), .ZN(n4887)
         );
  NOR2_X1 U5498 ( .A1(n4887), .A2(n6050), .ZN(n4423) );
  OAI21_X1 U5499 ( .B1(n5254), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4421), 
        .ZN(n4422) );
  OAI22_X1 U5500 ( .A1(n4423), .A2(n4422), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6052), .ZN(n4424) );
  OAI21_X1 U5501 ( .B1(n4886), .B2(n6050), .A(n4424), .ZN(U3461) );
  XNOR2_X1 U5502 ( .A(n2988), .B(n4425), .ZN(n4564) );
  NAND2_X1 U5503 ( .A1(n5988), .A2(n5986), .ZN(n6395) );
  NAND2_X1 U5504 ( .A1(n6395), .A2(n4426), .ZN(n4427) );
  MUX2_X1 U5505 ( .A(n4427), .B(n6391), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4431) );
  INV_X1 U5506 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6656) );
  OAI22_X1 U5507 ( .A1(n6434), .A2(n4428), .B1(n6656), .B2(n6435), .ZN(n4429)
         );
  INV_X1 U5508 ( .A(n4429), .ZN(n4430) );
  OAI211_X1 U5509 ( .C1(n4564), .C2(n6351), .A(n4431), .B(n4430), .ZN(U3017)
         );
  INV_X1 U5510 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4436) );
  OR2_X1 U5511 ( .A1(n4432), .A2(n4592), .ZN(n4433) );
  NAND2_X1 U5512 ( .A1(n6261), .A2(n5270), .ZN(n6250) );
  INV_X2 U5513 ( .A(n6263), .ZN(n6664) );
  NOR2_X4 U5514 ( .A1(n6261), .A2(n6664), .ZN(n6276) );
  AOI22_X1 U5515 ( .A1(n6664), .A2(UWORD_REG_14__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4435) );
  OAI21_X1 U5516 ( .B1(n4436), .B2(n6250), .A(n4435), .ZN(U2893) );
  AOI22_X1 U5517 ( .A1(n6664), .A2(UWORD_REG_0__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4437) );
  OAI21_X1 U5518 ( .B1(n4317), .B2(n6250), .A(n4437), .ZN(U2907) );
  INV_X1 U5519 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4439) );
  AOI22_X1 U5520 ( .A1(n6664), .A2(UWORD_REG_1__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4438) );
  OAI21_X1 U5521 ( .B1(n4439), .B2(n6250), .A(n4438), .ZN(U2906) );
  AOI22_X1 U5522 ( .A1(n6664), .A2(UWORD_REG_2__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4440) );
  OAI21_X1 U5523 ( .B1(n4321), .B2(n6250), .A(n4440), .ZN(U2905) );
  INV_X1 U5524 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4442) );
  AOI22_X1 U5525 ( .A1(n6664), .A2(UWORD_REG_3__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4441) );
  OAI21_X1 U5526 ( .B1(n4442), .B2(n6250), .A(n4441), .ZN(U2904) );
  INV_X1 U5527 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4444) );
  AOI22_X1 U5528 ( .A1(n6664), .A2(UWORD_REG_4__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4443) );
  OAI21_X1 U5529 ( .B1(n4444), .B2(n6250), .A(n4443), .ZN(U2903) );
  AOI22_X1 U5530 ( .A1(n6664), .A2(UWORD_REG_11__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4445) );
  OAI21_X1 U5531 ( .B1(n3862), .B2(n6250), .A(n4445), .ZN(U2896) );
  INV_X1 U5532 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4447) );
  AOI22_X1 U5533 ( .A1(n6664), .A2(UWORD_REG_6__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4446) );
  OAI21_X1 U5534 ( .B1(n4447), .B2(n6250), .A(n4446), .ZN(U2901) );
  AOI22_X1 U5535 ( .A1(n6664), .A2(UWORD_REG_7__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4448) );
  OAI21_X1 U5536 ( .B1(n4324), .B2(n6250), .A(n4448), .ZN(U2900) );
  INV_X1 U5537 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4450) );
  AOI22_X1 U5538 ( .A1(n6664), .A2(UWORD_REG_8__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4449) );
  OAI21_X1 U5539 ( .B1(n4450), .B2(n6250), .A(n4449), .ZN(U2899) );
  AOI22_X1 U5540 ( .A1(n6664), .A2(UWORD_REG_9__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4451) );
  OAI21_X1 U5541 ( .B1(n3825), .B2(n6250), .A(n4451), .ZN(U2898) );
  AOI22_X1 U5542 ( .A1(n6664), .A2(UWORD_REG_10__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4452) );
  OAI21_X1 U5543 ( .B1(n6282), .B2(n6250), .A(n4452), .ZN(U2897) );
  AOI22_X1 U5544 ( .A1(n6664), .A2(UWORD_REG_13__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4453) );
  OAI21_X1 U5545 ( .B1(n3906), .B2(n6250), .A(n4453), .ZN(U2894) );
  NAND2_X1 U5546 ( .A1(n4709), .A2(n4454), .ZN(n4608) );
  OAI21_X1 U5547 ( .B1(n4709), .B2(n4454), .A(n4608), .ZN(n5557) );
  INV_X1 U5548 ( .A(n4456), .ZN(n5560) );
  NAND2_X1 U5549 ( .A1(n4142), .A2(n5560), .ZN(n4458) );
  INV_X1 U5550 ( .A(n4457), .ZN(n4612) );
  AOI21_X1 U5551 ( .B1(n4459), .B2(n4458), .A(n4612), .ZN(n6421) );
  INV_X1 U5552 ( .A(n6243), .ZN(n5592) );
  AOI22_X1 U5553 ( .A1(n6239), .A2(n6421), .B1(EBX_REG_3__SCAN_IN), .B2(n5592), 
        .ZN(n4460) );
  OAI21_X1 U5554 ( .B1(n5557), .B2(n5609), .A(n4460), .ZN(U2856) );
  INV_X1 U5555 ( .A(n6391), .ZN(n4462) );
  INV_X1 U5556 ( .A(n5986), .ZN(n4461) );
  OAI22_X1 U5557 ( .A1(n3010), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(n4462), 
        .B2(n4461), .ZN(n4465) );
  AOI21_X1 U5558 ( .B1(n6422), .B2(n5577), .A(n4463), .ZN(n4464) );
  OAI211_X1 U5559 ( .C1(n4466), .C2(n6351), .A(n4465), .B(n4464), .ZN(U3018)
         );
  NOR2_X1 U5560 ( .A1(n4467), .A2(n5242), .ZN(n4469) );
  NAND2_X1 U5561 ( .A1(n4472), .A2(n4548), .ZN(n4473) );
  INV_X1 U5562 ( .A(n4473), .ZN(n4474) );
  INV_X1 U5563 ( .A(DATAI_0_), .ZN(n4490) );
  OAI222_X1 U5564 ( .A1(n5658), .A2(n5584), .B1(n4711), .B2(n4490), .C1(n6249), 
        .C2(n4312), .ZN(U2891) );
  INV_X1 U5565 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6729) );
  OAI222_X1 U5566 ( .A1(n5576), .A2(n5658), .B1(n4711), .B2(n4553), .C1(n6249), 
        .C2(n6729), .ZN(U2890) );
  INV_X1 U5567 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6822) );
  OAI222_X1 U5568 ( .A1(n5557), .A2(n5658), .B1(n4711), .B2(n4503), .C1(n6822), 
        .C2(n6249), .ZN(U2888) );
  XNOR2_X1 U5569 ( .A(n4608), .B(n4606), .ZN(n6331) );
  INV_X1 U5570 ( .A(n6331), .ZN(n6219) );
  INV_X1 U5571 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4475) );
  XNOR2_X1 U5572 ( .A(n4612), .B(n4611), .ZN(n6208) );
  OAI222_X1 U5573 ( .A1(n5609), .A2(n6219), .B1(n4475), .B2(n6243), .C1(n5608), 
        .C2(n6208), .ZN(U2855) );
  INV_X1 U5574 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6781) );
  OAI222_X1 U5575 ( .A1(n5658), .A2(n6219), .B1(n4711), .B2(n4512), .C1(n6249), 
        .C2(n6781), .ZN(U2887) );
  INV_X1 U5576 ( .A(n4476), .ZN(n4478) );
  AOI21_X1 U5577 ( .B1(n4478), .B2(n4477), .A(n4709), .ZN(n6341) );
  INV_X1 U5578 ( .A(n6341), .ZN(n4479) );
  INV_X1 U5579 ( .A(DATAI_2_), .ZN(n4526) );
  OAI222_X1 U5580 ( .A1(n4479), .A2(n5658), .B1(n4711), .B2(n4526), .C1(n6249), 
        .C2(n4327), .ZN(U2889) );
  INV_X1 U5581 ( .A(n6042), .ZN(n4481) );
  OAI21_X1 U5582 ( .B1(n5033), .B2(n4481), .A(n6666), .ZN(n4495) );
  NAND2_X1 U5583 ( .A1(n4483), .A2(n5568), .ZN(n4719) );
  INV_X1 U5584 ( .A(n4719), .ZN(n4485) );
  NAND2_X1 U5585 ( .A1(n4485), .A2(n5552), .ZN(n5093) );
  OR2_X1 U5586 ( .A1(n5093), .A2(n6490), .ZN(n4487) );
  INV_X1 U5587 ( .A(n4720), .ZN(n4486) );
  NAND2_X1 U5588 ( .A1(n4486), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6562) );
  NAND3_X1 U5589 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n4895), .ZN(n5084) );
  OAI22_X1 U5590 ( .A1(n4495), .A2(n4491), .B1(n5084), .B2(n6575), .ZN(n6567)
         );
  INV_X1 U5591 ( .A(n6567), .ZN(n4518) );
  NOR2_X1 U5592 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6670) );
  INV_X1 U5593 ( .A(n4602), .ZN(n4488) );
  OR2_X1 U5594 ( .A1(n6670), .A2(n4488), .ZN(n4489) );
  INV_X1 U5595 ( .A(n4491), .ZN(n4494) );
  NOR2_X1 U5596 ( .A1(n4986), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4492)
         );
  AOI21_X1 U5597 ( .B1(n5084), .B2(n6497), .A(n5038), .ZN(n4493) );
  OAI21_X1 U5598 ( .B1(n4495), .B2(n4494), .A(n4493), .ZN(n6569) );
  INV_X1 U5599 ( .A(DATAI_24_), .ZN(n4496) );
  NOR2_X1 U5600 ( .A1(n5779), .A2(n4496), .ZN(n6502) );
  INV_X1 U5601 ( .A(n6502), .ZN(n5119) );
  NOR2_X1 U5602 ( .A1(n6572), .A2(n5119), .ZN(n4501) );
  NAND2_X1 U5603 ( .A1(n6332), .A2(DATAI_16_), .ZN(n6495) );
  INV_X1 U5604 ( .A(n4921), .ZN(n4498) );
  AND2_X1 U5605 ( .A1(n4555), .A2(n5270), .ZN(n6469) );
  OAI22_X1 U5606 ( .A1(n6565), .A2(n6495), .B1(n6494), .B2(n6562), .ZN(n4500)
         );
  AOI211_X1 U5607 ( .C1(n6569), .C2(INSTQUEUE_REG_11__0__SCAN_IN), .A(n4501), 
        .B(n4500), .ZN(n4502) );
  OAI21_X1 U5608 ( .B1(n4518), .B2(n6505), .A(n4502), .ZN(U3108) );
  NAND2_X1 U5609 ( .A1(n6332), .A2(DATAI_27_), .ZN(n6512) );
  NOR2_X1 U5610 ( .A1(n6572), .A2(n6512), .ZN(n4505) );
  NAND2_X1 U5611 ( .A1(n6332), .A2(DATAI_19_), .ZN(n6489) );
  AND2_X1 U5612 ( .A1(n4555), .A2(n3283), .ZN(n6483) );
  OAI22_X1 U5613 ( .A1(n6565), .A2(n6489), .B1(n6511), .B2(n6562), .ZN(n4504)
         );
  AOI211_X1 U5614 ( .C1(n6569), .C2(INSTQUEUE_REG_11__3__SCAN_IN), .A(n4505), 
        .B(n4504), .ZN(n4506) );
  OAI21_X1 U5615 ( .B1(n4518), .B2(n6517), .A(n4506), .ZN(U3111) );
  NAND2_X1 U5616 ( .A1(n6332), .A2(DATAI_30_), .ZN(n6532) );
  NOR2_X1 U5617 ( .A1(n6572), .A2(n6532), .ZN(n4510) );
  INV_X1 U5618 ( .A(DATAI_22_), .ZN(n4507) );
  NOR2_X1 U5619 ( .A1(n5779), .A2(n4507), .ZN(n6534) );
  INV_X1 U5620 ( .A(n6534), .ZN(n6091) );
  AND2_X1 U5621 ( .A1(n4555), .A2(n4508), .ZN(n6459) );
  OAI22_X1 U5622 ( .A1(n6565), .A2(n6091), .B1(n6531), .B2(n6562), .ZN(n4509)
         );
  AOI211_X1 U5623 ( .C1(n6569), .C2(INSTQUEUE_REG_11__6__SCAN_IN), .A(n4510), 
        .B(n4509), .ZN(n4511) );
  OAI21_X1 U5624 ( .B1(n4518), .B2(n6537), .A(n4511), .ZN(U3114) );
  INV_X1 U5625 ( .A(DATAI_28_), .ZN(n4513) );
  NOR2_X1 U5626 ( .A1(n5779), .A2(n4513), .ZN(n6522) );
  INV_X1 U5627 ( .A(n6522), .ZN(n6455) );
  NOR2_X1 U5628 ( .A1(n6572), .A2(n6455), .ZN(n4516) );
  INV_X1 U5629 ( .A(DATAI_20_), .ZN(n4514) );
  NOR2_X1 U5630 ( .A1(n5779), .A2(n4514), .ZN(n6451) );
  INV_X1 U5631 ( .A(n6451), .ZN(n6519) );
  AND2_X1 U5632 ( .A1(n4555), .A2(n3271), .ZN(n6450) );
  OAI22_X1 U5633 ( .A1(n6565), .A2(n6519), .B1(n6518), .B2(n6562), .ZN(n4515)
         );
  AOI211_X1 U5634 ( .C1(n6569), .C2(INSTQUEUE_REG_11__4__SCAN_IN), .A(n4516), 
        .B(n4515), .ZN(n4517) );
  OAI21_X1 U5635 ( .B1(n4518), .B2(n6525), .A(n4517), .ZN(U3112) );
  NAND2_X1 U5636 ( .A1(n6332), .A2(DATAI_26_), .ZN(n6678) );
  AOI21_X1 U5637 ( .B1(n4659), .B2(n4480), .A(n5779), .ZN(n4521) );
  NOR2_X1 U5638 ( .A1(n6497), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5150) );
  NOR2_X1 U5639 ( .A1(n4483), .A2(n6039), .ZN(n4956) );
  INV_X1 U5640 ( .A(n4556), .ZN(n4520) );
  AOI21_X1 U5641 ( .B1(n5036), .B2(n4956), .A(n4520), .ZN(n4523) );
  OAI21_X1 U5642 ( .B1(n4521), .B2(n5150), .A(n4523), .ZN(n4522) );
  NAND2_X1 U5643 ( .A1(n4552), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4530)
         );
  NAND2_X1 U5644 ( .A1(n4659), .A2(n6054), .ZN(n4833) );
  NAND2_X1 U5645 ( .A1(n6332), .A2(DATAI_18_), .ZN(n6681) );
  INV_X1 U5646 ( .A(n6681), .ZN(n6447) );
  INV_X1 U5647 ( .A(n4523), .ZN(n4525) );
  AOI22_X1 U5648 ( .A1(n4525), .A2(n6666), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4524), .ZN(n4557) );
  OAI22_X1 U5649 ( .A1(n4557), .A2(n6682), .B1(n4556), .B2(n6676), .ZN(n4528)
         );
  AOI21_X1 U5650 ( .B1(n4874), .B2(n6447), .A(n4528), .ZN(n4529) );
  OAI211_X1 U5651 ( .C1(n4953), .C2(n6678), .A(n4530), .B(n4529), .ZN(U3142)
         );
  NAND2_X1 U5652 ( .A1(n4552), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4533)
         );
  INV_X1 U5653 ( .A(n6489), .ZN(n6514) );
  OAI22_X1 U5654 ( .A1(n4557), .A2(n6517), .B1(n4556), .B2(n6511), .ZN(n4531)
         );
  AOI21_X1 U5655 ( .B1(n4874), .B2(n6514), .A(n4531), .ZN(n4532) );
  OAI211_X1 U5656 ( .C1(n4953), .C2(n6512), .A(n4533), .B(n4532), .ZN(U3143)
         );
  NAND2_X1 U5657 ( .A1(n6332), .A2(DATAI_29_), .ZN(n6561) );
  NAND2_X1 U5658 ( .A1(n4552), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4537)
         );
  INV_X1 U5659 ( .A(DATAI_21_), .ZN(n4534) );
  NOR2_X1 U5660 ( .A1(n5779), .A2(n4534), .ZN(n6527) );
  INV_X1 U5661 ( .A(DATAI_5_), .ZN(n4615) );
  AND2_X1 U5662 ( .A1(n4555), .A2(n5610), .ZN(n6456) );
  OAI22_X1 U5663 ( .A1(n4557), .A2(n6530), .B1(n4556), .B2(n6555), .ZN(n4535)
         );
  AOI21_X1 U5664 ( .B1(n4874), .B2(n6527), .A(n4535), .ZN(n4536) );
  OAI211_X1 U5665 ( .C1(n4953), .C2(n6561), .A(n4537), .B(n4536), .ZN(U3145)
         );
  NAND2_X1 U5666 ( .A1(n4552), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4540)
         );
  INV_X1 U5667 ( .A(n6495), .ZN(n5117) );
  OAI22_X1 U5668 ( .A1(n4557), .A2(n6505), .B1(n4556), .B2(n6494), .ZN(n4538)
         );
  AOI21_X1 U5669 ( .B1(n4874), .B2(n5117), .A(n4538), .ZN(n4539) );
  OAI211_X1 U5670 ( .C1(n4953), .C2(n5119), .A(n4540), .B(n4539), .ZN(U3140)
         );
  NAND2_X1 U5671 ( .A1(n4552), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4543)
         );
  OAI22_X1 U5672 ( .A1(n4557), .A2(n6525), .B1(n4556), .B2(n6518), .ZN(n4541)
         );
  AOI21_X1 U5673 ( .B1(n4874), .B2(n6451), .A(n4541), .ZN(n4542) );
  OAI211_X1 U5674 ( .C1(n4953), .C2(n6455), .A(n4543), .B(n4542), .ZN(U3144)
         );
  NAND2_X1 U5675 ( .A1(n4552), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4546)
         );
  OAI22_X1 U5676 ( .A1(n4557), .A2(n6537), .B1(n4556), .B2(n6531), .ZN(n4544)
         );
  AOI21_X1 U5677 ( .B1(n4874), .B2(n6534), .A(n4544), .ZN(n4545) );
  OAI211_X1 U5678 ( .C1(n4953), .C2(n6532), .A(n4546), .B(n4545), .ZN(U3146)
         );
  NAND2_X1 U5679 ( .A1(n6332), .A2(DATAI_31_), .ZN(n6573) );
  NAND2_X1 U5680 ( .A1(n4552), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4551)
         );
  INV_X1 U5681 ( .A(DATAI_23_), .ZN(n4547) );
  NOR2_X1 U5682 ( .A1(n5779), .A2(n4547), .ZN(n6540) );
  INV_X1 U5683 ( .A(DATAI_7_), .ZN(n6750) );
  AND2_X1 U5684 ( .A1(n4555), .A2(n4548), .ZN(n5112) );
  OAI22_X1 U5685 ( .A1(n4557), .A2(n6543), .B1(n4556), .B2(n6563), .ZN(n4549)
         );
  AOI21_X1 U5686 ( .B1(n4874), .B2(n6540), .A(n4549), .ZN(n4550) );
  OAI211_X1 U5687 ( .C1(n4953), .C2(n6573), .A(n4551), .B(n4550), .ZN(U3147)
         );
  NAND2_X1 U5688 ( .A1(n6332), .A2(DATAI_25_), .ZN(n6550) );
  NAND2_X1 U5689 ( .A1(n4552), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4560)
         );
  NAND2_X1 U5690 ( .A1(n6332), .A2(DATAI_17_), .ZN(n6545) );
  INV_X1 U5691 ( .A(n6545), .ZN(n6507) );
  AND2_X1 U5692 ( .A1(n4555), .A2(n4554), .ZN(n6472) );
  OAI22_X1 U5693 ( .A1(n4557), .A2(n6510), .B1(n4556), .B2(n6544), .ZN(n4558)
         );
  AOI21_X1 U5694 ( .B1(n4874), .B2(n6507), .A(n4558), .ZN(n4559) );
  OAI211_X1 U5695 ( .C1(n4953), .C2(n6550), .A(n4560), .B(n4559), .ZN(U3141)
         );
  INV_X1 U5696 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5569) );
  OAI22_X1 U5697 ( .A1(n5833), .A2(n5569), .B1(n6435), .B2(n6656), .ZN(n4562)
         );
  NOR2_X1 U5698 ( .A1(n5576), .A2(n5779), .ZN(n4561) );
  AOI211_X1 U5699 ( .C1(n6312), .C2(n5569), .A(n4562), .B(n4561), .ZN(n4563)
         );
  OAI21_X1 U5700 ( .B1(n4564), .B2(n6316), .A(n4563), .ZN(U2985) );
  NAND2_X1 U5701 ( .A1(n6209), .A2(n4565), .ZN(n4566) );
  OAI21_X1 U5702 ( .B1(n4891), .B2(n4370), .A(n4566), .ZN(n4567) );
  NAND2_X1 U5703 ( .A1(n4567), .A2(n5254), .ZN(n4570) );
  INV_X1 U5704 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6105) );
  NAND2_X1 U5705 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6105), .ZN(n4572) );
  INV_X1 U5706 ( .A(n4572), .ZN(n4568) );
  NAND2_X1 U5707 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4568), .ZN(n4569) );
  NAND2_X1 U5708 ( .A1(n4570), .A2(n4569), .ZN(n4574) );
  INV_X1 U5709 ( .A(n4574), .ZN(n4600) );
  NOR2_X1 U5710 ( .A1(n4572), .A2(n4571), .ZN(n4573) );
  NOR2_X1 U5711 ( .A1(n4574), .A2(n4573), .ZN(n4599) );
  NAND2_X1 U5712 ( .A1(n5552), .A2(n4589), .ZN(n4588) );
  INV_X1 U5713 ( .A(n4575), .ZN(n4576) );
  OR2_X1 U5714 ( .A1(n4577), .A2(n4576), .ZN(n4595) );
  MUX2_X1 U5715 ( .A(n4578), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4402), 
        .Z(n4579) );
  XNOR2_X1 U5716 ( .A(n4580), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4584)
         );
  AOI21_X1 U5717 ( .B1(n4402), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4581), 
        .ZN(n4582) );
  NOR2_X1 U5718 ( .A1(n4583), .A2(n4582), .ZN(n6049) );
  OAI22_X1 U5719 ( .A1(n4592), .A2(n4584), .B1(n6049), .B2(n4590), .ZN(n4585)
         );
  AOI21_X1 U5720 ( .B1(n4595), .B2(n4586), .A(n4585), .ZN(n4587) );
  NAND2_X1 U5721 ( .A1(n4588), .A2(n4587), .ZN(n6047) );
  MUX2_X1 U5722 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6047), .S(n4891), 
        .Z(n4900) );
  INV_X1 U5723 ( .A(n4589), .ZN(n4597) );
  XNOR2_X1 U5724 ( .A(n4402), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4594)
         );
  XNOR2_X1 U5725 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4591) );
  OAI22_X1 U5726 ( .A1(n4592), .A2(n4591), .B1(n4590), .B2(n4594), .ZN(n4593)
         );
  AOI21_X1 U5727 ( .B1(n4595), .B2(n4594), .A(n4593), .ZN(n4596) );
  OAI21_X1 U5728 ( .B1(n4483), .B2(n4597), .A(n4596), .ZN(n5230) );
  MUX2_X1 U5729 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5230), .S(n4891), 
        .Z(n4896) );
  NAND3_X1 U5730 ( .A1(n4900), .A2(n4896), .A3(n5254), .ZN(n4598) );
  AOI21_X1 U5731 ( .B1(n4600), .B2(n4401), .A(n4915), .ZN(n4603) );
  OAI21_X1 U5732 ( .B1(n4603), .B2(FLUSH_REG_SCAN_IN), .A(n4920), .ZN(n4601)
         );
  NAND2_X1 U5733 ( .A1(n4601), .A2(n4926), .ZN(n6443) );
  NOR2_X1 U5734 ( .A1(n4603), .A2(n4602), .ZN(n6576) );
  NAND2_X1 U5735 ( .A1(n4986), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4662) );
  INV_X1 U5736 ( .A(n4662), .ZN(n6044) );
  OAI22_X1 U5737 ( .A1(n5043), .A2(n6497), .B1(n6044), .B2(n6490), .ZN(n4604)
         );
  OAI21_X1 U5738 ( .B1(n6576), .B2(n4604), .A(n6443), .ZN(n4605) );
  OAI21_X1 U5739 ( .B1(n6443), .B2(n5152), .A(n4605), .ZN(U3465) );
  INV_X1 U5740 ( .A(n4606), .ZN(n4607) );
  NOR2_X1 U5741 ( .A1(n4608), .A2(n4607), .ZN(n4609) );
  NAND2_X1 U5742 ( .A1(n4609), .A2(n4708), .ZN(n4700) );
  OAI21_X1 U5743 ( .B1(n4609), .B2(n4708), .A(n4700), .ZN(n5529) );
  INV_X1 U5744 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4614) );
  AOI21_X1 U5745 ( .B1(n4612), .B2(n4611), .A(n4610), .ZN(n4613) );
  OR2_X1 U5746 ( .A1(n4613), .A2(n4703), .ZN(n5537) );
  OAI222_X1 U5747 ( .A1(n5529), .A2(n5609), .B1(n6243), .B2(n4614), .C1(n5537), 
        .C2(n5608), .ZN(U2854) );
  INV_X1 U5748 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6271) );
  OAI222_X1 U5749 ( .A1(n5529), .A2(n5658), .B1(n4711), .B2(n4615), .C1(n6249), 
        .C2(n6271), .ZN(U2886) );
  AND2_X1 U5750 ( .A1(n4726), .A2(n4738), .ZN(n4616) );
  INV_X1 U5751 ( .A(n6043), .ZN(n4727) );
  INV_X1 U5752 ( .A(n5150), .ZN(n4617) );
  OAI21_X1 U5753 ( .B1(n4619), .B2(n6497), .A(n4617), .ZN(n4623) );
  NAND2_X1 U5754 ( .A1(n4483), .A2(n6039), .ZN(n6056) );
  NOR2_X1 U5755 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5035) );
  AND2_X1 U5756 ( .A1(n5035), .A2(n6811), .ZN(n4837) );
  AND2_X1 U5757 ( .A1(n4837), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4620)
         );
  AOI21_X1 U5758 ( .B1(n4834), .B2(n3552), .A(n4620), .ZN(n4622) );
  INV_X1 U5759 ( .A(n4622), .ZN(n4618) );
  INV_X1 U5760 ( .A(n4620), .ZN(n4645) );
  OAI22_X1 U5761 ( .A1(n4993), .A2(n6495), .B1(n6494), .B2(n4645), .ZN(n4621)
         );
  AOI21_X1 U5762 ( .B1(n6502), .B2(n4647), .A(n4621), .ZN(n4626) );
  NAND2_X1 U5763 ( .A1(n4623), .A2(n4622), .ZN(n4624) );
  NAND2_X1 U5764 ( .A1(n4648), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4625) );
  OAI211_X1 U5765 ( .C1(n4651), .C2(n6505), .A(n4626), .B(n4625), .ZN(U3028)
         );
  INV_X1 U5766 ( .A(n6561), .ZN(n6084) );
  INV_X1 U5767 ( .A(n6527), .ZN(n6556) );
  OAI22_X1 U5768 ( .A1(n4993), .A2(n6556), .B1(n6555), .B2(n4645), .ZN(n4627)
         );
  AOI21_X1 U5769 ( .B1(n6084), .B2(n4647), .A(n4627), .ZN(n4629) );
  NAND2_X1 U5770 ( .A1(n4648), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4628) );
  OAI211_X1 U5771 ( .C1(n4651), .C2(n6530), .A(n4629), .B(n4628), .ZN(U3033)
         );
  INV_X1 U5772 ( .A(n6512), .ZN(n6485) );
  OAI22_X1 U5773 ( .A1(n4993), .A2(n6489), .B1(n6511), .B2(n4645), .ZN(n4630)
         );
  AOI21_X1 U5774 ( .B1(n6485), .B2(n4647), .A(n4630), .ZN(n4632) );
  NAND2_X1 U5775 ( .A1(n4648), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4631) );
  OAI211_X1 U5776 ( .C1(n4651), .C2(n6517), .A(n4632), .B(n4631), .ZN(U3031)
         );
  INV_X1 U5777 ( .A(n6573), .ZN(n6096) );
  INV_X1 U5778 ( .A(n6540), .ZN(n6564) );
  OAI22_X1 U5779 ( .A1(n4993), .A2(n6564), .B1(n6563), .B2(n4645), .ZN(n4633)
         );
  AOI21_X1 U5780 ( .B1(n6096), .B2(n4647), .A(n4633), .ZN(n4635) );
  NAND2_X1 U5781 ( .A1(n4648), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4634) );
  OAI211_X1 U5782 ( .C1(n4651), .C2(n6543), .A(n4635), .B(n4634), .ZN(U3035)
         );
  INV_X1 U5783 ( .A(n6532), .ZN(n6088) );
  OAI22_X1 U5784 ( .A1(n4993), .A2(n6091), .B1(n6531), .B2(n4645), .ZN(n4636)
         );
  AOI21_X1 U5785 ( .B1(n6088), .B2(n4647), .A(n4636), .ZN(n4638) );
  NAND2_X1 U5786 ( .A1(n4648), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4637) );
  OAI211_X1 U5787 ( .C1(n4651), .C2(n6537), .A(n4638), .B(n4637), .ZN(U3034)
         );
  INV_X1 U5788 ( .A(n6678), .ZN(n6477) );
  OAI22_X1 U5789 ( .A1(n4993), .A2(n6681), .B1(n6676), .B2(n4645), .ZN(n4639)
         );
  AOI21_X1 U5790 ( .B1(n6477), .B2(n4647), .A(n4639), .ZN(n4641) );
  NAND2_X1 U5791 ( .A1(n4648), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4640) );
  OAI211_X1 U5792 ( .C1(n4651), .C2(n6682), .A(n4641), .B(n4640), .ZN(U3030)
         );
  OAI22_X1 U5793 ( .A1(n4993), .A2(n6519), .B1(n6518), .B2(n4645), .ZN(n4642)
         );
  AOI21_X1 U5794 ( .B1(n6522), .B2(n4647), .A(n4642), .ZN(n4644) );
  NAND2_X1 U5795 ( .A1(n4648), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4643) );
  OAI211_X1 U5796 ( .C1(n4651), .C2(n6525), .A(n4644), .B(n4643), .ZN(U3032)
         );
  INV_X1 U5797 ( .A(n6550), .ZN(n6473) );
  OAI22_X1 U5798 ( .A1(n4993), .A2(n6545), .B1(n6544), .B2(n4645), .ZN(n4646)
         );
  AOI21_X1 U5799 ( .B1(n6473), .B2(n4647), .A(n4646), .ZN(n4650) );
  NAND2_X1 U5800 ( .A1(n4648), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4649) );
  OAI211_X1 U5801 ( .C1(n4651), .C2(n6510), .A(n4650), .B(n4649), .ZN(U3029)
         );
  INV_X1 U5802 ( .A(n4654), .ZN(n6423) );
  NAND2_X1 U5803 ( .A1(n6423), .A2(n6340), .ZN(n4658) );
  INV_X1 U5804 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4655) );
  NOR2_X1 U5805 ( .A1(n6435), .A2(n4655), .ZN(n6420) );
  NOR2_X1 U5806 ( .A1(n6345), .A2(n5547), .ZN(n4656) );
  AOI211_X1 U5807 ( .C1(n6336), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6420), 
        .B(n4656), .ZN(n4657) );
  OAI211_X1 U5808 ( .C1(n5779), .C2(n5557), .A(n4658), .B(n4657), .ZN(U2983)
         );
  INV_X1 U5809 ( .A(n4726), .ZN(n4661) );
  NAND2_X1 U5810 ( .A1(n4670), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4668) );
  NAND2_X1 U5811 ( .A1(n6055), .A2(n6042), .ZN(n6498) );
  NAND3_X1 U5812 ( .A1(n4668), .A2(n5033), .A3(n6498), .ZN(n4718) );
  AOI222_X1 U5813 ( .A1(n4662), .A2(n5552), .B1(n4661), .B2(n5150), .C1(n4718), 
        .C2(n6666), .ZN(n4665) );
  INV_X1 U5814 ( .A(n6443), .ZN(n4664) );
  NAND2_X1 U5815 ( .A1(n4664), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4663) );
  OAI21_X1 U5816 ( .B1(n4665), .B2(n4664), .A(n4663), .ZN(U3462) );
  AND3_X1 U5817 ( .A1(n4889), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4758) );
  INV_X1 U5818 ( .A(n4483), .ZN(n5563) );
  NAND2_X1 U5819 ( .A1(n5563), .A2(n6039), .ZN(n5158) );
  INV_X1 U5820 ( .A(n5158), .ZN(n4762) );
  NAND2_X1 U5821 ( .A1(n4762), .A2(n5036), .ZN(n4666) );
  NAND2_X1 U5822 ( .A1(n4758), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4693) );
  AOI21_X1 U5823 ( .B1(n4666), .B2(n4693), .A(n6497), .ZN(n4667) );
  AOI21_X1 U5824 ( .B1(n4758), .B2(STATE2_REG_2__SCAN_IN), .A(n4667), .ZN(
        n4698) );
  NOR2_X1 U5825 ( .A1(n4668), .A2(n6497), .ZN(n4669) );
  NAND2_X1 U5826 ( .A1(n4692), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4673)
         );
  OAI22_X1 U5827 ( .A1(n4985), .A2(n6091), .B1(n6531), .B2(n4693), .ZN(n4671)
         );
  AOI21_X1 U5828 ( .B1(n6088), .B2(n4695), .A(n4671), .ZN(n4672) );
  OAI211_X1 U5829 ( .C1(n4698), .C2(n6537), .A(n4673), .B(n4672), .ZN(U3130)
         );
  NAND2_X1 U5830 ( .A1(n4692), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4676)
         );
  OAI22_X1 U5831 ( .A1(n4985), .A2(n6556), .B1(n6555), .B2(n4693), .ZN(n4674)
         );
  AOI21_X1 U5832 ( .B1(n6084), .B2(n4695), .A(n4674), .ZN(n4675) );
  OAI211_X1 U5833 ( .C1(n4698), .C2(n6530), .A(n4676), .B(n4675), .ZN(U3129)
         );
  NAND2_X1 U5834 ( .A1(n4692), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4679)
         );
  OAI22_X1 U5835 ( .A1(n4985), .A2(n6564), .B1(n6563), .B2(n4693), .ZN(n4677)
         );
  AOI21_X1 U5836 ( .B1(n6096), .B2(n4695), .A(n4677), .ZN(n4678) );
  OAI211_X1 U5837 ( .C1(n4698), .C2(n6543), .A(n4679), .B(n4678), .ZN(U3131)
         );
  NAND2_X1 U5838 ( .A1(n4692), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4682)
         );
  OAI22_X1 U5839 ( .A1(n4985), .A2(n6681), .B1(n6676), .B2(n4693), .ZN(n4680)
         );
  AOI21_X1 U5840 ( .B1(n6477), .B2(n4695), .A(n4680), .ZN(n4681) );
  OAI211_X1 U5841 ( .C1(n4698), .C2(n6682), .A(n4682), .B(n4681), .ZN(U3126)
         );
  NAND2_X1 U5842 ( .A1(n4692), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4685)
         );
  OAI22_X1 U5843 ( .A1(n4985), .A2(n6545), .B1(n6544), .B2(n4693), .ZN(n4683)
         );
  AOI21_X1 U5844 ( .B1(n6473), .B2(n4695), .A(n4683), .ZN(n4684) );
  OAI211_X1 U5845 ( .C1(n4698), .C2(n6510), .A(n4685), .B(n4684), .ZN(U3125)
         );
  NAND2_X1 U5846 ( .A1(n4692), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4688)
         );
  OAI22_X1 U5847 ( .A1(n4985), .A2(n6489), .B1(n6511), .B2(n4693), .ZN(n4686)
         );
  AOI21_X1 U5848 ( .B1(n6485), .B2(n4695), .A(n4686), .ZN(n4687) );
  OAI211_X1 U5849 ( .C1(n4698), .C2(n6517), .A(n4688), .B(n4687), .ZN(U3127)
         );
  NAND2_X1 U5850 ( .A1(n4692), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4691)
         );
  OAI22_X1 U5851 ( .A1(n4985), .A2(n6519), .B1(n6518), .B2(n4693), .ZN(n4689)
         );
  AOI21_X1 U5852 ( .B1(n6522), .B2(n4695), .A(n4689), .ZN(n4690) );
  OAI211_X1 U5853 ( .C1(n4698), .C2(n6525), .A(n4691), .B(n4690), .ZN(U3128)
         );
  NAND2_X1 U5854 ( .A1(n4692), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4697)
         );
  OAI22_X1 U5855 ( .A1(n4985), .A2(n6495), .B1(n6494), .B2(n4693), .ZN(n4694)
         );
  AOI21_X1 U5856 ( .B1(n6502), .B2(n4695), .A(n4694), .ZN(n4696) );
  OAI211_X1 U5857 ( .C1(n4698), .C2(n6505), .A(n4697), .B(n4696), .ZN(U3124)
         );
  XNOR2_X1 U5858 ( .A(n4700), .B(n4699), .ZN(n6322) );
  INV_X1 U5859 ( .A(n6322), .ZN(n6200) );
  OR2_X1 U5860 ( .A1(n4703), .A2(n4702), .ZN(n4704) );
  AND2_X1 U5861 ( .A1(n4701), .A2(n4704), .ZN(n6397) );
  AOI22_X1 U5862 ( .A1(n6239), .A2(n6397), .B1(EBX_REG_6__SCAN_IN), .B2(n5592), 
        .ZN(n4705) );
  OAI21_X1 U5863 ( .B1(n6200), .B2(n5609), .A(n4705), .ZN(U2853) );
  OAI222_X1 U5864 ( .A1(n5658), .A2(n6200), .B1(n4711), .B2(n4706), .C1(n6249), 
        .C2(n3589), .ZN(U2885) );
  XOR2_X1 U5865 ( .A(n4707), .B(n4825), .Z(n5142) );
  INV_X1 U5866 ( .A(n5142), .ZN(n5528) );
  OAI222_X1 U5867 ( .A1(n5658), .A2(n5528), .B1(n4711), .B2(n6750), .C1(n6249), 
        .C2(n4319), .ZN(U2884) );
  INV_X1 U5868 ( .A(n4712), .ZN(n4714) );
  NAND2_X1 U5869 ( .A1(n4825), .A2(n4707), .ZN(n4713) );
  AOI21_X1 U5870 ( .B1(n4714), .B2(n4713), .A(n4792), .ZN(n5199) );
  INV_X1 U5871 ( .A(n5199), .ZN(n5515) );
  XNOR2_X1 U5872 ( .A(n4828), .B(n4830), .ZN(n6372) );
  AOI22_X1 U5873 ( .A1(n6239), .A2(n6372), .B1(EBX_REG_8__SCAN_IN), .B2(n5592), 
        .ZN(n4715) );
  OAI21_X1 U5874 ( .B1(n5515), .B2(n5609), .A(n4715), .ZN(U2851) );
  AOI22_X1 U5875 ( .A1(n6246), .A2(DATAI_8_), .B1(n5656), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4716) );
  OAI21_X1 U5876 ( .B1(n5515), .B2(n5658), .A(n4716), .ZN(U2883) );
  NAND2_X1 U5877 ( .A1(n4727), .A2(n6042), .ZN(n4717) );
  OAI21_X1 U5878 ( .B1(n4718), .B2(n4717), .A(n6666), .ZN(n4724) );
  NOR2_X1 U5879 ( .A1(n4720), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6460)
         );
  AOI21_X1 U5880 ( .B1(n4987), .B2(n3552), .A(n6460), .ZN(n4723) );
  INV_X1 U5881 ( .A(n4723), .ZN(n4722) );
  NAND3_X1 U5882 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6811), .A3(n4895), .ZN(n4989) );
  AOI21_X1 U5883 ( .B1(n4989), .B2(n6497), .A(n5038), .ZN(n4721) );
  INV_X1 U5884 ( .A(n6464), .ZN(n4732) );
  INV_X1 U5885 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6697) );
  OAI22_X1 U5886 ( .A1(n4724), .A2(n4723), .B1(n4989), .B2(n6575), .ZN(n6462)
         );
  NAND2_X1 U5887 ( .A1(n4726), .A2(n4922), .ZN(n4725) );
  AND2_X1 U5888 ( .A1(n4726), .A2(n6054), .ZN(n4728) );
  AOI22_X1 U5889 ( .A1(n6461), .A2(n6540), .B1(n6460), .B2(n5112), .ZN(n4729)
         );
  OAI21_X1 U5890 ( .B1(n6467), .B2(n6573), .A(n4729), .ZN(n4730) );
  AOI21_X1 U5891 ( .B1(n6462), .B2(n6568), .A(n4730), .ZN(n4731) );
  OAI21_X1 U5892 ( .B1(n4732), .B2(n6697), .A(n4731), .ZN(U3051) );
  NAND3_X1 U5893 ( .A1(n6055), .A2(STATEBS16_REG_SCAN_IN), .A3(n4738), .ZN(
        n4733) );
  NAND2_X1 U5894 ( .A1(n4733), .A2(n6666), .ZN(n4743) );
  INV_X1 U5895 ( .A(n4743), .ZN(n4736) );
  OR2_X1 U5896 ( .A1(n5158), .A2(n4734), .ZN(n5149) );
  NOR2_X1 U5897 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4735) );
  NAND2_X1 U5898 ( .A1(n4735), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4740) );
  OR2_X1 U5899 ( .A1(n4740), .A2(n5152), .ZN(n4778) );
  OAI21_X1 U5900 ( .B1(n5149), .B2(n6490), .A(n4778), .ZN(n4742) );
  INV_X1 U5901 ( .A(n4740), .ZN(n5153) );
  NOR2_X1 U5902 ( .A1(n4480), .A2(n5043), .ZN(n4737) );
  OAI22_X1 U5903 ( .A1(n5189), .A2(n6678), .B1(n6676), .B2(n4778), .ZN(n4739)
         );
  AOI21_X1 U5904 ( .B1(n6447), .B2(n6484), .A(n4739), .ZN(n4745) );
  AOI21_X1 U5905 ( .B1(n6497), .B2(n4740), .A(n5038), .ZN(n4741) );
  NAND2_X1 U5906 ( .A1(n4780), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4744) );
  OAI211_X1 U5907 ( .C1(n4783), .C2(n6682), .A(n4745), .B(n4744), .ZN(U3062)
         );
  OAI22_X1 U5908 ( .A1(n5189), .A2(n5119), .B1(n6494), .B2(n4778), .ZN(n4746)
         );
  AOI21_X1 U5909 ( .B1(n5117), .B2(n6484), .A(n4746), .ZN(n4748) );
  NAND2_X1 U5910 ( .A1(n4780), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4747) );
  OAI211_X1 U5911 ( .C1(n4783), .C2(n6505), .A(n4748), .B(n4747), .ZN(U3060)
         );
  OAI22_X1 U5912 ( .A1(n5189), .A2(n6512), .B1(n6511), .B2(n4778), .ZN(n4749)
         );
  AOI21_X1 U5913 ( .B1(n6514), .B2(n6484), .A(n4749), .ZN(n4751) );
  NAND2_X1 U5914 ( .A1(n4780), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4750) );
  OAI211_X1 U5915 ( .C1(n4783), .C2(n6517), .A(n4751), .B(n4750), .ZN(U3063)
         );
  OAI22_X1 U5916 ( .A1(n5189), .A2(n6550), .B1(n6544), .B2(n4778), .ZN(n4752)
         );
  AOI21_X1 U5917 ( .B1(n6507), .B2(n6484), .A(n4752), .ZN(n4754) );
  NAND2_X1 U5918 ( .A1(n4780), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4753) );
  OAI211_X1 U5919 ( .C1(n4783), .C2(n6510), .A(n4754), .B(n4753), .ZN(U3061)
         );
  OAI22_X1 U5920 ( .A1(n5189), .A2(n6455), .B1(n6518), .B2(n4778), .ZN(n4755)
         );
  AOI21_X1 U5921 ( .B1(n6451), .B2(n6484), .A(n4755), .ZN(n4757) );
  NAND2_X1 U5922 ( .A1(n4780), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4756) );
  OAI211_X1 U5923 ( .C1(n4783), .C2(n6525), .A(n4757), .B(n4756), .ZN(U3064)
         );
  AOI21_X1 U5924 ( .B1(n4823), .B2(n6565), .A(n6104), .ZN(n4761) );
  OAI21_X1 U5925 ( .B1(n5158), .B2(n4923), .A(n6666), .ZN(n4760) );
  NAND2_X1 U5926 ( .A1(n4758), .A2(n5152), .ZN(n4818) );
  NOR2_X1 U5927 ( .A1(n4763), .A2(n6575), .ZN(n5155) );
  INV_X1 U5928 ( .A(n5092), .ZN(n4994) );
  AOI21_X1 U5929 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4994), .A(n4926), .ZN(
        n4836) );
  OAI21_X1 U5930 ( .B1(n6065), .B2(n6575), .A(n4836), .ZN(n6059) );
  AOI211_X1 U5931 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4818), .A(n5155), .B(
        n6059), .ZN(n4759) );
  NAND2_X1 U5932 ( .A1(n4820), .A2(n6502), .ZN(n4769) );
  AND2_X1 U5933 ( .A1(n5552), .A2(n6666), .ZN(n6067) );
  NAND2_X1 U5934 ( .A1(n6067), .A2(n4762), .ZN(n4765) );
  NAND2_X1 U5935 ( .A1(n4763), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5086) );
  NOR2_X1 U5936 ( .A1(n5086), .A2(n4994), .ZN(n5161) );
  NAND2_X1 U5937 ( .A1(n5161), .A2(n6065), .ZN(n4764) );
  INV_X1 U5938 ( .A(n4817), .ZN(n4767) );
  INV_X1 U5939 ( .A(n4818), .ZN(n4766) );
  AOI22_X1 U5940 ( .A1(n4767), .A2(n6468), .B1(n6469), .B2(n4766), .ZN(n4768)
         );
  OAI211_X1 U5941 ( .C1(n4823), .C2(n6495), .A(n4769), .B(n4768), .ZN(n4770)
         );
  AOI21_X1 U5942 ( .B1(n4816), .B2(INSTQUEUE_REG_12__0__SCAN_IN), .A(n4770), 
        .ZN(n4771) );
  INV_X1 U5943 ( .A(n4771), .ZN(U3116) );
  OAI22_X1 U5944 ( .A1(n5189), .A2(n6532), .B1(n6531), .B2(n4778), .ZN(n4772)
         );
  AOI21_X1 U5945 ( .B1(n6534), .B2(n6484), .A(n4772), .ZN(n4774) );
  NAND2_X1 U5946 ( .A1(n4780), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4773) );
  OAI211_X1 U5947 ( .C1(n4783), .C2(n6537), .A(n4774), .B(n4773), .ZN(U3066)
         );
  OAI22_X1 U5948 ( .A1(n5189), .A2(n6561), .B1(n6555), .B2(n4778), .ZN(n4775)
         );
  AOI21_X1 U5949 ( .B1(n6527), .B2(n6484), .A(n4775), .ZN(n4777) );
  NAND2_X1 U5950 ( .A1(n4780), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4776) );
  OAI211_X1 U5951 ( .C1(n4783), .C2(n6530), .A(n4777), .B(n4776), .ZN(U3065)
         );
  OAI22_X1 U5952 ( .A1(n5189), .A2(n6573), .B1(n6563), .B2(n4778), .ZN(n4779)
         );
  AOI21_X1 U5953 ( .B1(n6540), .B2(n6484), .A(n4779), .ZN(n4782) );
  NAND2_X1 U5954 ( .A1(n4780), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4781) );
  OAI211_X1 U5955 ( .C1(n4783), .C2(n6543), .A(n4782), .B(n4781), .ZN(U3067)
         );
  INV_X1 U5956 ( .A(n6462), .ZN(n4790) );
  AOI22_X1 U5957 ( .A1(n6461), .A2(n5117), .B1(n6460), .B2(n6469), .ZN(n4784)
         );
  OAI21_X1 U5958 ( .B1(n5119), .B2(n6467), .A(n4784), .ZN(n4785) );
  AOI21_X1 U5959 ( .B1(n6464), .B2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4785), 
        .ZN(n4786) );
  OAI21_X1 U5960 ( .B1(n4790), .B2(n6505), .A(n4786), .ZN(U3044) );
  AOI22_X1 U5961 ( .A1(n6461), .A2(n6514), .B1(n6460), .B2(n6483), .ZN(n4787)
         );
  OAI21_X1 U5962 ( .B1(n6467), .B2(n6512), .A(n4787), .ZN(n4788) );
  AOI21_X1 U5963 ( .B1(n6464), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4788), 
        .ZN(n4789) );
  OAI21_X1 U5964 ( .B1(n4790), .B2(n6517), .A(n4789), .ZN(U3047) );
  NAND2_X1 U5965 ( .A1(n4792), .A2(n4791), .ZN(n5145) );
  OR2_X1 U5966 ( .A1(n4792), .A2(n4791), .ZN(n4793) );
  NAND2_X1 U5967 ( .A1(n5145), .A2(n4793), .ZN(n6187) );
  AOI22_X1 U5968 ( .A1(n6246), .A2(DATAI_9_), .B1(n5656), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4794) );
  OAI21_X1 U5969 ( .B1(n6187), .B2(n5658), .A(n4794), .ZN(U2882) );
  NAND2_X1 U5970 ( .A1(n4701), .A2(n4795), .ZN(n4796) );
  NAND2_X1 U5971 ( .A1(n4828), .A2(n4796), .ZN(n5516) );
  INV_X1 U5972 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4797) );
  OAI222_X1 U5973 ( .A1(n5516), .A2(n5608), .B1(n4797), .B2(n6243), .C1(n5609), 
        .C2(n5528), .ZN(U2852) );
  NAND2_X1 U5974 ( .A1(n4816), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4800)
         );
  OAI22_X1 U5975 ( .A1(n6676), .A2(n4818), .B1(n4817), .B2(n6682), .ZN(n4798)
         );
  AOI21_X1 U5976 ( .B1(n4820), .B2(n6477), .A(n4798), .ZN(n4799) );
  OAI211_X1 U5977 ( .C1(n4823), .C2(n6681), .A(n4800), .B(n4799), .ZN(U3118)
         );
  NAND2_X1 U5978 ( .A1(n4816), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4803)
         );
  OAI22_X1 U5979 ( .A1(n6555), .A2(n4818), .B1(n4817), .B2(n6530), .ZN(n4801)
         );
  AOI21_X1 U5980 ( .B1(n4820), .B2(n6084), .A(n4801), .ZN(n4802) );
  OAI211_X1 U5981 ( .C1(n4823), .C2(n6556), .A(n4803), .B(n4802), .ZN(U3121)
         );
  NAND2_X1 U5982 ( .A1(n4816), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4806)
         );
  OAI22_X1 U5983 ( .A1(n6518), .A2(n4818), .B1(n4817), .B2(n6525), .ZN(n4804)
         );
  AOI21_X1 U5984 ( .B1(n4820), .B2(n6522), .A(n4804), .ZN(n4805) );
  OAI211_X1 U5985 ( .C1(n4823), .C2(n6519), .A(n4806), .B(n4805), .ZN(U3120)
         );
  NAND2_X1 U5986 ( .A1(n4816), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4809)
         );
  OAI22_X1 U5987 ( .A1(n6531), .A2(n4818), .B1(n4817), .B2(n6537), .ZN(n4807)
         );
  AOI21_X1 U5988 ( .B1(n4820), .B2(n6088), .A(n4807), .ZN(n4808) );
  OAI211_X1 U5989 ( .C1(n4823), .C2(n6091), .A(n4809), .B(n4808), .ZN(U3122)
         );
  NAND2_X1 U5990 ( .A1(n4816), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4812)
         );
  OAI22_X1 U5991 ( .A1(n6563), .A2(n4818), .B1(n4817), .B2(n6543), .ZN(n4810)
         );
  AOI21_X1 U5992 ( .B1(n4820), .B2(n6096), .A(n4810), .ZN(n4811) );
  OAI211_X1 U5993 ( .C1(n4823), .C2(n6564), .A(n4812), .B(n4811), .ZN(U3123)
         );
  NAND2_X1 U5994 ( .A1(n4816), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4815)
         );
  OAI22_X1 U5995 ( .A1(n6544), .A2(n4818), .B1(n4817), .B2(n6510), .ZN(n4813)
         );
  AOI21_X1 U5996 ( .B1(n4820), .B2(n6473), .A(n4813), .ZN(n4814) );
  OAI211_X1 U5997 ( .C1(n4823), .C2(n6545), .A(n4815), .B(n4814), .ZN(U3117)
         );
  NAND2_X1 U5998 ( .A1(n4816), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4822)
         );
  OAI22_X1 U5999 ( .A1(n6511), .A2(n4818), .B1(n4817), .B2(n6517), .ZN(n4819)
         );
  AOI21_X1 U6000 ( .B1(n4820), .B2(n6485), .A(n4819), .ZN(n4821) );
  OAI211_X1 U6001 ( .C1(n4823), .C2(n6489), .A(n4822), .B(n4821), .ZN(U3119)
         );
  NAND2_X1 U6002 ( .A1(n4825), .A2(n4824), .ZN(n6174) );
  XNOR2_X1 U6003 ( .A(n6174), .B(n4826), .ZN(n5821) );
  INV_X1 U6004 ( .A(n5821), .ZN(n6160) );
  AOI22_X1 U6005 ( .A1(n6246), .A2(DATAI_12_), .B1(n5656), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4827) );
  OAI21_X1 U6006 ( .B1(n6160), .B2(n5658), .A(n4827), .ZN(U2879) );
  AOI21_X1 U6007 ( .B1(n3103), .B2(n4830), .A(n4829), .ZN(n4831) );
  OR2_X1 U6008 ( .A1(n4831), .A2(n5192), .ZN(n6359) );
  INV_X1 U6009 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4832) );
  OAI222_X1 U6010 ( .A1(n6359), .A2(n5608), .B1(n4832), .B2(n6243), .C1(n6187), 
        .C2(n5609), .ZN(U2850) );
  AOI21_X1 U6011 ( .B1(n4872), .B2(n4833), .A(n6104), .ZN(n4835) );
  NOR3_X1 U6012 ( .A1(n4835), .A2(n4834), .A3(n6497), .ZN(n4839) );
  INV_X1 U6013 ( .A(n6065), .ZN(n5160) );
  OAI21_X1 U6014 ( .B1(n6575), .B2(n5160), .A(n4836), .ZN(n5154) );
  AND2_X1 U6015 ( .A1(n4837), .A2(n5152), .ZN(n4869) );
  OAI21_X1 U6016 ( .B1(n4869), .B2(n4986), .A(n5086), .ZN(n4838) );
  NOR3_X2 U6017 ( .A1(n4839), .A2(n5154), .A3(n4838), .ZN(n4877) );
  INV_X1 U6018 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4845) );
  AND2_X1 U6019 ( .A1(n5155), .A2(n5092), .ZN(n6064) );
  NAND2_X1 U6020 ( .A1(n5160), .A2(n6064), .ZN(n4840) );
  OAI21_X1 U6021 ( .B1(n4841), .B2(n6497), .A(n4840), .ZN(n4870) );
  AOI22_X1 U6022 ( .A1(n6452), .A2(n4870), .B1(n6450), .B2(n4869), .ZN(n4842)
         );
  OAI21_X1 U6023 ( .B1(n4872), .B2(n6519), .A(n4842), .ZN(n4843) );
  AOI21_X1 U6024 ( .B1(n6522), .B2(n4874), .A(n4843), .ZN(n4844) );
  OAI21_X1 U6025 ( .B1(n4877), .B2(n4845), .A(n4844), .ZN(U3024) );
  INV_X1 U6026 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6731) );
  AOI22_X1 U6027 ( .A1(n6552), .A2(n4870), .B1(n6476), .B2(n4869), .ZN(n4846)
         );
  OAI21_X1 U6028 ( .B1(n4872), .B2(n6681), .A(n4846), .ZN(n4847) );
  AOI21_X1 U6029 ( .B1(n6477), .B2(n4874), .A(n4847), .ZN(n4848) );
  OAI21_X1 U6030 ( .B1(n4877), .B2(n6731), .A(n4848), .ZN(U3022) );
  INV_X1 U6031 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4852) );
  AOI22_X1 U6032 ( .A1(n6463), .A2(n4870), .B1(n6459), .B2(n4869), .ZN(n4849)
         );
  OAI21_X1 U6033 ( .B1(n4872), .B2(n6091), .A(n4849), .ZN(n4850) );
  AOI21_X1 U6034 ( .B1(n6088), .B2(n4874), .A(n4850), .ZN(n4851) );
  OAI21_X1 U6035 ( .B1(n4877), .B2(n4852), .A(n4851), .ZN(U3026) );
  INV_X1 U6036 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4856) );
  AOI22_X1 U6037 ( .A1(n6568), .A2(n4870), .B1(n5112), .B2(n4869), .ZN(n4853)
         );
  OAI21_X1 U6038 ( .B1(n4872), .B2(n6564), .A(n4853), .ZN(n4854) );
  AOI21_X1 U6039 ( .B1(n6096), .B2(n4874), .A(n4854), .ZN(n4855) );
  OAI21_X1 U6040 ( .B1(n4877), .B2(n4856), .A(n4855), .ZN(U3027) );
  INV_X1 U6041 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4860) );
  AOI22_X1 U6042 ( .A1(n6547), .A2(n4870), .B1(n6472), .B2(n4869), .ZN(n4857)
         );
  OAI21_X1 U6043 ( .B1(n4872), .B2(n6545), .A(n4857), .ZN(n4858) );
  AOI21_X1 U6044 ( .B1(n6473), .B2(n4874), .A(n4858), .ZN(n4859) );
  OAI21_X1 U6045 ( .B1(n4877), .B2(n4860), .A(n4859), .ZN(U3021) );
  INV_X1 U6046 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4864) );
  AOI22_X1 U6047 ( .A1(n6558), .A2(n4870), .B1(n6456), .B2(n4869), .ZN(n4861)
         );
  OAI21_X1 U6048 ( .B1(n4872), .B2(n6556), .A(n4861), .ZN(n4862) );
  AOI21_X1 U6049 ( .B1(n6084), .B2(n4874), .A(n4862), .ZN(n4863) );
  OAI21_X1 U6050 ( .B1(n4877), .B2(n4864), .A(n4863), .ZN(U3025) );
  INV_X1 U6051 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4868) );
  AOI22_X1 U6052 ( .A1(n6480), .A2(n4870), .B1(n6483), .B2(n4869), .ZN(n4865)
         );
  OAI21_X1 U6053 ( .B1(n4872), .B2(n6489), .A(n4865), .ZN(n4866) );
  AOI21_X1 U6054 ( .B1(n6485), .B2(n4874), .A(n4866), .ZN(n4867) );
  OAI21_X1 U6055 ( .B1(n4877), .B2(n4868), .A(n4867), .ZN(U3023) );
  INV_X1 U6056 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4876) );
  AOI22_X1 U6057 ( .A1(n6468), .A2(n4870), .B1(n6469), .B2(n4869), .ZN(n4871)
         );
  OAI21_X1 U6058 ( .B1(n4872), .B2(n6495), .A(n4871), .ZN(n4873) );
  AOI21_X1 U6059 ( .B1(n6502), .B2(n4874), .A(n4873), .ZN(n4875) );
  OAI21_X1 U6060 ( .B1(n4877), .B2(n4876), .A(n4875), .ZN(U3020) );
  OAI21_X1 U6061 ( .B1(n4880), .B2(n4879), .A(n4878), .ZN(n6402) );
  NAND2_X1 U6062 ( .A1(n3009), .A2(REIP_REG_5__SCAN_IN), .ZN(n6405) );
  OAI21_X1 U6063 ( .B1(n5833), .B2(n5535), .A(n6405), .ZN(n4882) );
  NOR2_X1 U6064 ( .A1(n5529), .A2(n5779), .ZN(n4881) );
  AOI211_X1 U6065 ( .C1(n6312), .C2(n5533), .A(n4882), .B(n4881), .ZN(n4883)
         );
  OAI21_X1 U6066 ( .B1(n6316), .B2(n6402), .A(n4883), .ZN(U2981) );
  NAND2_X1 U6067 ( .A1(n4884), .A2(n6104), .ZN(n5296) );
  INV_X1 U6068 ( .A(n5296), .ZN(n4885) );
  NAND2_X1 U6069 ( .A1(n5269), .A2(n4885), .ZN(n5278) );
  INV_X1 U6070 ( .A(n4896), .ZN(n4898) );
  NAND3_X1 U6071 ( .A1(n4887), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n4886), .ZN(n4888) );
  INV_X1 U6072 ( .A(n4888), .ZN(n4893) );
  AOI22_X1 U6073 ( .A1(n4891), .A2(n4890), .B1(n4889), .B2(n4888), .ZN(n4892)
         );
  AOI21_X1 U6074 ( .B1(n4893), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n4892), 
        .ZN(n4894) );
  OAI21_X1 U6075 ( .B1(n4896), .B2(n4895), .A(n4894), .ZN(n4897) );
  OAI21_X1 U6076 ( .B1(n4898), .B2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n4897), 
        .ZN(n4899) );
  AOI222_X1 U6077 ( .A1(n4900), .A2(n6811), .B1(n4900), .B2(n4899), .C1(n6811), 
        .C2(n4899), .ZN(n4905) );
  NOR3_X1 U6078 ( .A1(n5530), .A2(n5269), .A3(n4901), .ZN(n4902) );
  NOR2_X1 U6079 ( .A1(n4902), .A2(READY_N), .ZN(n6669) );
  NOR2_X1 U6080 ( .A1(n4903), .A2(n6669), .ZN(n5248) );
  OAI21_X1 U6081 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n5248), 
        .ZN(n4904) );
  OAI21_X1 U6082 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n4905), .A(n4904), 
        .ZN(n4917) );
  INV_X1 U6083 ( .A(n4301), .ZN(n4906) );
  NOR2_X1 U6084 ( .A1(n4907), .A2(n4906), .ZN(n4908) );
  MUX2_X1 U6085 ( .A(n4909), .B(n4908), .S(n6581), .Z(n4913) );
  NAND2_X1 U6086 ( .A1(n4911), .A2(n4910), .ZN(n4912) );
  AND2_X1 U6087 ( .A1(n4913), .A2(n4912), .ZN(n5247) );
  NAND3_X1 U6088 ( .A1(n4915), .A2(n5247), .A3(n4914), .ZN(n4916) );
  OAI22_X1 U6089 ( .A1(n6574), .A2(n6587), .B1(n6263), .B2(n4884), .ZN(n4918)
         );
  OAI21_X1 U6090 ( .B1(n5278), .B2(n4919), .A(n4918), .ZN(n6592) );
  INV_X1 U6091 ( .A(n4920), .ZN(n6596) );
  OAI211_X1 U6092 ( .C1(n6592), .C2(n4986), .A(n4921), .B(n6596), .ZN(U3453)
         );
  INV_X1 U6093 ( .A(n6679), .ZN(n6521) );
  OAI21_X1 U6094 ( .B1(n6521), .B2(n6484), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4924) );
  NAND2_X1 U6095 ( .A1(n4956), .A2(n4923), .ZN(n6491) );
  NAND3_X1 U6096 ( .A1(n4924), .A2(n6666), .A3(n6491), .ZN(n4929) );
  AND2_X1 U6097 ( .A1(n5092), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4925) );
  NAND2_X1 U6098 ( .A1(n6500), .A2(n5152), .ZN(n4930) );
  AOI21_X1 U6099 ( .B1(n4930), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4928) );
  INV_X1 U6100 ( .A(n5155), .ZN(n4927) );
  NAND4_X1 U6101 ( .A1(n4929), .A2(n5088), .A3(n4928), .A4(n4927), .ZN(n6486)
         );
  NAND2_X1 U6102 ( .A1(n6484), .A2(n6096), .ZN(n4934) );
  INV_X1 U6103 ( .A(n4930), .ZN(n6482) );
  INV_X1 U6104 ( .A(n5552), .ZN(n6057) );
  NAND3_X1 U6105 ( .A1(n6057), .A2(n4956), .A3(n6666), .ZN(n4932) );
  INV_X1 U6106 ( .A(n5086), .ZN(n6060) );
  NAND3_X1 U6107 ( .A1(n6060), .A2(n4994), .A3(n6811), .ZN(n4931) );
  NAND2_X1 U6108 ( .A1(n4932), .A2(n4931), .ZN(n6481) );
  AOI22_X1 U6109 ( .A1(n5112), .A2(n6482), .B1(n6481), .B2(n6568), .ZN(n4933)
         );
  OAI211_X1 U6110 ( .C1(n6679), .C2(n6564), .A(n4934), .B(n4933), .ZN(n4935)
         );
  AOI21_X1 U6111 ( .B1(n6486), .B2(INSTQUEUE_REG_6__7__SCAN_IN), .A(n4935), 
        .ZN(n4936) );
  INV_X1 U6112 ( .A(n4936), .ZN(U3075) );
  NAND2_X1 U6113 ( .A1(n6484), .A2(n6088), .ZN(n4938) );
  AOI22_X1 U6114 ( .A1(n6459), .A2(n6482), .B1(n6481), .B2(n6463), .ZN(n4937)
         );
  OAI211_X1 U6115 ( .C1(n6679), .C2(n6091), .A(n4938), .B(n4937), .ZN(n4939)
         );
  AOI21_X1 U6116 ( .B1(n6486), .B2(INSTQUEUE_REG_6__6__SCAN_IN), .A(n4939), 
        .ZN(n4940) );
  INV_X1 U6117 ( .A(n4940), .ZN(U3074) );
  NAND2_X1 U6118 ( .A1(n6484), .A2(n6522), .ZN(n4942) );
  AOI22_X1 U6119 ( .A1(n6450), .A2(n6482), .B1(n6481), .B2(n6452), .ZN(n4941)
         );
  OAI211_X1 U6120 ( .C1(n6679), .C2(n6519), .A(n4942), .B(n4941), .ZN(n4943)
         );
  AOI21_X1 U6121 ( .B1(n6486), .B2(INSTQUEUE_REG_6__4__SCAN_IN), .A(n4943), 
        .ZN(n4944) );
  INV_X1 U6122 ( .A(n4944), .ZN(U3072) );
  NAND2_X1 U6123 ( .A1(n6484), .A2(n6084), .ZN(n4946) );
  AOI22_X1 U6124 ( .A1(n6456), .A2(n6482), .B1(n6481), .B2(n6558), .ZN(n4945)
         );
  OAI211_X1 U6125 ( .C1(n6679), .C2(n6556), .A(n4946), .B(n4945), .ZN(n4947)
         );
  AOI21_X1 U6126 ( .B1(n6486), .B2(INSTQUEUE_REG_6__5__SCAN_IN), .A(n4947), 
        .ZN(n4948) );
  INV_X1 U6127 ( .A(n4948), .ZN(U3073) );
  AOI21_X1 U6128 ( .B1(n4985), .B2(n4953), .A(n6104), .ZN(n4949) );
  NOR3_X1 U6129 ( .A1(n4949), .A2(n4956), .A3(n6497), .ZN(n4952) );
  INV_X1 U6130 ( .A(n5088), .ZN(n4990) );
  NOR2_X1 U6131 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4950), .ZN(n4954)
         );
  OAI21_X1 U6132 ( .B1(n4986), .B2(n4954), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n4951) );
  NAND2_X1 U6133 ( .A1(n4978), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4959)
         );
  INV_X1 U6134 ( .A(n4954), .ZN(n4980) );
  NOR3_X1 U6135 ( .A1(n5086), .A2(n5092), .A3(n6811), .ZN(n4955) );
  AOI21_X1 U6136 ( .B1(n6067), .B2(n4956), .A(n4955), .ZN(n4979) );
  OAI22_X1 U6137 ( .A1(n6676), .A2(n4980), .B1(n4979), .B2(n6682), .ZN(n4957)
         );
  AOI21_X1 U6138 ( .B1(n4982), .B2(n6447), .A(n4957), .ZN(n4958) );
  OAI211_X1 U6139 ( .C1(n4985), .C2(n6678), .A(n4959), .B(n4958), .ZN(U3134)
         );
  NAND2_X1 U6140 ( .A1(n4978), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4962)
         );
  OAI22_X1 U6141 ( .A1(n6511), .A2(n4980), .B1(n4979), .B2(n6517), .ZN(n4960)
         );
  AOI21_X1 U6142 ( .B1(n4982), .B2(n6514), .A(n4960), .ZN(n4961) );
  OAI211_X1 U6143 ( .C1(n4985), .C2(n6512), .A(n4962), .B(n4961), .ZN(U3135)
         );
  NAND2_X1 U6144 ( .A1(n4978), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4965)
         );
  OAI22_X1 U6145 ( .A1(n6563), .A2(n4980), .B1(n4979), .B2(n6543), .ZN(n4963)
         );
  AOI21_X1 U6146 ( .B1(n4982), .B2(n6540), .A(n4963), .ZN(n4964) );
  OAI211_X1 U6147 ( .C1(n4985), .C2(n6573), .A(n4965), .B(n4964), .ZN(U3139)
         );
  NAND2_X1 U6148 ( .A1(n4978), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4968)
         );
  OAI22_X1 U6149 ( .A1(n6531), .A2(n4980), .B1(n4979), .B2(n6537), .ZN(n4966)
         );
  AOI21_X1 U6150 ( .B1(n4982), .B2(n6534), .A(n4966), .ZN(n4967) );
  OAI211_X1 U6151 ( .C1(n4985), .C2(n6532), .A(n4968), .B(n4967), .ZN(U3138)
         );
  NAND2_X1 U6152 ( .A1(n4978), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4971)
         );
  OAI22_X1 U6153 ( .A1(n6518), .A2(n4980), .B1(n4979), .B2(n6525), .ZN(n4969)
         );
  AOI21_X1 U6154 ( .B1(n4982), .B2(n6451), .A(n4969), .ZN(n4970) );
  OAI211_X1 U6155 ( .C1(n4985), .C2(n6455), .A(n4971), .B(n4970), .ZN(U3136)
         );
  NAND2_X1 U6156 ( .A1(n4978), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4974)
         );
  OAI22_X1 U6157 ( .A1(n6494), .A2(n4980), .B1(n4979), .B2(n6505), .ZN(n4972)
         );
  AOI21_X1 U6158 ( .B1(n4982), .B2(n5117), .A(n4972), .ZN(n4973) );
  OAI211_X1 U6159 ( .C1(n4985), .C2(n5119), .A(n4974), .B(n4973), .ZN(U3132)
         );
  NAND2_X1 U6160 ( .A1(n4978), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4977)
         );
  OAI22_X1 U6161 ( .A1(n6544), .A2(n4980), .B1(n4979), .B2(n6510), .ZN(n4975)
         );
  AOI21_X1 U6162 ( .B1(n4982), .B2(n6507), .A(n4975), .ZN(n4976) );
  OAI211_X1 U6163 ( .C1(n4985), .C2(n6550), .A(n4977), .B(n4976), .ZN(U3133)
         );
  NAND2_X1 U6164 ( .A1(n4978), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4984)
         );
  OAI22_X1 U6165 ( .A1(n6555), .A2(n4980), .B1(n4979), .B2(n6530), .ZN(n4981)
         );
  AOI21_X1 U6166 ( .B1(n4982), .B2(n6527), .A(n4981), .ZN(n4983) );
  OAI211_X1 U6167 ( .C1(n4985), .C2(n6561), .A(n4984), .B(n4983), .ZN(U3137)
         );
  AOI21_X1 U6168 ( .B1(n4993), .B2(n6467), .A(n5150), .ZN(n4988) );
  OAI21_X1 U6169 ( .B1(n4988), .B2(n4987), .A(n4986), .ZN(n4992) );
  NOR2_X1 U6170 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4989), .ZN(n5025)
         );
  INV_X1 U6171 ( .A(n5025), .ZN(n4991) );
  INV_X1 U6172 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5000) );
  NAND3_X1 U6173 ( .A1(n5155), .A2(n4994), .A3(n6811), .ZN(n4995) );
  OAI21_X1 U6174 ( .B1(n4996), .B2(n6497), .A(n4995), .ZN(n5026) );
  AOI22_X1 U6175 ( .A1(n6452), .A2(n5026), .B1(n6450), .B2(n5025), .ZN(n4997)
         );
  OAI21_X1 U6176 ( .B1(n6467), .B2(n6519), .A(n4997), .ZN(n4998) );
  AOI21_X1 U6177 ( .B1(n5029), .B2(n6522), .A(n4998), .ZN(n4999) );
  OAI21_X1 U6178 ( .B1(n5032), .B2(n5000), .A(n4999), .ZN(U3040) );
  INV_X1 U6179 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5004) );
  AOI22_X1 U6180 ( .A1(n6552), .A2(n5026), .B1(n6476), .B2(n5025), .ZN(n5001)
         );
  OAI21_X1 U6181 ( .B1(n6467), .B2(n6681), .A(n5001), .ZN(n5002) );
  AOI21_X1 U6182 ( .B1(n5029), .B2(n6477), .A(n5002), .ZN(n5003) );
  OAI21_X1 U6183 ( .B1(n5032), .B2(n5004), .A(n5003), .ZN(U3038) );
  INV_X1 U6184 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5008) );
  AOI22_X1 U6185 ( .A1(n6547), .A2(n5026), .B1(n6472), .B2(n5025), .ZN(n5005)
         );
  OAI21_X1 U6186 ( .B1(n6467), .B2(n6545), .A(n5005), .ZN(n5006) );
  AOI21_X1 U6187 ( .B1(n5029), .B2(n6473), .A(n5006), .ZN(n5007) );
  OAI21_X1 U6188 ( .B1(n5032), .B2(n5008), .A(n5007), .ZN(U3037) );
  INV_X1 U6189 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5012) );
  AOI22_X1 U6190 ( .A1(n6568), .A2(n5026), .B1(n5112), .B2(n5025), .ZN(n5009)
         );
  OAI21_X1 U6191 ( .B1(n6467), .B2(n6564), .A(n5009), .ZN(n5010) );
  AOI21_X1 U6192 ( .B1(n5029), .B2(n6096), .A(n5010), .ZN(n5011) );
  OAI21_X1 U6193 ( .B1(n5032), .B2(n5012), .A(n5011), .ZN(U3043) );
  INV_X1 U6194 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5016) );
  AOI22_X1 U6195 ( .A1(n6558), .A2(n5026), .B1(n6456), .B2(n5025), .ZN(n5013)
         );
  OAI21_X1 U6196 ( .B1(n6467), .B2(n6556), .A(n5013), .ZN(n5014) );
  AOI21_X1 U6197 ( .B1(n5029), .B2(n6084), .A(n5014), .ZN(n5015) );
  OAI21_X1 U6198 ( .B1(n5032), .B2(n5016), .A(n5015), .ZN(U3041) );
  INV_X1 U6199 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5020) );
  AOI22_X1 U6200 ( .A1(n6480), .A2(n5026), .B1(n6483), .B2(n5025), .ZN(n5017)
         );
  OAI21_X1 U6201 ( .B1(n6467), .B2(n6489), .A(n5017), .ZN(n5018) );
  AOI21_X1 U6202 ( .B1(n5029), .B2(n6485), .A(n5018), .ZN(n5019) );
  OAI21_X1 U6203 ( .B1(n5032), .B2(n5020), .A(n5019), .ZN(U3039) );
  INV_X1 U6204 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5024) );
  AOI22_X1 U6205 ( .A1(n6463), .A2(n5026), .B1(n6459), .B2(n5025), .ZN(n5021)
         );
  OAI21_X1 U6206 ( .B1(n6467), .B2(n6091), .A(n5021), .ZN(n5022) );
  AOI21_X1 U6207 ( .B1(n5029), .B2(n6088), .A(n5022), .ZN(n5023) );
  OAI21_X1 U6208 ( .B1(n5032), .B2(n5024), .A(n5023), .ZN(U3042) );
  INV_X1 U6209 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U6210 ( .A1(n6468), .A2(n5026), .B1(n6469), .B2(n5025), .ZN(n5027)
         );
  OAI21_X1 U6211 ( .B1(n6467), .B2(n6495), .A(n5027), .ZN(n5028) );
  AOI21_X1 U6212 ( .B1(n6502), .B2(n5029), .A(n5028), .ZN(n5030) );
  OAI21_X1 U6213 ( .B1(n5032), .B2(n5031), .A(n5030), .ZN(U3036) );
  INV_X1 U6214 ( .A(n5045), .ZN(n5034) );
  AOI21_X1 U6215 ( .B1(n5034), .B2(n6666), .A(n5150), .ZN(n5042) );
  INV_X1 U6216 ( .A(n5042), .ZN(n5040) );
  INV_X1 U6217 ( .A(n6056), .ZN(n6066) );
  NAND2_X1 U6218 ( .A1(n5035), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6058) );
  NOR2_X1 U6219 ( .A1(n6058), .A2(n5152), .ZN(n5074) );
  AOI21_X1 U6220 ( .B1(n5036), .B2(n6066), .A(n5074), .ZN(n5041) );
  INV_X1 U6221 ( .A(n6058), .ZN(n5037) );
  NOR2_X1 U6222 ( .A1(n5037), .A2(n6666), .ZN(n5039) );
  INV_X1 U6223 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n5049) );
  OAI22_X1 U6224 ( .A1(n5042), .A2(n5041), .B1(n6575), .B2(n6058), .ZN(n5077)
         );
  AOI22_X1 U6225 ( .A1(n5095), .A2(n6507), .B1(n6472), .B2(n5074), .ZN(n5046)
         );
  OAI21_X1 U6226 ( .B1(n6550), .B2(n6099), .A(n5046), .ZN(n5047) );
  AOI21_X1 U6227 ( .B1(n5077), .B2(n6547), .A(n5047), .ZN(n5048) );
  OAI21_X1 U6228 ( .B1(n5080), .B2(n5049), .A(n5048), .ZN(U3093) );
  INV_X1 U6229 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n5053) );
  AOI22_X1 U6230 ( .A1(n5095), .A2(n5117), .B1(n6469), .B2(n5074), .ZN(n5050)
         );
  OAI21_X1 U6231 ( .B1(n5119), .B2(n6099), .A(n5050), .ZN(n5051) );
  AOI21_X1 U6232 ( .B1(n5077), .B2(n6468), .A(n5051), .ZN(n5052) );
  OAI21_X1 U6233 ( .B1(n5080), .B2(n5053), .A(n5052), .ZN(U3092) );
  INV_X1 U6234 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n5057) );
  AOI22_X1 U6235 ( .A1(n5095), .A2(n6514), .B1(n6483), .B2(n5074), .ZN(n5054)
         );
  OAI21_X1 U6236 ( .B1(n6512), .B2(n6099), .A(n5054), .ZN(n5055) );
  AOI21_X1 U6237 ( .B1(n5077), .B2(n6480), .A(n5055), .ZN(n5056) );
  OAI21_X1 U6238 ( .B1(n5080), .B2(n5057), .A(n5056), .ZN(U3095) );
  INV_X1 U6239 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n5061) );
  AOI22_X1 U6240 ( .A1(n5095), .A2(n6451), .B1(n6450), .B2(n5074), .ZN(n5058)
         );
  OAI21_X1 U6241 ( .B1(n6455), .B2(n6099), .A(n5058), .ZN(n5059) );
  AOI21_X1 U6242 ( .B1(n5077), .B2(n6452), .A(n5059), .ZN(n5060) );
  OAI21_X1 U6243 ( .B1(n5080), .B2(n5061), .A(n5060), .ZN(U3096) );
  INV_X1 U6244 ( .A(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n5065) );
  AOI22_X1 U6245 ( .A1(n5095), .A2(n6540), .B1(n5112), .B2(n5074), .ZN(n5062)
         );
  OAI21_X1 U6246 ( .B1(n6573), .B2(n6099), .A(n5062), .ZN(n5063) );
  AOI21_X1 U6247 ( .B1(n5077), .B2(n6568), .A(n5063), .ZN(n5064) );
  OAI21_X1 U6248 ( .B1(n5080), .B2(n5065), .A(n5064), .ZN(U3099) );
  INV_X1 U6249 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n5069) );
  AOI22_X1 U6250 ( .A1(n5095), .A2(n6534), .B1(n6459), .B2(n5074), .ZN(n5066)
         );
  OAI21_X1 U6251 ( .B1(n6532), .B2(n6099), .A(n5066), .ZN(n5067) );
  AOI21_X1 U6252 ( .B1(n5077), .B2(n6463), .A(n5067), .ZN(n5068) );
  OAI21_X1 U6253 ( .B1(n5080), .B2(n5069), .A(n5068), .ZN(U3098) );
  INV_X1 U6254 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n5073) );
  AOI22_X1 U6255 ( .A1(n5095), .A2(n6447), .B1(n6476), .B2(n5074), .ZN(n5070)
         );
  OAI21_X1 U6256 ( .B1(n6678), .B2(n6099), .A(n5070), .ZN(n5071) );
  AOI21_X1 U6257 ( .B1(n5077), .B2(n6552), .A(n5071), .ZN(n5072) );
  OAI21_X1 U6258 ( .B1(n5080), .B2(n5073), .A(n5072), .ZN(U3094) );
  INV_X1 U6259 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n5079) );
  AOI22_X1 U6260 ( .A1(n5095), .A2(n6527), .B1(n6456), .B2(n5074), .ZN(n5075)
         );
  OAI21_X1 U6261 ( .B1(n6561), .B2(n6099), .A(n5075), .ZN(n5076) );
  AOI21_X1 U6262 ( .B1(n5077), .B2(n6558), .A(n5076), .ZN(n5078) );
  OAI21_X1 U6263 ( .B1(n5080), .B2(n5079), .A(n5078), .ZN(U3097) );
  NAND2_X1 U6264 ( .A1(n6031), .A2(n5081), .ZN(n5082) );
  NAND2_X1 U6265 ( .A1(n6000), .A2(n5082), .ZN(n6166) );
  OAI222_X1 U6266 ( .A1(n5608), .A2(n6166), .B1(n6243), .B2(n6157), .C1(n5609), 
        .C2(n6160), .ZN(U2847) );
  OAI21_X1 U6267 ( .B1(n5095), .B2(n5128), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5083) );
  NAND2_X1 U6268 ( .A1(n5083), .A2(n6666), .ZN(n5094) );
  INV_X1 U6269 ( .A(n5094), .ZN(n5090) );
  NOR2_X1 U6270 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5084), .ZN(n5127)
         );
  INV_X1 U6271 ( .A(n5127), .ZN(n5085) );
  AOI22_X1 U6272 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6811), .B1(
        STATE2_REG_3__SCAN_IN), .B2(n5085), .ZN(n5087) );
  NAND3_X1 U6273 ( .A1(n5088), .A2(n5087), .A3(n5086), .ZN(n5089) );
  INV_X1 U6274 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6275 ( .A1(n5155), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5091) );
  AOI22_X1 U6276 ( .A1(n5128), .A2(n6447), .B1(n5127), .B2(n6476), .ZN(n5096)
         );
  OAI21_X1 U6277 ( .B1(n5130), .B2(n6678), .A(n5096), .ZN(n5097) );
  AOI21_X1 U6278 ( .B1(n5132), .B2(n6552), .A(n5097), .ZN(n5098) );
  OAI21_X1 U6279 ( .B1(n5135), .B2(n5099), .A(n5098), .ZN(U3102) );
  INV_X1 U6280 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5103) );
  AOI22_X1 U6281 ( .A1(n5128), .A2(n6514), .B1(n6483), .B2(n5127), .ZN(n5100)
         );
  OAI21_X1 U6282 ( .B1(n5130), .B2(n6512), .A(n5100), .ZN(n5101) );
  AOI21_X1 U6283 ( .B1(n5132), .B2(n6480), .A(n5101), .ZN(n5102) );
  OAI21_X1 U6284 ( .B1(n5135), .B2(n5103), .A(n5102), .ZN(U3103) );
  INV_X1 U6285 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5107) );
  AOI22_X1 U6286 ( .A1(n5128), .A2(n6527), .B1(n5127), .B2(n6456), .ZN(n5104)
         );
  OAI21_X1 U6287 ( .B1(n5130), .B2(n6561), .A(n5104), .ZN(n5105) );
  AOI21_X1 U6288 ( .B1(n5132), .B2(n6558), .A(n5105), .ZN(n5106) );
  OAI21_X1 U6289 ( .B1(n5135), .B2(n5107), .A(n5106), .ZN(U3105) );
  INV_X1 U6290 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5111) );
  AOI22_X1 U6291 ( .A1(n5128), .A2(n6534), .B1(n5127), .B2(n6459), .ZN(n5108)
         );
  OAI21_X1 U6292 ( .B1(n5130), .B2(n6532), .A(n5108), .ZN(n5109) );
  AOI21_X1 U6293 ( .B1(n5132), .B2(n6463), .A(n5109), .ZN(n5110) );
  OAI21_X1 U6294 ( .B1(n5135), .B2(n5111), .A(n5110), .ZN(U3106) );
  INV_X1 U6295 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5116) );
  AOI22_X1 U6296 ( .A1(n5128), .A2(n6540), .B1(n5112), .B2(n5127), .ZN(n5113)
         );
  OAI21_X1 U6297 ( .B1(n5130), .B2(n6573), .A(n5113), .ZN(n5114) );
  AOI21_X1 U6298 ( .B1(n5132), .B2(n6568), .A(n5114), .ZN(n5115) );
  OAI21_X1 U6299 ( .B1(n5135), .B2(n5116), .A(n5115), .ZN(U3107) );
  INV_X1 U6300 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5122) );
  AOI22_X1 U6301 ( .A1(n5128), .A2(n5117), .B1(n6469), .B2(n5127), .ZN(n5118)
         );
  OAI21_X1 U6302 ( .B1(n5119), .B2(n5130), .A(n5118), .ZN(n5120) );
  AOI21_X1 U6303 ( .B1(n5132), .B2(n6468), .A(n5120), .ZN(n5121) );
  OAI21_X1 U6304 ( .B1(n5135), .B2(n5122), .A(n5121), .ZN(U3100) );
  INV_X1 U6305 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5126) );
  AOI22_X1 U6306 ( .A1(n5128), .A2(n6507), .B1(n5127), .B2(n6472), .ZN(n5123)
         );
  OAI21_X1 U6307 ( .B1(n5130), .B2(n6550), .A(n5123), .ZN(n5124) );
  AOI21_X1 U6308 ( .B1(n5132), .B2(n6547), .A(n5124), .ZN(n5125) );
  OAI21_X1 U6309 ( .B1(n5135), .B2(n5126), .A(n5125), .ZN(U3101) );
  INV_X1 U6310 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5134) );
  AOI22_X1 U6311 ( .A1(n5128), .A2(n6451), .B1(n5127), .B2(n6450), .ZN(n5129)
         );
  OAI21_X1 U6312 ( .B1(n5130), .B2(n6455), .A(n5129), .ZN(n5131) );
  AOI21_X1 U6313 ( .B1(n5132), .B2(n6452), .A(n5131), .ZN(n5133) );
  OAI21_X1 U6314 ( .B1(n5135), .B2(n5134), .A(n5133), .ZN(U3104) );
  OAI21_X1 U6315 ( .B1(n5138), .B2(n5137), .A(n5136), .ZN(n6381) );
  INV_X1 U6316 ( .A(n5517), .ZN(n5140) );
  NAND2_X1 U6317 ( .A1(n3009), .A2(REIP_REG_7__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U6318 ( .A1(n6336), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5139)
         );
  OAI211_X1 U6319 ( .C1(n6345), .C2(n5140), .A(n6378), .B(n5139), .ZN(n5141)
         );
  AOI21_X1 U6320 ( .B1(n5142), .B2(n6332), .A(n5141), .ZN(n5143) );
  OAI21_X1 U6321 ( .B1(n6381), .B2(n6316), .A(n5143), .ZN(U2979) );
  INV_X1 U6322 ( .A(n5144), .ZN(n5146) );
  NOR2_X1 U6323 ( .A1(n5145), .A2(n5146), .ZN(n6176) );
  AOI21_X1 U6324 ( .B1(n5146), .B2(n5145), .A(n6176), .ZN(n5827) );
  INV_X1 U6325 ( .A(n5827), .ZN(n5501) );
  AOI22_X1 U6326 ( .A1(n6246), .A2(DATAI_10_), .B1(n5656), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5147) );
  OAI21_X1 U6327 ( .B1(n5501), .B2(n5658), .A(n5147), .ZN(U2881) );
  INV_X1 U6328 ( .A(n5189), .ZN(n5148) );
  NOR3_X1 U6329 ( .A1(n5148), .A2(n6461), .A3(n6497), .ZN(n5151) );
  OAI21_X1 U6330 ( .B1(n5151), .B2(n5150), .A(n5149), .ZN(n5157) );
  NAND2_X1 U6331 ( .A1(n5153), .A2(n5152), .ZN(n5184) );
  AOI211_X1 U6332 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5184), .A(n5155), .B(
        n5154), .ZN(n5156) );
  NAND2_X1 U6333 ( .A1(n5183), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5164) );
  NOR3_X1 U6334 ( .A1(n5158), .A2(n5552), .A3(n6497), .ZN(n5159) );
  AOI21_X1 U6335 ( .B1(n5161), .B2(n5160), .A(n5159), .ZN(n5185) );
  OAI22_X1 U6336 ( .A1(n5185), .A2(n6510), .B1(n6544), .B2(n5184), .ZN(n5162)
         );
  AOI21_X1 U6337 ( .B1(n6461), .B2(n6473), .A(n5162), .ZN(n5163) );
  OAI211_X1 U6338 ( .C1(n5189), .C2(n6545), .A(n5164), .B(n5163), .ZN(U3053)
         );
  NAND2_X1 U6339 ( .A1(n5183), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5167) );
  OAI22_X1 U6340 ( .A1(n5185), .A2(n6505), .B1(n6494), .B2(n5184), .ZN(n5165)
         );
  AOI21_X1 U6341 ( .B1(n6461), .B2(n6502), .A(n5165), .ZN(n5166) );
  OAI211_X1 U6342 ( .C1(n5189), .C2(n6495), .A(n5167), .B(n5166), .ZN(U3052)
         );
  NAND2_X1 U6343 ( .A1(n5183), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5170) );
  OAI22_X1 U6344 ( .A1(n5185), .A2(n6517), .B1(n6511), .B2(n5184), .ZN(n5168)
         );
  AOI21_X1 U6345 ( .B1(n6461), .B2(n6485), .A(n5168), .ZN(n5169) );
  OAI211_X1 U6346 ( .C1(n5189), .C2(n6489), .A(n5170), .B(n5169), .ZN(U3055)
         );
  NAND2_X1 U6347 ( .A1(n5183), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5173) );
  OAI22_X1 U6348 ( .A1(n5185), .A2(n6530), .B1(n6555), .B2(n5184), .ZN(n5171)
         );
  AOI21_X1 U6349 ( .B1(n6461), .B2(n6084), .A(n5171), .ZN(n5172) );
  OAI211_X1 U6350 ( .C1(n5189), .C2(n6556), .A(n5173), .B(n5172), .ZN(U3057)
         );
  NAND2_X1 U6351 ( .A1(n5183), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5176) );
  OAI22_X1 U6352 ( .A1(n5185), .A2(n6537), .B1(n6531), .B2(n5184), .ZN(n5174)
         );
  AOI21_X1 U6353 ( .B1(n6461), .B2(n6088), .A(n5174), .ZN(n5175) );
  OAI211_X1 U6354 ( .C1(n5189), .C2(n6091), .A(n5176), .B(n5175), .ZN(U3058)
         );
  NAND2_X1 U6355 ( .A1(n5183), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5179) );
  OAI22_X1 U6356 ( .A1(n5185), .A2(n6525), .B1(n6518), .B2(n5184), .ZN(n5177)
         );
  AOI21_X1 U6357 ( .B1(n6461), .B2(n6522), .A(n5177), .ZN(n5178) );
  OAI211_X1 U6358 ( .C1(n5189), .C2(n6519), .A(n5179), .B(n5178), .ZN(U3056)
         );
  NAND2_X1 U6359 ( .A1(n5183), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5182) );
  OAI22_X1 U6360 ( .A1(n5185), .A2(n6682), .B1(n6676), .B2(n5184), .ZN(n5180)
         );
  AOI21_X1 U6361 ( .B1(n6461), .B2(n6477), .A(n5180), .ZN(n5181) );
  OAI211_X1 U6362 ( .C1(n5189), .C2(n6681), .A(n5182), .B(n5181), .ZN(U3054)
         );
  NAND2_X1 U6363 ( .A1(n5183), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5188) );
  OAI22_X1 U6364 ( .A1(n5185), .A2(n6543), .B1(n6563), .B2(n5184), .ZN(n5186)
         );
  AOI21_X1 U6365 ( .B1(n6461), .B2(n6096), .A(n5186), .ZN(n5187) );
  OAI211_X1 U6366 ( .C1(n5189), .C2(n6564), .A(n5188), .B(n5187), .ZN(U3059)
         );
  INV_X1 U6367 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5193) );
  INV_X1 U6368 ( .A(n6029), .ZN(n5190) );
  OAI21_X1 U6369 ( .B1(n5192), .B2(n5191), .A(n5190), .ZN(n6352) );
  OAI222_X1 U6370 ( .A1(n5501), .A2(n5609), .B1(n6243), .B2(n5193), .C1(n6352), 
        .C2(n5608), .ZN(U2849) );
  OAI21_X1 U6371 ( .B1(n5196), .B2(n5195), .A(n5194), .ZN(n6373) );
  NAND2_X1 U6372 ( .A1(n3009), .A2(REIP_REG_8__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U6373 ( .A1(n6336), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5197)
         );
  OAI211_X1 U6374 ( .C1(n6345), .C2(n5507), .A(n6370), .B(n5197), .ZN(n5198)
         );
  AOI21_X1 U6375 ( .B1(n5199), .B2(n6332), .A(n5198), .ZN(n5200) );
  OAI21_X1 U6376 ( .B1(n6373), .B2(n6316), .A(n5200), .ZN(U2978) );
  INV_X1 U6377 ( .A(n5201), .ZN(n5205) );
  AOI21_X1 U6378 ( .B1(n5202), .B2(n5407), .A(n5203), .ZN(n5204) );
  NOR2_X1 U6379 ( .A1(n5205), .A2(n5204), .ZN(n5395) );
  AOI21_X1 U6380 ( .B1(n6336), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5206), 
        .ZN(n5207) );
  OAI21_X1 U6381 ( .B1(n5399), .B2(n6345), .A(n5207), .ZN(n5208) );
  AOI21_X1 U6382 ( .B1(n5395), .B2(n6332), .A(n5208), .ZN(n5209) );
  OAI21_X1 U6383 ( .B1(n5210), .B2(n6316), .A(n5209), .ZN(U2964) );
  NAND2_X1 U6384 ( .A1(n5684), .A2(n5211), .ZN(n5667) );
  INV_X1 U6385 ( .A(n5213), .ZN(n5847) );
  INV_X1 U6386 ( .A(n5709), .ZN(n5214) );
  NAND2_X1 U6387 ( .A1(n6395), .A2(n5214), .ZN(n5215) );
  INV_X1 U6388 ( .A(n6428), .ZN(n5218) );
  AOI21_X1 U6389 ( .B1(n5218), .B2(n6432), .A(n5217), .ZN(n5219) );
  OAI21_X1 U6390 ( .B1(n5962), .B2(n5220), .A(n5890), .ZN(n5869) );
  AOI21_X1 U6391 ( .B1(n6395), .B2(n5847), .A(n5869), .ZN(n5846) );
  OAI21_X1 U6392 ( .B1(n5962), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5846), 
        .ZN(n5837) );
  INV_X1 U6393 ( .A(n5221), .ZN(n5872) );
  NAND2_X1 U6394 ( .A1(n5872), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5222) );
  NOR2_X1 U6395 ( .A1(n5902), .A2(n5222), .ZN(n5878) );
  NAND2_X1 U6396 ( .A1(n5878), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U6397 ( .A1(n3009), .A2(REIP_REG_30__SCAN_IN), .ZN(n5660) );
  OAI21_X1 U6398 ( .B1(n5840), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5660), 
        .ZN(n5224) );
  INV_X1 U6399 ( .A(n5224), .ZN(n5225) );
  NAND2_X1 U6400 ( .A1(n4402), .A2(n5234), .ZN(n5228) );
  OAI22_X1 U6401 ( .A1(n6048), .A2(n5228), .B1(n5227), .B2(n5226), .ZN(n5229)
         );
  AOI21_X1 U6402 ( .B1(n5231), .B2(n5230), .A(n5229), .ZN(n5237) );
  INV_X1 U6403 ( .A(n6048), .ZN(n5233) );
  AOI21_X1 U6404 ( .B1(n5233), .B2(n5232), .A(n5236), .ZN(n5235) );
  OAI22_X1 U6405 ( .A1(n5237), .A2(n5236), .B1(n5235), .B2(n5234), .ZN(U3459)
         );
  NAND2_X1 U6406 ( .A1(n5250), .A2(n5238), .ZN(n5241) );
  AOI22_X1 U6407 ( .A1(n5650), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5656), .ZN(n5240) );
  NAND2_X1 U6408 ( .A1(n5241), .A2(n5240), .ZN(U2860) );
  OR2_X1 U6409 ( .A1(n5441), .A2(READREQUEST_REG_SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6410 ( .A1(n5242), .A2(n4212), .ZN(n5245) );
  MUX2_X1 U6411 ( .A(n5246), .B(n5245), .S(n6668), .Z(U3474) );
  INV_X1 U6412 ( .A(n5247), .ZN(n5249) );
  NOR2_X1 U6413 ( .A1(n5248), .A2(n6587), .ZN(n6106) );
  MUX2_X1 U6414 ( .A(MORE_REG_SCAN_IN), .B(n5249), .S(n6106), .Z(U3471) );
  INV_X1 U6415 ( .A(n5250), .ZN(n5294) );
  NAND2_X1 U6416 ( .A1(n6670), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6580) );
  OR2_X1 U6417 ( .A1(n6580), .A2(n6579), .ZN(n6577) );
  NAND2_X1 U6418 ( .A1(n5252), .A2(n5251), .ZN(n6589) );
  NAND3_X1 U6419 ( .A1(n6435), .A2(n6577), .A3(n6589), .ZN(n5253) );
  INV_X1 U6420 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5587) );
  MUX2_X1 U6421 ( .A(EBX_REG_29__SCAN_IN), .B(n3137), .S(n5418), .Z(n5256) );
  AOI21_X1 U6422 ( .B1(n5257), .B2(n5587), .A(n5256), .ZN(n5312) );
  NAND2_X1 U6423 ( .A1(n5312), .A2(n5258), .ZN(n5259) );
  OAI22_X1 U6424 ( .A1(n5262), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5267), .ZN(n5263) );
  INV_X1 U6425 ( .A(n5263), .ZN(n5264) );
  NAND2_X1 U6426 ( .A1(n5296), .A2(EBX_REG_31__SCAN_IN), .ZN(n5266) );
  NOR2_X1 U6427 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  AND3_X1 U6428 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6429 ( .A1(n5270), .A2(n5269), .ZN(n5271) );
  AOI21_X1 U6430 ( .B1(n5267), .B2(n5271), .A(n5296), .ZN(n5272) );
  NAND2_X2 U6431 ( .A1(n5545), .A2(n5272), .ZN(n6150) );
  NAND2_X1 U6432 ( .A1(n6150), .A2(n6151), .ZN(n5582) );
  INV_X1 U6433 ( .A(n5582), .ZN(n5553) );
  INV_X1 U6434 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6626) );
  INV_X1 U6435 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6828) );
  INV_X1 U6436 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6623) );
  INV_X1 U6437 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6618) );
  INV_X1 U6438 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6612) );
  INV_X1 U6439 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6610) );
  INV_X1 U6440 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6606) );
  INV_X1 U6441 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6603) );
  NOR3_X1 U6442 ( .A1(n6656), .A2(n4655), .A3(n6603), .ZN(n6206) );
  NAND2_X1 U6443 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6206), .ZN(n5538) );
  NOR2_X1 U6444 ( .A1(n6606), .A2(n5538), .ZN(n6196) );
  NAND2_X1 U6445 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6196), .ZN(n5500) );
  NOR3_X1 U6446 ( .A1(n6612), .A2(n6610), .A3(n5500), .ZN(n5510) );
  NAND3_X1 U6447 ( .A1(n5510), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n6167) );
  NOR2_X1 U6448 ( .A1(n6618), .A2(n6167), .ZN(n6149) );
  NAND3_X1 U6449 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        n6149), .ZN(n6130) );
  NOR2_X1 U6450 ( .A1(n6623), .A2(n6130), .ZN(n5280) );
  NAND2_X1 U6451 ( .A1(n5280), .A2(n6151), .ZN(n5493) );
  NOR3_X1 U6452 ( .A1(n6626), .A2(n6828), .A3(n5493), .ZN(n5273) );
  NAND2_X1 U6453 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5273), .ZN(n5274) );
  NAND2_X1 U6454 ( .A1(n5582), .A2(n5274), .ZN(n5470) );
  INV_X1 U6455 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6629) );
  NAND2_X1 U6456 ( .A1(n6207), .A2(n6629), .ZN(n5275) );
  NAND2_X1 U6457 ( .A1(n5470), .A2(n5275), .ZN(n5457) );
  NAND2_X1 U6458 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_20__SCAN_IN), .ZN(
        n5283) );
  AND2_X1 U6459 ( .A1(n5582), .A2(n5283), .ZN(n5276) );
  OR2_X2 U6460 ( .A1(n5457), .A2(n5276), .ZN(n5423) );
  AND3_X1 U6461 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5284) );
  NOR2_X1 U6462 ( .A1(n6150), .A2(n5284), .ZN(n5277) );
  NOR2_X1 U6463 ( .A1(n5423), .A2(n5277), .ZN(n5387) );
  OAI21_X1 U6464 ( .B1(n5285), .B2(n5553), .A(n5387), .ZN(n5353) );
  INV_X1 U6465 ( .A(n5353), .ZN(n5343) );
  AND2_X1 U6466 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5286) );
  NOR2_X1 U6467 ( .A1(n5353), .A2(n6207), .ZN(n5305) );
  AOI21_X1 U6468 ( .B1(n5343), .B2(n5286), .A(n5305), .ZN(n5328) );
  INV_X1 U6469 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6646) );
  NOR2_X1 U6470 ( .A1(n5328), .A2(n6646), .ZN(n5306) );
  AOI211_X1 U6471 ( .C1(n5306), .C2(REIP_REG_30__SCAN_IN), .A(n5305), .B(n6650), .ZN(n5292) );
  AND2_X1 U6472 ( .A1(n5279), .A2(n5278), .ZN(n5295) );
  NAND3_X1 U6473 ( .A1(n5545), .A2(EBX_REG_31__SCAN_IN), .A3(n5295), .ZN(n5289) );
  INV_X1 U6474 ( .A(n5280), .ZN(n5281) );
  NOR2_X1 U6475 ( .A1(n6828), .A2(n5492), .ZN(n5488) );
  NAND2_X1 U6476 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5488), .ZN(n5471) );
  INV_X1 U6477 ( .A(n5471), .ZN(n5282) );
  NAND2_X1 U6478 ( .A1(n5456), .A2(REIP_REG_18__SCAN_IN), .ZN(n5424) );
  NOR2_X1 U6479 ( .A1(n5424), .A2(n5283), .ZN(n5408) );
  AND2_X1 U6480 ( .A1(n5408), .A2(n5284), .ZN(n5352) );
  NAND2_X1 U6481 ( .A1(n5352), .A2(n5285), .ZN(n5339) );
  INV_X1 U6482 ( .A(n5286), .ZN(n5287) );
  NOR2_X1 U6483 ( .A1(n5339), .A2(n5287), .ZN(n5316) );
  NAND4_X1 U6484 ( .A1(n5316), .A2(REIP_REG_29__SCAN_IN), .A3(
        REIP_REG_30__SCAN_IN), .A4(n6650), .ZN(n5288) );
  OAI211_X1 U6485 ( .C1(n5290), .C2(n6143), .A(n5289), .B(n5288), .ZN(n5291)
         );
  AOI211_X1 U6486 ( .C1(n5843), .C2(n6211), .A(n5292), .B(n5291), .ZN(n5293)
         );
  OAI21_X1 U6487 ( .B1(n5294), .B2(n6199), .A(n5293), .ZN(U2796) );
  NAND2_X1 U6488 ( .A1(n5663), .A2(n6190), .ZN(n5310) );
  INV_X1 U6489 ( .A(n5295), .ZN(n5298) );
  INV_X1 U6490 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5585) );
  NAND3_X1 U6491 ( .A1(n5270), .A2(n5585), .A3(n5296), .ZN(n5297) );
  NAND2_X1 U6492 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  NOR2_X1 U6493 ( .A1(n6646), .A2(REIP_REG_30__SCAN_IN), .ZN(n5302) );
  AOI22_X1 U6494 ( .A1(n6214), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .B1(n5316), 
        .B2(n5302), .ZN(n5303) );
  OAI21_X1 U6495 ( .B1(n5661), .B2(n6217), .A(n5303), .ZN(n5308) );
  INV_X1 U6496 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5304) );
  NOR3_X1 U6497 ( .A1(n5306), .A2(n5305), .A3(n5304), .ZN(n5307) );
  AOI211_X1 U6498 ( .C1(EBX_REG_30__SCAN_IN), .C2(n6222), .A(n5308), .B(n5307), 
        .ZN(n5309) );
  OAI211_X1 U6499 ( .C1(n6184), .C2(n5311), .A(n5310), .B(n5309), .ZN(U2797)
         );
  XNOR2_X1 U6500 ( .A(n5322), .B(n5312), .ZN(n5851) );
  NAND2_X1 U6501 ( .A1(n5672), .A2(n6190), .ZN(n5320) );
  OAI22_X1 U6502 ( .A1(n6217), .A2(n5670), .B1(n6827), .B2(n6143), .ZN(n5318)
         );
  MUX2_X1 U6503 ( .A(n5316), .B(n5328), .S(REIP_REG_29__SCAN_IN), .Z(n5317) );
  AOI211_X1 U6504 ( .C1(EBX_REG_29__SCAN_IN), .C2(n6222), .A(n5318), .B(n5317), 
        .ZN(n5319) );
  OAI211_X1 U6505 ( .C1(n6184), .C2(n5851), .A(n5320), .B(n5319), .ZN(U2798)
         );
  AND2_X1 U6506 ( .A1(n5338), .A2(n5321), .ZN(n5323) );
  INV_X1 U6507 ( .A(n5682), .ZN(n5326) );
  NAND2_X1 U6508 ( .A1(n5326), .A2(n6190), .ZN(n5333) );
  OAI22_X1 U6509 ( .A1(n6217), .A2(n5674), .B1(n5327), .B2(n6143), .ZN(n5331)
         );
  INV_X1 U6510 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6808) );
  NOR2_X1 U6511 ( .A1(n5339), .A2(n6808), .ZN(n5329) );
  MUX2_X1 U6512 ( .A(n5329), .B(n5328), .S(REIP_REG_28__SCAN_IN), .Z(n5330) );
  AOI211_X1 U6513 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6222), .A(n5331), .B(n5330), 
        .ZN(n5332) );
  OAI211_X1 U6514 ( .C1(n6184), .C2(n5857), .A(n5333), .B(n5332), .ZN(U2799)
         );
  AOI21_X1 U6515 ( .B1(n5335), .B2(n5347), .A(n5324), .ZN(n5690) );
  INV_X1 U6516 ( .A(n5690), .ZN(n5623) );
  NAND2_X1 U6517 ( .A1(n5351), .A2(n5336), .ZN(n5337) );
  AND2_X1 U6518 ( .A1(n5338), .A2(n5337), .ZN(n5864) );
  OAI22_X1 U6519 ( .A1(n6143), .A2(n5688), .B1(REIP_REG_27__SCAN_IN), .B2(
        n5339), .ZN(n5340) );
  AOI21_X1 U6520 ( .B1(n5686), .B2(n6189), .A(n5340), .ZN(n5342) );
  NAND2_X1 U6521 ( .A1(n6222), .A2(EBX_REG_27__SCAN_IN), .ZN(n5341) );
  OAI211_X1 U6522 ( .C1(n5343), .C2(n6808), .A(n5342), .B(n5341), .ZN(n5344)
         );
  AOI21_X1 U6523 ( .B1(n5864), .B2(n6211), .A(n5344), .ZN(n5345) );
  OAI21_X1 U6524 ( .B1(n5623), .B2(n6199), .A(n5345), .ZN(U2800) );
  OR2_X1 U6525 ( .A1(n5364), .A2(n5349), .ZN(n5350) );
  NAND2_X1 U6526 ( .A1(n5351), .A2(n5350), .ZN(n5874) );
  INV_X1 U6527 ( .A(n5874), .ZN(n5358) );
  INV_X1 U6528 ( .A(n5352), .ZN(n5377) );
  INV_X1 U6529 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6784) );
  INV_X1 U6530 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6638) );
  NOR3_X1 U6531 ( .A1(n5377), .A2(n6784), .A3(n6638), .ZN(n5354) );
  OAI21_X1 U6532 ( .B1(REIP_REG_26__SCAN_IN), .B2(n5354), .A(n5353), .ZN(n5356) );
  AOI22_X1 U6533 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6214), .B1(n6189), 
        .B2(n5699), .ZN(n5355) );
  OAI211_X1 U6534 ( .C1(n6714), .C2(n6171), .A(n5356), .B(n5355), .ZN(n5357)
         );
  AOI21_X1 U6535 ( .B1(n5358), .B2(n6211), .A(n5357), .ZN(n5359) );
  OAI21_X1 U6536 ( .B1(n5697), .B2(n6199), .A(n5359), .ZN(U2801) );
  AOI21_X1 U6537 ( .B1(n5362), .B2(n5360), .A(n5361), .ZN(n5363) );
  INV_X1 U6538 ( .A(n5363), .ZN(n5708) );
  AOI21_X1 U6539 ( .B1(n3099), .B2(n5365), .A(n5364), .ZN(n5886) );
  XNOR2_X1 U6540 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .ZN(
        n5366) );
  OAI22_X1 U6541 ( .A1(n6143), .A2(n5700), .B1(n5377), .B2(n5366), .ZN(n5367)
         );
  AOI21_X1 U6542 ( .B1(n5702), .B2(n6189), .A(n5367), .ZN(n5369) );
  NAND2_X1 U6543 ( .A1(n6222), .A2(EBX_REG_25__SCAN_IN), .ZN(n5368) );
  OAI211_X1 U6544 ( .C1(n5387), .C2(n6638), .A(n5369), .B(n5368), .ZN(n5370)
         );
  AOI21_X1 U6545 ( .B1(n5886), .B2(n6211), .A(n5370), .ZN(n5371) );
  OAI21_X1 U6546 ( .B1(n5708), .B2(n6199), .A(n5371), .ZN(U2802) );
  OAI21_X1 U6547 ( .B1(n5372), .B2(n5373), .A(n5360), .ZN(n5714) );
  AND2_X1 U6548 ( .A1(n5386), .A2(n5374), .ZN(n5375) );
  NOR2_X1 U6549 ( .A1(n5376), .A2(n5375), .ZN(n5895) );
  OAI22_X1 U6550 ( .A1(n6143), .A2(n5713), .B1(REIP_REG_24__SCAN_IN), .B2(
        n5377), .ZN(n5378) );
  AOI21_X1 U6551 ( .B1(n5717), .B2(n6189), .A(n5378), .ZN(n5380) );
  NAND2_X1 U6552 ( .A1(n6222), .A2(EBX_REG_24__SCAN_IN), .ZN(n5379) );
  OAI211_X1 U6553 ( .C1(n5387), .C2(n6784), .A(n5380), .B(n5379), .ZN(n5381)
         );
  AOI21_X1 U6554 ( .B1(n5895), .B2(n6211), .A(n5381), .ZN(n5382) );
  OAI21_X1 U6555 ( .B1(n5714), .B2(n6199), .A(n5382), .ZN(U2803) );
  AOI21_X1 U6556 ( .B1(n5383), .B2(n5201), .A(n5372), .ZN(n5726) );
  INV_X1 U6557 ( .A(n5726), .ZN(n5632) );
  NAND2_X1 U6558 ( .A1(n4263), .A2(n5384), .ZN(n5385) );
  NAND2_X1 U6559 ( .A1(n5386), .A2(n5385), .ZN(n5899) );
  INV_X1 U6560 ( .A(n5899), .ZN(n5393) );
  INV_X1 U6561 ( .A(REIP_REG_23__SCAN_IN), .ZN(n5389) );
  NAND3_X1 U6562 ( .A1(n5408), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5388) );
  AOI21_X1 U6563 ( .B1(n5389), .B2(n5388), .A(n5387), .ZN(n5392) );
  INV_X1 U6564 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6719) );
  AOI22_X1 U6565 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n6214), .B1(n6189), 
        .B2(n5722), .ZN(n5390) );
  OAI21_X1 U6566 ( .B1(n6171), .B2(n6719), .A(n5390), .ZN(n5391) );
  AOI211_X1 U6567 ( .C1(n5393), .C2(n6211), .A(n5392), .B(n5391), .ZN(n5394)
         );
  OAI21_X1 U6568 ( .B1(n5632), .B2(n6199), .A(n5394), .ZN(U2804) );
  INV_X1 U6569 ( .A(n5395), .ZN(n5635) );
  NAND2_X1 U6570 ( .A1(n6222), .A2(EBX_REG_22__SCAN_IN), .ZN(n5398) );
  XOR2_X1 U6571 ( .A(REIP_REG_22__SCAN_IN), .B(REIP_REG_21__SCAN_IN), .Z(n5396) );
  AOI22_X1 U6572 ( .A1(n6214), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .B1(n5408), 
        .B2(n5396), .ZN(n5397) );
  OAI211_X1 U6573 ( .C1(n6217), .C2(n5399), .A(n5398), .B(n5397), .ZN(n5400)
         );
  AOI21_X1 U6574 ( .B1(n5423), .B2(REIP_REG_22__SCAN_IN), .A(n5400), .ZN(n5402) );
  NAND2_X1 U6575 ( .A1(n5593), .A2(n6211), .ZN(n5401) );
  OAI211_X1 U6576 ( .C1(n5635), .C2(n6199), .A(n5402), .B(n5401), .ZN(U2805)
         );
  NOR2_X1 U6577 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  OR2_X1 U6578 ( .A1(n5406), .A2(n5405), .ZN(n5910) );
  XOR2_X1 U6579 ( .A(n5407), .B(n5202), .Z(n5734) );
  NAND2_X1 U6580 ( .A1(n5734), .A2(n6190), .ZN(n5415) );
  NAND2_X1 U6581 ( .A1(n6222), .A2(EBX_REG_21__SCAN_IN), .ZN(n5412) );
  INV_X1 U6582 ( .A(n5408), .ZN(n5409) );
  OAI22_X1 U6583 ( .A1(n6143), .A2(n6745), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5409), .ZN(n5410) );
  INV_X1 U6584 ( .A(n5410), .ZN(n5411) );
  OAI211_X1 U6585 ( .C1(n6217), .C2(n5732), .A(n5412), .B(n5411), .ZN(n5413)
         );
  AOI21_X1 U6586 ( .B1(n5423), .B2(REIP_REG_21__SCAN_IN), .A(n5413), .ZN(n5414) );
  OAI211_X1 U6587 ( .C1(n5910), .C2(n6184), .A(n5415), .B(n5414), .ZN(U2806)
         );
  INV_X1 U6588 ( .A(n5416), .ZN(n5433) );
  MUX2_X1 U6589 ( .A(n5433), .B(n5418), .S(n5417), .Z(n5420) );
  XNOR2_X1 U6590 ( .A(n5420), .B(n5419), .ZN(n5925) );
  NOR2_X1 U6591 ( .A1(n5437), .A2(n5421), .ZN(n5422) );
  OR2_X1 U6592 ( .A1(n5202), .A2(n5422), .ZN(n5641) );
  INV_X1 U6593 ( .A(n5641), .ZN(n5743) );
  NAND2_X1 U6594 ( .A1(n5743), .A2(n6190), .ZN(n5430) );
  OAI22_X1 U6595 ( .A1(n6217), .A2(n5739), .B1(n5740), .B2(n6143), .ZN(n5428)
         );
  INV_X1 U6596 ( .A(n5423), .ZN(n5426) );
  INV_X1 U6597 ( .A(n5424), .ZN(n5440) );
  AOI21_X1 U6598 ( .B1(n5440), .B2(REIP_REG_19__SCAN_IN), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5425) );
  NOR2_X1 U6599 ( .A1(n5426), .A2(n5425), .ZN(n5427) );
  AOI211_X1 U6600 ( .C1(n6222), .C2(EBX_REG_20__SCAN_IN), .A(n5428), .B(n5427), 
        .ZN(n5429) );
  OAI211_X1 U6601 ( .C1(n5925), .C2(n6184), .A(n5430), .B(n5429), .ZN(U2807)
         );
  MUX2_X1 U6602 ( .A(n5433), .B(n5432), .S(n4110), .Z(n5448) );
  OR2_X1 U6603 ( .A1(n5431), .A2(n5448), .ZN(n5449) );
  XNOR2_X1 U6604 ( .A(n5449), .B(n5434), .ZN(n5933) );
  INV_X1 U6605 ( .A(n5436), .ZN(n5453) );
  INV_X1 U6606 ( .A(n5753), .ZN(n5438) );
  NAND2_X1 U6607 ( .A1(n5438), .A2(n6190), .ZN(n5447) );
  AOI22_X1 U6608 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n6214), .B1(n6189), 
        .B2(n5750), .ZN(n5444) );
  NAND2_X1 U6609 ( .A1(n6222), .A2(EBX_REG_19__SCAN_IN), .ZN(n5443) );
  INV_X1 U6610 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6611 ( .A1(n5440), .A2(n5439), .ZN(n5442) );
  NAND2_X1 U6612 ( .A1(n6151), .A2(n5441), .ZN(n6197) );
  NAND4_X1 U6613 ( .A1(n5444), .A2(n5443), .A3(n5442), .A4(n6197), .ZN(n5445)
         );
  AOI21_X1 U6614 ( .B1(n5457), .B2(REIP_REG_19__SCAN_IN), .A(n5445), .ZN(n5446) );
  OAI211_X1 U6615 ( .C1(n5933), .C2(n6184), .A(n5447), .B(n5446), .ZN(U2808)
         );
  INV_X1 U6616 ( .A(n5431), .ZN(n5451) );
  INV_X1 U6617 ( .A(n5448), .ZN(n5450) );
  OAI21_X1 U6618 ( .B1(n5451), .B2(n5450), .A(n5449), .ZN(n5944) );
  AOI21_X1 U6619 ( .B1(n5454), .B2(n5467), .A(n5453), .ZN(n5764) );
  NAND2_X1 U6620 ( .A1(n5764), .A2(n6190), .ZN(n5463) );
  NAND2_X1 U6621 ( .A1(n6189), .A2(n5760), .ZN(n5455) );
  OAI211_X1 U6622 ( .C1(n6143), .C2(n5762), .A(n5455), .B(n6197), .ZN(n5461)
         );
  INV_X1 U6623 ( .A(n5456), .ZN(n5459) );
  INV_X1 U6624 ( .A(n5457), .ZN(n5458) );
  AOI21_X1 U6625 ( .B1(n6629), .B2(n5459), .A(n5458), .ZN(n5460) );
  AOI211_X1 U6626 ( .C1(EBX_REG_18__SCAN_IN), .C2(n6222), .A(n5461), .B(n5460), 
        .ZN(n5462) );
  OAI211_X1 U6627 ( .C1(n6184), .C2(n5944), .A(n5463), .B(n5462), .ZN(U2809)
         );
  OR2_X1 U6628 ( .A1(n5484), .A2(n5464), .ZN(n5465) );
  NAND2_X1 U6629 ( .A1(n5431), .A2(n5465), .ZN(n5951) );
  OAI21_X1 U6630 ( .B1(n5466), .B2(n5468), .A(n5467), .ZN(n5778) );
  INV_X1 U6631 ( .A(n5778), .ZN(n5469) );
  NAND2_X1 U6632 ( .A1(n5469), .A2(n6190), .ZN(n5480) );
  INV_X1 U6633 ( .A(n5470), .ZN(n5478) );
  INV_X1 U6634 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U6635 ( .A1(n5773), .A2(n5471), .ZN(n5477) );
  NAND2_X1 U6636 ( .A1(n6222), .A2(EBX_REG_17__SCAN_IN), .ZN(n5475) );
  OAI21_X1 U6637 ( .B1(n6143), .B2(n5472), .A(n6197), .ZN(n5473) );
  INV_X1 U6638 ( .A(n5473), .ZN(n5474) );
  OAI211_X1 U6639 ( .C1(n6217), .C2(n5774), .A(n5475), .B(n5474), .ZN(n5476)
         );
  AOI21_X1 U6640 ( .B1(n5478), .B2(n5477), .A(n5476), .ZN(n5479) );
  OAI211_X1 U6641 ( .C1(n5951), .C2(n6184), .A(n5480), .B(n5479), .ZN(U2810)
         );
  NOR2_X1 U6642 ( .A1(n5481), .A2(n5482), .ZN(n5483) );
  OR2_X1 U6643 ( .A1(n5484), .A2(n5483), .ZN(n5964) );
  OR2_X1 U6644 ( .A1(n5485), .A2(n5654), .ZN(n5486) );
  AOI21_X1 U6645 ( .B1(n5487), .B2(n5486), .A(n5466), .ZN(n5787) );
  NAND2_X1 U6646 ( .A1(n5787), .A2(n6190), .ZN(n5497) );
  INV_X1 U6647 ( .A(n5488), .ZN(n5491) );
  INV_X1 U6648 ( .A(n5785), .ZN(n5489) );
  AOI22_X1 U6649 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n6214), .B1(n6189), 
        .B2(n5489), .ZN(n5490) );
  OAI211_X1 U6650 ( .C1(REIP_REG_16__SCAN_IN), .C2(n5491), .A(n5490), .B(n6197), .ZN(n5495) );
  OR2_X1 U6651 ( .A1(n5492), .A2(REIP_REG_15__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U6652 ( .A1(n5582), .A2(n5493), .ZN(n6132) );
  AOI21_X1 U6653 ( .B1(n6122), .B2(n6132), .A(n6626), .ZN(n5494) );
  AOI211_X1 U6654 ( .C1(EBX_REG_16__SCAN_IN), .C2(n6222), .A(n5495), .B(n5494), 
        .ZN(n5496) );
  OAI211_X1 U6655 ( .C1(n5964), .C2(n6184), .A(n5497), .B(n5496), .ZN(U2811)
         );
  INV_X1 U6656 ( .A(n6197), .ZN(n6212) );
  AOI21_X1 U6657 ( .B1(n6214), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6212), 
        .ZN(n5499) );
  OAI21_X1 U6658 ( .B1(n6150), .B2(n5510), .A(n6151), .ZN(n6186) );
  AOI22_X1 U6659 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6222), .B1(
        REIP_REG_10__SCAN_IN), .B2(n6186), .ZN(n5498) );
  OAI211_X1 U6660 ( .C1(n6184), .C2(n6352), .A(n5499), .B(n5498), .ZN(n5504)
         );
  INV_X1 U6661 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6616) );
  INV_X1 U6662 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6614) );
  OR2_X1 U6663 ( .A1(n6150), .A2(n5500), .ZN(n5523) );
  NOR2_X1 U6664 ( .A1(n5523), .A2(n6610), .ZN(n5512) );
  NAND2_X1 U6665 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5512), .ZN(n6194) );
  AOI221_X1 U6666 ( .B1(REIP_REG_10__SCAN_IN), .B2(REIP_REG_9__SCAN_IN), .C1(
        n6616), .C2(n6614), .A(n6194), .ZN(n5503) );
  OAI22_X1 U6667 ( .A1(n5501), .A2(n6199), .B1(n5825), .B2(n6217), .ZN(n5502)
         );
  OR3_X1 U6668 ( .A1(n5504), .A2(n5503), .A3(n5502), .ZN(U2817) );
  AOI22_X1 U6669 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6214), .B1(n6211), 
        .B2(n6372), .ZN(n5505) );
  OAI211_X1 U6670 ( .C1(n6171), .C2(n5506), .A(n5505), .B(n6197), .ZN(n5509)
         );
  NOR2_X1 U6671 ( .A1(n6217), .A2(n5507), .ZN(n5508) );
  AOI211_X1 U6672 ( .C1(REIP_REG_8__SCAN_IN), .C2(n6186), .A(n5509), .B(n5508), 
        .ZN(n5514) );
  INV_X1 U6673 ( .A(n5510), .ZN(n5511) );
  NAND2_X1 U6674 ( .A1(n5512), .A2(n5511), .ZN(n5513) );
  OAI211_X1 U6675 ( .C1(n5515), .C2(n6199), .A(n5514), .B(n5513), .ZN(U2819)
         );
  INV_X1 U6676 ( .A(n5516), .ZN(n6380) );
  AOI22_X1 U6677 ( .A1(n6211), .A2(n6380), .B1(n6222), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5522) );
  NAND2_X1 U6678 ( .A1(n6189), .A2(n5517), .ZN(n5518) );
  OAI211_X1 U6679 ( .C1(n5519), .C2(n6143), .A(n5518), .B(n6197), .ZN(n5520)
         );
  INV_X1 U6680 ( .A(n5520), .ZN(n5521) );
  OAI211_X1 U6681 ( .C1(REIP_REG_7__SCAN_IN), .C2(n5523), .A(n5522), .B(n5521), 
        .ZN(n5524) );
  INV_X1 U6682 ( .A(n5524), .ZN(n5527) );
  NOR2_X1 U6683 ( .A1(n6150), .A2(REIP_REG_6__SCAN_IN), .ZN(n6195) );
  OR2_X1 U6684 ( .A1(n6150), .A2(n6196), .ZN(n5525) );
  NAND2_X1 U6685 ( .A1(n5525), .A2(n6151), .ZN(n6203) );
  OAI21_X1 U6686 ( .B1(n6195), .B2(n6203), .A(REIP_REG_7__SCAN_IN), .ZN(n5526)
         );
  OAI211_X1 U6687 ( .C1(n5528), .C2(n6199), .A(n5527), .B(n5526), .ZN(U2820)
         );
  INV_X1 U6688 ( .A(n5529), .ZN(n5532) );
  NAND2_X1 U6689 ( .A1(n5545), .A2(n5530), .ZN(n5531) );
  NAND2_X1 U6690 ( .A1(n5531), .A2(n6199), .ZN(n5558) );
  NAND2_X1 U6691 ( .A1(n5532), .A2(n5558), .ZN(n5543) );
  NAND2_X1 U6692 ( .A1(n6189), .A2(n5533), .ZN(n5534) );
  OAI211_X1 U6693 ( .C1(n5535), .C2(n6143), .A(n5534), .B(n6197), .ZN(n5536)
         );
  INV_X1 U6694 ( .A(n5536), .ZN(n5542) );
  INV_X1 U6695 ( .A(n5537), .ZN(n6403) );
  AOI22_X1 U6696 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6222), .B1(n6211), .B2(n6403), 
        .ZN(n5541) );
  OAI21_X1 U6697 ( .B1(n6150), .B2(n5538), .A(n6606), .ZN(n5539) );
  NAND2_X1 U6698 ( .A1(n6203), .A2(n5539), .ZN(n5540) );
  NAND4_X1 U6699 ( .A1(n5543), .A2(n5542), .A3(n5541), .A4(n5540), .ZN(U2822)
         );
  AND2_X1 U6700 ( .A1(n5545), .A2(n5544), .ZN(n6210) );
  OAI22_X1 U6701 ( .A1(n6217), .A2(n5547), .B1(n5546), .B2(n6143), .ZN(n5551)
         );
  INV_X1 U6702 ( .A(n6421), .ZN(n5549) );
  INV_X1 U6703 ( .A(EBX_REG_3__SCAN_IN), .ZN(n5548) );
  OAI22_X1 U6704 ( .A1(n6184), .A2(n5549), .B1(n6171), .B2(n5548), .ZN(n5550)
         );
  AOI211_X1 U6705 ( .C1(n6210), .C2(n5552), .A(n5551), .B(n5550), .ZN(n5556)
         );
  AOI21_X1 U6706 ( .B1(n6151), .B2(REIP_REG_1__SCAN_IN), .A(n5553), .ZN(n5554)
         );
  NOR2_X1 U6707 ( .A1(n5554), .A2(n6603), .ZN(n5567) );
  OAI21_X1 U6708 ( .B1(n6150), .B2(n6206), .A(n6151), .ZN(n6213) );
  OAI21_X1 U6709 ( .B1(n5567), .B2(REIP_REG_3__SCAN_IN), .A(n6213), .ZN(n5555)
         );
  OAI211_X1 U6710 ( .C1(n5557), .C2(n6218), .A(n5556), .B(n5555), .ZN(U2824)
         );
  AOI21_X1 U6711 ( .B1(n6207), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U6712 ( .A1(n6341), .A2(n5558), .ZN(n5565) );
  INV_X1 U6713 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5559) );
  OAI22_X1 U6714 ( .A1(n6217), .A2(n6344), .B1(n5559), .B2(n6143), .ZN(n5562)
         );
  XNOR2_X1 U6715 ( .A(n4455), .B(n5560), .ZN(n6238) );
  INV_X1 U6716 ( .A(n6238), .ZN(n6433) );
  OAI22_X1 U6717 ( .A1(n6242), .A2(n6171), .B1(n6184), .B2(n6433), .ZN(n5561)
         );
  AOI211_X1 U6718 ( .C1(n5563), .C2(n6210), .A(n5562), .B(n5561), .ZN(n5564)
         );
  OAI211_X1 U6719 ( .C1(n5567), .C2(n5566), .A(n5565), .B(n5564), .ZN(U2825)
         );
  AOI22_X1 U6720 ( .A1(EBX_REG_1__SCAN_IN), .A2(n6222), .B1(n6211), .B2(n4377), 
        .ZN(n5574) );
  AOI22_X1 U6721 ( .A1(n6207), .A2(n6656), .B1(n6210), .B2(n5568), .ZN(n5573)
         );
  OAI22_X1 U6722 ( .A1(n6143), .A2(n5569), .B1(n6151), .B2(n6656), .ZN(n5570)
         );
  INV_X1 U6723 ( .A(n5570), .ZN(n5572) );
  NAND2_X1 U6724 ( .A1(n6189), .A2(n5569), .ZN(n5571) );
  AND4_X1 U6725 ( .A1(n5574), .A2(n5573), .A3(n5572), .A4(n5571), .ZN(n5575)
         );
  OAI21_X1 U6726 ( .B1(n6218), .B2(n5576), .A(n5575), .ZN(U2826) );
  INV_X1 U6727 ( .A(n6210), .ZN(n5580) );
  AOI22_X1 U6728 ( .A1(EBX_REG_0__SCAN_IN), .A2(n6222), .B1(n6211), .B2(n5577), 
        .ZN(n5579) );
  OAI21_X1 U6729 ( .B1(n6214), .B2(n6189), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5578) );
  OAI211_X1 U6730 ( .C1(n5580), .C2(n6490), .A(n5579), .B(n5578), .ZN(n5581)
         );
  AOI21_X1 U6731 ( .B1(n5582), .B2(REIP_REG_0__SCAN_IN), .A(n5581), .ZN(n5583)
         );
  OAI21_X1 U6732 ( .B1(n6218), .B2(n5584), .A(n5583), .ZN(U2827) );
  INV_X1 U6733 ( .A(n5843), .ZN(n5586) );
  OAI22_X1 U6734 ( .A1(n5586), .A2(n5608), .B1(n6243), .B2(n5585), .ZN(U2828)
         );
  INV_X1 U6735 ( .A(n5672), .ZN(n5618) );
  OAI222_X1 U6736 ( .A1(n5609), .A2(n5618), .B1(n5587), .B2(n6243), .C1(n5851), 
        .C2(n5608), .ZN(U2830) );
  OAI222_X1 U6737 ( .A1(n5609), .A2(n5682), .B1(n5588), .B2(n6243), .C1(n5857), 
        .C2(n5608), .ZN(U2831) );
  AOI22_X1 U6738 ( .A1(n5864), .A2(n6239), .B1(EBX_REG_27__SCAN_IN), .B2(n5592), .ZN(n5589) );
  OAI21_X1 U6739 ( .B1(n5623), .B2(n5609), .A(n5589), .ZN(U2832) );
  OAI222_X1 U6740 ( .A1(n5609), .A2(n5697), .B1(n6714), .B2(n6243), .C1(n5874), 
        .C2(n5608), .ZN(U2833) );
  AOI22_X1 U6741 ( .A1(n5886), .A2(n6239), .B1(EBX_REG_25__SCAN_IN), .B2(n5592), .ZN(n5590) );
  OAI21_X1 U6742 ( .B1(n5708), .B2(n5609), .A(n5590), .ZN(U2834) );
  AOI22_X1 U6743 ( .A1(n5895), .A2(n6239), .B1(EBX_REG_24__SCAN_IN), .B2(n5592), .ZN(n5591) );
  OAI21_X1 U6744 ( .B1(n5714), .B2(n5609), .A(n5591), .ZN(U2835) );
  OAI222_X1 U6745 ( .A1(n5609), .A2(n5632), .B1(n6719), .B2(n6243), .C1(n5899), 
        .C2(n5608), .ZN(U2836) );
  AOI22_X1 U6746 ( .A1(n5593), .A2(n6239), .B1(EBX_REG_22__SCAN_IN), .B2(n5592), .ZN(n5594) );
  OAI21_X1 U6747 ( .B1(n5635), .B2(n5609), .A(n5594), .ZN(U2837) );
  INV_X1 U6748 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5595) );
  INV_X1 U6749 ( .A(n5734), .ZN(n5638) );
  OAI222_X1 U6750 ( .A1(n5910), .A2(n5608), .B1(n5595), .B2(n6243), .C1(n5609), 
        .C2(n5638), .ZN(U2838) );
  INV_X1 U6751 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5596) );
  OAI222_X1 U6752 ( .A1(n5641), .A2(n5609), .B1(n5596), .B2(n6243), .C1(n5608), 
        .C2(n5925), .ZN(U2839) );
  OAI222_X1 U6753 ( .A1(n5753), .A2(n5609), .B1(n5597), .B2(n6243), .C1(n5608), 
        .C2(n5933), .ZN(U2840) );
  INV_X1 U6754 ( .A(n5764), .ZN(n5646) );
  OAI222_X1 U6755 ( .A1(n5609), .A2(n5646), .B1(n5598), .B2(n6243), .C1(n5944), 
        .C2(n5608), .ZN(U2841) );
  OAI22_X1 U6756 ( .A1(n5951), .A2(n5608), .B1(n5599), .B2(n6243), .ZN(n5600)
         );
  INV_X1 U6757 ( .A(n5600), .ZN(n5601) );
  OAI21_X1 U6758 ( .B1(n5778), .B2(n5609), .A(n5601), .ZN(U2842) );
  INV_X1 U6759 ( .A(n5787), .ZN(n5653) );
  INV_X1 U6760 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5602) );
  OAI222_X1 U6761 ( .A1(n5653), .A2(n5609), .B1(n5602), .B2(n6243), .C1(n5964), 
        .C2(n5608), .ZN(U2843) );
  OR2_X1 U6762 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  NAND2_X1 U6763 ( .A1(n5485), .A2(n5605), .ZN(n6137) );
  AND2_X1 U6764 ( .A1(n6002), .A2(n5606), .ZN(n5607) );
  OR2_X1 U6765 ( .A1(n5607), .A2(n5973), .ZN(n6141) );
  OAI222_X1 U6766 ( .A1(n6137), .A2(n5609), .B1(n6243), .B2(n4172), .C1(n6141), 
        .C2(n5608), .ZN(U2845) );
  NOR3_X1 U6767 ( .A1(n5656), .A2(n5611), .A3(n5610), .ZN(n5612) );
  AOI22_X1 U6768 ( .A1(n5649), .A2(DATAI_14_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5656), .ZN(n5614) );
  NAND2_X1 U6769 ( .A1(n5650), .A2(DATAI_30_), .ZN(n5613) );
  OAI211_X1 U6770 ( .C1(n5615), .C2(n5658), .A(n5614), .B(n5613), .ZN(U2861)
         );
  AOI22_X1 U6771 ( .A1(n5649), .A2(DATAI_13_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n5656), .ZN(n5617) );
  NAND2_X1 U6772 ( .A1(n5650), .A2(DATAI_29_), .ZN(n5616) );
  OAI211_X1 U6773 ( .C1(n5618), .C2(n5658), .A(n5617), .B(n5616), .ZN(U2862)
         );
  AOI22_X1 U6774 ( .A1(n5649), .A2(DATAI_12_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5656), .ZN(n5620) );
  NAND2_X1 U6775 ( .A1(n5650), .A2(DATAI_28_), .ZN(n5619) );
  OAI211_X1 U6776 ( .C1(n5682), .C2(n5658), .A(n5620), .B(n5619), .ZN(U2863)
         );
  AOI22_X1 U6777 ( .A1(n5649), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5656), .ZN(n5622) );
  NAND2_X1 U6778 ( .A1(n5650), .A2(DATAI_27_), .ZN(n5621) );
  OAI211_X1 U6779 ( .C1(n5623), .C2(n5658), .A(n5622), .B(n5621), .ZN(U2864)
         );
  AOI22_X1 U6780 ( .A1(n5649), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5656), .ZN(n5625) );
  NAND2_X1 U6781 ( .A1(n5650), .A2(DATAI_26_), .ZN(n5624) );
  OAI211_X1 U6782 ( .C1(n5697), .C2(n5658), .A(n5625), .B(n5624), .ZN(U2865)
         );
  AOI22_X1 U6783 ( .A1(n5649), .A2(DATAI_9_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n5656), .ZN(n5627) );
  NAND2_X1 U6784 ( .A1(n5650), .A2(DATAI_25_), .ZN(n5626) );
  OAI211_X1 U6785 ( .C1(n5708), .C2(n5658), .A(n5627), .B(n5626), .ZN(U2866)
         );
  AOI22_X1 U6786 ( .A1(n5649), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n5656), .ZN(n5629) );
  NAND2_X1 U6787 ( .A1(n5650), .A2(DATAI_24_), .ZN(n5628) );
  OAI211_X1 U6788 ( .C1(n5714), .C2(n5658), .A(n5629), .B(n5628), .ZN(U2867)
         );
  AOI22_X1 U6789 ( .A1(n5649), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n5656), .ZN(n5631) );
  NAND2_X1 U6790 ( .A1(n5650), .A2(DATAI_23_), .ZN(n5630) );
  OAI211_X1 U6791 ( .C1(n5632), .C2(n5658), .A(n5631), .B(n5630), .ZN(U2868)
         );
  AOI22_X1 U6792 ( .A1(n5649), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n5656), .ZN(n5634) );
  NAND2_X1 U6793 ( .A1(n5650), .A2(DATAI_22_), .ZN(n5633) );
  OAI211_X1 U6794 ( .C1(n5635), .C2(n5658), .A(n5634), .B(n5633), .ZN(U2869)
         );
  AOI22_X1 U6795 ( .A1(n5649), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n5656), .ZN(n5637) );
  NAND2_X1 U6796 ( .A1(n5650), .A2(DATAI_21_), .ZN(n5636) );
  OAI211_X1 U6797 ( .C1(n5638), .C2(n5658), .A(n5637), .B(n5636), .ZN(U2870)
         );
  AOI22_X1 U6798 ( .A1(n5649), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n5656), .ZN(n5640) );
  NAND2_X1 U6799 ( .A1(n5650), .A2(DATAI_20_), .ZN(n5639) );
  OAI211_X1 U6800 ( .C1(n5641), .C2(n5658), .A(n5640), .B(n5639), .ZN(U2871)
         );
  AOI22_X1 U6801 ( .A1(n5649), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n5656), .ZN(n5643) );
  NAND2_X1 U6802 ( .A1(n5650), .A2(DATAI_19_), .ZN(n5642) );
  OAI211_X1 U6803 ( .C1(n5753), .C2(n5658), .A(n5643), .B(n5642), .ZN(U2872)
         );
  AOI22_X1 U6804 ( .A1(n5649), .A2(DATAI_2_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n5656), .ZN(n5645) );
  NAND2_X1 U6805 ( .A1(n5650), .A2(DATAI_18_), .ZN(n5644) );
  OAI211_X1 U6806 ( .C1(n5646), .C2(n5658), .A(n5645), .B(n5644), .ZN(U2873)
         );
  AOI22_X1 U6807 ( .A1(n5649), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n5656), .ZN(n5648) );
  NAND2_X1 U6808 ( .A1(n5650), .A2(DATAI_17_), .ZN(n5647) );
  OAI211_X1 U6809 ( .C1(n5778), .C2(n5658), .A(n5648), .B(n5647), .ZN(U2874)
         );
  AOI22_X1 U6810 ( .A1(n5649), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n5656), .ZN(n5652) );
  NAND2_X1 U6811 ( .A1(n5650), .A2(DATAI_16_), .ZN(n5651) );
  OAI211_X1 U6812 ( .C1(n5653), .C2(n5658), .A(n5652), .B(n5651), .ZN(U2875)
         );
  XNOR2_X1 U6813 ( .A(n5485), .B(n5654), .ZN(n6227) );
  AOI22_X1 U6814 ( .A1(n6246), .A2(DATAI_15_), .B1(n5656), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5655) );
  OAI21_X1 U6815 ( .B1(n6227), .B2(n5658), .A(n5655), .ZN(U2876) );
  AOI22_X1 U6816 ( .A1(n6246), .A2(DATAI_14_), .B1(n5656), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5657) );
  OAI21_X1 U6817 ( .B1(n6137), .B2(n5658), .A(n5657), .ZN(U2877) );
  NAND2_X1 U6818 ( .A1(n6336), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5659)
         );
  OAI211_X1 U6819 ( .C1(n6345), .C2(n5661), .A(n5660), .B(n5659), .ZN(n5662)
         );
  AOI21_X1 U6820 ( .B1(n5663), .B2(n6332), .A(n5662), .ZN(n5664) );
  OAI21_X1 U6821 ( .B1(n5665), .B2(n6316), .A(n5664), .ZN(U2956) );
  NAND2_X1 U6822 ( .A1(n5667), .A2(n5666), .ZN(n5668) );
  XNOR2_X1 U6823 ( .A(n5668), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5855)
         );
  NOR2_X1 U6824 ( .A1(n6435), .A2(n6646), .ZN(n5849) );
  AOI21_X1 U6825 ( .B1(n6336), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5849), 
        .ZN(n5669) );
  OAI21_X1 U6826 ( .B1(n6345), .B2(n5670), .A(n5669), .ZN(n5671) );
  AOI21_X1 U6827 ( .B1(n5672), .B2(n6332), .A(n5671), .ZN(n5673) );
  OAI21_X1 U6828 ( .B1(n5855), .B2(n6316), .A(n5673), .ZN(U2957) );
  INV_X1 U6829 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6642) );
  NOR2_X1 U6830 ( .A1(n6435), .A2(n6642), .ZN(n5859) );
  NOR2_X1 U6831 ( .A1(n6345), .A2(n5674), .ZN(n5675) );
  AOI211_X1 U6832 ( .C1(PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n6336), .A(n5859), 
        .B(n5675), .ZN(n5681) );
  INV_X1 U6833 ( .A(n5693), .ZN(n5676) );
  INV_X1 U6834 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6775) );
  NAND3_X1 U6835 ( .A1(n5705), .A2(n5676), .A3(n6775), .ZN(n5683) );
  AOI22_X1 U6836 ( .A1(n5677), .A2(n5683), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5877), .ZN(n5679) );
  XNOR2_X1 U6837 ( .A(n5679), .B(n5678), .ZN(n5856) );
  NAND2_X1 U6838 ( .A1(n5856), .A2(n6340), .ZN(n5680) );
  OAI211_X1 U6839 ( .C1(n5682), .C2(n5779), .A(n5681), .B(n5680), .ZN(U2958)
         );
  NAND2_X1 U6840 ( .A1(n6025), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5692) );
  OAI21_X1 U6841 ( .B1(n5684), .B2(n5692), .A(n5683), .ZN(n5685) );
  XNOR2_X1 U6842 ( .A(n5685), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5871)
         );
  NAND2_X1 U6843 ( .A1(n6312), .A2(n5686), .ZN(n5687) );
  NAND2_X1 U6844 ( .A1(n3009), .A2(REIP_REG_27__SCAN_IN), .ZN(n5865) );
  OAI211_X1 U6845 ( .C1(n5688), .C2(n5833), .A(n5687), .B(n5865), .ZN(n5689)
         );
  AOI21_X1 U6846 ( .B1(n5690), .B2(n6332), .A(n5689), .ZN(n5691) );
  OAI21_X1 U6847 ( .B1(n5871), .B2(n6316), .A(n5691), .ZN(U2959) );
  NAND2_X1 U6848 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  XNOR2_X1 U6849 ( .A(n5695), .B(n5694), .ZN(n5880) );
  NAND2_X1 U6850 ( .A1(n3009), .A2(REIP_REG_26__SCAN_IN), .ZN(n5873) );
  OAI21_X1 U6851 ( .B1(n5833), .B2(n5696), .A(n5873), .ZN(n5698) );
  NAND2_X1 U6852 ( .A1(n3009), .A2(REIP_REG_25__SCAN_IN), .ZN(n5882) );
  OAI21_X1 U6853 ( .B1(n5833), .B2(n5700), .A(n5882), .ZN(n5701) );
  AOI21_X1 U6854 ( .B1(n6312), .B2(n5702), .A(n5701), .ZN(n5707) );
  OAI21_X1 U6855 ( .B1(n5705), .B2(n5704), .A(n5703), .ZN(n5881) );
  NAND2_X1 U6856 ( .A1(n5881), .A2(n6340), .ZN(n5706) );
  OAI211_X1 U6857 ( .C1(n5708), .C2(n5779), .A(n5707), .B(n5706), .ZN(U2961)
         );
  NAND2_X1 U6858 ( .A1(n5728), .A2(n2983), .ZN(n5711) );
  NAND4_X1 U6859 ( .A1(n5730), .A2(n5709), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n5781), .ZN(n5710) );
  NAND2_X1 U6860 ( .A1(n5711), .A2(n5710), .ZN(n5712) );
  XNOR2_X1 U6861 ( .A(n5712), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5897)
         );
  NAND2_X1 U6862 ( .A1(n3009), .A2(REIP_REG_24__SCAN_IN), .ZN(n5889) );
  OAI21_X1 U6863 ( .B1(n5833), .B2(n5713), .A(n5889), .ZN(n5716) );
  NOR2_X1 U6864 ( .A1(n5714), .A2(n5779), .ZN(n5715) );
  AOI211_X1 U6865 ( .C1(n5717), .C2(n6312), .A(n5716), .B(n5715), .ZN(n5718)
         );
  OAI21_X1 U6866 ( .B1(n5897), .B2(n6316), .A(n5718), .ZN(U2962) );
  AOI22_X1 U6867 ( .A1(n5728), .A2(n5719), .B1(n5746), .B2(n5900), .ZN(n5721)
         );
  XNOR2_X1 U6868 ( .A(n5721), .B(n5720), .ZN(n5907) );
  NAND2_X1 U6869 ( .A1(n6312), .A2(n5722), .ZN(n5723) );
  NAND2_X1 U6870 ( .A1(n3009), .A2(REIP_REG_23__SCAN_IN), .ZN(n5898) );
  OAI211_X1 U6871 ( .C1(n5724), .C2(n5833), .A(n5723), .B(n5898), .ZN(n5725)
         );
  AOI21_X1 U6872 ( .B1(n5726), .B2(n6332), .A(n5725), .ZN(n5727) );
  OAI21_X1 U6873 ( .B1(n5907), .B2(n6316), .A(n5727), .ZN(U2963) );
  AOI21_X1 U6874 ( .B1(n5730), .B2(n5729), .A(n5728), .ZN(n5915) );
  INV_X1 U6875 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6633) );
  NOR2_X1 U6876 ( .A1(n6435), .A2(n6633), .ZN(n5908) );
  AOI21_X1 U6877 ( .B1(n6336), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5908), 
        .ZN(n5731) );
  OAI21_X1 U6878 ( .B1(n5732), .B2(n6345), .A(n5731), .ZN(n5733) );
  AOI21_X1 U6879 ( .B1(n5734), .B2(n6332), .A(n5733), .ZN(n5735) );
  OAI21_X1 U6880 ( .B1(n5915), .B2(n6316), .A(n5735), .ZN(U2965) );
  XNOR2_X1 U6881 ( .A(n6025), .B(n5736), .ZN(n5737) );
  XNOR2_X1 U6882 ( .A(n5738), .B(n5737), .ZN(n5928) );
  INV_X1 U6883 ( .A(n5739), .ZN(n5742) );
  NAND2_X1 U6884 ( .A1(n3009), .A2(REIP_REG_20__SCAN_IN), .ZN(n5923) );
  OAI21_X1 U6885 ( .B1(n5833), .B2(n5740), .A(n5923), .ZN(n5741) );
  AOI21_X1 U6886 ( .B1(n6312), .B2(n5742), .A(n5741), .ZN(n5745) );
  NAND2_X1 U6887 ( .A1(n5743), .A2(n6332), .ZN(n5744) );
  OAI211_X1 U6888 ( .C1(n5928), .C2(n6316), .A(n5745), .B(n5744), .ZN(U2966)
         );
  INV_X1 U6889 ( .A(n5746), .ZN(n5931) );
  NAND2_X1 U6890 ( .A1(n2971), .A2(n5747), .ZN(n5930) );
  NAND3_X1 U6891 ( .A1(n5931), .A2(n6340), .A3(n5930), .ZN(n5752) );
  NAND2_X1 U6892 ( .A1(n3009), .A2(REIP_REG_19__SCAN_IN), .ZN(n5932) );
  OAI21_X1 U6893 ( .B1(n5833), .B2(n5748), .A(n5932), .ZN(n5749) );
  AOI21_X1 U6894 ( .B1(n6312), .B2(n5750), .A(n5749), .ZN(n5751) );
  OAI211_X1 U6895 ( .C1(n5779), .C2(n5753), .A(n5752), .B(n5751), .ZN(U2967)
         );
  AOI21_X1 U6896 ( .B1(n5756), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n5755), 
        .ZN(n5791) );
  XNOR2_X1 U6897 ( .A(n6025), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5790)
         );
  INV_X1 U6898 ( .A(n5789), .ZN(n5758) );
  NOR2_X1 U6899 ( .A1(n5781), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5780)
         );
  NAND3_X1 U6900 ( .A1(n5758), .A2(n5780), .A3(n5957), .ZN(n5770) );
  NAND2_X1 U6901 ( .A1(n5766), .A2(n5770), .ZN(n5759) );
  XNOR2_X1 U6902 ( .A(n5759), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5948)
         );
  NAND2_X1 U6903 ( .A1(n6312), .A2(n5760), .ZN(n5761) );
  NAND2_X1 U6904 ( .A1(n3009), .A2(REIP_REG_18__SCAN_IN), .ZN(n5942) );
  OAI211_X1 U6905 ( .C1(n5833), .C2(n5762), .A(n5761), .B(n5942), .ZN(n5763)
         );
  AOI21_X1 U6906 ( .B1(n5764), .B2(n6332), .A(n5763), .ZN(n5765) );
  OAI21_X1 U6907 ( .B1(n5948), .B2(n6316), .A(n5765), .ZN(U2968) );
  NAND2_X1 U6908 ( .A1(n5756), .A2(n5957), .ZN(n5768) );
  INV_X1 U6909 ( .A(n5780), .ZN(n5767) );
  AOI22_X1 U6910 ( .A1(n5769), .A2(n5768), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5767), .ZN(n5771) );
  OAI21_X1 U6911 ( .B1(n5772), .B2(n5771), .A(n5770), .ZN(n5950) );
  NAND2_X1 U6912 ( .A1(n5950), .A2(n6340), .ZN(n5777) );
  NOR2_X1 U6913 ( .A1(n6435), .A2(n5773), .ZN(n5952) );
  NOR2_X1 U6914 ( .A1(n6345), .A2(n5774), .ZN(n5775) );
  AOI211_X1 U6915 ( .C1(n6336), .C2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n5952), 
        .B(n5775), .ZN(n5776) );
  AOI21_X1 U6916 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n5781), .A(n5780), 
        .ZN(n5782) );
  XNOR2_X1 U6917 ( .A(n5783), .B(n5782), .ZN(n5970) );
  NAND2_X1 U6918 ( .A1(n3009), .A2(REIP_REG_16__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U6919 ( .A1(n6336), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5784)
         );
  OAI211_X1 U6920 ( .C1(n6345), .C2(n5785), .A(n5963), .B(n5784), .ZN(n5786)
         );
  AOI21_X1 U6921 ( .B1(n5787), .B2(n6332), .A(n5786), .ZN(n5788) );
  OAI21_X1 U6922 ( .B1(n5970), .B2(n6316), .A(n5788), .ZN(U2970) );
  OAI21_X1 U6923 ( .B1(n5791), .B2(n5790), .A(n5789), .ZN(n5971) );
  NAND2_X1 U6924 ( .A1(n5971), .A2(n6340), .ZN(n5794) );
  NAND2_X1 U6925 ( .A1(n3009), .A2(REIP_REG_15__SCAN_IN), .ZN(n5975) );
  OAI21_X1 U6926 ( .B1(n5833), .B2(n6757), .A(n5975), .ZN(n5792) );
  AOI21_X1 U6927 ( .B1(n6312), .B2(n6127), .A(n5792), .ZN(n5793) );
  OAI211_X1 U6928 ( .C1(n6227), .C2(n5779), .A(n5794), .B(n5793), .ZN(U2971)
         );
  XNOR2_X1 U6929 ( .A(n6025), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5796)
         );
  XNOR2_X1 U6930 ( .A(n5795), .B(n5796), .ZN(n5998) );
  NAND2_X1 U6931 ( .A1(n5998), .A2(n6340), .ZN(n5799) );
  NOR2_X1 U6932 ( .A1(n6435), .A2(n6623), .ZN(n5991) );
  NOR2_X1 U6933 ( .A1(n6345), .A2(n6136), .ZN(n5797) );
  AOI211_X1 U6934 ( .C1(n6336), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5991), 
        .B(n5797), .ZN(n5798) );
  OAI211_X1 U6935 ( .C1(n5779), .C2(n6137), .A(n5799), .B(n5798), .ZN(U2972)
         );
  XOR2_X1 U6936 ( .A(n5800), .B(n5801), .Z(n6012) );
  INV_X1 U6937 ( .A(n5802), .ZN(n5803) );
  AOI21_X1 U6938 ( .B1(n5805), .B2(n5804), .A(n5803), .ZN(n6244) );
  NAND2_X1 U6939 ( .A1(n3009), .A2(REIP_REG_13__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U6940 ( .A1(n6336), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5806)
         );
  OAI211_X1 U6941 ( .C1(n6345), .C2(n6155), .A(n6007), .B(n5806), .ZN(n5807)
         );
  AOI21_X1 U6942 ( .B1(n6244), .B2(n6332), .A(n5807), .ZN(n5808) );
  OAI21_X1 U6943 ( .B1(n6012), .B2(n6316), .A(n5808), .ZN(U2973) );
  OAI21_X1 U6944 ( .B1(n5781), .B2(n5810), .A(n5809), .ZN(n5817) );
  INV_X1 U6945 ( .A(n5811), .ZN(n5815) );
  NAND2_X1 U6946 ( .A1(n5815), .A2(n5812), .ZN(n6024) );
  OAI21_X1 U6947 ( .B1(n6024), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5756), 
        .ZN(n5813) );
  OAI21_X1 U6948 ( .B1(n5815), .B2(n5814), .A(n5813), .ZN(n5816) );
  XOR2_X1 U6949 ( .A(n5817), .B(n5816), .Z(n6023) );
  INV_X1 U6950 ( .A(n6162), .ZN(n5819) );
  NAND2_X1 U6951 ( .A1(n3009), .A2(REIP_REG_12__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U6952 ( .A1(n6336), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5818)
         );
  OAI211_X1 U6953 ( .C1(n6345), .C2(n5819), .A(n6013), .B(n5818), .ZN(n5820)
         );
  AOI21_X1 U6954 ( .B1(n5821), .B2(n6332), .A(n5820), .ZN(n5822) );
  OAI21_X1 U6955 ( .B1(n6023), .B2(n6316), .A(n5822), .ZN(U2974) );
  XNOR2_X1 U6956 ( .A(n6025), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5823)
         );
  XNOR2_X1 U6957 ( .A(n5811), .B(n5823), .ZN(n6350) );
  AOI22_X1 U6958 ( .A1(n6336), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n3009), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5824) );
  OAI21_X1 U6959 ( .B1(n5825), .B2(n6345), .A(n5824), .ZN(n5826) );
  AOI21_X1 U6960 ( .B1(n5827), .B2(n6332), .A(n5826), .ZN(n5828) );
  OAI21_X1 U6961 ( .B1(n6350), .B2(n6316), .A(n5828), .ZN(U2976) );
  NAND2_X1 U6962 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  XNOR2_X1 U6963 ( .A(n5829), .B(n5832), .ZN(n6364) );
  NAND2_X1 U6964 ( .A1(n6364), .A2(n6340), .ZN(n5836) );
  NAND2_X1 U6965 ( .A1(n3009), .A2(REIP_REG_9__SCAN_IN), .ZN(n6360) );
  OAI21_X1 U6966 ( .B1(n5833), .B2(n6181), .A(n6360), .ZN(n5834) );
  AOI21_X1 U6967 ( .B1(n6312), .B2(n6188), .A(n5834), .ZN(n5835) );
  OAI211_X1 U6968 ( .C1(n5779), .C2(n6187), .A(n5836), .B(n5835), .ZN(U2977)
         );
  NOR3_X1 U6969 ( .A1(n5840), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5839), 
        .ZN(n5841) );
  NAND2_X1 U6970 ( .A1(n5843), .A2(n6422), .ZN(n5844) );
  INV_X1 U6971 ( .A(n5846), .ZN(n5850) );
  NOR3_X1 U6972 ( .A1(n5863), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5847), 
        .ZN(n5848) );
  AOI211_X1 U6973 ( .C1(n5850), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5849), .B(n5848), .ZN(n5854) );
  INV_X1 U6974 ( .A(n5851), .ZN(n5852) );
  NAND2_X1 U6975 ( .A1(n5852), .A2(n6422), .ZN(n5853) );
  OAI211_X1 U6976 ( .C1(n5855), .C2(n6351), .A(n5854), .B(n5853), .ZN(U2989)
         );
  XNOR2_X1 U6977 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U6978 ( .A1(n5856), .A2(n6438), .ZN(n5861) );
  NOR2_X1 U6979 ( .A1(n5857), .A2(n6434), .ZN(n5858) );
  AOI211_X1 U6980 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5869), .A(n5859), .B(n5858), .ZN(n5860) );
  OAI211_X1 U6981 ( .C1(n5863), .C2(n5862), .A(n5861), .B(n5860), .ZN(U2990)
         );
  NOR2_X1 U6982 ( .A1(n5863), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5868)
         );
  INV_X1 U6983 ( .A(n5864), .ZN(n5866) );
  OAI21_X1 U6984 ( .B1(n5866), .B2(n6434), .A(n5865), .ZN(n5867) );
  AOI211_X1 U6985 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5869), .A(n5868), .B(n5867), .ZN(n5870) );
  OAI21_X1 U6986 ( .B1(n5871), .B2(n6351), .A(n5870), .ZN(U2991) );
  NAND3_X1 U6987 ( .A1(n5935), .A2(n5872), .A3(n6775), .ZN(n5883) );
  AOI21_X1 U6988 ( .B1(n5883), .B2(n5890), .A(n5877), .ZN(n5876) );
  OAI21_X1 U6989 ( .B1(n5874), .B2(n6434), .A(n5873), .ZN(n5875) );
  AOI211_X1 U6990 ( .C1(n5878), .C2(n5877), .A(n5876), .B(n5875), .ZN(n5879)
         );
  OAI21_X1 U6991 ( .B1(n5880), .B2(n6351), .A(n5879), .ZN(U2992) );
  NAND2_X1 U6992 ( .A1(n5881), .A2(n6438), .ZN(n5888) );
  INV_X1 U6993 ( .A(n5882), .ZN(n5885) );
  INV_X1 U6994 ( .A(n5883), .ZN(n5884) );
  AOI211_X1 U6995 ( .C1(n5886), .C2(n6422), .A(n5885), .B(n5884), .ZN(n5887)
         );
  OAI211_X1 U6996 ( .C1(n5890), .C2(n6775), .A(n5888), .B(n5887), .ZN(U2993)
         );
  INV_X1 U6997 ( .A(n5889), .ZN(n5894) );
  NAND3_X1 U6998 ( .A1(n5935), .A2(n5900), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5891) );
  AOI21_X1 U6999 ( .B1(n5892), .B2(n5891), .A(n5890), .ZN(n5893) );
  AOI211_X1 U7000 ( .C1(n6422), .C2(n5895), .A(n5894), .B(n5893), .ZN(n5896)
         );
  OAI21_X1 U7001 ( .B1(n5897), .B2(n6351), .A(n5896), .ZN(U2994) );
  OAI21_X1 U7002 ( .B1(n5899), .B2(n6434), .A(n5898), .ZN(n5904) );
  INV_X1 U7003 ( .A(n5900), .ZN(n5901) );
  NOR3_X1 U7004 ( .A1(n5902), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5901), 
        .ZN(n5903) );
  AOI211_X1 U7005 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5905), .A(n5904), .B(n5903), .ZN(n5906) );
  OAI21_X1 U7006 ( .B1(n5907), .B2(n6351), .A(n5906), .ZN(U2995) );
  INV_X1 U7007 ( .A(n5908), .ZN(n5909) );
  OAI21_X1 U7008 ( .B1(n5910), .B2(n6434), .A(n5909), .ZN(n5912) );
  AOI211_X1 U7009 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5913), .A(n5912), .B(n5911), .ZN(n5914) );
  OAI21_X1 U7010 ( .B1(n5915), .B2(n6351), .A(n5914), .ZN(U2997) );
  NAND2_X1 U7011 ( .A1(n5941), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5916) );
  OAI21_X1 U7012 ( .B1(n5983), .B2(n5916), .A(n6346), .ZN(n5918) );
  NAND2_X1 U7013 ( .A1(n5918), .A2(n5917), .ZN(n5949) );
  NOR2_X1 U7014 ( .A1(n6014), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5919)
         );
  OR2_X1 U7015 ( .A1(n5949), .A2(n5919), .ZN(n5946) );
  INV_X1 U7016 ( .A(n5946), .ZN(n5920) );
  OAI21_X1 U7017 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5962), .A(n5920), 
        .ZN(n5929) );
  NAND3_X1 U7018 ( .A1(n5935), .A2(n5922), .A3(n5921), .ZN(n5924) );
  OAI211_X1 U7019 ( .C1(n6434), .C2(n5925), .A(n5924), .B(n5923), .ZN(n5926)
         );
  AOI21_X1 U7020 ( .B1(INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n5929), .A(n5926), 
        .ZN(n5927) );
  OAI21_X1 U7021 ( .B1(n5928), .B2(n6351), .A(n5927), .ZN(U2998) );
  INV_X1 U7022 ( .A(n5929), .ZN(n5939) );
  NAND3_X1 U7023 ( .A1(n5931), .A2(n6438), .A3(n5930), .ZN(n5937) );
  OAI21_X1 U7024 ( .B1(n5933), .B2(n6434), .A(n5932), .ZN(n5934) );
  AOI21_X1 U7025 ( .B1(n5935), .B2(n5938), .A(n5934), .ZN(n5936) );
  OAI211_X1 U7026 ( .C1(n5939), .C2(n5938), .A(n5937), .B(n5936), .ZN(U2999)
         );
  NAND4_X1 U7027 ( .A1(n6036), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5941), .A4(n5940), .ZN(n5943) );
  OAI211_X1 U7028 ( .C1(n6434), .C2(n5944), .A(n5943), .B(n5942), .ZN(n5945)
         );
  AOI21_X1 U7029 ( .B1(n5946), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5945), 
        .ZN(n5947) );
  OAI21_X1 U7030 ( .B1(n5948), .B2(n6351), .A(n5947), .ZN(U3000) );
  INV_X1 U7031 ( .A(n5949), .ZN(n5958) );
  NAND2_X1 U7032 ( .A1(n5950), .A2(n6438), .ZN(n5956) );
  NOR2_X1 U7033 ( .A1(n5951), .A2(n6434), .ZN(n5953) );
  AOI211_X1 U7034 ( .C1(n5954), .C2(n5957), .A(n5953), .B(n5952), .ZN(n5955)
         );
  NAND2_X1 U7035 ( .A1(n6387), .A2(n5959), .ZN(n5960) );
  OAI21_X1 U7036 ( .B1(n5965), .B2(n5962), .A(n6033), .ZN(n5979) );
  OAI21_X1 U7037 ( .B1(n5964), .B2(n6434), .A(n5963), .ZN(n5968) );
  NAND2_X1 U7038 ( .A1(n6036), .A2(n5965), .ZN(n5977) );
  XNOR2_X1 U7039 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5966) );
  NOR2_X1 U7040 ( .A1(n5977), .A2(n5966), .ZN(n5967) );
  AOI211_X1 U7041 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n5979), .A(n5968), .B(n5967), .ZN(n5969) );
  OAI21_X1 U7042 ( .B1(n5970), .B2(n6351), .A(n5969), .ZN(U3002) );
  INV_X1 U7043 ( .A(n5971), .ZN(n5981) );
  NOR2_X1 U7044 ( .A1(n5973), .A2(n5972), .ZN(n5974) );
  OR2_X1 U7045 ( .A1(n5481), .A2(n5974), .ZN(n6226) );
  INV_X1 U7046 ( .A(n6226), .ZN(n6126) );
  NAND2_X1 U7047 ( .A1(n6126), .A2(n6422), .ZN(n5976) );
  OAI211_X1 U7048 ( .C1(n5977), .C2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5976), .B(n5975), .ZN(n5978) );
  AOI21_X1 U7049 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5979), .A(n5978), 
        .ZN(n5980) );
  OAI21_X1 U7050 ( .B1(n5981), .B2(n6351), .A(n5980), .ZN(U3003) );
  AOI21_X1 U7051 ( .B1(n6036), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5996) );
  AOI21_X1 U7052 ( .B1(n5983), .B2(n5982), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5985) );
  INV_X1 U7053 ( .A(n6015), .ZN(n6006) );
  OAI21_X1 U7054 ( .B1(n5985), .B2(n5984), .A(n6006), .ZN(n5995) );
  NOR2_X1 U7055 ( .A1(n6015), .A2(n6005), .ZN(n5987) );
  OAI22_X1 U7056 ( .A1(n5988), .A2(n6006), .B1(n5987), .B2(n5986), .ZN(n5989)
         );
  INV_X1 U7057 ( .A(n5989), .ZN(n5990) );
  NAND2_X1 U7058 ( .A1(n6033), .A2(n5990), .ZN(n6010) );
  NAND2_X1 U7059 ( .A1(n6010), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5994) );
  INV_X1 U7060 ( .A(n6141), .ZN(n5992) );
  AOI21_X1 U7061 ( .B1(n5992), .B2(n6422), .A(n5991), .ZN(n5993) );
  OAI211_X1 U7062 ( .C1(n5996), .C2(n5995), .A(n5994), .B(n5993), .ZN(n5997)
         );
  AOI21_X1 U7063 ( .B1(n5998), .B2(n6438), .A(n5997), .ZN(n5999) );
  INV_X1 U7064 ( .A(n5999), .ZN(U3004) );
  INV_X1 U7065 ( .A(n6000), .ZN(n6004) );
  INV_X1 U7066 ( .A(n6001), .ZN(n6003) );
  OAI21_X1 U7067 ( .B1(n6004), .B2(n6003), .A(n6002), .ZN(n6231) );
  NAND3_X1 U7068 ( .A1(n6036), .A2(n6006), .A3(n6005), .ZN(n6008) );
  OAI211_X1 U7069 ( .C1(n6434), .C2(n6231), .A(n6008), .B(n6007), .ZN(n6009)
         );
  AOI21_X1 U7070 ( .B1(n6010), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n6009), 
        .ZN(n6011) );
  OAI21_X1 U7071 ( .B1(n6012), .B2(n6351), .A(n6011), .ZN(U3005) );
  INV_X1 U7072 ( .A(n6166), .ZN(n6021) );
  INV_X1 U7073 ( .A(n6013), .ZN(n6020) );
  INV_X1 U7074 ( .A(n6014), .ZN(n6016) );
  INV_X1 U7075 ( .A(n6432), .ZN(n6390) );
  OAI21_X1 U7076 ( .B1(n6016), .B2(n6390), .A(n6015), .ZN(n6018) );
  AOI21_X1 U7077 ( .B1(n6036), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6017) );
  AOI21_X1 U7078 ( .B1(n6033), .B2(n6018), .A(n6017), .ZN(n6019) );
  AOI211_X1 U7079 ( .C1(n6422), .C2(n6021), .A(n6020), .B(n6019), .ZN(n6022)
         );
  OAI21_X1 U7080 ( .B1(n6023), .B2(n6351), .A(n6022), .ZN(U3006) );
  AOI22_X1 U7081 ( .A1(n6024), .A2(n5756), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5811), .ZN(n6027) );
  XNOR2_X1 U7082 ( .A(n6025), .B(n6037), .ZN(n6026) );
  XNOR2_X1 U7083 ( .A(n6027), .B(n6026), .ZN(n6317) );
  OR2_X1 U7084 ( .A1(n6029), .A2(n6028), .ZN(n6030) );
  AND2_X1 U7085 ( .A1(n6031), .A2(n6030), .ZN(n6235) );
  INV_X1 U7086 ( .A(n6235), .ZN(n6032) );
  NAND2_X1 U7087 ( .A1(n3009), .A2(REIP_REG_11__SCAN_IN), .ZN(n6309) );
  OAI21_X1 U7088 ( .B1(n6032), .B2(n6434), .A(n6309), .ZN(n6035) );
  NOR2_X1 U7089 ( .A1(n6033), .A2(n6037), .ZN(n6034) );
  AOI211_X1 U7090 ( .C1(n6037), .C2(n6036), .A(n6035), .B(n6034), .ZN(n6038)
         );
  OAI21_X1 U7091 ( .B1(n6317), .B2(n6351), .A(n6038), .ZN(U3007) );
  OAI21_X1 U7092 ( .B1(n4480), .B2(STATEBS16_REG_SCAN_IN), .A(n6666), .ZN(
        n6040) );
  OAI22_X1 U7093 ( .A1(n6040), .A2(n6042), .B1(n6044), .B2(n6039), .ZN(n6041)
         );
  MUX2_X1 U7094 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n6041), .S(n6443), 
        .Z(U3464) );
  XNOR2_X1 U7095 ( .A(n6043), .B(n6042), .ZN(n6045) );
  OAI22_X1 U7096 ( .A1(n6045), .A2(n6497), .B1(n6044), .B2(n4483), .ZN(n6046)
         );
  MUX2_X1 U7097 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n6046), .S(n6443), 
        .Z(U3463) );
  INV_X1 U7098 ( .A(n6047), .ZN(n6051) );
  OAI22_X1 U7099 ( .A1(n6051), .A2(n6050), .B1(n6049), .B2(n6048), .ZN(n6053)
         );
  MUX2_X1 U7100 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6053), .S(n6052), 
        .Z(U3456) );
  NAND2_X1 U7101 ( .A1(n6055), .A2(n6054), .ZN(n6680) );
  AOI21_X1 U7102 ( .B1(n6099), .B2(n6680), .A(n6104), .ZN(n6063) );
  OAI21_X1 U7103 ( .B1(n6057), .B2(n6056), .A(n6666), .ZN(n6062) );
  OR2_X1 U7104 ( .A1(n6058), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6094)
         );
  AOI211_X1 U7105 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6094), .A(n6060), .B(
        n6059), .ZN(n6061) );
  NAND2_X1 U7106 ( .A1(n6092), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6070) );
  AOI22_X1 U7107 ( .A1(n6067), .A2(n6066), .B1(n6065), .B2(n6064), .ZN(n6093)
         );
  OAI22_X1 U7108 ( .A1(n6494), .A2(n6094), .B1(n6093), .B2(n6505), .ZN(n6068)
         );
  AOI21_X1 U7109 ( .B1(n6539), .B2(n6502), .A(n6068), .ZN(n6069) );
  OAI211_X1 U7110 ( .C1(n6099), .C2(n6495), .A(n6070), .B(n6069), .ZN(U3084)
         );
  NAND2_X1 U7111 ( .A1(n6092), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6073) );
  OAI22_X1 U7112 ( .A1(n6544), .A2(n6094), .B1(n6093), .B2(n6510), .ZN(n6071)
         );
  AOI21_X1 U7113 ( .B1(n6539), .B2(n6473), .A(n6071), .ZN(n6072) );
  OAI211_X1 U7114 ( .C1(n6099), .C2(n6545), .A(n6073), .B(n6072), .ZN(U3085)
         );
  NAND2_X1 U7115 ( .A1(n6092), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6076) );
  OAI22_X1 U7116 ( .A1(n6676), .A2(n6094), .B1(n6093), .B2(n6682), .ZN(n6074)
         );
  AOI21_X1 U7117 ( .B1(n6539), .B2(n6477), .A(n6074), .ZN(n6075) );
  OAI211_X1 U7118 ( .C1(n6099), .C2(n6681), .A(n6076), .B(n6075), .ZN(U3086)
         );
  NAND2_X1 U7119 ( .A1(n6092), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6079) );
  OAI22_X1 U7120 ( .A1(n6511), .A2(n6094), .B1(n6093), .B2(n6517), .ZN(n6077)
         );
  AOI21_X1 U7121 ( .B1(n6539), .B2(n6485), .A(n6077), .ZN(n6078) );
  OAI211_X1 U7122 ( .C1(n6099), .C2(n6489), .A(n6079), .B(n6078), .ZN(U3087)
         );
  NAND2_X1 U7123 ( .A1(n6092), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6082) );
  OAI22_X1 U7124 ( .A1(n6518), .A2(n6094), .B1(n6093), .B2(n6525), .ZN(n6080)
         );
  AOI21_X1 U7125 ( .B1(n6539), .B2(n6522), .A(n6080), .ZN(n6081) );
  OAI211_X1 U7126 ( .C1(n6099), .C2(n6519), .A(n6082), .B(n6081), .ZN(U3088)
         );
  NAND2_X1 U7127 ( .A1(n6092), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6086) );
  OAI22_X1 U7128 ( .A1(n6555), .A2(n6094), .B1(n6093), .B2(n6530), .ZN(n6083)
         );
  AOI21_X1 U7129 ( .B1(n6539), .B2(n6084), .A(n6083), .ZN(n6085) );
  OAI211_X1 U7130 ( .C1(n6099), .C2(n6556), .A(n6086), .B(n6085), .ZN(U3089)
         );
  NAND2_X1 U7131 ( .A1(n6092), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6090) );
  OAI22_X1 U7132 ( .A1(n6531), .A2(n6094), .B1(n6093), .B2(n6537), .ZN(n6087)
         );
  AOI21_X1 U7133 ( .B1(n6539), .B2(n6088), .A(n6087), .ZN(n6089) );
  OAI211_X1 U7134 ( .C1(n6099), .C2(n6091), .A(n6090), .B(n6089), .ZN(U3090)
         );
  NAND2_X1 U7135 ( .A1(n6092), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6098) );
  OAI22_X1 U7136 ( .A1(n6563), .A2(n6094), .B1(n6093), .B2(n6543), .ZN(n6095)
         );
  AOI21_X1 U7137 ( .B1(n6539), .B2(n6096), .A(n6095), .ZN(n6097) );
  OAI211_X1 U7138 ( .C1(n6099), .C2(n6564), .A(n6098), .B(n6097), .ZN(U3091)
         );
  AND2_X1 U7139 ( .A1(n6276), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7140 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6809) );
  AOI221_X2 U7141 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_0__SCAN_IN), .C1(
        n6100), .C2(STATE_REG_0__SCAN_IN), .A(n6675), .ZN(n6654) );
  OAI21_X1 U7142 ( .B1(n6809), .B2(n6101), .A(n6652), .ZN(U2789) );
  NOR2_X1 U7143 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6103) );
  OAI21_X1 U7144 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6103), .A(n6663), .ZN(n6102)
         );
  OAI21_X1 U7145 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6663), .A(n6102), .ZN(
        U2791) );
  OAI21_X1 U7146 ( .B1(BS16_N), .B2(n6103), .A(n6654), .ZN(n6653) );
  OAI21_X1 U7147 ( .B1(n6654), .B2(n6104), .A(n6653), .ZN(U2792) );
  OAI21_X1 U7148 ( .B1(n6106), .B2(n6105), .A(n6316), .ZN(U2793) );
  NOR4_X1 U7149 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n6116) );
  NOR4_X1 U7150 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6115) );
  INV_X1 U7151 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6736) );
  INV_X1 U7152 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6761) );
  INV_X1 U7153 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6760) );
  INV_X1 U7154 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6785) );
  NAND4_X1 U7155 ( .A1(n6736), .A2(n6761), .A3(n6760), .A4(n6785), .ZN(n6113)
         );
  INV_X1 U7156 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6776) );
  INV_X1 U7157 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6717) );
  INV_X1 U7158 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n6722) );
  INV_X1 U7159 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6728) );
  OAI211_X1 U7160 ( .C1(n6776), .C2(n6717), .A(n6722), .B(n6728), .ZN(n6112)
         );
  NOR4_X1 U7161 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6110) );
  NOR4_X1 U7162 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6109) );
  NOR4_X1 U7163 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6108) );
  NOR4_X1 U7164 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n6107) );
  NAND4_X1 U7165 ( .A1(n6110), .A2(n6109), .A3(n6108), .A4(n6107), .ZN(n6111)
         );
  NOR3_X1 U7166 ( .A1(n6113), .A2(n6112), .A3(n6111), .ZN(n6114) );
  NAND3_X1 U7167 ( .A1(n6116), .A2(n6115), .A3(n6114), .ZN(n6660) );
  INV_X1 U7168 ( .A(n6660), .ZN(n6658) );
  NOR3_X1 U7169 ( .A1(DATAWIDTH_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(REIP_REG_0__SCAN_IN), .ZN(n6119) );
  NOR2_X1 U7170 ( .A1(n6660), .A2(REIP_REG_1__SCAN_IN), .ZN(n6659) );
  INV_X1 U7171 ( .A(n6659), .ZN(n6117) );
  OAI22_X1 U7172 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(n6658), .B1(n6119), 
        .B2(n6117), .ZN(n6118) );
  INV_X1 U7173 ( .A(n6118), .ZN(U2794) );
  AOI21_X1 U7174 ( .B1(n6656), .B2(n6717), .A(n6119), .ZN(n6120) );
  INV_X1 U7175 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6748) );
  AOI22_X1 U7176 ( .A1(n6658), .A2(n6120), .B1(n6748), .B2(n6660), .ZN(U2795)
         );
  INV_X1 U7177 ( .A(n6132), .ZN(n6125) );
  AOI21_X1 U7178 ( .B1(n6214), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6212), 
        .ZN(n6121) );
  OAI211_X1 U7179 ( .C1(n6171), .C2(n6230), .A(n6122), .B(n6121), .ZN(n6124)
         );
  NOR2_X1 U7180 ( .A1(n6227), .A2(n6199), .ZN(n6123) );
  AOI211_X1 U7181 ( .C1(REIP_REG_15__SCAN_IN), .C2(n6125), .A(n6124), .B(n6123), .ZN(n6129) );
  AOI22_X1 U7182 ( .A1(n6127), .A2(n6189), .B1(n6211), .B2(n6126), .ZN(n6128)
         );
  NAND2_X1 U7183 ( .A1(n6129), .A2(n6128), .ZN(U2812) );
  INV_X1 U7184 ( .A(n6130), .ZN(n6131) );
  AOI21_X1 U7185 ( .B1(n6207), .B2(n6131), .A(REIP_REG_14__SCAN_IN), .ZN(n6133) );
  NOR2_X1 U7186 ( .A1(n6133), .A2(n6132), .ZN(n6135) );
  OAI21_X1 U7187 ( .B1(n6143), .B2(n6812), .A(n6197), .ZN(n6134) );
  AOI211_X1 U7188 ( .C1(n6222), .C2(EBX_REG_14__SCAN_IN), .A(n6135), .B(n6134), 
        .ZN(n6140) );
  OAI22_X1 U7189 ( .A1(n6137), .A2(n6199), .B1(n6136), .B2(n6217), .ZN(n6138)
         );
  INV_X1 U7190 ( .A(n6138), .ZN(n6139) );
  OAI211_X1 U7191 ( .C1(n6184), .C2(n6141), .A(n6140), .B(n6139), .ZN(U2813)
         );
  NAND2_X1 U7192 ( .A1(n6207), .A2(n6149), .ZN(n6148) );
  INV_X1 U7193 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6620) );
  NOR3_X1 U7194 ( .A1(n6148), .A2(REIP_REG_13__SCAN_IN), .A3(n6620), .ZN(n6147) );
  INV_X1 U7195 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6142) );
  OAI21_X1 U7196 ( .B1(n6143), .B2(n6142), .A(n6197), .ZN(n6144) );
  AOI21_X1 U7197 ( .B1(n6222), .B2(EBX_REG_13__SCAN_IN), .A(n6144), .ZN(n6145)
         );
  OAI21_X1 U7198 ( .B1(n6184), .B2(n6231), .A(n6145), .ZN(n6146) );
  AOI211_X1 U7199 ( .C1(n6244), .C2(n6190), .A(n6147), .B(n6146), .ZN(n6154)
         );
  NOR2_X1 U7200 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6148), .ZN(n6163) );
  NOR2_X1 U7201 ( .A1(n6150), .A2(n6149), .ZN(n6168) );
  INV_X1 U7202 ( .A(n6168), .ZN(n6152) );
  NAND2_X1 U7203 ( .A1(n6152), .A2(n6151), .ZN(n6173) );
  OAI21_X1 U7204 ( .B1(n6163), .B2(n6173), .A(REIP_REG_13__SCAN_IN), .ZN(n6153) );
  OAI211_X1 U7205 ( .C1(n6217), .C2(n6155), .A(n6154), .B(n6153), .ZN(U2814)
         );
  AOI21_X1 U7206 ( .B1(n6214), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6212), 
        .ZN(n6156) );
  OAI21_X1 U7207 ( .B1(n6171), .B2(n6157), .A(n6156), .ZN(n6158) );
  AOI21_X1 U7208 ( .B1(n6173), .B2(REIP_REG_12__SCAN_IN), .A(n6158), .ZN(n6159) );
  OAI21_X1 U7209 ( .B1(n6160), .B2(n6199), .A(n6159), .ZN(n6161) );
  AOI21_X1 U7210 ( .B1(n6162), .B2(n6189), .A(n6161), .ZN(n6165) );
  INV_X1 U7211 ( .A(n6163), .ZN(n6164) );
  OAI211_X1 U7212 ( .C1(n6166), .C2(n6184), .A(n6165), .B(n6164), .ZN(U2815)
         );
  INV_X1 U7213 ( .A(n6167), .ZN(n6169) );
  AOI22_X1 U7214 ( .A1(n6211), .A2(n6235), .B1(n6169), .B2(n6168), .ZN(n6180)
         );
  OAI22_X1 U7215 ( .A1(n6171), .A2(n6237), .B1(n6170), .B2(n6143), .ZN(n6172)
         );
  AOI211_X1 U7216 ( .C1(REIP_REG_11__SCAN_IN), .C2(n6173), .A(n6212), .B(n6172), .ZN(n6179) );
  OAI21_X1 U7217 ( .B1(n6176), .B2(n6175), .A(n6174), .ZN(n6177) );
  INV_X1 U7218 ( .A(n6177), .ZN(n6313) );
  AOI22_X1 U7219 ( .A1(n6313), .A2(n6190), .B1(n6189), .B2(n6311), .ZN(n6178)
         );
  NAND3_X1 U7220 ( .A1(n6180), .A2(n6179), .A3(n6178), .ZN(U2816) );
  OAI21_X1 U7221 ( .B1(n6143), .B2(n6181), .A(n6197), .ZN(n6182) );
  AOI21_X1 U7222 ( .B1(n6222), .B2(EBX_REG_9__SCAN_IN), .A(n6182), .ZN(n6183)
         );
  OAI21_X1 U7223 ( .B1(n6184), .B2(n6359), .A(n6183), .ZN(n6185) );
  AOI21_X1 U7224 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6186), .A(n6185), .ZN(n6193)
         );
  INV_X1 U7225 ( .A(n6187), .ZN(n6191) );
  AOI22_X1 U7226 ( .A1(n6191), .A2(n6190), .B1(n6189), .B2(n6188), .ZN(n6192)
         );
  OAI211_X1 U7227 ( .C1(REIP_REG_9__SCAN_IN), .C2(n6194), .A(n6193), .B(n6192), 
        .ZN(U2818) );
  AOI22_X1 U7228 ( .A1(n6211), .A2(n6397), .B1(n6196), .B2(n6195), .ZN(n6205)
         );
  NAND2_X1 U7229 ( .A1(n6222), .A2(EBX_REG_6__SCAN_IN), .ZN(n6198) );
  OAI211_X1 U7230 ( .C1(n3583), .C2(n6143), .A(n6198), .B(n6197), .ZN(n6202)
         );
  NOR2_X1 U7231 ( .A1(n6200), .A2(n6199), .ZN(n6201) );
  AOI211_X1 U7232 ( .C1(REIP_REG_6__SCAN_IN), .C2(n6203), .A(n6202), .B(n6201), 
        .ZN(n6204) );
  OAI211_X1 U7233 ( .C1(n6325), .C2(n6217), .A(n6205), .B(n6204), .ZN(U2821)
         );
  NAND2_X1 U7234 ( .A1(n6207), .A2(n6206), .ZN(n6225) );
  INV_X1 U7235 ( .A(n6208), .ZN(n6410) );
  AOI22_X1 U7236 ( .A1(n6211), .A2(n6410), .B1(n6210), .B2(n6209), .ZN(n6224)
         );
  AOI21_X1 U7237 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6213), .A(n6212), .ZN(n6216)
         );
  NAND2_X1 U7238 ( .A1(n6214), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6215)
         );
  OAI211_X1 U7239 ( .C1(n6217), .C2(n6335), .A(n6216), .B(n6215), .ZN(n6221)
         );
  NOR2_X1 U7240 ( .A1(n6219), .A2(n6218), .ZN(n6220) );
  AOI211_X1 U7241 ( .C1(n6222), .C2(EBX_REG_4__SCAN_IN), .A(n6221), .B(n6220), 
        .ZN(n6223) );
  OAI211_X1 U7242 ( .C1(REIP_REG_4__SCAN_IN), .C2(n6225), .A(n6224), .B(n6223), 
        .ZN(U2823) );
  OAI22_X1 U7243 ( .A1(n6227), .A2(n5609), .B1(n5608), .B2(n6226), .ZN(n6228)
         );
  INV_X1 U7244 ( .A(n6228), .ZN(n6229) );
  OAI21_X1 U7245 ( .B1(n6243), .B2(n6230), .A(n6229), .ZN(U2844) );
  INV_X1 U7246 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6234) );
  INV_X1 U7247 ( .A(n6231), .ZN(n6232) );
  AOI22_X1 U7248 ( .A1(n6244), .A2(n6240), .B1(n6239), .B2(n6232), .ZN(n6233)
         );
  OAI21_X1 U7249 ( .B1(n6243), .B2(n6234), .A(n6233), .ZN(U2846) );
  AOI22_X1 U7250 ( .A1(n6313), .A2(n6240), .B1(n6239), .B2(n6235), .ZN(n6236)
         );
  OAI21_X1 U7251 ( .B1(n6243), .B2(n6237), .A(n6236), .ZN(U2848) );
  AOI22_X1 U7252 ( .A1(n6341), .A2(n6240), .B1(n6239), .B2(n6238), .ZN(n6241)
         );
  OAI21_X1 U7253 ( .B1(n6243), .B2(n6242), .A(n6241), .ZN(U2857) );
  INV_X1 U7254 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6824) );
  AOI22_X1 U7255 ( .A1(n6244), .A2(n6247), .B1(DATAI_13_), .B2(n6246), .ZN(
        n6245) );
  OAI21_X1 U7256 ( .B1(n6824), .B2(n6249), .A(n6245), .ZN(U2878) );
  INV_X1 U7257 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U7258 ( .A1(n6313), .A2(n6247), .B1(DATAI_11_), .B2(n6246), .ZN(
        n6248) );
  OAI21_X1 U7259 ( .B1(n6743), .B2(n6249), .A(n6248), .ZN(U2880) );
  INV_X1 U7260 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6797) );
  INV_X1 U7261 ( .A(n6250), .ZN(n6252) );
  AOI22_X1 U7262 ( .A1(n6276), .A2(DATAO_REG_28__SCAN_IN), .B1(n6252), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6251) );
  OAI21_X1 U7263 ( .B1(n6263), .B2(n6797), .A(n6251), .ZN(U2895) );
  INV_X1 U7264 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n6805) );
  INV_X1 U7265 ( .A(n6276), .ZN(n6254) );
  AOI22_X1 U7266 ( .A1(n6252), .A2(EAX_REG_21__SCAN_IN), .B1(
        UWORD_REG_5__SCAN_IN), .B2(n6664), .ZN(n6253) );
  OAI21_X1 U7267 ( .B1(n6805), .B2(n6254), .A(n6253), .ZN(U2902) );
  INV_X1 U7268 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6308) );
  AOI22_X1 U7269 ( .A1(n6664), .A2(LWORD_REG_15__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6255) );
  OAI21_X1 U7270 ( .B1(n6308), .B2(n6278), .A(n6255), .ZN(U2908) );
  INV_X1 U7271 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6257) );
  AOI22_X1 U7272 ( .A1(n6664), .A2(LWORD_REG_14__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6256) );
  OAI21_X1 U7273 ( .B1(n6257), .B2(n6278), .A(n6256), .ZN(U2909) );
  AOI22_X1 U7274 ( .A1(n6664), .A2(LWORD_REG_13__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6258) );
  OAI21_X1 U7275 ( .B1(n6824), .B2(n6278), .A(n6258), .ZN(U2910) );
  INV_X1 U7276 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6782) );
  AOI22_X1 U7277 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6261), .B1(n6276), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7278 ( .B1(n6263), .B2(n6782), .A(n6259), .ZN(U2911) );
  AOI22_X1 U7279 ( .A1(n6664), .A2(LWORD_REG_11__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6260) );
  OAI21_X1 U7280 ( .B1(n6743), .B2(n6278), .A(n6260), .ZN(U2912) );
  INV_X1 U7281 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6764) );
  AOI22_X1 U7282 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6261), .B1(n6276), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6262) );
  OAI21_X1 U7283 ( .B1(n6263), .B2(n6764), .A(n6262), .ZN(U2913) );
  INV_X1 U7284 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6265) );
  AOI22_X1 U7285 ( .A1(n6664), .A2(LWORD_REG_9__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6264) );
  OAI21_X1 U7286 ( .B1(n6265), .B2(n6278), .A(n6264), .ZN(U2914) );
  INV_X1 U7287 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6267) );
  AOI22_X1 U7288 ( .A1(n6664), .A2(LWORD_REG_8__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6266) );
  OAI21_X1 U7289 ( .B1(n6267), .B2(n6278), .A(n6266), .ZN(U2915) );
  AOI22_X1 U7290 ( .A1(n6664), .A2(LWORD_REG_7__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6268) );
  OAI21_X1 U7291 ( .B1(n4319), .B2(n6278), .A(n6268), .ZN(U2916) );
  AOI22_X1 U7292 ( .A1(n6664), .A2(LWORD_REG_6__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6269) );
  OAI21_X1 U7293 ( .B1(n3589), .B2(n6278), .A(n6269), .ZN(U2917) );
  AOI22_X1 U7294 ( .A1(n6664), .A2(LWORD_REG_5__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6270) );
  OAI21_X1 U7295 ( .B1(n6271), .B2(n6278), .A(n6270), .ZN(U2918) );
  AOI22_X1 U7296 ( .A1(n6664), .A2(LWORD_REG_4__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6272) );
  OAI21_X1 U7297 ( .B1(n6781), .B2(n6278), .A(n6272), .ZN(U2919) );
  AOI22_X1 U7298 ( .A1(n6664), .A2(LWORD_REG_3__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6273) );
  OAI21_X1 U7299 ( .B1(n6822), .B2(n6278), .A(n6273), .ZN(U2920) );
  AOI22_X1 U7300 ( .A1(n6664), .A2(LWORD_REG_2__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6274) );
  OAI21_X1 U7301 ( .B1(n4327), .B2(n6278), .A(n6274), .ZN(U2921) );
  AOI22_X1 U7302 ( .A1(n6664), .A2(LWORD_REG_1__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6275) );
  OAI21_X1 U7303 ( .B1(n6729), .B2(n6278), .A(n6275), .ZN(U2922) );
  AOI22_X1 U7304 ( .A1(n6664), .A2(LWORD_REG_0__SCAN_IN), .B1(n6276), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6277) );
  OAI21_X1 U7305 ( .B1(n4312), .B2(n6278), .A(n6277), .ZN(U2923) );
  AOI22_X1 U7306 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6301), .B1(n6305), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7307 ( .A1(n6304), .A2(DATAI_9_), .ZN(n6290) );
  NAND2_X1 U7308 ( .A1(n6279), .A2(n6290), .ZN(U2933) );
  INV_X1 U7309 ( .A(DATAI_10_), .ZN(n6280) );
  NOR2_X1 U7310 ( .A1(n6287), .A2(n6280), .ZN(n6292) );
  AOI21_X1 U7311 ( .B1(n6305), .B2(UWORD_REG_10__SCAN_IN), .A(n6292), .ZN(
        n6281) );
  OAI21_X1 U7312 ( .B1(n6282), .B2(n6307), .A(n6281), .ZN(U2934) );
  AOI22_X1 U7313 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6301), .B1(n6305), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7314 ( .A1(n6304), .A2(DATAI_11_), .ZN(n6294) );
  NAND2_X1 U7315 ( .A1(n6283), .A2(n6294), .ZN(U2935) );
  INV_X1 U7316 ( .A(DATAI_12_), .ZN(n6284) );
  NOR2_X1 U7317 ( .A1(n6287), .A2(n6284), .ZN(n6296) );
  AOI21_X1 U7318 ( .B1(n6301), .B2(EAX_REG_28__SCAN_IN), .A(n6296), .ZN(n6285)
         );
  OAI21_X1 U7319 ( .B1(n6797), .B2(n6298), .A(n6285), .ZN(U2936) );
  INV_X1 U7320 ( .A(DATAI_13_), .ZN(n6286) );
  NOR2_X1 U7321 ( .A1(n6287), .A2(n6286), .ZN(n6299) );
  AOI21_X1 U7322 ( .B1(n6305), .B2(UWORD_REG_13__SCAN_IN), .A(n6299), .ZN(
        n6288) );
  OAI21_X1 U7323 ( .B1(n3906), .B2(n6307), .A(n6288), .ZN(U2937) );
  AOI22_X1 U7324 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6301), .B1(n6305), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7325 ( .A1(n6304), .A2(DATAI_14_), .ZN(n6302) );
  NAND2_X1 U7326 ( .A1(n6289), .A2(n6302), .ZN(U2938) );
  AOI22_X1 U7327 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6301), .B1(n6305), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U7328 ( .A1(n6291), .A2(n6290), .ZN(U2948) );
  AOI21_X1 U7329 ( .B1(n6301), .B2(EAX_REG_10__SCAN_IN), .A(n6292), .ZN(n6293)
         );
  OAI21_X1 U7330 ( .B1(n6764), .B2(n6298), .A(n6293), .ZN(U2949) );
  AOI22_X1 U7331 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6301), .B1(n6305), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7332 ( .A1(n6295), .A2(n6294), .ZN(U2950) );
  AOI21_X1 U7333 ( .B1(n6301), .B2(EAX_REG_12__SCAN_IN), .A(n6296), .ZN(n6297)
         );
  OAI21_X1 U7334 ( .B1(n6782), .B2(n6298), .A(n6297), .ZN(U2951) );
  AOI21_X1 U7335 ( .B1(n6305), .B2(LWORD_REG_13__SCAN_IN), .A(n6299), .ZN(
        n6300) );
  OAI21_X1 U7336 ( .B1(n6824), .B2(n6307), .A(n6300), .ZN(U2952) );
  AOI22_X1 U7337 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6301), .B1(n6305), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7338 ( .A1(n6303), .A2(n6302), .ZN(U2953) );
  AOI22_X1 U7339 ( .A1(n6305), .A2(LWORD_REG_15__SCAN_IN), .B1(n6304), .B2(
        DATAI_15_), .ZN(n6306) );
  OAI21_X1 U7340 ( .B1(n6308), .B2(n6307), .A(n6306), .ZN(U2954) );
  INV_X1 U7341 ( .A(n6309), .ZN(n6310) );
  AOI21_X1 U7342 ( .B1(n6336), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6310), 
        .ZN(n6315) );
  AOI22_X1 U7343 ( .A1(n6313), .A2(n6332), .B1(n6312), .B2(n6311), .ZN(n6314)
         );
  OAI211_X1 U7344 ( .C1(n6317), .C2(n6316), .A(n6315), .B(n6314), .ZN(U2975)
         );
  AOI22_X1 U7345 ( .A1(n6336), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n3009), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6324) );
  OAI21_X1 U7346 ( .B1(n6320), .B2(n6319), .A(n6318), .ZN(n6321) );
  INV_X1 U7347 ( .A(n6321), .ZN(n6396) );
  AOI22_X1 U7348 ( .A1(n6396), .A2(n6340), .B1(n6332), .B2(n6322), .ZN(n6323)
         );
  OAI211_X1 U7349 ( .C1(n6345), .C2(n6325), .A(n6324), .B(n6323), .ZN(U2980)
         );
  INV_X1 U7350 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6326) );
  NOR2_X1 U7351 ( .A1(n6435), .A2(n6326), .ZN(n6409) );
  AOI21_X1 U7352 ( .B1(n6336), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6409), 
        .ZN(n6334) );
  OAI21_X1 U7353 ( .B1(n6329), .B2(n6328), .A(n6327), .ZN(n6330) );
  INV_X1 U7354 ( .A(n6330), .ZN(n6414) );
  AOI22_X1 U7355 ( .A1(n6414), .A2(n6340), .B1(n6332), .B2(n6331), .ZN(n6333)
         );
  OAI211_X1 U7356 ( .C1(n6345), .C2(n6335), .A(n6334), .B(n6333), .ZN(U2982)
         );
  AOI22_X1 U7357 ( .A1(n6336), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n3009), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6343) );
  XNOR2_X1 U7358 ( .A(n6337), .B(n6388), .ZN(n6338) );
  XNOR2_X1 U7359 ( .A(n6339), .B(n6338), .ZN(n6439) );
  AOI22_X1 U7360 ( .A1(n6341), .A2(n6332), .B1(n6340), .B2(n6439), .ZN(n6342)
         );
  OAI211_X1 U7361 ( .C1(n6345), .C2(n6344), .A(n6343), .B(n6342), .ZN(U2984)
         );
  INV_X1 U7362 ( .A(n6346), .ZN(n6412) );
  INV_X1 U7363 ( .A(n6387), .ZN(n6348) );
  OAI22_X1 U7364 ( .A1(n6349), .A2(n6412), .B1(n6348), .B2(n6347), .ZN(n6382)
         );
  AOI21_X1 U7365 ( .B1(n6369), .B2(n6395), .A(n6382), .ZN(n6368) );
  OAI222_X1 U7366 ( .A1(n6352), .A2(n6434), .B1(n6351), .B2(n6350), .C1(n6435), 
        .C2(n6616), .ZN(n6353) );
  INV_X1 U7367 ( .A(n6353), .ZN(n6358) );
  INV_X1 U7368 ( .A(n6413), .ZN(n6354) );
  NAND3_X1 U7369 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6428), .ZN(n6392) );
  NAND2_X1 U7370 ( .A1(n6355), .A2(n6419), .ZN(n6386) );
  NOR2_X1 U7371 ( .A1(n6369), .A2(n6386), .ZN(n6363) );
  OAI211_X1 U7372 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6363), .B(n6356), .ZN(n6357) );
  OAI211_X1 U7373 ( .C1(n6368), .C2(n5812), .A(n6358), .B(n6357), .ZN(U3008)
         );
  INV_X1 U7374 ( .A(n6359), .ZN(n6362) );
  INV_X1 U7375 ( .A(n6360), .ZN(n6361) );
  AOI21_X1 U7376 ( .B1(n6422), .B2(n6362), .A(n6361), .ZN(n6366) );
  AOI22_X1 U7377 ( .A1(n6364), .A2(n6438), .B1(n6363), .B2(n6367), .ZN(n6365)
         );
  OAI211_X1 U7378 ( .C1(n6368), .C2(n6367), .A(n6366), .B(n6365), .ZN(U3009)
         );
  OAI21_X1 U7379 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6369), .ZN(n6377) );
  INV_X1 U7380 ( .A(n6370), .ZN(n6371) );
  AOI21_X1 U7381 ( .B1(n6422), .B2(n6372), .A(n6371), .ZN(n6376) );
  INV_X1 U7382 ( .A(n6373), .ZN(n6374) );
  AOI22_X1 U7383 ( .A1(n6374), .A2(n6438), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n6382), .ZN(n6375) );
  OAI211_X1 U7384 ( .C1(n6386), .C2(n6377), .A(n6376), .B(n6375), .ZN(U3010)
         );
  INV_X1 U7385 ( .A(n6378), .ZN(n6379) );
  AOI21_X1 U7386 ( .B1(n6422), .B2(n6380), .A(n6379), .ZN(n6385) );
  INV_X1 U7387 ( .A(n6381), .ZN(n6383) );
  AOI22_X1 U7388 ( .A1(n6383), .A2(n6438), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6382), .ZN(n6384) );
  OAI211_X1 U7389 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6386), .A(n6385), 
        .B(n6384), .ZN(U3011) );
  NAND3_X1 U7390 ( .A1(n6401), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6419), 
        .ZN(n6400) );
  OAI21_X1 U7391 ( .B1(n6389), .B2(n6388), .A(n6387), .ZN(n6411) );
  OAI21_X1 U7392 ( .B1(n6391), .B2(n6390), .A(n6411), .ZN(n6437) );
  NOR2_X1 U7393 ( .A1(n6429), .A2(n6742), .ZN(n6393) );
  OAI22_X1 U7394 ( .A1(n6393), .A2(n6432), .B1(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .B2(n6392), .ZN(n6394) );
  AOI211_X1 U7395 ( .C1(n6415), .C2(n6395), .A(n6437), .B(n6394), .ZN(n6408)
         );
  AOI222_X1 U7396 ( .A1(REIP_REG_6__SCAN_IN), .A2(n3009), .B1(n6422), .B2(
        n6397), .C1(n6438), .C2(n6396), .ZN(n6398) );
  OAI221_X1 U7397 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6400), .C1(n6399), .C2(n6408), .A(n6398), .ZN(U3012) );
  AOI21_X1 U7398 ( .B1(n6401), .B2(n6419), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6407) );
  INV_X1 U7399 ( .A(n6402), .ZN(n6404) );
  AOI22_X1 U7400 ( .A1(n6404), .A2(n6438), .B1(n6422), .B2(n6403), .ZN(n6406)
         );
  OAI211_X1 U7401 ( .C1(n6408), .C2(n6407), .A(n6406), .B(n6405), .ZN(U3013)
         );
  AOI21_X1 U7402 ( .B1(n6422), .B2(n6410), .A(n6409), .ZN(n6418) );
  OAI21_X1 U7403 ( .B1(n6413), .B2(n6412), .A(n6411), .ZN(n6424) );
  AOI22_X1 U7404 ( .A1(n6424), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n6438), 
        .B2(n6414), .ZN(n6417) );
  OAI211_X1 U7405 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6419), .B(n6415), .ZN(n6416) );
  NAND3_X1 U7406 ( .A1(n6418), .A2(n6417), .A3(n6416), .ZN(U3014) );
  INV_X1 U7407 ( .A(n6419), .ZN(n6427) );
  AOI21_X1 U7408 ( .B1(n6422), .B2(n6421), .A(n6420), .ZN(n6426) );
  AOI22_X1 U7409 ( .A1(n6424), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n6438), 
        .B2(n6423), .ZN(n6425) );
  OAI211_X1 U7410 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n6427), .A(n6426), 
        .B(n6425), .ZN(U3015) );
  NAND2_X1 U7411 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6428), .ZN(n6442)
         );
  AOI21_X1 U7412 ( .B1(n6430), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6429), 
        .ZN(n6431) );
  OAI222_X1 U7413 ( .A1(n6435), .A2(n6603), .B1(n6434), .B2(n6433), .C1(n6432), 
        .C2(n6431), .ZN(n6436) );
  INV_X1 U7414 ( .A(n6436), .ZN(n6441) );
  AOI22_X1 U7415 ( .A1(n6439), .A2(n6438), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6437), .ZN(n6440) );
  OAI211_X1 U7416 ( .C1(INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n6442), .A(n6441), 
        .B(n6440), .ZN(U3016) );
  NOR2_X1 U7417 ( .A1(n6444), .A2(n6443), .ZN(U3019) );
  AOI22_X1 U7418 ( .A1(n6461), .A2(n6507), .B1(n6460), .B2(n6472), .ZN(n6446)
         );
  AOI22_X1 U7419 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6464), .B1(n6547), 
        .B2(n6462), .ZN(n6445) );
  OAI211_X1 U7420 ( .C1(n6467), .C2(n6550), .A(n6446), .B(n6445), .ZN(U3045)
         );
  AOI22_X1 U7421 ( .A1(n6461), .A2(n6447), .B1(n6460), .B2(n6476), .ZN(n6449)
         );
  AOI22_X1 U7422 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6464), .B1(n6552), 
        .B2(n6462), .ZN(n6448) );
  OAI211_X1 U7423 ( .C1(n6467), .C2(n6678), .A(n6449), .B(n6448), .ZN(U3046)
         );
  AOI22_X1 U7424 ( .A1(n6461), .A2(n6451), .B1(n6460), .B2(n6450), .ZN(n6454)
         );
  AOI22_X1 U7425 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6464), .B1(n6452), 
        .B2(n6462), .ZN(n6453) );
  OAI211_X1 U7426 ( .C1(n6467), .C2(n6455), .A(n6454), .B(n6453), .ZN(U3048)
         );
  AOI22_X1 U7427 ( .A1(n6461), .A2(n6527), .B1(n6460), .B2(n6456), .ZN(n6458)
         );
  AOI22_X1 U7428 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6464), .B1(n6558), 
        .B2(n6462), .ZN(n6457) );
  OAI211_X1 U7429 ( .C1(n6467), .C2(n6561), .A(n6458), .B(n6457), .ZN(U3049)
         );
  AOI22_X1 U7430 ( .A1(n6461), .A2(n6534), .B1(n6460), .B2(n6459), .ZN(n6466)
         );
  AOI22_X1 U7431 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6464), .B1(n6463), 
        .B2(n6462), .ZN(n6465) );
  OAI211_X1 U7432 ( .C1(n6467), .C2(n6532), .A(n6466), .B(n6465), .ZN(U3050)
         );
  AOI22_X1 U7433 ( .A1(n6469), .A2(n6482), .B1(n6481), .B2(n6468), .ZN(n6471)
         );
  AOI22_X1 U7434 ( .A1(n6486), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6502), 
        .B2(n6484), .ZN(n6470) );
  OAI211_X1 U7435 ( .C1(n6495), .C2(n6679), .A(n6471), .B(n6470), .ZN(U3068)
         );
  AOI22_X1 U7436 ( .A1(n6472), .A2(n6482), .B1(n6481), .B2(n6547), .ZN(n6475)
         );
  AOI22_X1 U7437 ( .A1(n6486), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6473), 
        .B2(n6484), .ZN(n6474) );
  OAI211_X1 U7438 ( .C1(n6545), .C2(n6679), .A(n6475), .B(n6474), .ZN(U3069)
         );
  AOI22_X1 U7439 ( .A1(n6476), .A2(n6482), .B1(n6481), .B2(n6552), .ZN(n6479)
         );
  AOI22_X1 U7440 ( .A1(n6486), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6477), 
        .B2(n6484), .ZN(n6478) );
  OAI211_X1 U7441 ( .C1(n6681), .C2(n6679), .A(n6479), .B(n6478), .ZN(U3070)
         );
  AOI22_X1 U7442 ( .A1(n6483), .A2(n6482), .B1(n6481), .B2(n6480), .ZN(n6488)
         );
  AOI22_X1 U7443 ( .A1(n6486), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6485), 
        .B2(n6484), .ZN(n6487) );
  OAI211_X1 U7444 ( .C1(n6489), .C2(n6679), .A(n6488), .B(n6487), .ZN(U3071)
         );
  OAI21_X1 U7445 ( .B1(n6491), .B2(n6490), .A(n6677), .ZN(n6492) );
  AND2_X1 U7446 ( .A1(n6492), .A2(n6666), .ZN(n6493) );
  OAI22_X1 U7447 ( .A1(n6680), .A2(n6495), .B1(n6677), .B2(n6494), .ZN(n6496)
         );
  INV_X1 U7448 ( .A(n6496), .ZN(n6504) );
  NOR2_X1 U7449 ( .A1(n6498), .A2(n6497), .ZN(n6501) );
  AOI22_X1 U7450 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6686), .B1(n6502), 
        .B2(n6521), .ZN(n6503) );
  OAI211_X1 U7451 ( .C1(n6683), .C2(n6505), .A(n6504), .B(n6503), .ZN(U3076)
         );
  OAI22_X1 U7452 ( .A1(n6679), .A2(n6550), .B1(n6677), .B2(n6544), .ZN(n6506)
         );
  INV_X1 U7453 ( .A(n6506), .ZN(n6509) );
  AOI22_X1 U7454 ( .A1(n6686), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n6507), 
        .B2(n6539), .ZN(n6508) );
  OAI211_X1 U7455 ( .C1(n6683), .C2(n6510), .A(n6509), .B(n6508), .ZN(U3077)
         );
  OAI22_X1 U7456 ( .A1(n6679), .A2(n6512), .B1(n6677), .B2(n6511), .ZN(n6513)
         );
  INV_X1 U7457 ( .A(n6513), .ZN(n6516) );
  AOI22_X1 U7458 ( .A1(n6686), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n6514), 
        .B2(n6539), .ZN(n6515) );
  OAI211_X1 U7459 ( .C1(n6683), .C2(n6517), .A(n6516), .B(n6515), .ZN(U3079)
         );
  OAI22_X1 U7460 ( .A1(n6680), .A2(n6519), .B1(n6677), .B2(n6518), .ZN(n6520)
         );
  INV_X1 U7461 ( .A(n6520), .ZN(n6524) );
  AOI22_X1 U7462 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6686), .B1(n6522), 
        .B2(n6521), .ZN(n6523) );
  OAI211_X1 U7463 ( .C1(n6683), .C2(n6525), .A(n6524), .B(n6523), .ZN(U3080)
         );
  OAI22_X1 U7464 ( .A1(n6679), .A2(n6561), .B1(n6677), .B2(n6555), .ZN(n6526)
         );
  INV_X1 U7465 ( .A(n6526), .ZN(n6529) );
  AOI22_X1 U7466 ( .A1(n6686), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n6527), 
        .B2(n6539), .ZN(n6528) );
  OAI211_X1 U7467 ( .C1(n6683), .C2(n6530), .A(n6529), .B(n6528), .ZN(U3081)
         );
  OAI22_X1 U7468 ( .A1(n6679), .A2(n6532), .B1(n6677), .B2(n6531), .ZN(n6533)
         );
  INV_X1 U7469 ( .A(n6533), .ZN(n6536) );
  AOI22_X1 U7470 ( .A1(n6686), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n6534), 
        .B2(n6539), .ZN(n6535) );
  OAI211_X1 U7471 ( .C1(n6683), .C2(n6537), .A(n6536), .B(n6535), .ZN(U3082)
         );
  OAI22_X1 U7472 ( .A1(n6679), .A2(n6573), .B1(n6677), .B2(n6563), .ZN(n6538)
         );
  INV_X1 U7473 ( .A(n6538), .ZN(n6542) );
  AOI22_X1 U7474 ( .A1(n6686), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n6540), 
        .B2(n6539), .ZN(n6541) );
  OAI211_X1 U7475 ( .C1(n6683), .C2(n6543), .A(n6542), .B(n6541), .ZN(U3083)
         );
  OAI22_X1 U7476 ( .A1(n6565), .A2(n6545), .B1(n6544), .B2(n6562), .ZN(n6546)
         );
  INV_X1 U7477 ( .A(n6546), .ZN(n6549) );
  AOI22_X1 U7478 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6569), .B1(n6547), 
        .B2(n6567), .ZN(n6548) );
  OAI211_X1 U7479 ( .C1(n6550), .C2(n6572), .A(n6549), .B(n6548), .ZN(U3109)
         );
  OAI22_X1 U7480 ( .A1(n6565), .A2(n6681), .B1(n6676), .B2(n6562), .ZN(n6551)
         );
  INV_X1 U7481 ( .A(n6551), .ZN(n6554) );
  AOI22_X1 U7482 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6569), .B1(n6552), 
        .B2(n6567), .ZN(n6553) );
  OAI211_X1 U7483 ( .C1(n6678), .C2(n6572), .A(n6554), .B(n6553), .ZN(U3110)
         );
  OAI22_X1 U7484 ( .A1(n6565), .A2(n6556), .B1(n6555), .B2(n6562), .ZN(n6557)
         );
  INV_X1 U7485 ( .A(n6557), .ZN(n6560) );
  AOI22_X1 U7486 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6569), .B1(n6558), 
        .B2(n6567), .ZN(n6559) );
  OAI211_X1 U7487 ( .C1(n6561), .C2(n6572), .A(n6560), .B(n6559), .ZN(U3113)
         );
  OAI22_X1 U7488 ( .A1(n6565), .A2(n6564), .B1(n6563), .B2(n6562), .ZN(n6566)
         );
  INV_X1 U7489 ( .A(n6566), .ZN(n6571) );
  AOI22_X1 U7490 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6569), .B1(n6568), 
        .B2(n6567), .ZN(n6570) );
  OAI211_X1 U7491 ( .C1(n6573), .C2(n6572), .A(n6571), .B(n6570), .ZN(U3115)
         );
  INV_X1 U7492 ( .A(n6574), .ZN(n6584) );
  NAND2_X1 U7493 ( .A1(n6575), .A2(READY_N), .ZN(n6595) );
  NAND2_X1 U7494 ( .A1(n6592), .A2(n6595), .ZN(n6585) );
  OAI21_X1 U7495 ( .B1(n6585), .B2(n6576), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6578) );
  AND2_X1 U7496 ( .A1(n6578), .A2(n6577), .ZN(n6583) );
  OAI211_X1 U7497 ( .C1(n6581), .C2(n6580), .A(n6579), .B(n6592), .ZN(n6582)
         );
  OAI211_X1 U7498 ( .C1(n6584), .C2(n6587), .A(n6583), .B(n6582), .ZN(U3148)
         );
  NOR2_X1 U7499 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6600) );
  INV_X1 U7500 ( .A(n6600), .ZN(n6586) );
  NAND3_X1 U7501 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6586), .A3(n6585), .ZN(
        n6594) );
  OAI21_X1 U7502 ( .B1(n6588), .B2(READY_N), .A(n6587), .ZN(n6591) );
  INV_X1 U7503 ( .A(n6589), .ZN(n6590) );
  AOI21_X1 U7504 ( .B1(n6592), .B2(n6591), .A(n6590), .ZN(n6593) );
  NAND2_X1 U7505 ( .A1(n6594), .A2(n6593), .ZN(U3149) );
  INV_X1 U7506 ( .A(n6670), .ZN(n6597) );
  NAND3_X1 U7507 ( .A1(n6597), .A2(n6596), .A3(n6595), .ZN(n6599) );
  OAI21_X1 U7508 ( .B1(n6600), .B2(n6599), .A(n6598), .ZN(U3150) );
  AND2_X1 U7509 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6652), .ZN(U3151) );
  AND2_X1 U7510 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6652), .ZN(U3152) );
  NOR2_X1 U7511 ( .A1(n6654), .A2(n6722), .ZN(U3153) );
  NOR2_X1 U7512 ( .A1(n6654), .A2(n6785), .ZN(U3154) );
  AND2_X1 U7513 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6652), .ZN(U3155) );
  AND2_X1 U7514 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6652), .ZN(U3156) );
  INV_X1 U7515 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6806) );
  NOR2_X1 U7516 ( .A1(n6654), .A2(n6806), .ZN(U3157) );
  AND2_X1 U7517 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6652), .ZN(U3158) );
  NOR2_X1 U7518 ( .A1(n6654), .A2(n6736), .ZN(U3159) );
  AND2_X1 U7519 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6652), .ZN(U3160) );
  AND2_X1 U7520 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6652), .ZN(U3161) );
  AND2_X1 U7521 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6652), .ZN(U3162) );
  AND2_X1 U7522 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6652), .ZN(U3163) );
  AND2_X1 U7523 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6652), .ZN(U3164) );
  AND2_X1 U7524 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6652), .ZN(U3165) );
  AND2_X1 U7525 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6652), .ZN(U3166) );
  AND2_X1 U7526 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6652), .ZN(U3167) );
  AND2_X1 U7527 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6652), .ZN(U3168) );
  AND2_X1 U7528 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6652), .ZN(U3169) );
  AND2_X1 U7529 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6652), .ZN(U3170) );
  AND2_X1 U7530 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6652), .ZN(U3171) );
  NOR2_X1 U7531 ( .A1(n6654), .A2(n6728), .ZN(U3172) );
  AND2_X1 U7532 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6652), .ZN(U3173) );
  NOR2_X1 U7533 ( .A1(n6654), .A2(n6760), .ZN(U3174) );
  AND2_X1 U7534 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6652), .ZN(U3175) );
  AND2_X1 U7535 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6652), .ZN(U3176) );
  NOR2_X1 U7536 ( .A1(n6654), .A2(n6761), .ZN(U3177) );
  AND2_X1 U7537 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6652), .ZN(U3178) );
  AND2_X1 U7538 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6652), .ZN(U3179) );
  AND2_X1 U7539 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6652), .ZN(U3180) );
  NAND2_X1 U7540 ( .A1(n6675), .A2(n6601), .ZN(n6649) );
  NOR2_X2 U7541 ( .A1(n6601), .A2(n6663), .ZN(n6647) );
  AOI22_X1 U7542 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6663), .ZN(n6602) );
  OAI21_X1 U7543 ( .B1(n6603), .B2(n6649), .A(n6602), .ZN(U3184) );
  AOI22_X1 U7544 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6663), .ZN(n6604) );
  OAI21_X1 U7545 ( .B1(n4655), .B2(n6649), .A(n6604), .ZN(U3185) );
  INV_X1 U7546 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6747) );
  OAI222_X1 U7547 ( .A1(n6645), .A2(n4655), .B1(n6747), .B2(n6675), .C1(n6326), 
        .C2(n6649), .ZN(U3186) );
  AOI22_X1 U7548 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6663), .ZN(n6605) );
  OAI21_X1 U7549 ( .B1(n6606), .B2(n6649), .A(n6605), .ZN(U3187) );
  INV_X1 U7550 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6608) );
  AOI22_X1 U7551 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6663), .ZN(n6607) );
  OAI21_X1 U7552 ( .B1(n6608), .B2(n6649), .A(n6607), .ZN(U3188) );
  AOI22_X1 U7553 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6663), .ZN(n6609) );
  OAI21_X1 U7554 ( .B1(n6610), .B2(n6649), .A(n6609), .ZN(U3189) );
  AOI22_X1 U7555 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6663), .ZN(n6611) );
  OAI21_X1 U7556 ( .B1(n6612), .B2(n6649), .A(n6611), .ZN(U3190) );
  AOI22_X1 U7557 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6663), .ZN(n6613) );
  OAI21_X1 U7558 ( .B1(n6614), .B2(n6649), .A(n6613), .ZN(U3191) );
  AOI22_X1 U7559 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6663), .ZN(n6615) );
  OAI21_X1 U7560 ( .B1(n6616), .B2(n6649), .A(n6615), .ZN(U3192) );
  AOI22_X1 U7561 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6663), .ZN(n6617) );
  OAI21_X1 U7562 ( .B1(n6618), .B2(n6649), .A(n6617), .ZN(U3193) );
  INV_X1 U7563 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6763) );
  OAI222_X1 U7564 ( .A1(n6645), .A2(n6618), .B1(n6763), .B2(n6675), .C1(n6620), 
        .C2(n6649), .ZN(U3194) );
  INV_X1 U7565 ( .A(n6649), .ZN(n6643) );
  AOI22_X1 U7566 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6663), .ZN(n6619) );
  OAI21_X1 U7567 ( .B1(n6620), .B2(n6645), .A(n6619), .ZN(U3195) );
  AOI22_X1 U7568 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6663), .ZN(n6621) );
  OAI21_X1 U7569 ( .B1(n6623), .B2(n6649), .A(n6621), .ZN(U3196) );
  AOI22_X1 U7570 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6663), .ZN(n6622) );
  OAI21_X1 U7571 ( .B1(n6623), .B2(n6645), .A(n6622), .ZN(U3197) );
  AOI22_X1 U7572 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6663), .ZN(n6624) );
  OAI21_X1 U7573 ( .B1(n6828), .B2(n6645), .A(n6624), .ZN(U3198) );
  AOI22_X1 U7574 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6663), .ZN(n6625) );
  OAI21_X1 U7575 ( .B1(n6626), .B2(n6645), .A(n6625), .ZN(U3199) );
  AOI22_X1 U7576 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6663), .ZN(n6627) );
  OAI21_X1 U7577 ( .B1(n6629), .B2(n6649), .A(n6627), .ZN(U3200) );
  AOI22_X1 U7578 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6663), .ZN(n6628) );
  OAI21_X1 U7579 ( .B1(n6629), .B2(n6645), .A(n6628), .ZN(U3201) );
  INV_X1 U7580 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6793) );
  AOI22_X1 U7581 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6663), .ZN(n6630) );
  OAI21_X1 U7582 ( .B1(n6793), .B2(n6649), .A(n6630), .ZN(U3202) );
  AOI22_X1 U7583 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6663), .ZN(n6631) );
  OAI21_X1 U7584 ( .B1(n6793), .B2(n6645), .A(n6631), .ZN(U3203) );
  AOI22_X1 U7585 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6663), .ZN(n6632) );
  OAI21_X1 U7586 ( .B1(n6633), .B2(n6645), .A(n6632), .ZN(U3204) );
  AOI22_X1 U7587 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6663), .ZN(n6634) );
  OAI21_X1 U7588 ( .B1(n6635), .B2(n6645), .A(n6634), .ZN(U3205) );
  AOI22_X1 U7589 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6663), .ZN(n6636) );
  OAI21_X1 U7590 ( .B1(n6784), .B2(n6649), .A(n6636), .ZN(U3206) );
  INV_X1 U7591 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6821) );
  OAI222_X1 U7592 ( .A1(n6649), .A2(n6638), .B1(n6821), .B2(n6675), .C1(n6784), 
        .C2(n6645), .ZN(U3207) );
  AOI22_X1 U7593 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6663), .ZN(n6637) );
  OAI21_X1 U7594 ( .B1(n6638), .B2(n6645), .A(n6637), .ZN(U3208) );
  INV_X1 U7595 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6640) );
  AOI22_X1 U7596 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6663), .ZN(n6639) );
  OAI21_X1 U7597 ( .B1(n6640), .B2(n6645), .A(n6639), .ZN(U3209) );
  AOI22_X1 U7598 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6663), .ZN(n6641) );
  OAI21_X1 U7599 ( .B1(n6808), .B2(n6645), .A(n6641), .ZN(U3210) );
  INV_X1 U7600 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6713) );
  OAI222_X1 U7601 ( .A1(n6645), .A2(n6642), .B1(n6713), .B2(n6675), .C1(n6646), 
        .C2(n6649), .ZN(U3211) );
  AOI22_X1 U7602 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6643), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6663), .ZN(n6644) );
  OAI21_X1 U7603 ( .B1(n6646), .B2(n6645), .A(n6644), .ZN(U3212) );
  AOI22_X1 U7604 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6647), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6663), .ZN(n6648) );
  OAI21_X1 U7605 ( .B1(n6650), .B2(n6649), .A(n6648), .ZN(U3213) );
  MUX2_X1 U7606 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6675), .Z(U3445) );
  MUX2_X1 U7607 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6675), .Z(U3446) );
  MUX2_X1 U7608 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6675), .Z(U3447) );
  MUX2_X1 U7609 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6675), .Z(U3448) );
  INV_X1 U7610 ( .A(n6653), .ZN(n6651) );
  AOI21_X1 U7611 ( .B1(n6776), .B2(n6652), .A(n6651), .ZN(U3451) );
  OAI21_X1 U7612 ( .B1(n6654), .B2(n6717), .A(n6653), .ZN(U3452) );
  NOR2_X1 U7613 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(n6717), .ZN(n6704) );
  AOI21_X1 U7614 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(n6704), .ZN(n6655) );
  OAI22_X1 U7615 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6656), .B1(
        REIP_REG_1__SCAN_IN), .B2(n6655), .ZN(n6657) );
  INV_X1 U7616 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6790) );
  AOI22_X1 U7617 ( .A1(n6658), .A2(n6657), .B1(n6790), .B2(n6660), .ZN(U3468)
         );
  INV_X1 U7618 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6661) );
  AOI22_X1 U7619 ( .A1(n6661), .A2(n6660), .B1(n4386), .B2(n6659), .ZN(U3469)
         );
  NAND2_X1 U7620 ( .A1(n6663), .A2(W_R_N_REG_SCAN_IN), .ZN(n6662) );
  OAI21_X1 U7621 ( .B1(n6663), .B2(READREQUEST_REG_SCAN_IN), .A(n6662), .ZN(
        U3470) );
  AND2_X1 U7622 ( .A1(n6664), .A2(n4884), .ZN(n6665) );
  NOR4_X1 U7623 ( .A1(n6668), .A2(n6667), .A3(n6666), .A4(n6665), .ZN(n6674)
         );
  OAI211_X1 U7624 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3963), .A(n6669), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6671) );
  AOI21_X1 U7625 ( .B1(n6671), .B2(STATE2_REG_0__SCAN_IN), .A(n6670), .ZN(
        n6673) );
  NAND2_X1 U7626 ( .A1(n6674), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6672) );
  OAI21_X1 U7627 ( .B1(n6674), .B2(n6673), .A(n6672), .ZN(U3472) );
  MUX2_X1 U7628 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6675), .Z(U3473) );
  OAI22_X1 U7629 ( .A1(n6679), .A2(n6678), .B1(n6677), .B2(n6676), .ZN(n6685)
         );
  OAI22_X1 U7630 ( .A1(n6683), .A2(n6682), .B1(n6681), .B2(n6680), .ZN(n6684)
         );
  AOI211_X1 U7631 ( .C1(INSTQUEUE_REG_7__2__SCAN_IN), .C2(n6686), .A(n6685), 
        .B(n6684), .ZN(n6842) );
  NAND4_X1 U7632 ( .A1(EBX_REG_23__SCAN_IN), .A2(ADDRESS_REG_27__SCAN_IN), 
        .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(n6714), .ZN(n6696) );
  NAND4_X1 U7633 ( .A1(EAX_REG_1__SCAN_IN), .A2(D_C_N_REG_SCAN_IN), .A3(
        DATAWIDTH_REG_10__SCAN_IN), .A4(n6734), .ZN(n6695) );
  NOR3_X1 U7634 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(EAX_REG_11__SCAN_IN), .A3(LWORD_REG_5__SCAN_IN), .ZN(n6688) );
  NOR3_X1 U7635 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        BYTEENABLE_REG_3__SCAN_IN), .A3(ADDRESS_REG_2__SCAN_IN), .ZN(n6687) );
  NAND4_X1 U7636 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6688), .A3(
        MEMORYFETCH_REG_SCAN_IN), .A4(n6687), .ZN(n6694) );
  NOR4_X1 U7637 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n4172), .A3(n6775), .A4(
        n6781), .ZN(n6692) );
  NOR4_X1 U7638 ( .A1(EAX_REG_29__SCAN_IN), .A2(EAX_REG_3__SCAN_IN), .A3(
        ADDRESS_REG_23__SCAN_IN), .A4(n5548), .ZN(n6691) );
  NOR4_X1 U7639 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(n6824), .A4(n6828), .ZN(n6690) );
  NOR4_X1 U7640 ( .A1(n6808), .A2(n6805), .A3(n6809), .A4(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6689) );
  NAND4_X1 U7641 ( .A1(n6692), .A2(n6691), .A3(n6690), .A4(n6689), .ZN(n6693)
         );
  NOR4_X1 U7642 ( .A1(n6696), .A2(n6695), .A3(n6694), .A4(n6693), .ZN(n6840)
         );
  INV_X1 U7643 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6699) );
  INV_X1 U7644 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6698) );
  NOR4_X1 U7645 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(
        INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6705) );
  INV_X1 U7646 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6702) );
  NOR4_X1 U7647 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .A3(n6731), .A4(n6811), .ZN(n6700) );
  INV_X1 U7648 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6732) );
  NAND4_X1 U7649 ( .A1(n6825), .A2(n5000), .A3(n6700), .A4(n6732), .ZN(n6701)
         );
  NOR4_X1 U7650 ( .A1(n6702), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .A3(
        INSTQUEUE_REG_0__4__SCAN_IN), .A4(n6701), .ZN(n6703) );
  NAND3_X1 U7651 ( .A1(n6705), .A2(n6704), .A3(n6703), .ZN(n6711) );
  NOR4_X1 U7652 ( .A1(EBX_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), .A3(
        n6757), .A4(n6750), .ZN(n6709) );
  NOR4_X1 U7653 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(LWORD_REG_10__SCAN_IN), 
        .A3(ADDRESS_REG_10__SCAN_IN), .A4(REIP_REG_0__SCAN_IN), .ZN(n6708) );
  NOR4_X1 U7654 ( .A1(DATAI_8_), .A2(BYTEENABLE_REG_2__SCAN_IN), .A3(n6793), 
        .A4(n6791), .ZN(n6707) );
  INV_X1 U7655 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6796) );
  NOR4_X1 U7656 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n6784), .A3(n6796), .A4(
        n6785), .ZN(n6706) );
  NAND4_X1 U7657 ( .A1(n6709), .A2(n6708), .A3(n6707), .A4(n6706), .ZN(n6710)
         );
  NOR2_X1 U7658 ( .A1(n6711), .A2(n6710), .ZN(n6839) );
  AOI22_X1 U7659 ( .A1(n6714), .A2(keyinput12), .B1(keyinput48), .B2(n6713), 
        .ZN(n6712) );
  OAI221_X1 U7660 ( .B1(n6714), .B2(keyinput12), .C1(n6713), .C2(keyinput48), 
        .A(n6712), .ZN(n6726) );
  INV_X1 U7661 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6716) );
  AOI22_X1 U7662 ( .A1(n6717), .A2(keyinput36), .B1(n6716), .B2(keyinput10), 
        .ZN(n6715) );
  OAI221_X1 U7663 ( .B1(n6717), .B2(keyinput36), .C1(n6716), .C2(keyinput10), 
        .A(n6715), .ZN(n6725) );
  AOI22_X1 U7664 ( .A1(n6699), .A2(keyinput3), .B1(keyinput51), .B2(n6719), 
        .ZN(n6718) );
  OAI221_X1 U7665 ( .B1(n6699), .B2(keyinput3), .C1(n6719), .C2(keyinput51), 
        .A(n6718), .ZN(n6724) );
  INV_X1 U7666 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6721) );
  AOI22_X1 U7667 ( .A1(n6722), .A2(keyinput34), .B1(keyinput27), .B2(n6721), 
        .ZN(n6720) );
  OAI221_X1 U7668 ( .B1(n6722), .B2(keyinput34), .C1(n6721), .C2(keyinput27), 
        .A(n6720), .ZN(n6723) );
  NOR4_X1 U7669 ( .A1(n6726), .A2(n6725), .A3(n6724), .A4(n6723), .ZN(n6773)
         );
  AOI22_X1 U7670 ( .A1(n6729), .A2(keyinput60), .B1(keyinput41), .B2(n6728), 
        .ZN(n6727) );
  OAI221_X1 U7671 ( .B1(n6729), .B2(keyinput60), .C1(n6728), .C2(keyinput41), 
        .A(n6727), .ZN(n6740) );
  AOI22_X1 U7672 ( .A1(n6732), .A2(keyinput63), .B1(keyinput19), .B2(n6731), 
        .ZN(n6730) );
  OAI221_X1 U7673 ( .B1(n6732), .B2(keyinput63), .C1(n6731), .C2(keyinput19), 
        .A(n6730), .ZN(n6739) );
  AOI22_X1 U7674 ( .A1(n6734), .A2(keyinput28), .B1(n5000), .B2(keyinput9), 
        .ZN(n6733) );
  OAI221_X1 U7675 ( .B1(n6734), .B2(keyinput28), .C1(n5000), .C2(keyinput9), 
        .A(n6733), .ZN(n6738) );
  AOI22_X1 U7676 ( .A1(n6702), .A2(keyinput49), .B1(keyinput32), .B2(n6736), 
        .ZN(n6735) );
  OAI221_X1 U7677 ( .B1(n6702), .B2(keyinput49), .C1(n6736), .C2(keyinput32), 
        .A(n6735), .ZN(n6737) );
  NOR4_X1 U7678 ( .A1(n6740), .A2(n6739), .A3(n6738), .A4(n6737), .ZN(n6772)
         );
  AOI22_X1 U7679 ( .A1(n6743), .A2(keyinput11), .B1(n6742), .B2(keyinput38), 
        .ZN(n6741) );
  OAI221_X1 U7680 ( .B1(n6743), .B2(keyinput11), .C1(n6742), .C2(keyinput38), 
        .A(n6741), .ZN(n6755) );
  AOI22_X1 U7681 ( .A1(n4355), .A2(keyinput50), .B1(n6745), .B2(keyinput21), 
        .ZN(n6744) );
  OAI221_X1 U7682 ( .B1(n4355), .B2(keyinput50), .C1(n6745), .C2(keyinput21), 
        .A(n6744), .ZN(n6754) );
  AOI22_X1 U7683 ( .A1(n6748), .A2(keyinput52), .B1(keyinput45), .B2(n6747), 
        .ZN(n6746) );
  OAI221_X1 U7684 ( .B1(n6748), .B2(keyinput52), .C1(n6747), .C2(keyinput45), 
        .A(n6746), .ZN(n6753) );
  AOI22_X1 U7685 ( .A1(n6751), .A2(keyinput46), .B1(n6750), .B2(keyinput0), 
        .ZN(n6749) );
  OAI221_X1 U7686 ( .B1(n6751), .B2(keyinput46), .C1(n6750), .C2(keyinput0), 
        .A(n6749), .ZN(n6752) );
  NOR4_X1 U7687 ( .A1(n6755), .A2(n6754), .A3(n6753), .A4(n6752), .ZN(n6771)
         );
  AOI22_X1 U7688 ( .A1(n6758), .A2(keyinput40), .B1(keyinput53), .B2(n6757), 
        .ZN(n6756) );
  OAI221_X1 U7689 ( .B1(n6758), .B2(keyinput40), .C1(n6757), .C2(keyinput53), 
        .A(n6756), .ZN(n6769) );
  AOI22_X1 U7690 ( .A1(n6761), .A2(keyinput39), .B1(keyinput56), .B2(n6760), 
        .ZN(n6759) );
  OAI221_X1 U7691 ( .B1(n6761), .B2(keyinput39), .C1(n6760), .C2(keyinput56), 
        .A(n6759), .ZN(n6768) );
  AOI22_X1 U7692 ( .A1(n6764), .A2(keyinput14), .B1(keyinput24), .B2(n6763), 
        .ZN(n6762) );
  OAI221_X1 U7693 ( .B1(n6764), .B2(keyinput14), .C1(n6763), .C2(keyinput24), 
        .A(n6762), .ZN(n6767) );
  AOI22_X1 U7694 ( .A1(n6697), .A2(keyinput26), .B1(keyinput7), .B2(n4386), 
        .ZN(n6765) );
  OAI221_X1 U7695 ( .B1(n6697), .B2(keyinput26), .C1(n4386), .C2(keyinput7), 
        .A(n6765), .ZN(n6766) );
  NOR4_X1 U7696 ( .A1(n6769), .A2(n6768), .A3(n6767), .A4(n6766), .ZN(n6770)
         );
  NAND4_X1 U7697 ( .A1(n6773), .A2(n6772), .A3(n6771), .A4(n6770), .ZN(n6838)
         );
  AOI22_X1 U7698 ( .A1(n4172), .A2(keyinput33), .B1(n6775), .B2(keyinput4), 
        .ZN(n6774) );
  OAI221_X1 U7699 ( .B1(n4172), .B2(keyinput33), .C1(n6775), .C2(keyinput4), 
        .A(n6774), .ZN(n6779) );
  XNOR2_X1 U7700 ( .A(n6776), .B(keyinput25), .ZN(n6778) );
  XOR2_X1 U7701 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .B(keyinput1), .Z(n6777) );
  OR3_X1 U7702 ( .A1(n6779), .A2(n6778), .A3(n6777), .ZN(n6788) );
  AOI22_X1 U7703 ( .A1(n6782), .A2(keyinput31), .B1(n6781), .B2(keyinput8), 
        .ZN(n6780) );
  OAI221_X1 U7704 ( .B1(n6782), .B2(keyinput31), .C1(n6781), .C2(keyinput8), 
        .A(n6780), .ZN(n6787) );
  AOI22_X1 U7705 ( .A1(n6785), .A2(keyinput6), .B1(n6784), .B2(keyinput29), 
        .ZN(n6783) );
  OAI221_X1 U7706 ( .B1(n6785), .B2(keyinput6), .C1(n6784), .C2(keyinput29), 
        .A(n6783), .ZN(n6786) );
  NOR3_X1 U7707 ( .A1(n6788), .A2(n6787), .A3(n6786), .ZN(n6836) );
  AOI22_X1 U7708 ( .A1(n6791), .A2(keyinput57), .B1(keyinput54), .B2(n6790), 
        .ZN(n6789) );
  OAI221_X1 U7709 ( .B1(n6791), .B2(keyinput57), .C1(n6790), .C2(keyinput54), 
        .A(n6789), .ZN(n6803) );
  AOI22_X1 U7710 ( .A1(n6794), .A2(keyinput59), .B1(n6793), .B2(keyinput23), 
        .ZN(n6792) );
  OAI221_X1 U7711 ( .B1(n6794), .B2(keyinput59), .C1(n6793), .C2(keyinput23), 
        .A(n6792), .ZN(n6802) );
  AOI22_X1 U7712 ( .A1(n6797), .A2(keyinput20), .B1(n6796), .B2(keyinput42), 
        .ZN(n6795) );
  OAI221_X1 U7713 ( .B1(n6797), .B2(keyinput20), .C1(n6796), .C2(keyinput42), 
        .A(n6795), .ZN(n6801) );
  XNOR2_X1 U7714 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .B(keyinput44), .ZN(n6799)
         );
  XNOR2_X1 U7715 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .B(keyinput18), .ZN(n6798) );
  NAND2_X1 U7716 ( .A1(n6799), .A2(n6798), .ZN(n6800) );
  NOR4_X1 U7717 ( .A1(n6803), .A2(n6802), .A3(n6801), .A4(n6800), .ZN(n6835)
         );
  AOI22_X1 U7718 ( .A1(n6806), .A2(keyinput30), .B1(keyinput13), .B2(n6805), 
        .ZN(n6804) );
  OAI221_X1 U7719 ( .B1(n6806), .B2(keyinput30), .C1(n6805), .C2(keyinput13), 
        .A(n6804), .ZN(n6818) );
  AOI22_X1 U7720 ( .A1(n6809), .A2(keyinput2), .B1(n6808), .B2(keyinput55), 
        .ZN(n6807) );
  OAI221_X1 U7721 ( .B1(n6809), .B2(keyinput2), .C1(n6808), .C2(keyinput55), 
        .A(n6807), .ZN(n6817) );
  AOI22_X1 U7722 ( .A1(n6812), .A2(keyinput35), .B1(n6811), .B2(keyinput15), 
        .ZN(n6810) );
  OAI221_X1 U7723 ( .B1(n6812), .B2(keyinput35), .C1(n6811), .C2(keyinput15), 
        .A(n6810), .ZN(n6816) );
  XOR2_X1 U7724 ( .A(n6698), .B(keyinput5), .Z(n6814) );
  XNOR2_X1 U7725 ( .A(STATE2_REG_3__SCAN_IN), .B(keyinput43), .ZN(n6813) );
  NAND2_X1 U7726 ( .A1(n6814), .A2(n6813), .ZN(n6815) );
  NOR4_X1 U7727 ( .A1(n6818), .A2(n6817), .A3(n6816), .A4(n6815), .ZN(n6834)
         );
  AOI22_X1 U7728 ( .A1(n5548), .A2(keyinput47), .B1(keyinput37), .B2(n3906), 
        .ZN(n6819) );
  OAI221_X1 U7729 ( .B1(n5548), .B2(keyinput47), .C1(n3906), .C2(keyinput37), 
        .A(n6819), .ZN(n6832) );
  AOI22_X1 U7730 ( .A1(n6822), .A2(keyinput58), .B1(keyinput62), .B2(n6821), 
        .ZN(n6820) );
  OAI221_X1 U7731 ( .B1(n6822), .B2(keyinput58), .C1(n6821), .C2(keyinput62), 
        .A(n6820), .ZN(n6831) );
  AOI22_X1 U7732 ( .A1(n6825), .A2(keyinput61), .B1(keyinput22), .B2(n6824), 
        .ZN(n6823) );
  OAI221_X1 U7733 ( .B1(n6825), .B2(keyinput61), .C1(n6824), .C2(keyinput22), 
        .A(n6823), .ZN(n6830) );
  AOI22_X1 U7734 ( .A1(n6828), .A2(keyinput16), .B1(n6827), .B2(keyinput17), 
        .ZN(n6826) );
  OAI221_X1 U7735 ( .B1(n6828), .B2(keyinput16), .C1(n6827), .C2(keyinput17), 
        .A(n6826), .ZN(n6829) );
  NOR4_X1 U7736 ( .A1(n6832), .A2(n6831), .A3(n6830), .A4(n6829), .ZN(n6833)
         );
  NAND4_X1 U7737 ( .A1(n6836), .A2(n6835), .A3(n6834), .A4(n6833), .ZN(n6837)
         );
  AOI211_X1 U7738 ( .C1(n6840), .C2(n6839), .A(n6838), .B(n6837), .ZN(n6841)
         );
  XNOR2_X1 U7739 ( .A(n6842), .B(n6841), .ZN(U3078) );
  CLKBUF_X1 U3653 ( .A(n3348), .Z(n3304) );
  CLKBUF_X1 U4310 ( .A(n3947), .Z(n5043) );
endmodule

