

module b15_C_AntiSAT_k_128_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736;

  OR2_X1 U34450 ( .A1(n3574), .A2(n3573), .ZN(n5743) );
  CLKBUF_X2 U34470 ( .A(n4477), .Z(n3033) );
  NAND2_X2 U34480 ( .A1(n4115), .A2(n3208), .ZN(n4163) );
  CLKBUF_X2 U3449 ( .A(n3168), .Z(n4038) );
  CLKBUF_X1 U3450 ( .A(n3159), .Z(n4013) );
  CLKBUF_X1 U34510 ( .A(n3241), .Z(n3938) );
  CLKBUF_X2 U34520 ( .A(n3198), .Z(n4060) );
  AND2_X1 U34530 ( .A1(n3279), .A2(n3231), .ZN(n3277) );
  AND2_X1 U3454 ( .A1(n3103), .A2(n4386), .ZN(n3242) );
  NOR2_X1 U34550 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3101) );
  AOI21_X1 U34560 ( .B1(n5018), .B2(n5231), .A(n5232), .ZN(n5069) );
  OR2_X1 U3458 ( .A1(n3223), .A2(n4116), .ZN(n4250) );
  INV_X2 U34590 ( .A(n5691), .ZN(n5467) );
  INV_X1 U34600 ( .A(n4328), .ZN(n5100) );
  NAND2_X1 U34610 ( .A1(n3900), .A2(n3899), .ZN(n4094) );
  OR2_X1 U34620 ( .A1(n3747), .A2(n4935), .ZN(n5231) );
  AND2_X1 U34630 ( .A1(n5454), .A2(n5455), .ZN(n5695) );
  NAND2_X1 U34640 ( .A1(n4898), .A2(n4936), .ZN(n4935) );
  INV_X1 U34650 ( .A(n5499), .ZN(n5941) );
  AOI211_X1 U3466 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5121), .A(n5112), .B(n5111), .ZN(n5113) );
  XOR2_X1 U3467 ( .A(n5107), .B(n5106), .Z(n5505) );
  NOR2_X2 U34680 ( .A1(n4445), .A2(n4131), .ZN(n4449) );
  NAND2_X2 U34690 ( .A1(n5430), .A2(n5429), .ZN(n5428) );
  AOI21_X2 U34700 ( .B1(n5434), .B2(n4088), .A(n3082), .ZN(n5430) );
  NAND2_X2 U34710 ( .A1(n3203), .A2(n3090), .ZN(n3224) );
  INV_X2 U34720 ( .A(n3205), .ZN(n3230) );
  AND2_X4 U34730 ( .A1(n3102), .A2(n4536), .ZN(n3241) );
  OAI21_X2 U34740 ( .B1(n5142), .B2(n5143), .A(n5125), .ZN(n5376) );
  INV_X2 U3475 ( .A(n5776), .ZN(n5848) );
  INV_X2 U3476 ( .A(n5691), .ZN(n5436) );
  CLKBUF_X1 U3477 ( .A(n4479), .Z(n3031) );
  CLKBUF_X1 U3478 ( .A(n3606), .Z(n3029) );
  AND3_X1 U3479 ( .A1(n3229), .A2(n3207), .A3(n3280), .ZN(n3218) );
  OR2_X1 U3480 ( .A1(n3210), .A2(n4115), .ZN(n3229) );
  INV_X1 U3481 ( .A(n3231), .ZN(n4115) );
  OR2_X2 U3482 ( .A1(n3117), .A2(n3116), .ZN(n3191) );
  AND4_X1 U3483 ( .A1(n3125), .A2(n3124), .A3(n3123), .A4(n3122), .ZN(n3136)
         );
  CLKBUF_X2 U3484 ( .A(n3181), .Z(n4043) );
  BUF_X2 U3485 ( .A(n3030), .Z(n4000) );
  BUF_X2 U3486 ( .A(n3166), .Z(n3027) );
  AND2_X2 U3487 ( .A1(n3100), .A2(n3103), .ZN(n3165) );
  AND2_X2 U3488 ( .A1(n3100), .A2(n3101), .ZN(n3167) );
  AND2_X2 U3489 ( .A1(n3103), .A2(n3102), .ZN(n3159) );
  AND2_X2 U3490 ( .A1(n3101), .A2(n3102), .ZN(n3166) );
  INV_X2 U3491 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3095) );
  OR2_X1 U3492 ( .A1(n3469), .A2(n3468), .ZN(n3485) );
  NAND2_X1 U3493 ( .A1(n3271), .A2(n3270), .ZN(n3314) );
  CLKBUF_X1 U3494 ( .A(n4241), .Z(n3013) );
  OR2_X1 U3495 ( .A1(n3532), .A2(n3210), .ZN(n3086) );
  INV_X2 U3496 ( .A(n3224), .ZN(n3279) );
  INV_X2 U3497 ( .A(n3220), .ZN(n3189) );
  NAND2_X2 U3498 ( .A1(n3148), .A2(n3147), .ZN(n3209) );
  INV_X2 U3499 ( .A(n3208), .ZN(n2998) );
  CLKBUF_X2 U3500 ( .A(n3167), .Z(n4037) );
  BUF_X2 U3501 ( .A(n3164), .Z(n3932) );
  CLKBUF_X2 U3502 ( .A(n3182), .Z(n4018) );
  BUF_X2 U3503 ( .A(n3247), .Z(n4036) );
  CLKBUF_X2 U3504 ( .A(n3380), .Z(n3401) );
  BUF_X2 U3505 ( .A(n3169), .Z(n3901) );
  AND2_X1 U3506 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4536) );
  NOR2_X1 U3507 ( .A1(n3521), .A2(n3520), .ZN(n3522) );
  AOI21_X1 U3508 ( .B1(n5520), .B2(n5375), .A(n5374), .ZN(n5527) );
  AOI21_X1 U3509 ( .B1(n4091), .B2(n5421), .A(n4090), .ZN(n4092) );
  NAND2_X1 U3510 ( .A1(n5393), .A2(n3513), .ZN(n5371) );
  AND2_X1 U3511 ( .A1(n5383), .A2(n5500), .ZN(n3520) );
  AND2_X1 U3512 ( .A1(n5369), .A2(n3518), .ZN(n5383) );
  OAI21_X1 U3513 ( .B1(n3070), .B2(n5279), .A(n3035), .ZN(n5654) );
  AND2_X1 U3514 ( .A1(n5016), .A2(n3059), .ZN(n3058) );
  NAND3_X1 U3515 ( .A1(n4553), .A2(n4552), .A3(n4459), .ZN(n4462) );
  NAND2_X2 U3516 ( .A1(n5858), .A2(n4827), .ZN(n5785) );
  AND3_X2 U3517 ( .A1(n4457), .A2(n4441), .A3(n4447), .ZN(n4553) );
  XNOR2_X1 U3518 ( .A(n3485), .B(n3472), .ZN(n3648) );
  AND2_X2 U3519 ( .A1(n3485), .A2(n3484), .ZN(n5691) );
  NAND2_X1 U3520 ( .A1(n3597), .A2(n3596), .ZN(n4457) );
  XNOR2_X1 U3521 ( .A(n3469), .B(n3458), .ZN(n3635) );
  NOR2_X2 U3522 ( .A1(n6181), .A2(n6227), .ZN(n5004) );
  OR2_X1 U3523 ( .A1(n3617), .A2(n3616), .ZN(n4443) );
  INV_X1 U3524 ( .A(n3590), .ZN(n4638) );
  AND2_X1 U3525 ( .A1(n4325), .A2(n4324), .ZN(n3616) );
  AOI21_X1 U3526 ( .B1(n4432), .B2(n4433), .A(n3362), .ZN(n5938) );
  NAND2_X1 U3527 ( .A1(n3604), .A2(n3603), .ZN(n4325) );
  NAND2_X1 U3528 ( .A1(n3360), .A2(n3359), .ZN(n4432) );
  XNOR2_X1 U3529 ( .A(n3422), .B(n3085), .ZN(n3620) );
  AND2_X1 U3530 ( .A1(n5221), .A2(n3017), .ZN(n5294) );
  OR2_X1 U3531 ( .A1(n3393), .A2(n4637), .ZN(n3422) );
  NOR2_X1 U3532 ( .A1(n5078), .A2(n5780), .ZN(n5225) );
  BUF_X1 U3533 ( .A(n3598), .Z(n4476) );
  XNOR2_X1 U3535 ( .A(n3368), .B(n3337), .ZN(n3598) );
  NAND2_X2 U3536 ( .A1(n5357), .A2(n4573), .ZN(n5361) );
  NAND2_X1 U3537 ( .A1(n4159), .A2(n4158), .ZN(n5237) );
  NOR2_X1 U3538 ( .A1(n4750), .A2(n5313), .ZN(n6360) );
  NOR2_X1 U3539 ( .A1(n4750), .A2(n3230), .ZN(n6352) );
  NOR2_X1 U3540 ( .A1(n4750), .A2(n3176), .ZN(n6346) );
  NOR2_X1 U3541 ( .A1(n4750), .A2(n3206), .ZN(n6340) );
  NOR2_X1 U3542 ( .A1(n4750), .A2(n4115), .ZN(n6334) );
  NOR2_X1 U3543 ( .A1(n4750), .A2(n3279), .ZN(n6328) );
  NOR2_X1 U3544 ( .A1(n4750), .A2(n3189), .ZN(n6322) );
  NOR2_X1 U3545 ( .A1(n4750), .A2(n2998), .ZN(n6307) );
  AOI21_X1 U3546 ( .B1(n4479), .B2(n6414), .A(n3392), .ZN(n4637) );
  NAND2_X1 U3547 ( .A1(n6526), .A2(n4844), .ZN(n5833) );
  NOR2_X2 U3548 ( .A1(n5743), .A2(n6418), .ZN(n4409) );
  AND2_X1 U3549 ( .A1(n3015), .A2(n3016), .ZN(n4836) );
  OAI22_X1 U3550 ( .A1(n4480), .A2(STATE2_REG_0__SCAN_IN), .B1(n3395), .B2(
        n3379), .ZN(n3336) );
  NOR2_X1 U3551 ( .A1(n4561), .A2(n4559), .ZN(n3015) );
  NAND2_X1 U3552 ( .A1(n3341), .A2(n3345), .ZN(n4970) );
  NAND2_X1 U3553 ( .A1(n4378), .A2(n6414), .ZN(n3303) );
  INV_X1 U3554 ( .A(n3314), .ZN(n3291) );
  NOR2_X1 U3555 ( .A1(n3227), .A2(n4254), .ZN(n3238) );
  OAI21_X1 U3556 ( .B1(n3204), .B2(n3578), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3212) );
  INV_X1 U3557 ( .A(n4835), .ZN(n2999) );
  NOR2_X1 U3558 ( .A1(n3265), .A2(n6414), .ZN(n3481) );
  AND2_X1 U3559 ( .A1(n3138), .A2(n4107), .ZN(n3190) );
  INV_X1 U3560 ( .A(n3532), .ZN(n3560) );
  NAND2_X1 U3561 ( .A1(n3379), .A2(n3378), .ZN(n3569) );
  INV_X1 U3562 ( .A(n4246), .ZN(n5745) );
  INV_X1 U3563 ( .A(n4107), .ZN(n4882) );
  INV_X1 U3564 ( .A(n4251), .ZN(n5296) );
  NAND2_X1 U3565 ( .A1(n4328), .A2(n4251), .ZN(n4197) );
  NAND2_X1 U3566 ( .A1(n2998), .A2(n3189), .ZN(n4246) );
  AND2_X2 U3567 ( .A1(n4831), .A2(n3208), .ZN(n4328) );
  NAND2_X1 U3568 ( .A1(n3253), .A2(n3094), .ZN(n3487) );
  BUF_X4 U3569 ( .A(n4116), .Z(n4251) );
  OR2_X1 U3570 ( .A1(n3208), .A2(n6414), .ZN(n3378) );
  NAND2_X2 U3571 ( .A1(n3231), .A2(n3220), .ZN(n4116) );
  OR2_X1 U3572 ( .A1(n3263), .A2(n3262), .ZN(n3355) );
  INV_X2 U3573 ( .A(n3209), .ZN(n3206) );
  NOR2_X1 U3574 ( .A1(n5499), .A2(n4744), .ZN(n6355) );
  NOR2_X1 U3575 ( .A1(n5499), .A2(n4488), .ZN(n6348) );
  OR2_X2 U3576 ( .A1(n3175), .A2(n3174), .ZN(n3205) );
  AND4_X1 U3577 ( .A1(n3099), .A2(n3098), .A3(n3097), .A4(n3096), .ZN(n3037)
         );
  AND4_X1 U3578 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n3148)
         );
  AND4_X1 U3579 ( .A1(n3197), .A2(n3196), .A3(n3195), .A4(n3194), .ZN(n3203)
         );
  AND4_X1 U3580 ( .A1(n3121), .A2(n3120), .A3(n3119), .A4(n3118), .ZN(n3137)
         );
  AOI22_X1 U3581 ( .A1(n3247), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3140) );
  AND4_X1 U3582 ( .A1(n3146), .A2(n3145), .A3(n3144), .A4(n3143), .ZN(n3147)
         );
  AND4_X1 U3583 ( .A1(n3129), .A2(n3128), .A3(n3127), .A4(n3126), .ZN(n3135)
         );
  AND4_X1 U3584 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n3134)
         );
  BUF_X4 U3585 ( .A(n3165), .Z(n4019) );
  OR2_X2 U3586 ( .A1(n6425), .A2(n6305), .ZN(n5499) );
  BUF_X2 U3587 ( .A(n3406), .Z(n3937) );
  BUF_X2 U3588 ( .A(n3165), .Z(n3028) );
  AND2_X1 U3589 ( .A1(n3100), .A2(n4536), .ZN(n3164) );
  AND2_X2 U3590 ( .A1(n4515), .A2(n3100), .ZN(n3030) );
  AND2_X2 U3591 ( .A1(n4515), .A2(n4386), .ZN(n3380) );
  CLKBUF_X1 U3592 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n6645) );
  NAND2_X1 U3593 ( .A1(n3501), .A2(n3003), .ZN(n3000) );
  AND2_X2 U3594 ( .A1(n3000), .A2(n3001), .ZN(n5441) );
  OR2_X1 U3595 ( .A1(n3002), .A2(n3041), .ZN(n3001) );
  INV_X1 U3596 ( .A(n3506), .ZN(n3002) );
  AND2_X1 U3597 ( .A1(n3500), .A2(n3506), .ZN(n3003) );
  NAND2_X1 U3598 ( .A1(n3303), .A2(n3302), .ZN(n3004) );
  NAND3_X1 U3600 ( .A1(n3212), .A2(n3211), .A3(n3086), .ZN(n3318) );
  OAI21_X2 U3601 ( .B1(n3590), .B2(n3482), .A(n3398), .ZN(n3399) );
  AOI21_X1 U3602 ( .B1(n5018), .B2(n5231), .A(n5232), .ZN(n3006) );
  AOI21_X1 U3603 ( .B1(n5018), .B2(n5231), .A(n5232), .ZN(n3007) );
  AND2_X2 U3604 ( .A1(n5260), .A2(n3008), .ZN(n5141) );
  AND2_X1 U3605 ( .A1(n5261), .A2(n3009), .ZN(n3008) );
  INV_X1 U3606 ( .A(n5156), .ZN(n3009) );
  NAND2_X1 U3607 ( .A1(n3011), .A2(n5921), .ZN(n3010) );
  CLKBUF_X1 U3608 ( .A(n5919), .Z(n3011) );
  AND2_X1 U3609 ( .A1(n3286), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3012) );
  CLKBUF_X1 U3610 ( .A(n5476), .Z(n3014) );
  NAND2_X1 U3611 ( .A1(n4102), .A2(n5745), .ZN(n4241) );
  AND2_X1 U3612 ( .A1(n2999), .A2(n4656), .ZN(n3016) );
  AND2_X1 U3613 ( .A1(n4172), .A2(n3018), .ZN(n3017) );
  INV_X1 U3614 ( .A(n5181), .ZN(n3018) );
  AND2_X1 U3615 ( .A1(n5289), .A2(n4189), .ZN(n5276) );
  CLKBUF_X1 U3616 ( .A(n5910), .Z(n3019) );
  BUF_X1 U3617 ( .A(n3316), .Z(n3020) );
  NAND3_X1 U3618 ( .A1(n3216), .A2(n3280), .A3(n3206), .ZN(n3021) );
  NAND3_X1 U3619 ( .A1(n3216), .A2(n3280), .A3(n3206), .ZN(n3022) );
  OR2_X2 U3620 ( .A1(n3188), .A2(n3187), .ZN(n3280) );
  AND2_X1 U3621 ( .A1(n3100), .A2(n4536), .ZN(n3023) );
  NOR2_X2 U3622 ( .A1(n3278), .A2(n4103), .ZN(n4232) );
  AND2_X2 U3623 ( .A1(n3095), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3100)
         );
  AOI21_X1 U3624 ( .B1(n3005), .B2(n6645), .A(n3322), .ZN(n3370) );
  AND2_X1 U3625 ( .A1(n4515), .A2(n4386), .ZN(n3024) );
  AND2_X1 U3626 ( .A1(n4515), .A2(n4386), .ZN(n3025) );
  AND2_X1 U3627 ( .A1(n3103), .A2(n3102), .ZN(n3026) );
  AND2_X1 U3628 ( .A1(n3366), .A2(n3365), .ZN(n5928) );
  OR2_X2 U3629 ( .A1(n3158), .A2(n3157), .ZN(n3231) );
  AND2_X2 U3630 ( .A1(n3230), .A2(n3191), .ZN(n3210) );
  NAND2_X2 U3631 ( .A1(n3205), .A2(n3176), .ZN(n3216) );
  NAND2_X2 U3632 ( .A1(n3316), .A2(n3290), .ZN(n3313) );
  NAND2_X2 U3633 ( .A1(n3037), .A2(n3091), .ZN(n3220) );
  AND2_X4 U3634 ( .A1(n3102), .A2(n4515), .ZN(n3182) );
  NAND2_X2 U3635 ( .A1(n4923), .A2(n4922), .ZN(n4958) );
  NAND2_X2 U3636 ( .A1(n3494), .A2(n3493), .ZN(n4923) );
  NAND2_X2 U3637 ( .A1(n3619), .A2(n3618), .ZN(n4441) );
  NAND2_X1 U3638 ( .A1(n3206), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3379) );
  INV_X2 U3639 ( .A(n3191), .ZN(n3176) );
  AND2_X2 U3640 ( .A1(n3218), .A2(n3217), .ZN(n4102) );
  OAI21_X2 U3641 ( .B1(n5484), .B2(n5486), .A(n5485), .ZN(n5476) );
  OAI21_X2 U3642 ( .B1(n5051), .B2(n3057), .A(n3055), .ZN(n5484) );
  AND2_X2 U3643 ( .A1(n4854), .A2(n4900), .ZN(n4898) );
  NOR2_X2 U3644 ( .A1(n4555), .A2(n3077), .ZN(n4854) );
  OAI21_X4 U3645 ( .B1(n4958), .B2(n3498), .A(n3497), .ZN(n5051) );
  NOR2_X2 U3646 ( .A1(n4094), .A2(n3067), .ZN(n5260) );
  XNOR2_X1 U3647 ( .A(n3271), .B(n3240), .ZN(n3606) );
  AND2_X2 U3648 ( .A1(n5141), .A2(n3073), .ZN(n5126) );
  AND2_X2 U3649 ( .A1(n4391), .A2(n3103), .ZN(n3168) );
  XNOR2_X2 U3650 ( .A(n3291), .B(n3313), .ZN(n4378) );
  NAND2_X2 U3651 ( .A1(n3746), .A2(n3745), .ZN(n5018) );
  XNOR2_X1 U3652 ( .A(n3306), .B(n3354), .ZN(n4477) );
  AND2_X1 U3653 ( .A1(n4515), .A2(n4391), .ZN(n3034) );
  AND2_X1 U3654 ( .A1(n4515), .A2(n4391), .ZN(n3247) );
  AND2_X1 U3655 ( .A1(n3512), .A2(n5519), .ZN(n3513) );
  NAND2_X1 U3656 ( .A1(n5166), .A2(n3070), .ZN(n3069) );
  INV_X1 U3657 ( .A(n5280), .ZN(n3899) );
  NOR2_X1 U3658 ( .A1(n4385), .A2(n6414), .ZN(n4071) );
  INV_X1 U3659 ( .A(n5442), .ZN(n4087) );
  CLKBUF_X1 U3660 ( .A(n4237), .Z(n4238) );
  INV_X2 U3661 ( .A(n3792), .ZN(n4082) );
  AOI21_X1 U3662 ( .B1(n3047), .B2(n3050), .A(n3045), .ZN(n3044) );
  NAND2_X1 U3663 ( .A1(n5441), .A2(n3047), .ZN(n3046) );
  INV_X1 U3664 ( .A(n5400), .ZN(n3045) );
  AOI21_X1 U3665 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6414), .A(n3564), 
        .ZN(n3572) );
  NAND2_X1 U3666 ( .A1(n4232), .A2(n3092), .ZN(n6407) );
  AND2_X1 U3667 ( .A1(n4246), .A2(n3531), .ZN(n3552) );
  AND2_X1 U3668 ( .A1(n3208), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3538) );
  AND2_X1 U3669 ( .A1(n3457), .A2(n3456), .ZN(n3468) );
  OR2_X1 U3670 ( .A1(n3301), .A2(n3300), .ZN(n3356) );
  NAND2_X1 U3671 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4538), .ZN(n3567) );
  OR2_X1 U3672 ( .A1(n3566), .A2(n3567), .ZN(n4228) );
  NAND2_X1 U3673 ( .A1(n3538), .A2(n3209), .ZN(n3532) );
  AND2_X1 U3674 ( .A1(n3216), .A2(n3280), .ZN(n3192) );
  NAND2_X1 U3675 ( .A1(n2998), .A2(n3220), .ZN(n4107) );
  NOR2_X1 U3676 ( .A1(n5127), .A2(n3074), .ZN(n3073) );
  INV_X1 U3677 ( .A(n5143), .ZN(n3074) );
  NOR2_X1 U3678 ( .A1(n3042), .A2(n3064), .ZN(n3063) );
  INV_X1 U3679 ( .A(n5291), .ZN(n3064) );
  NAND2_X1 U3680 ( .A1(n3079), .A2(n4769), .ZN(n3078) );
  INV_X1 U3681 ( .A(n4655), .ZN(n3079) );
  NOR2_X2 U3682 ( .A1(n3205), .A2(n6303), .ZN(n3827) );
  AND2_X1 U3683 ( .A1(n4153), .A2(n4152), .ZN(n4902) );
  AND2_X1 U3684 ( .A1(n3191), .A2(n4831), .ZN(n3523) );
  INV_X1 U3685 ( .A(n3523), .ZN(n3482) );
  INV_X1 U3686 ( .A(n3356), .ZN(n3310) );
  OR2_X1 U3687 ( .A1(n3576), .A2(n3575), .ZN(n4385) );
  AND4_X1 U3688 ( .A1(n3230), .A2(n2998), .A3(n3209), .A4(n3280), .ZN(n3232)
         );
  INV_X1 U3689 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U3690 ( .A1(n3377), .A2(n3376), .ZN(n6059) );
  AND2_X1 U3691 ( .A1(n4238), .A2(n6528), .ZN(n4298) );
  AND2_X1 U3692 ( .A1(n6303), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4081) );
  INV_X1 U3693 ( .A(n3073), .ZN(n3072) );
  NAND2_X1 U3694 ( .A1(n4031), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4076)
         );
  NAND2_X1 U3695 ( .A1(n3068), .A2(n5266), .ZN(n3067) );
  INV_X1 U3696 ( .A(n3069), .ZN(n3068) );
  OR2_X1 U3697 ( .A1(n5672), .A2(n4074), .ZN(n3881) );
  AOI21_X1 U3698 ( .B1(n3058), .B2(n3056), .A(n3036), .ZN(n3055) );
  INV_X1 U3699 ( .A(n3058), .ZN(n3057) );
  XNOR2_X1 U3700 ( .A(n5436), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5400)
         );
  AOI21_X1 U3701 ( .B1(n3040), .B2(n5436), .A(n3048), .ZN(n3047) );
  NOR2_X1 U3702 ( .A1(n5444), .A2(n3049), .ZN(n3048) );
  INV_X1 U3703 ( .A(n3087), .ZN(n3049) );
  NOR2_X1 U3704 ( .A1(n5436), .A2(n3087), .ZN(n3050) );
  NAND2_X1 U3705 ( .A1(n5467), .A2(n5435), .ZN(n4088) );
  OR2_X1 U3706 ( .A1(n5436), .A2(n3505), .ZN(n3506) );
  OR2_X1 U3707 ( .A1(n5726), .A2(n5719), .ZN(n5586) );
  NAND2_X1 U3708 ( .A1(n4277), .A2(n6396), .ZN(n5721) );
  OR2_X1 U3709 ( .A1(n5586), .A2(n6016), .ZN(n4605) );
  OR2_X1 U3710 ( .A1(n5726), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4434)
         );
  INV_X1 U3711 ( .A(n3270), .ZN(n3240) );
  AND2_X1 U3712 ( .A1(n4580), .A2(n6028), .ZN(n6026) );
  NAND2_X1 U3713 ( .A1(n4476), .A2(n4637), .ZN(n6119) );
  NOR2_X1 U3714 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4475), .ZN(n4743) );
  INV_X1 U3715 ( .A(n6314), .ZN(n6222) );
  INV_X1 U3716 ( .A(n4970), .ZN(n6260) );
  INV_X2 U3717 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6303) );
  NOR2_X1 U3718 ( .A1(n5118), .A2(n5309), .ZN(n4211) );
  NAND2_X1 U3719 ( .A1(n4113), .A2(n4566), .ZN(n5305) );
  INV_X1 U3720 ( .A(n5305), .ZN(n5311) );
  AND2_X1 U3721 ( .A1(n5357), .A2(n3281), .ZN(n5353) );
  INV_X1 U3722 ( .A(n5357), .ZN(n5352) );
  AND2_X1 U3723 ( .A1(n4411), .A2(n4838), .ZN(n5871) );
  INV_X1 U3724 ( .A(n5908), .ZN(n5902) );
  XNOR2_X1 U3725 ( .A(n5126), .B(n3076), .ZN(n5115) );
  XNOR2_X1 U3726 ( .A(n4216), .B(n3514), .ZN(n5089) );
  OAI21_X1 U3727 ( .B1(n4215), .B2(n3515), .A(n4214), .ZN(n4216) );
  INV_X1 U3728 ( .A(n5362), .ZN(n4215) );
  AND2_X1 U3729 ( .A1(n4277), .A2(n4245), .ZN(n6021) );
  AND2_X1 U3730 ( .A1(n4277), .A2(n4249), .ZN(n6010) );
  INV_X1 U3731 ( .A(n6021), .ZN(n5623) );
  INV_X1 U3732 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U3733 ( .A1(n3435), .A2(n3434), .ZN(n3444) );
  OR2_X1 U3734 ( .A1(n3455), .A2(n3454), .ZN(n3474) );
  OR2_X1 U3735 ( .A1(n3412), .A2(n3411), .ZN(n3460) );
  OR2_X1 U3736 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  AOI21_X1 U3737 ( .B1(n3318), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3289), 
        .ZN(n3287) );
  AOI22_X1 U3738 ( .A1(n3380), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3023), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U3739 ( .A1(n3167), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3111) );
  AND2_X1 U3740 ( .A1(n4229), .A2(n4228), .ZN(n4293) );
  AOI22_X1 U3741 ( .A1(n3169), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3170) );
  OR2_X1 U3742 ( .A1(n3975), .A2(n3974), .ZN(n3994) );
  INV_X1 U3743 ( .A(n4071), .ZN(n4052) );
  AND2_X1 U3744 ( .A1(n3797), .A2(n5217), .ZN(n5189) );
  NOR2_X1 U3745 ( .A1(n3815), .A2(n5080), .ZN(n3780) );
  NAND2_X1 U3746 ( .A1(n5053), .A2(n5052), .ZN(n3059) );
  INV_X1 U3747 ( .A(n5444), .ZN(n3051) );
  NOR2_X1 U3748 ( .A1(n3503), .A2(n3066), .ZN(n3065) );
  AND2_X1 U3749 ( .A1(n5467), .A2(n5457), .ZN(n3503) );
  INV_X1 U3750 ( .A(n3502), .ZN(n3066) );
  INV_X1 U3751 ( .A(n5478), .ZN(n3500) );
  INV_X1 U3752 ( .A(n3333), .ZN(n3395) );
  OR2_X1 U3753 ( .A1(n3578), .A2(n3577), .ZN(n4242) );
  OR2_X1 U3754 ( .A1(n3379), .A2(n3310), .ZN(n3302) );
  AND2_X1 U3755 ( .A1(n3568), .A2(n3567), .ZN(n4222) );
  OR2_X1 U3756 ( .A1(n3566), .A2(n3565), .ZN(n3568) );
  AND2_X1 U3757 ( .A1(n6025), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3565)
         );
  OAI22_X1 U3758 ( .A1(n3563), .A2(n3562), .B1(n3561), .B2(n4228), .ZN(n3564)
         );
  INV_X1 U3759 ( .A(n3561), .ZN(n3570) );
  AND2_X1 U3760 ( .A1(n6185), .A2(n3321), .ZN(n4485) );
  AOI21_X1 U3761 ( .B1(n6424), .B2(n4544), .A(n5047), .ZN(n4475) );
  INV_X1 U3762 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6702) );
  AND2_X1 U3763 ( .A1(n6391), .A2(n6393), .ZN(n5744) );
  AND2_X1 U3764 ( .A1(n4102), .A2(n2998), .ZN(n6391) );
  INV_X1 U3765 ( .A(n4293), .ZN(n6393) );
  INV_X1 U3766 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5147) );
  INV_X1 U3767 ( .A(n5028), .ZN(n4159) );
  AND2_X1 U3768 ( .A1(n4161), .A2(n4160), .ZN(n5236) );
  OR2_X1 U3769 ( .A1(n3972), .A2(n3987), .ZN(n3992) );
  NOR2_X1 U3770 ( .A1(n3928), .A2(n4095), .ZN(n3947) );
  AND2_X1 U3771 ( .A1(n3949), .A2(n3948), .ZN(n3950) );
  NAND2_X1 U3772 ( .A1(n3879), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3896)
         );
  NOR2_X1 U3773 ( .A1(n5284), .A2(n3061), .ZN(n3060) );
  INV_X1 U3774 ( .A(n3063), .ZN(n3061) );
  AND2_X1 U3775 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n3584), .ZN(n3846)
         );
  INV_X1 U3776 ( .A(n3812), .ZN(n3584) );
  NAND2_X1 U3777 ( .A1(n3846), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3862)
         );
  AND2_X1 U3778 ( .A1(n3780), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3777)
         );
  AND2_X1 U3779 ( .A1(n3762), .A2(n3761), .ZN(n5232) );
  NAND2_X1 U3780 ( .A1(n3714), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3730)
         );
  INV_X1 U3781 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3731) );
  CLKBUF_X1 U3782 ( .A(n4898), .Z(n4899) );
  OR2_X1 U3783 ( .A1(n3666), .A2(n4846), .ZN(n3682) );
  NOR2_X1 U3784 ( .A1(n6711), .A2(n3682), .ZN(n3709) );
  OR2_X1 U3785 ( .A1(n3078), .A2(n3698), .ZN(n3077) );
  NAND2_X1 U3786 ( .A1(n3651), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3666)
         );
  INV_X1 U3787 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4846) );
  INV_X1 U3788 ( .A(n3643), .ZN(n3651) );
  NOR2_X1 U3789 ( .A1(n3636), .A2(n3583), .ZN(n3644) );
  INV_X1 U3790 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3583) );
  CLKBUF_X1 U3791 ( .A(n4555), .Z(n4556) );
  NOR2_X1 U3792 ( .A1(n4242), .A2(n3223), .ZN(n6389) );
  NOR2_X1 U3793 ( .A1(n5391), .A2(n3517), .ZN(n3518) );
  AND2_X1 U3794 ( .A1(n4196), .A2(n4195), .ZN(n5262) );
  NOR2_X2 U3795 ( .A1(n5270), .A2(n5262), .ZN(n5264) );
  INV_X1 U3796 ( .A(n4183), .ZN(n4184) );
  NOR2_X2 U3797 ( .A1(n5287), .A2(n5286), .ZN(n5289) );
  INV_X1 U3798 ( .A(n5434), .ZN(n5445) );
  NOR2_X1 U3799 ( .A1(n3483), .A2(n3482), .ZN(n3484) );
  INV_X1 U3800 ( .A(n4605), .ZN(n5615) );
  NAND2_X1 U3801 ( .A1(n4138), .A2(n4137), .ZN(n4551) );
  OR2_X1 U3802 ( .A1(n6510), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3587) );
  AND2_X1 U3803 ( .A1(n4277), .A2(n4263), .ZN(n5719) );
  AND2_X1 U3804 ( .A1(n4277), .A2(n6373), .ZN(n5726) );
  AND2_X1 U3805 ( .A1(n3266), .A2(n3265), .ZN(n3267) );
  OAI211_X1 U3806 ( .C1(n3310), .C2(n3378), .A(n3309), .B(n3308), .ZN(n3354)
         );
  OR3_X1 U3807 ( .A1(n4312), .A2(n4568), .A3(n4311), .ZN(n6375) );
  OR2_X1 U3808 ( .A1(n3031), .A2(n4704), .ZN(n4666) );
  OR2_X1 U3809 ( .A1(n3031), .A2(n4972), .ZN(n6030) );
  OR2_X1 U3810 ( .A1(n3033), .A2(n6260), .ZN(n6066) );
  AND2_X1 U3811 ( .A1(n4973), .A2(n3031), .ZN(n6184) );
  OR2_X1 U3812 ( .A1(n3033), .A2(n4970), .ZN(n6227) );
  OR2_X1 U3813 ( .A1(n4481), .A2(n6120), .ZN(n6301) );
  OR2_X1 U3814 ( .A1(n6228), .A2(n4579), .ZN(n6309) );
  NOR2_X2 U3815 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6317) );
  OR3_X1 U3816 ( .A1(n6501), .A2(STATE2_REG_0__SCAN_IN), .A3(n4475), .ZN(n4750) );
  NAND2_X1 U3817 ( .A1(n6526), .A2(n4833), .ZN(n5849) );
  OR3_X1 U3818 ( .A1(n6526), .A2(n4825), .A3(n6420), .ZN(n5858) );
  AND2_X1 U3819 ( .A1(n5858), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5843) );
  INV_X1 U3820 ( .A(n5849), .ZN(n5832) );
  INV_X1 U3821 ( .A(n5309), .ZN(n5306) );
  OR2_X1 U3822 ( .A1(n5353), .A2(n5354), .ZN(n5072) );
  NAND2_X1 U3823 ( .A1(n4570), .A2(n4569), .ZN(n5357) );
  OAI21_X1 U3824 ( .B1(n4568), .B2(n4567), .A(n4566), .ZN(n4569) );
  INV_X1 U3825 ( .A(n5072), .ZN(n5359) );
  NAND2_X1 U3826 ( .A1(n4409), .A2(n4297), .ZN(n5908) );
  INV_X1 U3827 ( .A(n4570), .ZN(n5906) );
  XNOR2_X1 U3828 ( .A(n3586), .B(n3585), .ZN(n4828) );
  OR2_X1 U3829 ( .A1(n4076), .A2(n5117), .ZN(n3586) );
  XNOR2_X1 U3830 ( .A(n3075), .B(n4083), .ZN(n5314) );
  NOR2_X1 U3831 ( .A1(n3076), .A2(n3072), .ZN(n3071) );
  INV_X1 U3832 ( .A(n5652), .ZN(n4097) );
  OR2_X1 U3833 ( .A1(n5654), .A2(n5499), .ZN(n4099) );
  INV_X1 U3834 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5424) );
  INV_X1 U3835 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5690) );
  INV_X1 U3836 ( .A(n5936), .ZN(n5492) );
  CLKBUF_X1 U3837 ( .A(n4891), .Z(n4892) );
  INV_X1 U3838 ( .A(n5753), .ZN(n5940) );
  INV_X1 U3839 ( .A(n5946), .ZN(n5494) );
  OAI21_X1 U3840 ( .B1(n5441), .B2(n3050), .A(n3047), .ZN(n5401) );
  NAND2_X1 U3841 ( .A1(n5418), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5409) );
  XNOR2_X1 U3842 ( .A(n4092), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5558)
         );
  NAND2_X1 U3843 ( .A1(n4271), .A2(n4270), .ZN(n5571) );
  OR2_X1 U3844 ( .A1(n6013), .A2(n4282), .ZN(n4271) );
  INV_X1 U3845 ( .A(n5294), .ZN(n5295) );
  INV_X1 U3846 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5596) );
  INV_X1 U3847 ( .A(n6010), .ZN(n5967) );
  CLKBUF_X1 U3848 ( .A(n5911), .Z(n5912) );
  CLKBUF_X1 U3849 ( .A(n4599), .Z(n4600) );
  CLKBUF_X1 U3850 ( .A(n4602), .Z(n4603) );
  INV_X1 U3851 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6216) );
  INV_X1 U3852 ( .A(n6317), .ZN(n6305) );
  INV_X1 U3853 ( .A(n4378), .ZN(n6120) );
  CLKBUF_X1 U3854 ( .A(n4480), .Z(n4481) );
  INV_X1 U3855 ( .A(n4476), .ZN(n6028) );
  INV_X1 U3856 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6025) );
  OAI21_X1 U3857 ( .B1(n4542), .B2(n6499), .A(n4669), .ZN(n6024) );
  NOR2_X1 U3858 ( .A1(n6501), .A2(n5743), .ZN(n5047) );
  NAND2_X1 U3859 ( .A1(n4826), .A2(n6501), .ZN(n6510) );
  NOR2_X1 U3860 ( .A1(n4665), .A2(n6260), .ZN(n4762) );
  OAI21_X1 U3861 ( .B1(n4673), .B2(n4671), .A(n4670), .ZN(n4761) );
  OAI21_X1 U3862 ( .B1(n6036), .B2(n6033), .A(n6032), .ZN(n6054) );
  OR3_X1 U3863 ( .A1(n6065), .A2(n6064), .A3(n6063), .ZN(n6086) );
  INV_X1 U3864 ( .A(n6147), .ZN(n6174) );
  OAI21_X1 U3865 ( .B1(n6159), .B2(n6158), .A(n6157), .ZN(n6177) );
  INV_X1 U3866 ( .A(n4819), .ZN(n4810) );
  OR2_X1 U3867 ( .A1(n6119), .A2(n4703), .ZN(n6154) );
  NOR2_X1 U3868 ( .A1(n6181), .A2(n6118), .ZN(n6208) );
  OAI21_X1 U3869 ( .B1(n6193), .B2(n6192), .A(n6191), .ZN(n6211) );
  NOR2_X1 U3870 ( .A1(n5499), .A2(n4498), .ZN(n6270) );
  NOR2_X1 U3871 ( .A1(n5499), .A2(n4731), .ZN(n6284) );
  INV_X1 U3872 ( .A(n6231), .ZN(n6308) );
  INV_X1 U3873 ( .A(n6235), .ZN(n6323) );
  INV_X1 U3874 ( .A(n6238), .ZN(n6329) );
  INV_X1 U3875 ( .A(n6241), .ZN(n6335) );
  INV_X1 U3876 ( .A(n6244), .ZN(n6341) );
  INV_X1 U3877 ( .A(n6248), .ZN(n6347) );
  INV_X1 U3878 ( .A(n6252), .ZN(n6353) );
  OR2_X1 U3879 ( .A1(n6309), .A2(n6260), .ZN(n6369) );
  INV_X1 U3880 ( .A(n6358), .ZN(n6364) );
  INV_X1 U3881 ( .A(n6258), .ZN(n6363) );
  INV_X1 U3882 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U3883 ( .A1(n6411), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U3884 ( .A1(n6303), .A2(n4826), .ZN(n6424) );
  INV_X1 U3885 ( .A(READY_N), .ZN(n6528) );
  NOR2_X1 U3886 ( .A1(n4211), .A2(n4210), .ZN(n4212) );
  NOR2_X1 U3887 ( .A1(n5311), .A2(n4209), .ZN(n4210) );
  NOR2_X1 U3888 ( .A1(n4291), .A2(n4290), .ZN(n4292) );
  INV_X1 U3889 ( .A(n4289), .ZN(n4290) );
  INV_X1 U3890 ( .A(n4274), .ZN(n4291) );
  AND2_X2 U3891 ( .A1(n3189), .A2(n3208), .ZN(n3092) );
  OR2_X1 U3892 ( .A1(n4094), .A2(n4093), .ZN(n3035) );
  NAND2_X1 U3893 ( .A1(n5260), .A2(n5261), .ZN(n5155) );
  OR2_X1 U3894 ( .A1(n4555), .A2(n3078), .ZN(n4767) );
  NOR2_X1 U3895 ( .A1(n5177), .A2(n3042), .ZN(n5178) );
  AND2_X1 U3896 ( .A1(n5467), .A2(n3499), .ZN(n3036) );
  NOR2_X1 U3897 ( .A1(n4094), .A2(n3069), .ZN(n5167) );
  NAND2_X1 U3898 ( .A1(n3062), .A2(n3063), .ZN(n5283) );
  NAND2_X1 U3899 ( .A1(n5441), .A2(n5444), .ZN(n4086) );
  AND2_X1 U3900 ( .A1(n5456), .A2(n3065), .ZN(n5454) );
  NAND2_X1 U3901 ( .A1(n3206), .A2(n3191), .ZN(n3223) );
  NAND2_X1 U3902 ( .A1(n5456), .A2(n3502), .ZN(n5466) );
  AND2_X1 U3903 ( .A1(n4836), .A2(n4149), .ZN(n3038) );
  OR2_X1 U3904 ( .A1(n3289), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3039)
         );
  NAND2_X1 U3905 ( .A1(n3606), .A2(n6414), .ZN(n3341) );
  NAND2_X1 U3906 ( .A1(n3046), .A2(n3044), .ZN(n5369) );
  NAND2_X1 U3907 ( .A1(n3280), .A2(n3205), .ZN(n4571) );
  NOR2_X1 U3908 ( .A1(n4555), .A2(n4655), .ZN(n4654) );
  INV_X1 U3909 ( .A(n4093), .ZN(n3070) );
  NAND2_X1 U3910 ( .A1(n5911), .A2(n3480), .ZN(n4867) );
  OR2_X1 U3911 ( .A1(n3051), .A2(n3510), .ZN(n3040) );
  AND2_X1 U3912 ( .A1(n3065), .A2(n3084), .ZN(n3041) );
  INV_X1 U3913 ( .A(n5052), .ZN(n3056) );
  NAND2_X1 U3914 ( .A1(n3848), .A2(n3847), .ZN(n3042) );
  OAI33_X1 U3915 ( .A1(n6263), .A2(n6265), .A3(n6262), .B1(n6301), .B2(n6305), 
        .B3(n6261), .ZN(n3043) );
  INV_X1 U3916 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6265) );
  INV_X1 U3917 ( .A(n3031), .ZN(n6261) );
  AND2_X2 U3918 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4386) );
  OAI211_X1 U3919 ( .C1(n4869), .C2(n3054), .A(n3052), .B(n3492), .ZN(n3494)
         );
  NAND2_X1 U3920 ( .A1(n5911), .A2(n3053), .ZN(n3052) );
  AND2_X1 U3921 ( .A1(n3491), .A2(n3480), .ZN(n3053) );
  INV_X1 U3922 ( .A(n3491), .ZN(n3054) );
  NAND2_X1 U3923 ( .A1(n4868), .A2(n3491), .ZN(n4914) );
  NAND2_X1 U3924 ( .A1(n4867), .A2(n4869), .ZN(n4868) );
  OAI21_X1 U3925 ( .B1(n5051), .B2(n5053), .A(n5052), .ZN(n5015) );
  NAND2_X1 U3926 ( .A1(n3062), .A2(n3060), .ZN(n5278) );
  INV_X2 U3927 ( .A(n5177), .ZN(n3062) );
  NAND2_X1 U3928 ( .A1(n3501), .A2(n3500), .ZN(n5456) );
  NAND2_X1 U3929 ( .A1(n5141), .A2(n5143), .ZN(n5125) );
  AND2_X1 U3930 ( .A1(n5141), .A2(n3071), .ZN(n3075) );
  INV_X1 U3931 ( .A(n4101), .ZN(n3076) );
  NAND2_X1 U3932 ( .A1(n5383), .A2(n5520), .ZN(n5362) );
  NAND2_X1 U3933 ( .A1(n3394), .A2(n3422), .ZN(n3590) );
  INV_X1 U3934 ( .A(n4557), .ZN(n3649) );
  AND2_X2 U3935 ( .A1(n5753), .A2(n3579), .ZN(n5936) );
  AND4_X1 U3936 ( .A1(n5411), .A2(n5573), .A3(n5596), .A4(n5435), .ZN(n3080)
         );
  OR2_X1 U3937 ( .A1(n5691), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3081)
         );
  AND2_X1 U3938 ( .A1(n5691), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3082)
         );
  OR2_X1 U3939 ( .A1(n5691), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3083)
         );
  OR2_X1 U3940 ( .A1(n5691), .A2(n3504), .ZN(n3084) );
  NAND2_X1 U3941 ( .A1(n3414), .A2(n3413), .ZN(n3085) );
  XNOR2_X1 U3942 ( .A(n4935), .B(n3747), .ZN(n5017) );
  AND2_X1 U3943 ( .A1(n3080), .A2(n3511), .ZN(n3087) );
  NAND2_X1 U3944 ( .A1(n5369), .A2(n3083), .ZN(n5393) );
  OR2_X2 U3945 ( .A1(n5305), .A2(n5313), .ZN(n5312) );
  INV_X1 U3946 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5080) );
  INV_X1 U3947 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4095) );
  AND2_X1 U3948 ( .A1(n5218), .A2(n5189), .ZN(n3088) );
  AND2_X1 U3949 ( .A1(n4099), .A2(n4098), .ZN(n3089) );
  INV_X1 U3950 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6711) );
  INV_X1 U3951 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3514) );
  AND4_X1 U3952 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3090)
         );
  INV_X1 U3953 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4538) );
  INV_X1 U3954 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3515) );
  INV_X1 U3955 ( .A(n4550), .ZN(n4137) );
  AND4_X1 U3956 ( .A1(n3107), .A2(n3106), .A3(n3105), .A4(n3104), .ZN(n3091)
         );
  NAND2_X1 U3957 ( .A1(n4449), .A2(n4450), .ZN(n4549) );
  INV_X1 U3958 ( .A(n4549), .ZN(n4138) );
  OR2_X1 U3959 ( .A1(n5102), .A2(n5130), .ZN(n3093) );
  NOR2_X1 U3960 ( .A1(n3252), .A2(n3251), .ZN(n3094) );
  INV_X1 U3961 ( .A(n3536), .ZN(n3534) );
  OR2_X1 U3962 ( .A1(n3433), .A2(n3432), .ZN(n3459) );
  AND2_X1 U3963 ( .A1(n3923), .A2(n3924), .ZN(n3962) );
  AOI22_X1 U3964 ( .A1(n3159), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3030), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3161) );
  INV_X1 U3965 ( .A(n5020), .ZN(n3745) );
  OR2_X1 U3966 ( .A1(n3397), .A2(n6531), .ZN(n3398) );
  NAND2_X1 U3967 ( .A1(n3560), .A2(n3523), .ZN(n3561) );
  OR2_X1 U3968 ( .A1(n3390), .A2(n3389), .ZN(n3415) );
  INV_X1 U3969 ( .A(n4855), .ZN(n3698) );
  NOR2_X1 U3970 ( .A1(n4028), .A2(n5147), .ZN(n4031) );
  OR2_X1 U3971 ( .A1(n3896), .A2(n5424), .ZN(n3928) );
  NAND2_X1 U3972 ( .A1(n5313), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3792) );
  NOR2_X1 U3973 ( .A1(n5027), .A2(n5026), .ZN(n4158) );
  INV_X1 U3974 ( .A(n3370), .ZN(n3371) );
  AND2_X1 U3975 ( .A1(n3947), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3967)
         );
  INV_X1 U3976 ( .A(n4864), .ZN(n4149) );
  OR2_X1 U3977 ( .A1(n3992), .A2(n3991), .ZN(n4028) );
  NOR2_X1 U3978 ( .A1(n3862), .A2(n5690), .ZN(n3879) );
  NOR2_X1 U3979 ( .A1(n3730), .A2(n3731), .ZN(n3759) );
  NAND2_X1 U3980 ( .A1(n3515), .A2(n3514), .ZN(n3516) );
  AND2_X1 U3981 ( .A1(n4177), .A2(n4176), .ZN(n5181) );
  OR2_X1 U3982 ( .A1(n6391), .A2(n4106), .ZN(n4218) );
  INV_X1 U3983 ( .A(n3391), .ZN(n3392) );
  AND2_X1 U3984 ( .A1(n3272), .A2(n3320), .ZN(n4974) );
  INV_X1 U3985 ( .A(n4637), .ZN(n4478) );
  NAND2_X1 U3986 ( .A1(n3967), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3972)
         );
  AND2_X1 U3987 ( .A1(REIP_REG_8__SCAN_IN), .A2(n4907), .ZN(n4952) );
  AND2_X1 U3988 ( .A1(n4828), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4829) );
  AND2_X1 U3989 ( .A1(n4165), .A2(n4164), .ZN(n5074) );
  NAND2_X1 U3990 ( .A1(n4112), .A2(n4111), .ZN(n4113) );
  AND2_X1 U3991 ( .A1(n3864), .A2(n3863), .ZN(n5291) );
  NAND2_X1 U3992 ( .A1(n3759), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3815)
         );
  AND2_X1 U3993 ( .A1(n3709), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3714)
         );
  AND3_X1 U3994 ( .A1(n3679), .A2(n3678), .A3(n3677), .ZN(n3680) );
  NAND2_X1 U3995 ( .A1(n5371), .A2(n3515), .ZN(n4214) );
  INV_X1 U3996 ( .A(n5407), .ZN(n5408) );
  INV_X1 U3997 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U3998 ( .A1(n5586), .A2(n4434), .ZN(n6013) );
  NAND2_X1 U3999 ( .A1(n4236), .A2(n4235), .ZN(n4277) );
  AND2_X1 U4000 ( .A1(n4383), .A2(n4382), .ZN(n4532) );
  INV_X1 U4001 ( .A(n6051), .ZN(n4797) );
  AND2_X1 U4002 ( .A1(n6151), .A2(n6153), .ZN(n6155) );
  INV_X1 U4003 ( .A(n6208), .ZN(n5006) );
  NAND2_X1 U4004 ( .A1(n4638), .A2(n6028), .ZN(n6181) );
  OR2_X1 U4005 ( .A1(n6228), .A2(n6066), .ZN(n4746) );
  NAND2_X1 U4006 ( .A1(n5744), .A2(n4566), .ZN(n5090) );
  INV_X1 U4007 ( .A(n4510), .ZN(n6396) );
  NOR2_X1 U4008 ( .A1(n6476), .A2(n5682), .ZN(n5666) );
  NOR2_X1 U4009 ( .A1(n6551), .A2(n5212), .ZN(n5202) );
  NOR2_X1 U4010 ( .A1(n5833), .A2(n4906), .ZN(n5790) );
  NOR2_X1 U4011 ( .A1(n4828), .A2(n4826), .ZN(n4827) );
  AND2_X1 U4012 ( .A1(n5858), .A2(n4829), .ZN(n5776) );
  NAND2_X1 U4013 ( .A1(n5093), .A2(n5090), .ZN(n6526) );
  AND2_X1 U4014 ( .A1(n5264), .A2(n5158), .ZN(n5160) );
  AND2_X1 U4015 ( .A1(n5239), .A2(n5074), .ZN(n5221) );
  INV_X1 U4016 ( .A(n3280), .ZN(n5313) );
  AND2_X1 U4017 ( .A1(n5357), .A2(n4574), .ZN(n5354) );
  AND2_X1 U4018 ( .A1(n4572), .A2(n4571), .ZN(n4573) );
  NAND2_X1 U4019 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n4544) );
  OR2_X1 U4020 ( .A1(n4299), .A2(n3189), .ZN(n4570) );
  AND2_X1 U4021 ( .A1(n5908), .A2(n4299), .ZN(n5905) );
  NAND2_X1 U4022 ( .A1(n3777), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3812)
         );
  AND2_X1 U4023 ( .A1(n3007), .A2(n5071), .ZN(n5218) );
  INV_X1 U4024 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5411) );
  AND2_X1 U4025 ( .A1(n4284), .A2(n4283), .ZN(n5574) );
  INV_X1 U4026 ( .A(n5721), .ZN(n6016) );
  INV_X1 U4027 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4826) );
  INV_X1 U4028 ( .A(n6418), .ZN(n4566) );
  NAND2_X1 U4029 ( .A1(n4484), .A2(n4483), .ZN(n4786) );
  OAI21_X1 U4030 ( .B1(n4583), .B2(n4582), .A(n4981), .ZN(n4796) );
  AND2_X1 U4031 ( .A1(n6026), .A2(n4970), .ZN(n6051) );
  INV_X1 U4032 ( .A(n6154), .ZN(n6176) );
  OR2_X1 U4033 ( .A1(n4707), .A2(n4706), .ZN(n4809) );
  NOR2_X1 U4034 ( .A1(n6181), .A2(n6066), .ZN(n4819) );
  INV_X1 U4035 ( .A(n4979), .ZN(n5008) );
  NOR2_X1 U4036 ( .A1(n6181), .A2(n4703), .ZN(n6210) );
  INV_X1 U4037 ( .A(n4746), .ZN(n6253) );
  NOR2_X1 U4038 ( .A1(n5499), .A2(n4493), .ZN(n6324) );
  NOR2_X1 U4039 ( .A1(n5499), .A2(n4732), .ZN(n6342) );
  AND2_X1 U4040 ( .A1(n4826), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6411) );
  INV_X1 U4041 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6437) );
  INV_X1 U4042 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6429) );
  INV_X1 U4043 ( .A(n6494), .ZN(n6734) );
  INV_X1 U4044 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6446) );
  INV_X1 U4045 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5750) );
  INV_X1 U4046 ( .A(n5843), .ZN(n5821) );
  INV_X1 U4047 ( .A(n5831), .ZN(n5851) );
  INV_X1 U4048 ( .A(n5193), .ZN(n5253) );
  OR2_X1 U4049 ( .A1(n5305), .A2(n3280), .ZN(n5309) );
  INV_X1 U4050 ( .A(n5115), .ZN(n5319) );
  OR2_X1 U4051 ( .A1(n5260), .A2(n5267), .ZN(n5644) );
  OAI21_X1 U4052 ( .B1(n5191), .B2(n3088), .A(n5190), .ZN(n5452) );
  OR2_X1 U4053 ( .A1(n4854), .A2(n4856), .ZN(n5786) );
  OR2_X1 U4054 ( .A1(n3616), .A2(n4326), .ZN(n5846) );
  NAND2_X1 U4055 ( .A1(n5871), .A2(n3208), .ZN(n5859) );
  OR2_X1 U4056 ( .A1(n4544), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6405) );
  INV_X1 U4057 ( .A(n5871), .ZN(n5889) );
  INV_X1 U4058 ( .A(n5905), .ZN(n4377) );
  INV_X1 U4059 ( .A(n3589), .ZN(n4085) );
  OR2_X1 U4060 ( .A1(n5936), .A2(n3582), .ZN(n5946) );
  NAND2_X2 U4061 ( .A1(n4409), .A2(n6389), .ZN(n5753) );
  AND2_X1 U4062 ( .A1(n4285), .A2(n5574), .ZN(n5566) );
  OR2_X1 U4063 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4672), .ZN(n4792)
         );
  INV_X1 U4064 ( .A(n4667), .ZN(n4766) );
  INV_X1 U4065 ( .A(n4583), .ZN(n4803) );
  NAND2_X1 U4066 ( .A1(n6026), .A2(n6260), .ZN(n6089) );
  AOI22_X1 U4067 ( .A1(n6095), .A2(n6093), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6097), .ZN(n6117) );
  OR2_X1 U4068 ( .A1(n6119), .A2(n6118), .ZN(n6147) );
  INV_X1 U4069 ( .A(n6152), .ZN(n6180) );
  INV_X1 U4070 ( .A(n4702), .ZN(n4816) );
  INV_X1 U4071 ( .A(n6307), .ZN(n4726) );
  INV_X1 U4072 ( .A(n6346), .ZN(n4718) );
  AOI22_X1 U4073 ( .A1(n4978), .A2(n6184), .B1(n6264), .B2(n4975), .ZN(n5010)
         );
  AOI22_X1 U4074 ( .A1(n6188), .A2(n6192), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6189), .ZN(n6214) );
  AOI21_X1 U4075 ( .B1(n4621), .B2(n4620), .A(n4619), .ZN(n4755) );
  AOI22_X1 U4076 ( .A1(n6221), .A2(n6220), .B1(n6219), .B2(n6225), .ZN(n6259)
         );
  INV_X1 U4077 ( .A(n6330), .ZN(n6279) );
  INV_X1 U4078 ( .A(n6365), .ZN(n6299) );
  INV_X1 U4079 ( .A(n6245), .ZN(n6351) );
  INV_X1 U4080 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6501) );
  INV_X1 U4081 ( .A(n6498), .ZN(n6428) );
  NAND2_X1 U4082 ( .A1(n4221), .A2(n6437), .ZN(n6434) );
  INV_X1 U4083 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6456) );
  NOR2_X1 U4084 ( .A1(n6429), .A2(STATE_REG_0__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U4085 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6464), .ZN(n6494) );
  NAND2_X1 U4086 ( .A1(n4213), .A2(n4212), .ZN(U2829) );
  INV_X1 U4087 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3612) );
  AND2_X2 U4088 ( .A1(n3612), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4515)
         );
  NOR2_X2 U4089 ( .A1(n3095), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4391)
         );
  NOR2_X2 U4090 ( .A1(n3612), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3103)
         );
  AOI22_X1 U4091 ( .A1(n3034), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3099) );
  AOI22_X1 U4092 ( .A1(n3380), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3023), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3098) );
  NOR2_X4 U4093 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3102) );
  AOI22_X1 U4094 ( .A1(n3167), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3097) );
  AND2_X2 U4095 ( .A1(n3101), .A2(n4386), .ZN(n3169) );
  AOI22_X1 U4096 ( .A1(n3168), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3096) );
  AOI22_X1 U4097 ( .A1(n3030), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3107) );
  AND2_X2 U4098 ( .A1(n4391), .A2(n4536), .ZN(n3181) );
  AND2_X2 U4099 ( .A1(n4391), .A2(n3101), .ZN(n3406) );
  AOI22_X1 U4100 ( .A1(n3181), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3106) );
  AOI22_X1 U4101 ( .A1(n3182), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3105) );
  AND2_X2 U4102 ( .A1(n4536), .A2(n4386), .ZN(n3198) );
  AOI22_X1 U4103 ( .A1(n3242), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3104) );
  XNOR2_X1 U4104 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n4220) );
  NAND2_X1 U4105 ( .A1(n3189), .A2(n4220), .ZN(n3284) );
  AOI22_X1 U4106 ( .A1(n3168), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3110) );
  AOI22_X1 U4107 ( .A1(n3247), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3109) );
  AOI22_X1 U4108 ( .A1(n3024), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3164), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3108) );
  NAND4_X1 U4109 ( .A1(n3111), .A2(n3110), .A3(n3109), .A4(n3108), .ZN(n3117)
         );
  AOI22_X1 U4110 ( .A1(n3182), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4111 ( .A1(n3030), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3026), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U4112 ( .A1(n3181), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U4113 ( .A1(n3242), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3112) );
  NAND4_X1 U4114 ( .A1(n3115), .A2(n3114), .A3(n3113), .A4(n3112), .ZN(n3116)
         );
  NAND2_X1 U4115 ( .A1(n3284), .A2(n3176), .ZN(n3138) );
  NAND2_X1 U4116 ( .A1(n3030), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3121)
         );
  NAND2_X1 U4117 ( .A1(n3181), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3120)
         );
  NAND2_X1 U4118 ( .A1(n3167), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3119) );
  NAND2_X1 U4119 ( .A1(n3166), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3118) );
  NAND2_X1 U4120 ( .A1(n3034), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3125) );
  NAND2_X1 U4121 ( .A1(n4019), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3124) );
  NAND2_X1 U4122 ( .A1(n3168), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3123) );
  NAND2_X1 U4123 ( .A1(n3169), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3122) );
  NAND2_X1 U4124 ( .A1(n3182), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3129) );
  NAND2_X1 U4125 ( .A1(n3406), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3128) );
  NAND2_X1 U4126 ( .A1(n3159), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3127) );
  NAND2_X1 U4127 ( .A1(n3241), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3126)
         );
  NAND2_X1 U4128 ( .A1(n3025), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3133)
         );
  NAND2_X1 U4129 ( .A1(n3023), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3132)
         );
  NAND2_X1 U4130 ( .A1(n3242), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U4131 ( .A1(n3198), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3130)
         );
  NAND4_X4 U4132 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n3208)
         );
  AOI22_X1 U4133 ( .A1(n3167), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3142) );
  AOI22_X1 U4134 ( .A1(n3380), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3023), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U4135 ( .A1(n3168), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U4136 ( .A1(n3181), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4137 ( .A1(n3030), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4138 ( .A1(n3182), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U4139 ( .A1(n3242), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3143) );
  AOI22_X1 U4140 ( .A1(n3034), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4141 ( .A1(n3167), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U4142 ( .A1(n3168), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3149) );
  NAND4_X1 U4143 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n3158)
         );
  AOI22_X1 U4144 ( .A1(n3030), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4145 ( .A1(n3181), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4146 ( .A1(n3182), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4147 ( .A1(n3242), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3153) );
  NAND4_X1 U4148 ( .A1(n3156), .A2(n3155), .A3(n3154), .A4(n3153), .ZN(n3157)
         );
  AOI22_X1 U4149 ( .A1(n3182), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4150 ( .A1(n3181), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4151 ( .A1(n3242), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3160) );
  NAND4_X1 U4152 ( .A1(n3163), .A2(n3162), .A3(n3161), .A4(n3160), .ZN(n3175)
         );
  AOI22_X1 U4153 ( .A1(n3025), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3164), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4154 ( .A1(n3247), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4155 ( .A1(n3167), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3171) );
  NAND4_X1 U4156 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3174)
         );
  AOI22_X1 U4157 ( .A1(n3025), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3023), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4158 ( .A1(n3034), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4159 ( .A1(n3167), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4160 ( .A1(n3168), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3177) );
  NAND4_X1 U4161 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3188)
         );
  AOI22_X1 U4162 ( .A1(n3181), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4163 ( .A1(n3030), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3185) );
  AOI22_X1 U4164 ( .A1(n3182), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4165 ( .A1(n3242), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3183) );
  NAND4_X1 U4166 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(n3187)
         );
  NAND3_X1 U4167 ( .A1(n3216), .A2(n3280), .A3(n3206), .ZN(n4103) );
  NAND2_X1 U4168 ( .A1(n3021), .A2(n3092), .ZN(n3233) );
  NAND3_X1 U4169 ( .A1(n3190), .A2(n4250), .A3(n3233), .ZN(n3204) );
  NAND2_X1 U4170 ( .A1(n3210), .A2(n3206), .ZN(n3193) );
  AND2_X2 U4171 ( .A1(n3193), .A2(n3192), .ZN(n4252) );
  AOI22_X1 U4172 ( .A1(n3165), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3023), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4173 ( .A1(n3025), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3168), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3196) );
  AOI22_X1 U4174 ( .A1(n3181), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3195) );
  AOI22_X1 U4175 ( .A1(n3182), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4176 ( .A1(n3030), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3202) );
  AOI22_X1 U4177 ( .A1(n3167), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4178 ( .A1(n3034), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4179 ( .A1(n3242), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3199) );
  NAND2_X1 U4180 ( .A1(n4252), .A2(n3277), .ZN(n3578) );
  OAI211_X1 U4181 ( .C1(n3206), .C2(n3205), .A(n3279), .B(n3216), .ZN(n3207)
         );
  NAND2_X1 U4182 ( .A1(n3218), .A2(n3279), .ZN(n3219) );
  INV_X1 U4183 ( .A(n3378), .ZN(n3334) );
  NAND2_X1 U4184 ( .A1(n3219), .A2(n3334), .ZN(n3211) );
  NAND2_X1 U4185 ( .A1(n3318), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3215) );
  INV_X1 U4186 ( .A(n6411), .ZN(n3274) );
  INV_X1 U4187 ( .A(n3587), .ZN(n3273) );
  MUX2_X1 U4188 ( .A(n3274), .B(n3273), .S(n6216), .Z(n3213) );
  INV_X1 U4189 ( .A(n3213), .ZN(n3214) );
  NAND2_X1 U4190 ( .A1(n3215), .A2(n3214), .ZN(n3271) );
  AND3_X1 U4191 ( .A1(n3216), .A2(n3206), .A3(n3205), .ZN(n3217) );
  INV_X1 U4192 ( .A(n4102), .ZN(n3221) );
  NAND3_X1 U4193 ( .A1(n3221), .A2(n3219), .A3(n5745), .ZN(n4262) );
  OR2_X1 U4194 ( .A1(n6510), .A2(n6414), .ZN(n6419) );
  INV_X1 U4195 ( .A(n6419), .ZN(n3222) );
  NAND2_X1 U4196 ( .A1(n4250), .A2(n3222), .ZN(n3227) );
  NAND2_X1 U4197 ( .A1(n4882), .A2(n3223), .ZN(n3226) );
  NAND2_X1 U4198 ( .A1(n3224), .A2(n3208), .ZN(n3225) );
  NAND2_X1 U4199 ( .A1(n3226), .A2(n3225), .ZN(n4254) );
  INV_X1 U4200 ( .A(n3210), .ZN(n3576) );
  NAND2_X1 U4201 ( .A1(n3576), .A2(n3209), .ZN(n3228) );
  AOI21_X1 U4202 ( .B1(n4252), .B2(n3228), .A(n3189), .ZN(n3236) );
  NAND3_X1 U4203 ( .A1(n3229), .A2(n4246), .A3(n4116), .ZN(n3234) );
  NOR2_X1 U4204 ( .A1(n3224), .A2(n3231), .ZN(n4109) );
  NAND2_X1 U4205 ( .A1(n3232), .A2(n4109), .ZN(n4514) );
  NAND3_X1 U4206 ( .A1(n3234), .A2(n4514), .A3(n3233), .ZN(n3235) );
  NOR2_X1 U4207 ( .A1(n3236), .A2(n3235), .ZN(n3237) );
  AND2_X1 U4208 ( .A1(n3238), .A2(n3237), .ZN(n3239) );
  NAND2_X1 U4209 ( .A1(n4262), .A2(n3239), .ZN(n3270) );
  AOI22_X1 U4210 ( .A1(n4038), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4211 ( .A1(n4043), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3246) );
  AOI22_X1 U4212 ( .A1(n4000), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4213 ( .A1(n4018), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3244) );
  INV_X1 U4214 ( .A(n3242), .ZN(n4517) );
  AOI22_X1 U4215 ( .A1(n4055), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3243) );
  NAND4_X1 U4216 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(n3252)
         );
  AOI22_X1 U4217 ( .A1(n4036), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4218 ( .A1(n4037), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4219 ( .A1(n3380), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3248) );
  NAND3_X1 U4220 ( .A1(n3250), .A2(n3249), .A3(n3248), .ZN(n3251) );
  NOR2_X1 U4221 ( .A1(n3379), .A2(n3487), .ZN(n3307) );
  NAND2_X1 U4222 ( .A1(n3206), .A2(n3487), .ZN(n3265) );
  AOI22_X1 U4223 ( .A1(n4043), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4224 ( .A1(n4036), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4037), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4225 ( .A1(n4000), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4226 ( .A1(n4018), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3254) );
  NAND4_X1 U4227 ( .A1(n3257), .A2(n3256), .A3(n3255), .A4(n3254), .ZN(n3263)
         );
  AOI22_X1 U4228 ( .A1(n3380), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4229 ( .A1(n4019), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4230 ( .A1(n4038), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4231 ( .A1(n4013), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3258) );
  NAND4_X1 U4232 ( .A1(n3261), .A2(n3260), .A3(n3259), .A4(n3258), .ZN(n3262)
         );
  INV_X1 U4233 ( .A(n3355), .ZN(n3264) );
  MUX2_X1 U4234 ( .A(n3307), .B(n3481), .S(n3264), .Z(n3344) );
  NAND2_X1 U4235 ( .A1(n3560), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3268) );
  AOI21_X1 U4236 ( .B1(n2998), .B2(n3355), .A(n6414), .ZN(n3266) );
  NAND2_X1 U4237 ( .A1(n3268), .A2(n3267), .ZN(n3342) );
  AOI21_X1 U4238 ( .B1(n3344), .B2(n3342), .A(n3481), .ZN(n3269) );
  NAND2_X1 U4239 ( .A1(n3341), .A2(n3269), .ZN(n3305) );
  NAND2_X1 U4240 ( .A1(n4976), .A2(n6216), .ZN(n3272) );
  NAND2_X1 U4241 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4242 ( .A1(n3273), .A2(n4974), .ZN(n3276) );
  NAND2_X1 U4243 ( .A1(n3274), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U4244 ( .A1(n3276), .A2(n3275), .ZN(n3289) );
  NAND2_X1 U4245 ( .A1(n3277), .A2(n3176), .ZN(n3278) );
  AND2_X1 U4246 ( .A1(n4232), .A2(n3208), .ZN(n4237) );
  NAND3_X1 U4247 ( .A1(n3176), .A2(n3279), .A3(n4115), .ZN(n4247) );
  INV_X1 U4248 ( .A(n4247), .ZN(n3282) );
  INV_X1 U4249 ( .A(n4571), .ZN(n3281) );
  NAND2_X1 U4250 ( .A1(n3282), .A2(n3281), .ZN(n3283) );
  NOR2_X1 U4251 ( .A1(n3283), .A2(n4246), .ZN(n4239) );
  AOI21_X1 U4252 ( .B1(n4237), .B2(n3284), .A(n4239), .ZN(n3285) );
  NAND2_X1 U4253 ( .A1(n3285), .A2(n4241), .ZN(n3286) );
  NAND2_X1 U4254 ( .A1(n3286), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U4255 ( .A1(n3287), .A2(n3288), .ZN(n3316) );
  NAND2_X1 U4256 ( .A1(n3012), .A2(n3039), .ZN(n3290) );
  AOI22_X1 U4257 ( .A1(n4036), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4258 ( .A1(n3380), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4259 ( .A1(n4037), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4260 ( .A1(n4038), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3292) );
  NAND4_X1 U4261 ( .A1(n3295), .A2(n3294), .A3(n3293), .A4(n3292), .ZN(n3301)
         );
  AOI22_X1 U4262 ( .A1(n4043), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4263 ( .A1(n4000), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4264 ( .A1(n4018), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4265 ( .A1(n4055), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3296) );
  NAND4_X1 U4266 ( .A1(n3299), .A2(n3298), .A3(n3297), .A4(n3296), .ZN(n3300)
         );
  NAND2_X1 U4267 ( .A1(n3303), .A2(n3302), .ZN(n3304) );
  NAND2_X1 U4268 ( .A1(n3304), .A2(n3305), .ZN(n3311) );
  OAI21_X1 U4269 ( .B1(n3305), .B2(n3004), .A(n3311), .ZN(n3306) );
  INV_X1 U4270 ( .A(n3306), .ZN(n3353) );
  NAND2_X1 U4271 ( .A1(n3560), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3309) );
  INV_X1 U4272 ( .A(n3307), .ZN(n3308) );
  NAND2_X1 U4273 ( .A1(n3353), .A2(n3354), .ZN(n3312) );
  NAND2_X1 U4274 ( .A1(n3312), .A2(n3311), .ZN(n3368) );
  INV_X1 U4275 ( .A(n3313), .ZN(n3315) );
  NAND2_X1 U4276 ( .A1(n3315), .A2(n3314), .ZN(n3317) );
  NAND2_X1 U4277 ( .A1(n3317), .A2(n3020), .ZN(n3369) );
  INV_X1 U4278 ( .A(n3320), .ZN(n3319) );
  NAND2_X1 U4279 ( .A1(n3319), .A2(n6381), .ZN(n6185) );
  NAND2_X1 U4280 ( .A1(n3320), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3321) );
  OAI22_X1 U4281 ( .A1(n4485), .A2(n3587), .B1(n6411), .B2(n6381), .ZN(n3322)
         );
  XNOR2_X1 U4282 ( .A(n3369), .B(n3370), .ZN(n4480) );
  AOI22_X1 U4283 ( .A1(n4036), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4284 ( .A1(n3401), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4285 ( .A1(n4037), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4286 ( .A1(n4038), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3323) );
  NAND4_X1 U4287 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3332)
         );
  AOI22_X1 U4288 ( .A1(n4043), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4289 ( .A1(n4000), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3329) );
  INV_X1 U4290 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6689) );
  AOI22_X1 U4291 ( .A1(n4018), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3328) );
  INV_X2 U4292 ( .A(n4517), .ZN(n4055) );
  AOI22_X1 U4293 ( .A1(n4055), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3327) );
  NAND4_X1 U4294 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3331)
         );
  AOI22_X1 U4295 ( .A1(n3560), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3334), 
        .B2(n3333), .ZN(n3335) );
  XNOR2_X1 U4296 ( .A(n3336), .B(n3335), .ZN(n3367) );
  INV_X1 U4297 ( .A(n3367), .ZN(n3337) );
  NAND2_X1 U4298 ( .A1(n3598), .A2(n3523), .ZN(n3340) );
  NAND2_X1 U4299 ( .A1(n3355), .A2(n3356), .ZN(n3396) );
  XNOR2_X1 U4300 ( .A(n3396), .B(n3395), .ZN(n3338) );
  AND2_X1 U4301 ( .A1(n2998), .A2(n3231), .ZN(n3346) );
  AOI21_X1 U4302 ( .B1(n3338), .B2(n3092), .A(n3346), .ZN(n3339) );
  NAND2_X1 U4303 ( .A1(n3340), .A2(n3339), .ZN(n5937) );
  NAND2_X1 U4304 ( .A1(n5937), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3363)
         );
  INV_X1 U4305 ( .A(n3342), .ZN(n3343) );
  XNOR2_X1 U4306 ( .A(n3344), .B(n3343), .ZN(n3345) );
  OR2_X1 U4307 ( .A1(n4970), .A2(n3482), .ZN(n3350) );
  INV_X1 U4308 ( .A(n3092), .ZN(n6531) );
  INV_X1 U4309 ( .A(n3346), .ZN(n3347) );
  OAI21_X1 U4310 ( .B1(n6531), .B2(n3355), .A(n3347), .ZN(n3348) );
  INV_X1 U4311 ( .A(n3348), .ZN(n3349) );
  NAND2_X1 U4312 ( .A1(n3350), .A2(n3349), .ZN(n4394) );
  NAND2_X1 U4313 ( .A1(n4394), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3351)
         );
  INV_X1 U4314 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U4315 ( .A1(n3351), .A2(n6012), .ZN(n3352) );
  AND2_X1 U4316 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U4317 ( .A1(n4394), .A2(n6015), .ZN(n3361) );
  AND2_X1 U4318 ( .A1(n3352), .A2(n3361), .ZN(n4433) );
  NAND2_X1 U4319 ( .A1(n3033), .A2(n3523), .ZN(n3360) );
  OAI21_X1 U4320 ( .B1(n3356), .B2(n3355), .A(n3396), .ZN(n3357) );
  OAI211_X1 U4321 ( .C1(n3357), .C2(n6531), .A(n3277), .B(n3191), .ZN(n3358)
         );
  INV_X1 U4322 ( .A(n3358), .ZN(n3359) );
  INV_X1 U4323 ( .A(n3361), .ZN(n3362) );
  NAND2_X1 U4324 ( .A1(n3363), .A2(n5938), .ZN(n3366) );
  INV_X1 U4325 ( .A(n5937), .ZN(n3364) );
  NAND2_X1 U4326 ( .A1(n3364), .A2(n6669), .ZN(n3365) );
  NAND2_X1 U4327 ( .A1(n3368), .A2(n3367), .ZN(n3393) );
  INV_X1 U4328 ( .A(n3369), .ZN(n3372) );
  NAND2_X1 U4329 ( .A1(n3372), .A2(n3371), .ZN(n4314) );
  NAND2_X1 U4330 ( .A1(n3005), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3377) );
  NAND3_X1 U4331 ( .A1(n6265), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6156) );
  INV_X1 U4332 ( .A(n6156), .ZN(n3373) );
  NAND2_X1 U4333 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3373), .ZN(n6153) );
  NAND2_X1 U4334 ( .A1(n6265), .A2(n6153), .ZN(n3374) );
  NAND3_X1 U4335 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6304) );
  INV_X1 U4336 ( .A(n6304), .ZN(n6316) );
  NAND2_X1 U4337 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6316), .ZN(n6306) );
  NAND2_X1 U4338 ( .A1(n3374), .A2(n6306), .ZN(n4618) );
  OAI22_X1 U4339 ( .A1(n3587), .A2(n4618), .B1(n6411), .B2(n6265), .ZN(n3375)
         );
  INV_X1 U4340 ( .A(n3375), .ZN(n3376) );
  XNOR2_X1 U4341 ( .A(n4314), .B(n6059), .ZN(n4479) );
  AOI22_X1 U4342 ( .A1(n4018), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4343 ( .A1(n3401), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4344 ( .A1(n4000), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4345 ( .A1(n4019), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3381) );
  NAND4_X1 U4346 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3390)
         );
  AOI22_X1 U4347 ( .A1(n4036), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4037), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4348 ( .A1(n3937), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4349 ( .A1(n4055), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4350 ( .A1(n4038), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3385) );
  NAND4_X1 U4351 ( .A1(n3388), .A2(n3387), .A3(n3386), .A4(n3385), .ZN(n3389)
         );
  AOI22_X1 U4352 ( .A1(n3569), .A2(n3415), .B1(n3560), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3391) );
  NAND2_X1 U4353 ( .A1(n3393), .A2(n4637), .ZN(n3394) );
  NAND2_X1 U4354 ( .A1(n3396), .A2(n3395), .ZN(n3416) );
  XNOR2_X1 U4355 ( .A(n3416), .B(n3415), .ZN(n3397) );
  INV_X1 U4356 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6007) );
  XNOR2_X1 U4357 ( .A(n3399), .B(n6007), .ZN(n5929) );
  NAND2_X1 U4358 ( .A1(n5928), .A2(n5929), .ZN(n5931) );
  NAND2_X1 U4359 ( .A1(n3399), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3400)
         );
  NAND2_X1 U4360 ( .A1(n5931), .A2(n3400), .ZN(n4890) );
  AOI22_X1 U4361 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4036), .B1(n4019), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4362 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3401), .B1(n3932), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4363 ( .A1(n4037), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4364 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4038), .B1(n3901), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3402) );
  NAND4_X1 U4365 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(n3412)
         );
  AOI22_X1 U4366 ( .A1(n4043), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4367 ( .A1(n4000), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4368 ( .A1(n4018), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4369 ( .A1(n4055), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3407) );
  NAND4_X1 U4370 ( .A1(n3410), .A2(n3409), .A3(n3408), .A4(n3407), .ZN(n3411)
         );
  NAND2_X1 U4371 ( .A1(n3569), .A2(n3460), .ZN(n3414) );
  NAND2_X1 U4372 ( .A1(n3560), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3413) );
  NAND2_X1 U4373 ( .A1(n3620), .A2(n3523), .ZN(n3419) );
  NAND2_X1 U4374 ( .A1(n3416), .A2(n3415), .ZN(n3462) );
  XNOR2_X1 U4375 ( .A(n3462), .B(n3460), .ZN(n3417) );
  NAND2_X1 U4376 ( .A1(n3417), .A2(n3092), .ZN(n3418) );
  NAND2_X1 U4377 ( .A1(n3419), .A2(n3418), .ZN(n3420) );
  INV_X1 U4378 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5999) );
  XNOR2_X1 U4379 ( .A(n3420), .B(n5999), .ZN(n4893) );
  NAND2_X1 U4380 ( .A1(n4890), .A2(n4893), .ZN(n4891) );
  NAND2_X1 U4381 ( .A1(n3420), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3421)
         );
  NAND2_X1 U4382 ( .A1(n4891), .A2(n3421), .ZN(n5919) );
  INV_X1 U4383 ( .A(n3422), .ZN(n3423) );
  NAND2_X1 U4384 ( .A1(n3423), .A2(n3085), .ZN(n3443) );
  AOI22_X1 U4385 ( .A1(n4000), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4386 ( .A1(n3932), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4387 ( .A1(n4018), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4388 ( .A1(n4037), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3424) );
  NAND4_X1 U4389 ( .A1(n3427), .A2(n3426), .A3(n3425), .A4(n3424), .ZN(n3433)
         );
  AOI22_X1 U4390 ( .A1(n4036), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4391 ( .A1(n4043), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4392 ( .A1(n4055), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4393 ( .A1(n3401), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3428) );
  NAND4_X1 U4394 ( .A1(n3431), .A2(n3430), .A3(n3429), .A4(n3428), .ZN(n3432)
         );
  NAND2_X1 U4395 ( .A1(n3569), .A2(n3459), .ZN(n3435) );
  NAND2_X1 U4396 ( .A1(n3560), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3434) );
  XNOR2_X1 U4397 ( .A(n3443), .B(n3444), .ZN(n3629) );
  NAND2_X1 U4398 ( .A1(n3629), .A2(n3523), .ZN(n3440) );
  INV_X1 U4399 ( .A(n3460), .ZN(n3436) );
  OR2_X1 U4400 ( .A1(n3462), .A2(n3436), .ZN(n3437) );
  XNOR2_X1 U4401 ( .A(n3437), .B(n3459), .ZN(n3438) );
  NAND2_X1 U4402 ( .A1(n3438), .A2(n3092), .ZN(n3439) );
  NAND2_X1 U4403 ( .A1(n3440), .A2(n3439), .ZN(n3441) );
  INV_X1 U4404 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4265) );
  XNOR2_X1 U4405 ( .A(n3441), .B(n4265), .ZN(n5921) );
  NAND2_X1 U4406 ( .A1(n5919), .A2(n5921), .ZN(n5920) );
  NAND2_X1 U4407 ( .A1(n3441), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3442)
         );
  NAND2_X1 U4408 ( .A1(n5920), .A2(n3442), .ZN(n4599) );
  INV_X1 U4409 ( .A(n3443), .ZN(n3445) );
  NAND2_X1 U4410 ( .A1(n3445), .A2(n3444), .ZN(n3469) );
  AOI22_X1 U4411 ( .A1(n4036), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4412 ( .A1(n3401), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4413 ( .A1(n4037), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4414 ( .A1(n4038), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3446) );
  NAND4_X1 U4415 ( .A1(n3449), .A2(n3448), .A3(n3447), .A4(n3446), .ZN(n3455)
         );
  AOI22_X1 U4416 ( .A1(n4043), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4417 ( .A1(n4000), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4418 ( .A1(n4018), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4419 ( .A1(n4055), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3450) );
  NAND4_X1 U4420 ( .A1(n3453), .A2(n3452), .A3(n3451), .A4(n3450), .ZN(n3454)
         );
  NAND2_X1 U4421 ( .A1(n3569), .A2(n3474), .ZN(n3457) );
  NAND2_X1 U4422 ( .A1(n3560), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3456) );
  INV_X1 U4423 ( .A(n3468), .ZN(n3458) );
  NAND2_X1 U4424 ( .A1(n3635), .A2(n3523), .ZN(n3465) );
  NAND2_X1 U4425 ( .A1(n3460), .A2(n3459), .ZN(n3461) );
  OR2_X1 U4426 ( .A1(n3462), .A2(n3461), .ZN(n3473) );
  XNOR2_X1 U4427 ( .A(n3473), .B(n3474), .ZN(n3463) );
  NAND2_X1 U4428 ( .A1(n3463), .A2(n3092), .ZN(n3464) );
  NAND2_X1 U4429 ( .A1(n3465), .A2(n3464), .ZN(n3466) );
  INV_X1 U4430 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4607) );
  XNOR2_X1 U4431 ( .A(n3466), .B(n4607), .ZN(n4601) );
  NAND2_X1 U4432 ( .A1(n4599), .A2(n4601), .ZN(n4602) );
  NAND2_X1 U4433 ( .A1(n3466), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3467)
         );
  NAND2_X1 U4434 ( .A1(n4602), .A2(n3467), .ZN(n5910) );
  NAND2_X1 U4435 ( .A1(n3569), .A2(n3487), .ZN(n3471) );
  NAND2_X1 U4436 ( .A1(n3560), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3470) );
  NAND2_X1 U4437 ( .A1(n3471), .A2(n3470), .ZN(n3472) );
  NAND2_X1 U4438 ( .A1(n3648), .A2(n3523), .ZN(n3478) );
  INV_X1 U4439 ( .A(n3473), .ZN(n3475) );
  NAND2_X1 U4440 ( .A1(n3475), .A2(n3474), .ZN(n3486) );
  XNOR2_X1 U4441 ( .A(n3486), .B(n3487), .ZN(n3476) );
  NAND2_X1 U4442 ( .A1(n3476), .A2(n3092), .ZN(n3477) );
  NAND2_X1 U4443 ( .A1(n3478), .A2(n3477), .ZN(n3479) );
  INV_X1 U4444 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5978) );
  XNOR2_X1 U4445 ( .A(n3479), .B(n5978), .ZN(n5913) );
  NAND2_X1 U4446 ( .A1(n5910), .A2(n5913), .ZN(n5911) );
  NAND2_X1 U4447 ( .A1(n3479), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3480)
         );
  INV_X1 U4448 ( .A(n3481), .ZN(n3483) );
  INV_X1 U4449 ( .A(n3486), .ZN(n3488) );
  NAND3_X1 U4450 ( .A1(n3488), .A2(n3092), .A3(n3487), .ZN(n3489) );
  NAND2_X1 U4451 ( .A1(n5467), .A2(n3489), .ZN(n3490) );
  INV_X1 U4452 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5973) );
  XNOR2_X1 U4453 ( .A(n3490), .B(n5973), .ZN(n4869) );
  NAND2_X1 U4454 ( .A1(n3490), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3491)
         );
  INV_X1 U4455 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5963) );
  NAND2_X1 U4456 ( .A1(n5436), .A2(n5963), .ZN(n3492) );
  OR2_X1 U4457 ( .A1(n5436), .A2(n5963), .ZN(n3493) );
  INV_X1 U4458 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3495) );
  NAND2_X1 U4459 ( .A1(n5467), .A2(n3495), .ZN(n4922) );
  INV_X1 U4460 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5953) );
  AND2_X1 U4461 ( .A1(n5436), .A2(n5953), .ZN(n3498) );
  OR2_X1 U4462 ( .A1(n5436), .A2(n3495), .ZN(n4959) );
  OAI21_X1 U4463 ( .B1(n5953), .B2(n5436), .A(n4959), .ZN(n3496) );
  INV_X1 U4464 ( .A(n3496), .ZN(n3497) );
  INV_X1 U4465 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5060) );
  NOR2_X1 U4466 ( .A1(n5436), .A2(n5060), .ZN(n5053) );
  NAND2_X1 U4467 ( .A1(n5467), .A2(n5060), .ZN(n5052) );
  XNOR2_X1 U4468 ( .A(n5436), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5016)
         );
  INV_X1 U4469 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3499) );
  INV_X1 U4470 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6577) );
  AND2_X1 U4471 ( .A1(n5436), .A2(n6577), .ZN(n5486) );
  OR2_X1 U4472 ( .A1(n5436), .A2(n6577), .ZN(n5485) );
  INV_X1 U4473 ( .A(n5476), .ZN(n3501) );
  INV_X1 U4474 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5617) );
  XNOR2_X1 U4475 ( .A(n5436), .B(n5617), .ZN(n5478) );
  NAND2_X1 U4476 ( .A1(n5467), .A2(n5617), .ZN(n3502) );
  INV_X1 U4477 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U4478 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5589) );
  INV_X1 U4479 ( .A(n5589), .ZN(n3504) );
  NOR3_X1 U4480 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n3505) );
  NAND2_X1 U4481 ( .A1(n5436), .A2(n5596), .ZN(n5444) );
  NAND2_X1 U4482 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4089) );
  INV_X1 U4483 ( .A(n4089), .ZN(n3509) );
  NAND2_X1 U4484 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4286) );
  INV_X1 U4485 ( .A(n4286), .ZN(n3508) );
  INV_X1 U4486 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3507) );
  NAND3_X1 U4487 ( .A1(n3509), .A2(n3508), .A3(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3510) );
  INV_X1 U4488 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5573) );
  INV_X1 U4489 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5435) );
  AND2_X1 U4490 ( .A1(n3507), .A2(n6698), .ZN(n3511) );
  INV_X1 U4491 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U4492 ( .A1(n5691), .A2(n5539), .ZN(n5392) );
  INV_X1 U4493 ( .A(n5392), .ZN(n3512) );
  NOR2_X1 U4494 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5519) );
  NOR2_X1 U4495 ( .A1(n5371), .A2(n3516), .ZN(n3521) );
  NAND2_X1 U4496 ( .A1(n5436), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5391) );
  INV_X1 U4497 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U4498 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U4499 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3519) );
  NOR2_X1 U4500 ( .A1(n5510), .A2(n3519), .ZN(n5500) );
  INV_X1 U4501 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4390) );
  XNOR2_X1 U4502 ( .A(n3522), .B(n4390), .ZN(n5509) );
  NAND2_X1 U4503 ( .A1(n6216), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3536) );
  XNOR2_X1 U4504 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3535) );
  NAND2_X1 U4505 ( .A1(n3534), .A2(n3535), .ZN(n3525) );
  NAND2_X1 U4506 ( .A1(n4976), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3524) );
  NAND2_X1 U4507 ( .A1(n3525), .A2(n3524), .ZN(n3529) );
  XNOR2_X1 U4508 ( .A(n6645), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3530)
         );
  NAND2_X1 U4509 ( .A1(n3529), .A2(n3530), .ZN(n3527) );
  NAND2_X1 U4510 ( .A1(n6381), .A2(n6645), .ZN(n3526) );
  NAND2_X1 U4511 ( .A1(n3527), .A2(n3526), .ZN(n3557) );
  XNOR2_X1 U4512 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3556) );
  INV_X1 U4513 ( .A(n3556), .ZN(n3528) );
  XNOR2_X1 U4514 ( .A(n3557), .B(n3528), .ZN(n4225) );
  INV_X1 U4515 ( .A(n4225), .ZN(n3555) );
  XOR2_X1 U4516 ( .A(n3530), .B(n3529), .Z(n4224) );
  NAND2_X1 U4517 ( .A1(n3569), .A2(n4224), .ZN(n3551) );
  NAND2_X1 U4518 ( .A1(n3189), .A2(n3191), .ZN(n3531) );
  AND2_X1 U4519 ( .A1(n3551), .A2(n3552), .ZN(n3533) );
  OAI22_X1 U4520 ( .A1(n3533), .A2(n3555), .B1(n4224), .B2(n3532), .ZN(n3554)
         );
  INV_X1 U4521 ( .A(n3569), .ZN(n3542) );
  OAI21_X1 U4522 ( .B1(n3542), .B2(n3189), .A(n3191), .ZN(n3548) );
  XOR2_X1 U4523 ( .A(n3535), .B(n3534), .Z(n4223) );
  NOR2_X1 U4524 ( .A1(n3548), .A2(n4223), .ZN(n3543) );
  OAI21_X1 U4525 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6216), .A(n3536), 
        .ZN(n3541) );
  INV_X1 U4526 ( .A(n3541), .ZN(n3537) );
  NAND2_X1 U4527 ( .A1(n3223), .A2(n3537), .ZN(n3539) );
  NAND2_X1 U4528 ( .A1(n3539), .A2(n3538), .ZN(n3540) );
  AND2_X1 U4529 ( .A1(n3552), .A2(n3540), .ZN(n3544) );
  NOR4_X1 U4530 ( .A1(n3543), .A2(n3542), .A3(n3541), .A4(n3544), .ZN(n3547)
         );
  INV_X1 U4531 ( .A(n4223), .ZN(n3546) );
  INV_X1 U4532 ( .A(n3544), .ZN(n3545) );
  OAI22_X1 U4533 ( .A1(n3547), .A2(n3570), .B1(n3546), .B2(n3545), .ZN(n3550)
         );
  NAND3_X1 U4534 ( .A1(n3548), .A2(STATE2_REG_0__SCAN_IN), .A3(n4223), .ZN(
        n3549) );
  OAI211_X1 U4535 ( .C1(n3552), .C2(n3551), .A(n3550), .B(n3549), .ZN(n3553)
         );
  AOI22_X1 U4536 ( .A1(n3570), .A2(n3555), .B1(n3554), .B2(n3553), .ZN(n3563)
         );
  NAND2_X1 U4537 ( .A1(n3557), .A2(n3556), .ZN(n3559) );
  NAND2_X1 U4538 ( .A1(n6265), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3558) );
  NAND2_X1 U4539 ( .A1(n3559), .A2(n3558), .ZN(n3566) );
  NOR2_X1 U4540 ( .A1(n3560), .A2(n4228), .ZN(n3562) );
  NAND2_X1 U4541 ( .A1(n3569), .A2(n4222), .ZN(n3571) );
  AOI21_X1 U4542 ( .B1(n3572), .B2(n3571), .A(n3570), .ZN(n3574) );
  NOR2_X1 U4543 ( .A1(n3572), .A2(n4222), .ZN(n3573) );
  NAND2_X1 U4544 ( .A1(n3209), .A2(n3280), .ZN(n3575) );
  AND2_X1 U4545 ( .A1(n4385), .A2(n2998), .ZN(n3577) );
  NAND2_X1 U4546 ( .A1(n6305), .A2(n3587), .ZN(n6527) );
  NAND2_X1 U4547 ( .A1(n6527), .A2(n6414), .ZN(n3579) );
  NAND2_X1 U4548 ( .A1(n6414), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3581) );
  NAND2_X1 U4549 ( .A1(n5750), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3580) );
  NAND2_X1 U4550 ( .A1(n3581), .A2(n3580), .ZN(n4468) );
  INV_X1 U4551 ( .A(n4468), .ZN(n3582) );
  NAND2_X1 U4552 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3613) );
  NOR2_X1 U4553 ( .A1(n6702), .A2(n3613), .ZN(n3622) );
  NAND2_X1 U4554 ( .A1(n3622), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3621)
         );
  INV_X1 U4555 ( .A(n3621), .ZN(n3630) );
  NAND2_X1 U4556 ( .A1(n3630), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3636)
         );
  NAND2_X1 U4557 ( .A1(n3644), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3643)
         );
  INV_X1 U4558 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3987) );
  INV_X1 U4559 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3991) );
  INV_X1 U4560 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5117) );
  INV_X1 U4561 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3585) );
  NOR2_X4 U4562 ( .A1(n3587), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6000) );
  AND2_X1 U4563 ( .A1(n6000), .A2(REIP_REG_31__SCAN_IN), .ZN(n5503) );
  AOI21_X1 U4564 ( .B1(n5936), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5503), 
        .ZN(n3588) );
  OAI21_X1 U4565 ( .B1(n5946), .B2(n4828), .A(n3588), .ZN(n3589) );
  NAND2_X1 U4566 ( .A1(n4638), .A2(n3827), .ZN(n3597) );
  NAND2_X1 U4567 ( .A1(n3281), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3625) );
  INV_X1 U4568 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4523) );
  NOR2_X4 U4569 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4077) );
  INV_X1 U4570 ( .A(n3613), .ZN(n3592) );
  INV_X1 U4571 ( .A(n3622), .ZN(n3591) );
  OAI21_X1 U4572 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3592), .A(n3591), 
        .ZN(n5935) );
  AOI22_X1 U4573 ( .A1(n4077), .A2(n5935), .B1(n4081), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U4574 ( .A1(n4082), .A2(EAX_REG_3__SCAN_IN), .ZN(n3593) );
  OAI211_X1 U4575 ( .C1(n3625), .C2(n4523), .A(n3594), .B(n3593), .ZN(n3595)
         );
  INV_X1 U4576 ( .A(n3595), .ZN(n3596) );
  NAND2_X1 U4577 ( .A1(n4476), .A2(n3827), .ZN(n3599) );
  INV_X1 U4578 ( .A(n4081), .ZN(n3791) );
  NAND2_X1 U4579 ( .A1(n3599), .A2(n3791), .ZN(n3617) );
  NAND2_X1 U4580 ( .A1(n4477), .A2(n3827), .ZN(n3604) );
  AOI22_X1 U4581 ( .A1(n4082), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6303), .ZN(n3602) );
  INV_X1 U4582 ( .A(n3625), .ZN(n3600) );
  NAND2_X1 U4583 ( .A1(n3600), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3601) );
  AND2_X1 U4584 ( .A1(n3602), .A2(n3601), .ZN(n3603) );
  NAND2_X1 U4585 ( .A1(n4970), .A2(n3230), .ZN(n3605) );
  NAND2_X1 U4586 ( .A1(n3605), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U4587 ( .A1(n4082), .A2(EAX_REG_0__SCAN_IN), .ZN(n3608) );
  NAND2_X1 U4588 ( .A1(n6303), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3607)
         );
  OAI211_X1 U4589 ( .C1(n3625), .C2(n3095), .A(n3608), .B(n3607), .ZN(n3609)
         );
  AOI21_X1 U4590 ( .B1(n3029), .B2(n3827), .A(n3609), .ZN(n4406) );
  OR2_X1 U4591 ( .A1(n4405), .A2(n4406), .ZN(n4403) );
  INV_X1 U4592 ( .A(n4406), .ZN(n3610) );
  OR2_X1 U4593 ( .A1(n3610), .A2(n4074), .ZN(n3611) );
  NAND2_X1 U4594 ( .A1(n4403), .A2(n3611), .ZN(n4324) );
  OAI21_X1 U4595 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3613), .ZN(n5945) );
  AOI22_X1 U4596 ( .A1(n4081), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4077), 
        .B2(n5945), .ZN(n3615) );
  NAND2_X1 U4597 ( .A1(n4082), .A2(EAX_REG_2__SCAN_IN), .ZN(n3614) );
  OAI211_X1 U4598 ( .C1(n3625), .C2(n3612), .A(n3615), .B(n3614), .ZN(n4442)
         );
  NAND2_X1 U4599 ( .A1(n4443), .A2(n4442), .ZN(n3619) );
  NAND2_X1 U4600 ( .A1(n3617), .A2(n3616), .ZN(n3618) );
  NAND2_X1 U4601 ( .A1(n3620), .A2(n3827), .ZN(n3628) );
  OAI21_X1 U4602 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3622), .A(n3621), 
        .ZN(n5822) );
  NAND2_X1 U4603 ( .A1(n4082), .A2(EAX_REG_4__SCAN_IN), .ZN(n3624) );
  OAI21_X1 U4604 ( .B1(n5750), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6303), 
        .ZN(n3623) );
  OAI211_X1 U4605 ( .C1(n3625), .C2(n4538), .A(n3624), .B(n3623), .ZN(n3626)
         );
  OAI21_X1 U4606 ( .B1(n4074), .B2(n5822), .A(n3626), .ZN(n3627) );
  NAND2_X1 U4607 ( .A1(n3628), .A2(n3627), .ZN(n4447) );
  NAND2_X1 U4608 ( .A1(n3629), .A2(n3827), .ZN(n3634) );
  INV_X1 U4609 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5807) );
  OAI21_X1 U4610 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3630), .A(n3636), 
        .ZN(n5926) );
  NAND2_X1 U4611 ( .A1(n5926), .A2(n4077), .ZN(n3631) );
  OAI21_X1 U4612 ( .B1(n3791), .B2(n5807), .A(n3631), .ZN(n3632) );
  AOI21_X1 U4613 ( .B1(n4082), .B2(EAX_REG_5__SCAN_IN), .A(n3632), .ZN(n3633)
         );
  NAND2_X1 U4614 ( .A1(n3634), .A2(n3633), .ZN(n4552) );
  NAND2_X1 U4615 ( .A1(n3635), .A2(n3827), .ZN(n3642) );
  INV_X1 U4616 ( .A(n3636), .ZN(n3637) );
  XNOR2_X1 U4617 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3637), .ZN(n4943) );
  INV_X1 U4618 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3639) );
  OAI21_X1 U4619 ( .B1(n5750), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6303), 
        .ZN(n3638) );
  OAI21_X1 U4620 ( .B1(n3792), .B2(n3639), .A(n3638), .ZN(n3640) );
  OAI21_X1 U4621 ( .B1(n4943), .B2(n4074), .A(n3640), .ZN(n3641) );
  NAND2_X1 U4622 ( .A1(n3642), .A2(n3641), .ZN(n4459) );
  INV_X1 U4623 ( .A(n4462), .ZN(n3650) );
  INV_X1 U4624 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3646) );
  OAI21_X1 U4625 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n3644), .A(n3643), 
        .ZN(n5918) );
  AOI22_X1 U4626 ( .A1(n4077), .A2(n5918), .B1(n4081), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3645) );
  OAI21_X1 U4627 ( .B1(n3792), .B2(n3646), .A(n3645), .ZN(n3647) );
  AOI21_X1 U4628 ( .B1(n3648), .B2(n3827), .A(n3647), .ZN(n4557) );
  NAND2_X1 U4629 ( .A1(n3650), .A2(n3649), .ZN(n4555) );
  XNOR2_X1 U4630 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3651), .ZN(n4908) );
  AOI22_X1 U4631 ( .A1(n4018), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4632 ( .A1(n4037), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4633 ( .A1(n4036), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4634 ( .A1(n4000), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3652) );
  NAND4_X1 U4635 ( .A1(n3655), .A2(n3654), .A3(n3653), .A4(n3652), .ZN(n3661)
         );
  AOI22_X1 U4636 ( .A1(n4019), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3659) );
  AOI22_X1 U4637 ( .A1(n3401), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4638 ( .A1(n4043), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4639 ( .A1(n3937), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3656) );
  NAND4_X1 U4640 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(n3660)
         );
  OAI21_X1 U4641 ( .B1(n3661), .B2(n3660), .A(n3827), .ZN(n3664) );
  NAND2_X1 U4642 ( .A1(n4082), .A2(EAX_REG_8__SCAN_IN), .ZN(n3663) );
  NAND2_X1 U4643 ( .A1(n4081), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3662)
         );
  NAND3_X1 U4644 ( .A1(n3664), .A2(n3663), .A3(n3662), .ZN(n3665) );
  AOI21_X1 U4645 ( .B1(n4908), .B2(n4077), .A(n3665), .ZN(n4655) );
  XNOR2_X1 U4646 ( .A(n3666), .B(n4846), .ZN(n4917) );
  NAND2_X1 U4647 ( .A1(n4917), .A2(n4077), .ZN(n3681) );
  AOI22_X1 U4648 ( .A1(n3401), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4649 ( .A1(n4043), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4650 ( .A1(n4037), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4651 ( .A1(n4038), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3667) );
  NAND4_X1 U4652 ( .A1(n3670), .A2(n3669), .A3(n3668), .A4(n3667), .ZN(n3676)
         );
  AOI22_X1 U4653 ( .A1(n4036), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4654 ( .A1(n3937), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4655 ( .A1(n4018), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4656 ( .A1(n4000), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3671) );
  NAND4_X1 U4657 ( .A1(n3674), .A2(n3673), .A3(n3672), .A4(n3671), .ZN(n3675)
         );
  OAI21_X1 U4658 ( .B1(n3676), .B2(n3675), .A(n3827), .ZN(n3679) );
  NAND2_X1 U4659 ( .A1(n4082), .A2(EAX_REG_9__SCAN_IN), .ZN(n3678) );
  NAND2_X1 U4660 ( .A1(n4081), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3677)
         );
  NAND2_X1 U4661 ( .A1(n3681), .A2(n3680), .ZN(n4769) );
  AOI21_X1 U4662 ( .B1(n6711), .B2(n3682), .A(n3709), .ZN(n5783) );
  OR2_X1 U4663 ( .A1(n5783), .A2(n4074), .ZN(n3697) );
  AOI22_X1 U4664 ( .A1(n4018), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4665 ( .A1(n4036), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4037), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4666 ( .A1(n4043), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4667 ( .A1(n4055), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3683) );
  NAND4_X1 U4668 ( .A1(n3686), .A2(n3685), .A3(n3684), .A4(n3683), .ZN(n3692)
         );
  AOI22_X1 U4669 ( .A1(n3401), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4670 ( .A1(n4000), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4671 ( .A1(n4019), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4672 ( .A1(n4038), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3687) );
  NAND4_X1 U4673 ( .A1(n3690), .A2(n3689), .A3(n3688), .A4(n3687), .ZN(n3691)
         );
  OAI21_X1 U4674 ( .B1(n3692), .B2(n3691), .A(n3827), .ZN(n3695) );
  NAND2_X1 U4675 ( .A1(n4082), .A2(EAX_REG_10__SCAN_IN), .ZN(n3694) );
  NAND2_X1 U4676 ( .A1(n4081), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3693)
         );
  AND3_X1 U4677 ( .A1(n3695), .A2(n3694), .A3(n3693), .ZN(n3696) );
  NAND2_X1 U4678 ( .A1(n3697), .A2(n3696), .ZN(n4855) );
  AOI22_X1 U4679 ( .A1(n4043), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4680 ( .A1(n4037), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4681 ( .A1(n3401), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4682 ( .A1(n4038), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3699) );
  NAND4_X1 U4683 ( .A1(n3702), .A2(n3701), .A3(n3700), .A4(n3699), .ZN(n3708)
         );
  AOI22_X1 U4684 ( .A1(n4000), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4685 ( .A1(n4036), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4686 ( .A1(n4018), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4687 ( .A1(n4055), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3703) );
  NAND4_X1 U4688 ( .A1(n3706), .A2(n3705), .A3(n3704), .A4(n3703), .ZN(n3707)
         );
  NOR2_X1 U4689 ( .A1(n3708), .A2(n3707), .ZN(n3713) );
  INV_X1 U4690 ( .A(n3827), .ZN(n3712) );
  XNOR2_X1 U4691 ( .A(n3709), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4962)
         );
  NAND2_X1 U4692 ( .A1(n4962), .A2(n4077), .ZN(n3711) );
  AOI22_X1 U4693 ( .A1(n4082), .A2(EAX_REG_11__SCAN_IN), .B1(n4081), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3710) );
  OAI211_X1 U4694 ( .C1(n3713), .C2(n3712), .A(n3711), .B(n3710), .ZN(n4900)
         );
  XOR2_X1 U4695 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3714), .Z(n5777) );
  NAND2_X1 U4696 ( .A1(n5777), .A2(n4077), .ZN(n3717) );
  INV_X1 U4697 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4967) );
  OAI21_X1 U4698 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n5750), .A(n6303), 
        .ZN(n3715) );
  OAI21_X1 U4699 ( .B1(n3792), .B2(n4967), .A(n3715), .ZN(n3716) );
  NAND2_X1 U4700 ( .A1(n3717), .A2(n3716), .ZN(n3729) );
  AOI22_X1 U4701 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3028), .B1(n4037), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4702 ( .A1(n4036), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4703 ( .A1(n4043), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4704 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3401), .B1(n3901), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3718) );
  NAND4_X1 U4705 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), .ZN(n3727)
         );
  AOI22_X1 U4706 ( .A1(n4018), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4707 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4000), .B1(n4013), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4708 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4038), .B1(n3027), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4709 ( .A1(n4055), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3722) );
  NAND4_X1 U4710 ( .A1(n3725), .A2(n3724), .A3(n3723), .A4(n3722), .ZN(n3726)
         );
  OAI21_X1 U4711 ( .B1(n3727), .B2(n3726), .A(n3827), .ZN(n3728) );
  NAND2_X1 U4712 ( .A1(n3729), .A2(n3728), .ZN(n4936) );
  XNOR2_X1 U4713 ( .A(n3730), .B(n3731), .ZN(n5032) );
  INV_X1 U4714 ( .A(EAX_REG_13__SCAN_IN), .ZN(n3732) );
  OAI22_X1 U4715 ( .A1(n3792), .A2(n3732), .B1(n3791), .B2(n3731), .ZN(n3733)
         );
  AOI21_X1 U4716 ( .B1(n5032), .B2(n4077), .A(n3733), .ZN(n3747) );
  INV_X1 U4717 ( .A(n5017), .ZN(n3746) );
  AOI22_X1 U4718 ( .A1(n4018), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4037), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4719 ( .A1(n3932), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4720 ( .A1(n3401), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4721 ( .A1(n4036), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3734) );
  NAND4_X1 U4722 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), .ZN(n3743)
         );
  AOI22_X1 U4723 ( .A1(n3937), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4724 ( .A1(n4000), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4725 ( .A1(n4043), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4726 ( .A1(n4038), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3738) );
  NAND4_X1 U4727 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(n3742)
         );
  OR2_X1 U4728 ( .A1(n3743), .A2(n3742), .ZN(n3744) );
  NAND2_X1 U4729 ( .A1(n3827), .A2(n3744), .ZN(n5020) );
  INV_X1 U4730 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5358) );
  INV_X1 U4731 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5491) );
  OAI22_X1 U4732 ( .A1(n3792), .A2(n5358), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5491), .ZN(n3748) );
  NAND2_X1 U4733 ( .A1(n3748), .A2(n4074), .ZN(n3762) );
  AOI22_X1 U4734 ( .A1(n4043), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4735 ( .A1(n4019), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4736 ( .A1(n4037), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4737 ( .A1(n3937), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3749) );
  NAND4_X1 U4738 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3758)
         );
  AOI22_X1 U4739 ( .A1(n4000), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4740 ( .A1(n4036), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4741 ( .A1(n3027), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4742 ( .A1(n4038), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3753) );
  NAND4_X1 U4743 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3757)
         );
  OR2_X1 U4744 ( .A1(n3758), .A2(n3757), .ZN(n3760) );
  XNOR2_X1 U4745 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3759), .ZN(n5489)
         );
  AOI22_X1 U4746 ( .A1(n3827), .A2(n3760), .B1(n4077), .B2(n5489), .ZN(n3761)
         );
  AOI22_X1 U4747 ( .A1(n3182), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4748 ( .A1(n4000), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4749 ( .A1(n4036), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4750 ( .A1(n4038), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3763) );
  NAND4_X1 U4751 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3772)
         );
  AOI22_X1 U4752 ( .A1(n4037), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4753 ( .A1(n3401), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4754 ( .A1(n4043), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4755 ( .A1(n3027), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3767) );
  NAND4_X1 U4756 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n3771)
         );
  NOR2_X1 U4757 ( .A1(n3772), .A2(n3771), .ZN(n3776) );
  NAND2_X1 U4758 ( .A1(n6303), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3773)
         );
  NAND2_X1 U4759 ( .A1(n4074), .A2(n3773), .ZN(n3774) );
  AOI21_X1 U4760 ( .B1(n4082), .B2(EAX_REG_17__SCAN_IN), .A(n3774), .ZN(n3775)
         );
  OAI21_X1 U4761 ( .B1(n4052), .B2(n3776), .A(n3775), .ZN(n3779) );
  OAI21_X1 U4762 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3777), .A(n3812), 
        .ZN(n5700) );
  OR2_X1 U4763 ( .A1(n4074), .A2(n5700), .ZN(n3778) );
  NAND2_X1 U4764 ( .A1(n3779), .A2(n3778), .ZN(n5204) );
  INV_X1 U4765 ( .A(n5204), .ZN(n3797) );
  XNOR2_X1 U4766 ( .A(n3780), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5222)
         );
  NAND2_X1 U4767 ( .A1(n5222), .A2(n4077), .ZN(n3796) );
  AOI22_X1 U4768 ( .A1(n4036), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4769 ( .A1(n3932), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4770 ( .A1(n4037), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4771 ( .A1(n4043), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3781) );
  NAND4_X1 U4772 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3790)
         );
  AOI22_X1 U4773 ( .A1(n4018), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4774 ( .A1(n4055), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4775 ( .A1(n3401), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4776 ( .A1(n4000), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4777 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3789)
         );
  OR2_X1 U4778 ( .A1(n3790), .A2(n3789), .ZN(n3794) );
  INV_X1 U4779 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4301) );
  INV_X1 U4780 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5470) );
  OAI22_X1 U4781 ( .A1(n3792), .A2(n4301), .B1(n3791), .B2(n5470), .ZN(n3793)
         );
  AOI21_X1 U4782 ( .B1(n4071), .B2(n3794), .A(n3793), .ZN(n3795) );
  NAND2_X1 U4783 ( .A1(n3796), .A2(n3795), .ZN(n5217) );
  AOI22_X1 U4784 ( .A1(n4036), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4785 ( .A1(n3401), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4786 ( .A1(n4037), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4787 ( .A1(n4038), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3798) );
  NAND4_X1 U4788 ( .A1(n3801), .A2(n3800), .A3(n3799), .A4(n3798), .ZN(n3807)
         );
  AOI22_X1 U4789 ( .A1(n4043), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4790 ( .A1(n4000), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4791 ( .A1(n4018), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4792 ( .A1(n4055), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3802) );
  NAND4_X1 U4793 ( .A1(n3805), .A2(n3804), .A3(n3803), .A4(n3802), .ZN(n3806)
         );
  NOR2_X1 U4794 ( .A1(n3807), .A2(n3806), .ZN(n3811) );
  INV_X1 U4795 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3808) );
  AOI21_X1 U4796 ( .B1(n3808), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3809) );
  AOI21_X1 U4797 ( .B1(n4082), .B2(EAX_REG_18__SCAN_IN), .A(n3809), .ZN(n3810)
         );
  OAI21_X1 U4798 ( .B1(n4052), .B2(n3811), .A(n3810), .ZN(n3814) );
  XNOR2_X1 U4799 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3812), .ZN(n5451)
         );
  NAND2_X1 U4800 ( .A1(n5451), .A2(n4077), .ZN(n3813) );
  AND2_X1 U4801 ( .A1(n3814), .A2(n3813), .ZN(n5191) );
  AND2_X1 U4802 ( .A1(n5189), .A2(n5191), .ZN(n3830) );
  XOR2_X1 U4803 ( .A(n5080), .B(n3815), .Z(n5482) );
  AOI22_X1 U4804 ( .A1(n4037), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4805 ( .A1(n4036), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4806 ( .A1(n3182), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4807 ( .A1(n4043), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3816) );
  NAND4_X1 U4808 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3825)
         );
  AOI22_X1 U4809 ( .A1(n3937), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4810 ( .A1(n3932), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4811 ( .A1(n4000), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4812 ( .A1(n4038), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4813 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3824)
         );
  OR2_X1 U4814 ( .A1(n3825), .A2(n3824), .ZN(n3826) );
  AOI22_X1 U4815 ( .A1(n3827), .A2(n3826), .B1(n4081), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3829) );
  NAND2_X1 U4816 ( .A1(n4082), .A2(EAX_REG_15__SCAN_IN), .ZN(n3828) );
  OAI211_X1 U4817 ( .C1(n5482), .C2(n4074), .A(n3829), .B(n3828), .ZN(n5071)
         );
  AND2_X1 U4818 ( .A1(n3830), .A2(n5071), .ZN(n3831) );
  NAND2_X1 U4819 ( .A1(n5069), .A2(n3831), .ZN(n5177) );
  AOI22_X1 U4820 ( .A1(n4018), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4821 ( .A1(n4000), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4037), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4822 ( .A1(n4036), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3401), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4823 ( .A1(n4043), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3832) );
  NAND4_X1 U4824 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3841)
         );
  AOI22_X1 U4825 ( .A1(n3028), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4826 ( .A1(n4055), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4827 ( .A1(n4038), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4828 ( .A1(n3938), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3836) );
  NAND4_X1 U4829 ( .A1(n3839), .A2(n3838), .A3(n3837), .A4(n3836), .ZN(n3840)
         );
  NOR2_X1 U4830 ( .A1(n3841), .A2(n3840), .ZN(n3845) );
  NAND2_X1 U4831 ( .A1(n6303), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3842)
         );
  NAND2_X1 U4832 ( .A1(n4074), .A2(n3842), .ZN(n3843) );
  AOI21_X1 U4833 ( .B1(n4082), .B2(EAX_REG_19__SCAN_IN), .A(n3843), .ZN(n3844)
         );
  OAI21_X1 U4834 ( .B1(n4052), .B2(n3845), .A(n3844), .ZN(n3848) );
  OAI21_X1 U4835 ( .B1(n3846), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n3862), 
        .ZN(n5447) );
  OR2_X1 U4836 ( .A1(n5447), .A2(n4074), .ZN(n3847) );
  AOI22_X1 U4837 ( .A1(n4018), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4838 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4036), .B1(n3028), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4839 ( .A1(n4000), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4840 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4055), .B1(n3027), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3849) );
  NAND4_X1 U4841 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3858)
         );
  AOI22_X1 U4842 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n3932), .B1(n3401), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4843 ( .A1(n4037), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4844 ( .A1(n3937), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4845 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4038), .B1(n3901), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4846 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3857)
         );
  NOR2_X1 U4847 ( .A1(n3858), .A2(n3857), .ZN(n3861) );
  OAI21_X1 U4848 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5690), .A(n4074), .ZN(
        n3859) );
  AOI21_X1 U4849 ( .B1(n4082), .B2(EAX_REG_20__SCAN_IN), .A(n3859), .ZN(n3860)
         );
  OAI21_X1 U4850 ( .B1(n4052), .B2(n3861), .A(n3860), .ZN(n3864) );
  XNOR2_X1 U4851 ( .A(n3862), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5681)
         );
  NAND2_X1 U4852 ( .A1(n5681), .A2(n4077), .ZN(n3863) );
  AOI22_X1 U4853 ( .A1(n4037), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4854 ( .A1(n3401), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4855 ( .A1(n3937), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4856 ( .A1(n4055), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3865) );
  NAND4_X1 U4857 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3874)
         );
  AOI22_X1 U4858 ( .A1(n4018), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4859 ( .A1(n4000), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4860 ( .A1(n3028), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4861 ( .A1(n4036), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3869) );
  NAND4_X1 U4862 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3873)
         );
  NOR2_X1 U4863 ( .A1(n3874), .A2(n3873), .ZN(n3878) );
  NAND2_X1 U4864 ( .A1(n6303), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3875)
         );
  NAND2_X1 U4865 ( .A1(n4074), .A2(n3875), .ZN(n3876) );
  AOI21_X1 U4866 ( .B1(n4082), .B2(EAX_REG_21__SCAN_IN), .A(n3876), .ZN(n3877)
         );
  OAI21_X1 U4867 ( .B1(n4052), .B2(n3878), .A(n3877), .ZN(n3882) );
  OR2_X1 U4868 ( .A1(n3879), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3880)
         );
  NAND2_X1 U4869 ( .A1(n3896), .A2(n3880), .ZN(n5672) );
  NAND2_X1 U4870 ( .A1(n3882), .A2(n3881), .ZN(n5284) );
  INV_X1 U4871 ( .A(n5278), .ZN(n3900) );
  AOI22_X1 U4872 ( .A1(n4043), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4873 ( .A1(n4036), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4037), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4874 ( .A1(n4000), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4875 ( .A1(n3932), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3883) );
  NAND4_X1 U4876 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3892)
         );
  AOI22_X1 U4877 ( .A1(n3380), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4878 ( .A1(n3159), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4879 ( .A1(n4019), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4880 ( .A1(n3182), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3887) );
  NAND4_X1 U4881 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3891)
         );
  NOR2_X1 U4882 ( .A1(n3892), .A2(n3891), .ZN(n3895) );
  OAI21_X1 U4883 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5424), .A(n4074), .ZN(
        n3893) );
  AOI21_X1 U4884 ( .B1(n4082), .B2(EAX_REG_22__SCAN_IN), .A(n3893), .ZN(n3894)
         );
  OAI21_X1 U4885 ( .B1(n4052), .B2(n3895), .A(n3894), .ZN(n3898) );
  XNOR2_X1 U4886 ( .A(n3896), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5663)
         );
  NAND2_X1 U4887 ( .A1(n5663), .A2(n4077), .ZN(n3897) );
  NAND2_X1 U4888 ( .A1(n3898), .A2(n3897), .ZN(n5280) );
  AOI22_X1 U4889 ( .A1(n4036), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4890 ( .A1(n3401), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4891 ( .A1(n4037), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4892 ( .A1(n4038), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3902) );
  NAND4_X1 U4893 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3911)
         );
  AOI22_X1 U4894 ( .A1(n4043), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4895 ( .A1(n4000), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4896 ( .A1(n4018), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4897 ( .A1(n4055), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3906) );
  NAND4_X1 U4898 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(n3910)
         );
  OR2_X1 U4899 ( .A1(n3911), .A2(n3910), .ZN(n3924) );
  AOI22_X1 U4900 ( .A1(n4036), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4901 ( .A1(n3401), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4902 ( .A1(n4037), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4903 ( .A1(n4038), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3912) );
  NAND4_X1 U4904 ( .A1(n3915), .A2(n3914), .A3(n3913), .A4(n3912), .ZN(n3921)
         );
  AOI22_X1 U4905 ( .A1(n4043), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3919) );
  INV_X1 U4906 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6701) );
  AOI22_X1 U4907 ( .A1(n4000), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4908 ( .A1(n4018), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4909 ( .A1(n4055), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3916) );
  NAND4_X1 U4910 ( .A1(n3919), .A2(n3918), .A3(n3917), .A4(n3916), .ZN(n3920)
         );
  OR2_X1 U4911 ( .A1(n3921), .A2(n3920), .ZN(n3923) );
  INV_X1 U4912 ( .A(n3962), .ZN(n3922) );
  OAI21_X1 U4913 ( .B1(n3924), .B2(n3923), .A(n3922), .ZN(n3927) );
  OAI21_X1 U4914 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4095), .A(n4074), .ZN(
        n3925) );
  AOI21_X1 U4915 ( .B1(n4082), .B2(EAX_REG_23__SCAN_IN), .A(n3925), .ZN(n3926)
         );
  OAI21_X1 U4916 ( .B1(n4052), .B2(n3927), .A(n3926), .ZN(n3931) );
  AND2_X1 U4917 ( .A1(n3928), .A2(n4095), .ZN(n3929) );
  OR2_X1 U4918 ( .A1(n3929), .A2(n3947), .ZN(n5652) );
  NAND2_X1 U4919 ( .A1(n4097), .A2(n4077), .ZN(n3930) );
  NAND2_X1 U4920 ( .A1(n3931), .A2(n3930), .ZN(n4093) );
  AOI22_X1 U4921 ( .A1(n4036), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4922 ( .A1(n3401), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4923 ( .A1(n4037), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4924 ( .A1(n4038), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3933) );
  NAND4_X1 U4925 ( .A1(n3936), .A2(n3935), .A3(n3934), .A4(n3933), .ZN(n3944)
         );
  AOI22_X1 U4926 ( .A1(n4043), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4927 ( .A1(n4000), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4928 ( .A1(n3182), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4929 ( .A1(n4055), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3939) );
  NAND4_X1 U4930 ( .A1(n3942), .A2(n3941), .A3(n3940), .A4(n3939), .ZN(n3943)
         );
  OR2_X1 U4931 ( .A1(n3944), .A2(n3943), .ZN(n3963) );
  INV_X1 U4932 ( .A(n3963), .ZN(n3945) );
  XNOR2_X1 U4933 ( .A(n3962), .B(n3945), .ZN(n3946) );
  NAND2_X1 U4934 ( .A1(n4071), .A2(n3946), .ZN(n3951) );
  AOI22_X1 U4935 ( .A1(n4082), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4081), .ZN(n3949) );
  XNOR2_X1 U4936 ( .A(n3947), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5414)
         );
  NAND2_X1 U4937 ( .A1(n5414), .A2(n4077), .ZN(n3948) );
  NAND2_X1 U4938 ( .A1(n3951), .A2(n3950), .ZN(n5166) );
  AOI22_X1 U4939 ( .A1(n4036), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4940 ( .A1(n4000), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4941 ( .A1(n3401), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4942 ( .A1(n4043), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3952) );
  NAND4_X1 U4943 ( .A1(n3955), .A2(n3954), .A3(n3953), .A4(n3952), .ZN(n3961)
         );
  AOI22_X1 U4944 ( .A1(n3937), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4037), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4945 ( .A1(n4018), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4946 ( .A1(n3028), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4947 ( .A1(n4055), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3956) );
  NAND4_X1 U4948 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3960)
         );
  OR2_X1 U4949 ( .A1(n3961), .A2(n3960), .ZN(n3973) );
  NAND2_X1 U4950 ( .A1(n3963), .A2(n3962), .ZN(n3975) );
  XNOR2_X1 U4951 ( .A(n3973), .B(n3975), .ZN(n3964) );
  NAND2_X1 U4952 ( .A1(n4071), .A2(n3964), .ZN(n3971) );
  NAND2_X1 U4953 ( .A1(n6303), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3965)
         );
  NAND2_X1 U4954 ( .A1(n4074), .A2(n3965), .ZN(n3966) );
  AOI21_X1 U4955 ( .B1(n4082), .B2(EAX_REG_25__SCAN_IN), .A(n3966), .ZN(n3970)
         );
  OR2_X1 U4956 ( .A1(n3967), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3968)
         );
  NAND2_X1 U4957 ( .A1(n3972), .A2(n3968), .ZN(n5640) );
  NOR2_X1 U4958 ( .A1(n5640), .A2(n4074), .ZN(n3969) );
  AOI21_X1 U4959 ( .B1(n3971), .B2(n3970), .A(n3969), .ZN(n5266) );
  XNOR2_X1 U4960 ( .A(n3972), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5629)
         );
  INV_X1 U4961 ( .A(n3973), .ZN(n3974) );
  AOI22_X1 U4962 ( .A1(n3181), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4963 ( .A1(n4018), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4964 ( .A1(n4000), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4965 ( .A1(n4038), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U4966 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3985)
         );
  AOI22_X1 U4967 ( .A1(n4036), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4968 ( .A1(n3401), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4969 ( .A1(n4037), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4970 ( .A1(n4013), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3980) );
  NAND4_X1 U4971 ( .A1(n3983), .A2(n3982), .A3(n3981), .A4(n3980), .ZN(n3984)
         );
  NOR2_X1 U4972 ( .A1(n3985), .A2(n3984), .ZN(n3995) );
  XOR2_X1 U4973 ( .A(n3994), .B(n3995), .Z(n3989) );
  NAND2_X1 U4974 ( .A1(n4082), .A2(EAX_REG_26__SCAN_IN), .ZN(n3986) );
  OAI211_X1 U4975 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n3987), .A(n3986), .B(
        n4074), .ZN(n3988) );
  AOI21_X1 U4976 ( .B1(n3989), .B2(n4071), .A(n3988), .ZN(n3990) );
  AOI21_X1 U4977 ( .B1(n4077), .B2(n5629), .A(n3990), .ZN(n5261) );
  NAND2_X1 U4978 ( .A1(n3992), .A2(n3991), .ZN(n3993) );
  NAND2_X1 U4979 ( .A1(n4028), .A2(n3993), .ZN(n5387) );
  NOR2_X1 U4980 ( .A1(n3995), .A2(n3994), .ZN(n4012) );
  AOI22_X1 U4981 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4036), .B1(n4019), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4982 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3401), .B1(n3932), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4983 ( .A1(n4037), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4984 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4038), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3996) );
  NAND4_X1 U4985 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(n4006)
         );
  AOI22_X1 U4986 ( .A1(n3181), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4987 ( .A1(n4000), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4988 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3182), .B1(n3241), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4989 ( .A1(n4055), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U4990 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4005)
         );
  OR2_X1 U4991 ( .A1(n4006), .A2(n4005), .ZN(n4011) );
  XNOR2_X1 U4992 ( .A(n4012), .B(n4011), .ZN(n4009) );
  AOI21_X1 U4993 ( .B1(PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6303), .A(n4077), 
        .ZN(n4008) );
  NAND2_X1 U4994 ( .A1(n4082), .A2(EAX_REG_27__SCAN_IN), .ZN(n4007) );
  OAI211_X1 U4995 ( .C1(n4009), .C2(n4052), .A(n4008), .B(n4007), .ZN(n4010)
         );
  OAI21_X1 U4996 ( .B1(n4074), .B2(n5387), .A(n4010), .ZN(n5156) );
  NAND2_X1 U4997 ( .A1(n4012), .A2(n4011), .ZN(n4034) );
  AOI22_X1 U4998 ( .A1(n3937), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4999 ( .A1(n4037), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U5000 ( .A1(n4038), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U5001 ( .A1(n3159), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U5002 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4025)
         );
  AOI22_X1 U5003 ( .A1(n4018), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4043), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U5004 ( .A1(n4036), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4019), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U5005 ( .A1(n3401), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U5006 ( .A1(n4000), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4020) );
  NAND4_X1 U5007 ( .A1(n4023), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(n4024)
         );
  NOR2_X1 U5008 ( .A1(n4025), .A2(n4024), .ZN(n4035) );
  XOR2_X1 U5009 ( .A(n4034), .B(n4035), .Z(n4026) );
  NAND2_X1 U5010 ( .A1(n4026), .A2(n4071), .ZN(n4030) );
  AOI21_X1 U5011 ( .B1(n5147), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4027) );
  AOI21_X1 U5012 ( .B1(n4082), .B2(EAX_REG_28__SCAN_IN), .A(n4027), .ZN(n4029)
         );
  XNOR2_X1 U5013 ( .A(n4028), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5146)
         );
  AOI22_X1 U5014 ( .A1(n4030), .A2(n4029), .B1(n4077), .B2(n5146), .ZN(n5143)
         );
  INV_X1 U5015 ( .A(n4031), .ZN(n4032) );
  INV_X1 U5016 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U5017 ( .A1(n4032), .A2(n5134), .ZN(n4033) );
  NAND2_X1 U5018 ( .A1(n4076), .A2(n4033), .ZN(n5365) );
  NOR2_X1 U5019 ( .A1(n4035), .A2(n4034), .ZN(n4068) );
  AOI22_X1 U5020 ( .A1(n4036), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5021 ( .A1(n3380), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3932), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5022 ( .A1(n4037), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5023 ( .A1(n4038), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4039) );
  NAND4_X1 U5024 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4049)
         );
  AOI22_X1 U5025 ( .A1(n4043), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3937), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5026 ( .A1(n4000), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5027 ( .A1(n3182), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5028 ( .A1(n4055), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4044) );
  NAND4_X1 U5029 ( .A1(n4047), .A2(n4046), .A3(n4045), .A4(n4044), .ZN(n4048)
         );
  OR2_X1 U5030 ( .A1(n4049), .A2(n4048), .ZN(n4067) );
  XNOR2_X1 U5031 ( .A(n4068), .B(n4067), .ZN(n4053) );
  AOI21_X1 U5032 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6303), .A(n4077), 
        .ZN(n4051) );
  NAND2_X1 U5033 ( .A1(n4082), .A2(EAX_REG_29__SCAN_IN), .ZN(n4050) );
  OAI211_X1 U5034 ( .C1(n4053), .C2(n4052), .A(n4051), .B(n4050), .ZN(n4054)
         );
  OAI21_X1 U5035 ( .B1(n4074), .B2(n5365), .A(n4054), .ZN(n5127) );
  AOI22_X1 U5036 ( .A1(n3182), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5037 ( .A1(n4036), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4037), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5038 ( .A1(n3380), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4038), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5039 ( .A1(n4055), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4056) );
  NAND4_X1 U5040 ( .A1(n4059), .A2(n4058), .A3(n4057), .A4(n4056), .ZN(n4066)
         );
  AOI22_X1 U5041 ( .A1(n4000), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3159), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5042 ( .A1(n3937), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5043 ( .A1(n3932), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3901), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5044 ( .A1(n3028), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4060), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4061) );
  NAND4_X1 U5045 ( .A1(n4064), .A2(n4063), .A3(n4062), .A4(n4061), .ZN(n4065)
         );
  NOR2_X1 U5046 ( .A1(n4066), .A2(n4065), .ZN(n4070) );
  NAND2_X1 U5047 ( .A1(n4068), .A2(n4067), .ZN(n4069) );
  XOR2_X1 U5048 ( .A(n4070), .B(n4069), .Z(n4072) );
  NAND2_X1 U5049 ( .A1(n4072), .A2(n4071), .ZN(n4080) );
  NAND2_X1 U5050 ( .A1(n6303), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4073)
         );
  NAND2_X1 U5051 ( .A1(n4074), .A2(n4073), .ZN(n4075) );
  AOI21_X1 U5052 ( .B1(n4082), .B2(EAX_REG_30__SCAN_IN), .A(n4075), .ZN(n4079)
         );
  XNOR2_X1 U5053 ( .A(n4076), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5084)
         );
  AND2_X1 U5054 ( .A1(n5084), .A2(n4077), .ZN(n4078) );
  AOI21_X1 U5055 ( .B1(n4080), .B2(n4079), .A(n4078), .ZN(n4101) );
  AOI22_X1 U5056 ( .A1(n4082), .A2(EAX_REG_31__SCAN_IN), .B1(n4081), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4083) );
  AND2_X1 U5057 ( .A1(n6414), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4824) );
  NAND2_X1 U5058 ( .A1(n4824), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6425) );
  NAND2_X1 U5059 ( .A1(n5314), .A2(n5941), .ZN(n4084) );
  OAI211_X1 U5060 ( .C1(n5509), .C2(n5753), .A(n4084), .B(n4085), .ZN(U2955)
         );
  NOR2_X1 U5061 ( .A1(n5436), .A2(n5596), .ZN(n5442) );
  NAND2_X1 U5062 ( .A1(n4086), .A2(n4087), .ZN(n5434) );
  XNOR2_X1 U5063 ( .A(n5436), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5429)
         );
  INV_X1 U5064 ( .A(n5428), .ZN(n4091) );
  NOR2_X1 U5065 ( .A1(n5436), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5421)
         );
  NAND2_X1 U5066 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5419) );
  NOR3_X1 U5067 ( .A1(n4086), .A2(n4089), .A3(n5419), .ZN(n4090) );
  NAND2_X1 U5068 ( .A1(n5558), .A2(n5940), .ZN(n4100) );
  INV_X1 U5069 ( .A(n4094), .ZN(n5279) );
  NAND2_X1 U5070 ( .A1(n6000), .A2(REIP_REG_23__SCAN_IN), .ZN(n5560) );
  OAI21_X1 U5071 ( .B1(n5492), .B2(n4095), .A(n5560), .ZN(n4096) );
  AOI21_X1 U5072 ( .B1(n4097), .B2(n5494), .A(n4096), .ZN(n4098) );
  NAND2_X1 U5073 ( .A1(n4100), .A2(n3089), .ZN(U2963) );
  NAND2_X1 U5074 ( .A1(n3022), .A2(n3208), .ZN(n4104) );
  MUX2_X1 U5075 ( .A(n4104), .B(n6531), .S(n3210), .Z(n4260) );
  INV_X1 U5076 ( .A(n4260), .ZN(n4105) );
  NOR2_X1 U5077 ( .A1(n4105), .A2(n4242), .ZN(n4106) );
  NOR2_X1 U5078 ( .A1(n4385), .A2(n3189), .ZN(n4217) );
  OR2_X1 U5079 ( .A1(n4107), .A2(n3224), .ZN(n4309) );
  AND2_X1 U5080 ( .A1(n4217), .A2(n4309), .ZN(n4108) );
  NAND2_X1 U5081 ( .A1(n4218), .A2(n4108), .ZN(n4510) );
  NAND2_X1 U5082 ( .A1(n5743), .A2(n6396), .ZN(n4112) );
  INV_X1 U5083 ( .A(n3216), .ZN(n4110) );
  NOR2_X1 U5084 ( .A1(n3209), .A2(n3280), .ZN(n4563) );
  NAND4_X1 U5085 ( .A1(n4110), .A2(n4109), .A3(n4328), .A4(n4563), .ZN(n4111)
         );
  INV_X1 U5086 ( .A(n5312), .ZN(n4114) );
  NAND2_X1 U5087 ( .A1(n5115), .A2(n4114), .ZN(n4213) );
  NAND2_X1 U5088 ( .A1(n4163), .A2(n6012), .ZN(n4119) );
  INV_X1 U5089 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4117) );
  NAND2_X1 U5090 ( .A1(n4328), .A2(n4117), .ZN(n4118) );
  NAND3_X1 U5091 ( .A1(n4119), .A2(n4251), .A3(n4118), .ZN(n4121) );
  OR2_X1 U5092 ( .A1(n4251), .A2(EBX_REG_1__SCAN_IN), .ZN(n4120) );
  NAND2_X1 U5093 ( .A1(n4121), .A2(n4120), .ZN(n4124) );
  NAND2_X1 U5094 ( .A1(n4163), .A2(EBX_REG_0__SCAN_IN), .ZN(n4123) );
  INV_X1 U5095 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4407) );
  NAND2_X1 U5096 ( .A1(n4251), .A2(n4407), .ZN(n4122) );
  NAND2_X1 U5097 ( .A1(n4123), .A2(n4122), .ZN(n4398) );
  XNOR2_X1 U5098 ( .A(n4124), .B(n4398), .ZN(n4327) );
  NAND2_X1 U5099 ( .A1(n4327), .A2(n4328), .ZN(n4330) );
  INV_X1 U5100 ( .A(n4124), .ZN(n4125) );
  NAND2_X1 U5101 ( .A1(n4125), .A2(n4398), .ZN(n4126) );
  NAND2_X1 U5102 ( .A1(n4330), .A2(n4126), .ZN(n4445) );
  NAND2_X2 U5103 ( .A1(n4163), .A2(n4251), .ZN(n5101) );
  MUX2_X1 U5104 ( .A(n4197), .B(n4251), .S(EBX_REG_3__SCAN_IN), .Z(n4127) );
  OAI21_X1 U5105 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n5101), .A(n4127), 
        .ZN(n4128) );
  INV_X1 U5106 ( .A(n4128), .ZN(n4453) );
  MUX2_X1 U5107 ( .A(n4251), .B(n4163), .S(EBX_REG_2__SCAN_IN), .Z(n4130) );
  NAND2_X1 U5108 ( .A1(n5100), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4129)
         );
  NAND2_X1 U5109 ( .A1(n4130), .A2(n4129), .ZN(n4454) );
  NAND2_X1 U5110 ( .A1(n4453), .A2(n4454), .ZN(n4131) );
  NAND2_X1 U5111 ( .A1(n4163), .A2(n5999), .ZN(n4133) );
  INV_X1 U5112 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U5113 ( .A1(n4328), .A2(n5830), .ZN(n4132) );
  NAND3_X1 U5114 ( .A1(n4133), .A2(n4251), .A3(n4132), .ZN(n4135) );
  NAND2_X1 U5115 ( .A1(n5296), .A2(n5830), .ZN(n4134) );
  NAND2_X1 U5116 ( .A1(n4135), .A2(n4134), .ZN(n4450) );
  MUX2_X1 U5117 ( .A(n4197), .B(n4251), .S(EBX_REG_5__SCAN_IN), .Z(n4136) );
  OAI21_X1 U5118 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5101), .A(n4136), 
        .ZN(n4550) );
  MUX2_X1 U5119 ( .A(n4251), .B(n4163), .S(EBX_REG_6__SCAN_IN), .Z(n4140) );
  NAND2_X1 U5120 ( .A1(n5100), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4139)
         );
  AND2_X1 U5121 ( .A1(n4140), .A2(n4139), .ZN(n4464) );
  OR2_X2 U5122 ( .A1(n4551), .A2(n4464), .ZN(n4561) );
  MUX2_X1 U5123 ( .A(n4197), .B(n4251), .S(EBX_REG_7__SCAN_IN), .Z(n4141) );
  OAI21_X1 U5124 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5101), .A(n4141), 
        .ZN(n4559) );
  NOR2_X1 U5125 ( .A1(n4561), .A2(n4559), .ZN(n4657) );
  NAND2_X1 U5126 ( .A1(n4163), .A2(n5973), .ZN(n4143) );
  INV_X1 U5127 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4905) );
  NAND2_X1 U5128 ( .A1(n4328), .A2(n4905), .ZN(n4142) );
  NAND3_X1 U5129 ( .A1(n4143), .A2(n4251), .A3(n4142), .ZN(n4145) );
  NAND2_X1 U5130 ( .A1(n5296), .A2(n4905), .ZN(n4144) );
  NAND2_X1 U5131 ( .A1(n4145), .A2(n4144), .ZN(n4656) );
  NAND2_X1 U5132 ( .A1(n4657), .A2(n4656), .ZN(n4834) );
  MUX2_X1 U5133 ( .A(n4197), .B(n4251), .S(EBX_REG_9__SCAN_IN), .Z(n4146) );
  OAI21_X1 U5134 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5101), .A(n4146), 
        .ZN(n4835) );
  MUX2_X1 U5135 ( .A(n4251), .B(n4163), .S(EBX_REG_10__SCAN_IN), .Z(n4148) );
  NAND2_X1 U5136 ( .A1(n5100), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4147) );
  AND2_X1 U5137 ( .A1(n4148), .A2(n4147), .ZN(n4864) );
  INV_X1 U5138 ( .A(n4197), .ZN(n4166) );
  INV_X1 U5139 ( .A(EBX_REG_11__SCAN_IN), .ZN(n4150) );
  NAND2_X1 U5140 ( .A1(n4166), .A2(n4150), .ZN(n4153) );
  NAND2_X1 U5141 ( .A1(n4251), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4151) );
  OAI211_X1 U5142 ( .C1(n5100), .C2(EBX_REG_11__SCAN_IN), .A(n4163), .B(n4151), 
        .ZN(n4152) );
  NAND2_X1 U5143 ( .A1(n3038), .A2(n4902), .ZN(n5028) );
  MUX2_X1 U5144 ( .A(n4251), .B(n4163), .S(EBX_REG_12__SCAN_IN), .Z(n4155) );
  NAND2_X1 U5145 ( .A1(n5100), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4154) );
  NAND2_X1 U5146 ( .A1(n4155), .A2(n4154), .ZN(n4937) );
  INV_X1 U5147 ( .A(n4937), .ZN(n5027) );
  NAND2_X1 U5148 ( .A1(n4251), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4156) );
  OAI211_X1 U5149 ( .C1(n5100), .C2(EBX_REG_13__SCAN_IN), .A(n4163), .B(n4156), 
        .ZN(n4157) );
  OAI21_X1 U5150 ( .B1(n4197), .B2(EBX_REG_13__SCAN_IN), .A(n4157), .ZN(n5026)
         );
  MUX2_X1 U5151 ( .A(n4251), .B(n4163), .S(EBX_REG_14__SCAN_IN), .Z(n4161) );
  NAND2_X1 U5152 ( .A1(n5100), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4160) );
  NOR2_X2 U5153 ( .A1(n5237), .A2(n5236), .ZN(n5239) );
  INV_X1 U5154 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U5155 ( .A1(n4166), .A2(n5308), .ZN(n4165) );
  NAND2_X1 U5156 ( .A1(n4251), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4162) );
  OAI211_X1 U5157 ( .C1(n5100), .C2(EBX_REG_15__SCAN_IN), .A(n4163), .B(n4162), 
        .ZN(n4164) );
  INV_X1 U5158 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U5159 ( .A1(n4166), .A2(n5304), .ZN(n4169) );
  NAND2_X1 U5160 ( .A1(n4251), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4167) );
  OAI211_X1 U5161 ( .C1(n5100), .C2(EBX_REG_17__SCAN_IN), .A(n4163), .B(n4167), 
        .ZN(n4168) );
  AND2_X1 U5162 ( .A1(n4169), .A2(n4168), .ZN(n5205) );
  MUX2_X1 U5163 ( .A(n4251), .B(n4163), .S(EBX_REG_16__SCAN_IN), .Z(n4171) );
  NAND2_X1 U5164 ( .A1(n5100), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4170) );
  NAND2_X1 U5165 ( .A1(n4171), .A2(n4170), .ZN(n5219) );
  AND2_X1 U5166 ( .A1(n5205), .A2(n5219), .ZN(n4172) );
  NAND2_X1 U5167 ( .A1(n5221), .A2(n4172), .ZN(n5208) );
  NAND2_X1 U5168 ( .A1(n4163), .A2(n5596), .ZN(n4174) );
  INV_X1 U5169 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4175) );
  NAND2_X1 U5170 ( .A1(n4328), .A2(n4175), .ZN(n4173) );
  NAND3_X1 U5171 ( .A1(n4174), .A2(n4251), .A3(n4173), .ZN(n4177) );
  NAND2_X1 U5172 ( .A1(n5296), .A2(n4175), .ZN(n4176) );
  INV_X1 U5173 ( .A(n5101), .ZN(n4400) );
  NOR2_X1 U5174 ( .A1(n5100), .A2(EBX_REG_20__SCAN_IN), .ZN(n4178) );
  AOI21_X1 U5175 ( .B1(n4400), .B2(n5435), .A(n4178), .ZN(n5298) );
  OR2_X1 U5176 ( .A1(n5101), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4180)
         );
  INV_X1 U5177 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4179) );
  NAND2_X1 U5178 ( .A1(n4328), .A2(n4179), .ZN(n5180) );
  NAND2_X1 U5179 ( .A1(n4180), .A2(n5180), .ZN(n5293) );
  NAND2_X1 U5180 ( .A1(n5296), .A2(EBX_REG_20__SCAN_IN), .ZN(n4182) );
  NAND2_X1 U5181 ( .A1(n5293), .A2(n4251), .ZN(n4181) );
  OAI211_X1 U5182 ( .C1(n5298), .C2(n5293), .A(n4182), .B(n4181), .ZN(n4183)
         );
  NAND2_X1 U5183 ( .A1(n5294), .A2(n4184), .ZN(n5287) );
  MUX2_X1 U5184 ( .A(n4197), .B(n4251), .S(EBX_REG_21__SCAN_IN), .Z(n4185) );
  OAI21_X1 U5185 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5101), .A(n4185), 
        .ZN(n5286) );
  MUX2_X1 U5186 ( .A(n4197), .B(n4251), .S(EBX_REG_23__SCAN_IN), .Z(n4186) );
  OAI21_X1 U5187 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5101), .A(n4186), 
        .ZN(n5272) );
  MUX2_X1 U5188 ( .A(n4251), .B(n4163), .S(EBX_REG_22__SCAN_IN), .Z(n4188) );
  NAND2_X1 U5189 ( .A1(n5100), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4187) );
  NAND2_X1 U5190 ( .A1(n4188), .A2(n4187), .ZN(n5274) );
  INV_X1 U5191 ( .A(n5274), .ZN(n5281) );
  NOR2_X1 U5192 ( .A1(n5272), .A2(n5281), .ZN(n4189) );
  MUX2_X1 U5193 ( .A(n4251), .B(n4163), .S(EBX_REG_24__SCAN_IN), .Z(n4191) );
  NAND2_X1 U5194 ( .A1(n5100), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4190) );
  NAND2_X1 U5195 ( .A1(n4191), .A2(n4190), .ZN(n5171) );
  NAND2_X1 U5196 ( .A1(n5276), .A2(n5171), .ZN(n5170) );
  MUX2_X1 U5197 ( .A(n4197), .B(n4251), .S(EBX_REG_25__SCAN_IN), .Z(n4192) );
  OAI21_X1 U5198 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5101), .A(n4192), 
        .ZN(n5268) );
  OR2_X2 U5199 ( .A1(n5170), .A2(n5268), .ZN(n5270) );
  NAND2_X1 U5200 ( .A1(n4163), .A2(n5539), .ZN(n4194) );
  INV_X1 U5201 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U5202 ( .A1(n4328), .A2(n5639), .ZN(n4193) );
  NAND3_X1 U5203 ( .A1(n4194), .A2(n4251), .A3(n4193), .ZN(n4196) );
  NAND2_X1 U5204 ( .A1(n5296), .A2(n5639), .ZN(n4195) );
  MUX2_X1 U5205 ( .A(n4197), .B(n4251), .S(EBX_REG_27__SCAN_IN), .Z(n4198) );
  OAI21_X1 U5206 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5101), .A(n4198), 
        .ZN(n4199) );
  INV_X1 U5207 ( .A(n4199), .ZN(n5158) );
  INV_X1 U5208 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U5209 ( .A1(n4163), .A2(n5370), .ZN(n4201) );
  INV_X1 U5210 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U5211 ( .A1(n4328), .A2(n5256), .ZN(n4200) );
  NAND3_X1 U5212 ( .A1(n4201), .A2(n4251), .A3(n4200), .ZN(n4203) );
  NAND2_X1 U5213 ( .A1(n5296), .A2(n5256), .ZN(n4202) );
  NAND2_X1 U5214 ( .A1(n4203), .A2(n4202), .ZN(n5144) );
  NAND2_X2 U5215 ( .A1(n5160), .A2(n5144), .ZN(n5102) );
  INV_X1 U5216 ( .A(n5102), .ZN(n4205) );
  OAI22_X1 U5217 ( .A1(n5101), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n5100), .ZN(n5131) );
  NOR2_X2 U5218 ( .A1(n5102), .A2(n5131), .ZN(n4206) );
  INV_X1 U5219 ( .A(n4206), .ZN(n5103) );
  AOI22_X1 U5220 ( .A1(n5101), .A2(EBX_REG_30__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5100), .ZN(n5105) );
  INV_X1 U5221 ( .A(n5105), .ZN(n4204) );
  NOR2_X1 U5222 ( .A1(n4206), .A2(n5296), .ZN(n5104) );
  AOI211_X1 U5223 ( .C1(n4205), .C2(n5103), .A(n4204), .B(n5104), .ZN(n4208)
         );
  AOI211_X1 U5224 ( .C1(n5296), .C2(n5102), .A(n5105), .B(n4206), .ZN(n4207)
         );
  NOR2_X1 U5225 ( .A1(n4208), .A2(n4207), .ZN(n5118) );
  INV_X1 U5226 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4209) );
  INV_X1 U5227 ( .A(n5510), .ZN(n5520) );
  NAND2_X1 U5228 ( .A1(n5743), .A2(n4217), .ZN(n4219) );
  NAND2_X1 U5229 ( .A1(n4219), .A2(n4218), .ZN(n4312) );
  INV_X1 U5230 ( .A(n4220), .ZN(n4221) );
  NAND2_X1 U5231 ( .A1(n4831), .A2(n6434), .ZN(n4230) );
  INV_X1 U5232 ( .A(n4222), .ZN(n4227) );
  NAND3_X1 U5233 ( .A1(n4225), .A2(n4224), .A3(n4223), .ZN(n4226) );
  NAND2_X1 U5234 ( .A1(n4227), .A2(n4226), .ZN(n4229) );
  NOR2_X1 U5235 ( .A1(n4293), .A2(READY_N), .ZN(n4305) );
  AND3_X1 U5236 ( .A1(n4230), .A2(n4305), .A3(n3224), .ZN(n4231) );
  OAI21_X1 U5237 ( .B1(n4312), .B2(n4231), .A(n4566), .ZN(n4236) );
  NAND2_X1 U5238 ( .A1(n3189), .A2(n6434), .ZN(n4843) );
  NAND3_X1 U5239 ( .A1(n4232), .A2(n4843), .A3(n6528), .ZN(n4233) );
  NAND3_X1 U5240 ( .A1(n4233), .A2(n3208), .A3(n4571), .ZN(n4234) );
  NAND3_X1 U5241 ( .A1(n4409), .A2(n3279), .A3(n4234), .ZN(n4235) );
  INV_X1 U5242 ( .A(n6389), .ZN(n6400) );
  NAND2_X1 U5243 ( .A1(n4238), .A2(n4831), .ZN(n4307) );
  NAND2_X1 U5244 ( .A1(n4239), .A2(n3209), .ZN(n4240) );
  AND2_X1 U5245 ( .A1(n4307), .A2(n4240), .ZN(n4244) );
  INV_X1 U5246 ( .A(n4242), .ZN(n4243) );
  NAND2_X1 U5247 ( .A1(n4243), .A2(n5745), .ZN(n6388) );
  NAND4_X1 U5248 ( .A1(n6400), .A2(n4244), .A3(n3013), .A4(n6388), .ZN(n4245)
         );
  INV_X1 U5249 ( .A(n5118), .ZN(n4273) );
  NOR2_X1 U5250 ( .A1(n4247), .A2(n4246), .ZN(n4379) );
  NAND3_X1 U5251 ( .A1(n4379), .A2(n3206), .A3(n3281), .ZN(n4248) );
  NAND2_X1 U5252 ( .A1(n6407), .A2(n4248), .ZN(n4249) );
  AND2_X1 U5253 ( .A1(n6000), .A2(REIP_REG_30__SCAN_IN), .ZN(n5085) );
  AND2_X1 U5254 ( .A1(n4102), .A2(n4882), .ZN(n6373) );
  OR2_X1 U5255 ( .A1(n4252), .A2(n4251), .ZN(n4259) );
  AND2_X1 U5256 ( .A1(n4571), .A2(n3224), .ZN(n4253) );
  NOR2_X1 U5257 ( .A1(n4254), .A2(n4253), .ZN(n4258) );
  INV_X1 U5258 ( .A(n4309), .ZN(n4256) );
  INV_X1 U5259 ( .A(n3277), .ZN(n4255) );
  OAI21_X1 U5260 ( .B1(n4256), .B2(n5101), .A(n4255), .ZN(n4257) );
  AND4_X1 U5261 ( .A1(n4260), .A2(n4259), .A3(n4258), .A4(n4257), .ZN(n4261)
         );
  AND2_X1 U5262 ( .A1(n4262), .A2(n4261), .ZN(n4383) );
  OAI211_X1 U5263 ( .C1(n4250), .C2(n3208), .A(n4383), .B(n4514), .ZN(n4263)
         );
  NAND2_X1 U5264 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4264) );
  NOR2_X1 U5265 ( .A1(n5589), .A2(n4264), .ZN(n4269) );
  NAND2_X1 U5266 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5724) );
  NOR3_X1 U5267 ( .A1(n3499), .A2(n6577), .A3(n5724), .ZN(n5616) );
  AND2_X1 U5268 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5616), .ZN(n5712)
         );
  NAND2_X1 U5269 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5712), .ZN(n4268) );
  INV_X1 U5270 ( .A(n4268), .ZN(n5588) );
  NOR2_X1 U5271 ( .A1(n5978), .A2(n5973), .ZN(n5968) );
  INV_X1 U5272 ( .A(n5968), .ZN(n4926) );
  NAND2_X1 U5273 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4927) );
  NOR2_X1 U5274 ( .A1(n4926), .A2(n4927), .ZN(n4267) );
  NAND2_X1 U5275 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U5276 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5983) );
  NOR4_X1 U5277 ( .A1(n4265), .A2(n4607), .A3(n5995), .A4(n5983), .ZN(n4928)
         );
  NAND2_X1 U5278 ( .A1(n4267), .A2(n4928), .ZN(n5055) );
  INV_X1 U5279 ( .A(n5055), .ZN(n5725) );
  NAND2_X1 U5280 ( .A1(n5588), .A2(n5725), .ZN(n5584) );
  INV_X1 U5281 ( .A(n5584), .ZN(n4266) );
  NAND2_X1 U5282 ( .A1(n4269), .A2(n4266), .ZN(n4282) );
  AOI21_X1 U5283 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6011) );
  NOR2_X1 U5284 ( .A1(n6011), .A2(n5995), .ZN(n5980) );
  NAND2_X1 U5285 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5980), .ZN(n4606)
         );
  NOR2_X1 U5286 ( .A1(n4607), .A2(n4606), .ZN(n4929) );
  NAND2_X1 U5287 ( .A1(n4929), .A2(n4267), .ZN(n5720) );
  NOR2_X1 U5288 ( .A1(n5720), .A2(n4268), .ZN(n5581) );
  NAND2_X1 U5289 ( .A1(n5581), .A2(n4269), .ZN(n4279) );
  OR2_X1 U5290 ( .A1(n5721), .A2(n4279), .ZN(n4270) );
  AND2_X1 U5291 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4275) );
  NAND2_X1 U5292 ( .A1(n5571), .A2(n4275), .ZN(n5559) );
  NOR2_X1 U5293 ( .A1(n5559), .A2(n4286), .ZN(n5547) );
  AND2_X1 U5294 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U5295 ( .A1(n5547), .A2(n5538), .ZN(n5528) );
  NOR4_X1 U5296 ( .A1(n5528), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5510), 
        .A4(n3515), .ZN(n4272) );
  AOI211_X1 U5297 ( .C1(n4273), .C2(n6010), .A(n5085), .B(n4272), .ZN(n4274)
         );
  INV_X1 U5298 ( .A(n4275), .ZN(n4276) );
  NAND2_X1 U5299 ( .A1(n5571), .A2(n4276), .ZN(n4285) );
  INV_X1 U5300 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U5301 ( .A1(n5719), .A2(n6504), .ZN(n4278) );
  OR2_X1 U5302 ( .A1(n4277), .A2(n6000), .ZN(n4431) );
  NAND2_X1 U5303 ( .A1(n4278), .A2(n4431), .ZN(n5582) );
  INV_X1 U5304 ( .A(n4279), .ZN(n4280) );
  NOR2_X1 U5305 ( .A1(n5721), .A2(n4280), .ZN(n4281) );
  NOR2_X1 U5306 ( .A1(n5582), .A2(n4281), .ZN(n4284) );
  NAND2_X1 U5307 ( .A1(n5586), .A2(n4282), .ZN(n4283) );
  OAI21_X1 U5308 ( .B1(n5059), .B2(n6016), .A(n4286), .ZN(n4287) );
  NAND2_X1 U5309 ( .A1(n5566), .A2(n4287), .ZN(n5555) );
  INV_X1 U5310 ( .A(n5538), .ZN(n4288) );
  AOI21_X1 U5311 ( .B1(n4605), .B2(n4288), .A(n5555), .ZN(n5529) );
  OAI211_X1 U5312 ( .C1(n5520), .C2(n5615), .A(n5529), .B(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5515) );
  OAI211_X1 U5313 ( .C1(n5555), .C2(n4605), .A(n5515), .B(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4289) );
  OAI21_X1 U5314 ( .B1(n5089), .B2(n5623), .A(n4292), .ZN(U2988) );
  NAND2_X1 U5315 ( .A1(n4409), .A2(n4238), .ZN(n5093) );
  INV_X1 U5316 ( .A(n6526), .ZN(n4296) );
  OR2_X1 U5317 ( .A1(n3092), .A2(n4882), .ZN(n5751) );
  NAND2_X1 U5318 ( .A1(n6317), .A2(n4826), .ZN(n5091) );
  INV_X1 U5319 ( .A(n5091), .ZN(n4294) );
  OAI21_X1 U5320 ( .B1(READREQUEST_REG_SCAN_IN), .B2(n4294), .A(n4296), .ZN(
        n4295) );
  OAI21_X1 U5321 ( .B1(n4296), .B2(n5751), .A(n4295), .ZN(U3474) );
  INV_X1 U5322 ( .A(n6407), .ZN(n4297) );
  NAND2_X1 U5323 ( .A1(n4409), .A2(n4298), .ZN(n4299) );
  NAND2_X1 U5324 ( .A1(n5905), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4300) );
  INV_X1 U5325 ( .A(DATAI_0_), .ZN(n4611) );
  OR2_X1 U5326 ( .A1(n4570), .A2(n4611), .ZN(n4302) );
  OAI211_X1 U5327 ( .C1(n5908), .C2(n4301), .A(n4300), .B(n4302), .ZN(U2924)
         );
  INV_X1 U5328 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4304) );
  NAND2_X1 U5329 ( .A1(n5905), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4303) );
  OAI211_X1 U5330 ( .C1(n5908), .C2(n4304), .A(n4303), .B(n4302), .ZN(U2939)
         );
  INV_X1 U5331 ( .A(n4305), .ZN(n4306) );
  OAI22_X1 U5332 ( .A1(n5743), .A2(n6388), .B1(n4306), .B2(n3013), .ZN(n4568)
         );
  AOI21_X1 U5333 ( .B1(n4307), .B2(n6434), .A(READY_N), .ZN(n4308) );
  OAI21_X1 U5334 ( .B1(n6373), .B2(n4232), .A(n4308), .ZN(n4310) );
  OAI21_X1 U5335 ( .B1(n5743), .B2(n4310), .A(n4309), .ZN(n4311) );
  NOR2_X1 U5336 ( .A1(n6414), .A2(n4544), .ZN(n4541) );
  AOI22_X1 U5337 ( .A1(n6375), .A2(n4566), .B1(FLUSH_REG_SCAN_IN), .B2(n4541), 
        .ZN(n4318) );
  INV_X1 U5338 ( .A(n6059), .ZN(n4313) );
  OR2_X1 U5339 ( .A1(n4314), .A2(n4313), .ZN(n4315) );
  XNOR2_X1 U5340 ( .A(n4315), .B(n4538), .ZN(n4537) );
  INV_X1 U5341 ( .A(n4537), .ZN(n5814) );
  INV_X1 U5342 ( .A(n6510), .ZN(n5045) );
  INV_X1 U5343 ( .A(n3013), .ZN(n4316) );
  NAND3_X1 U5344 ( .A1(n5814), .A2(n5045), .A3(n4316), .ZN(n4317) );
  OAI21_X1 U5345 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6501), .A(n4318), .ZN(
        n6508) );
  OAI22_X1 U5346 ( .A1(n4318), .A2(n4317), .B1(n4538), .B2(n6508), .ZN(U3455)
         );
  INV_X1 U5347 ( .A(EAX_REG_2__SCAN_IN), .ZN(n4320) );
  NAND2_X1 U5348 ( .A1(n5906), .A2(DATAI_2_), .ZN(n4322) );
  NAND2_X1 U5349 ( .A1(n5905), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4319) );
  OAI211_X1 U5350 ( .C1(n5908), .C2(n4320), .A(n4322), .B(n4319), .ZN(U2941)
         );
  INV_X1 U5351 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4323) );
  NAND2_X1 U5352 ( .A1(n5905), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4321) );
  OAI211_X1 U5353 ( .C1(n5908), .C2(n4323), .A(n4322), .B(n4321), .ZN(U2926)
         );
  NOR2_X1 U5354 ( .A1(n4325), .A2(n4324), .ZN(n4326) );
  OR2_X1 U5355 ( .A1(n4327), .A2(n4328), .ZN(n4329) );
  NAND2_X1 U5356 ( .A1(n4330), .A2(n4329), .ZN(n4435) );
  AOI22_X1 U5357 ( .A1(n5306), .A2(n4435), .B1(EBX_REG_1__SCAN_IN), .B2(n5305), 
        .ZN(n4331) );
  OAI21_X1 U5358 ( .B1(n5312), .B2(n5846), .A(n4331), .ZN(U2858) );
  INV_X1 U5359 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4333) );
  INV_X1 U5360 ( .A(DATAI_7_), .ZN(n4575) );
  NOR2_X1 U5361 ( .A1(n4570), .A2(n4575), .ZN(n4342) );
  AOI21_X1 U5362 ( .B1(n5902), .B2(EAX_REG_23__SCAN_IN), .A(n4342), .ZN(n4332)
         );
  OAI21_X1 U5363 ( .B1(n4377), .B2(n4333), .A(n4332), .ZN(U2931) );
  INV_X1 U5364 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n4335) );
  INV_X1 U5365 ( .A(DATAI_1_), .ZN(n4614) );
  NOR2_X1 U5366 ( .A1(n4570), .A2(n4614), .ZN(n4360) );
  AOI21_X1 U5367 ( .B1(n5902), .B2(EAX_REG_1__SCAN_IN), .A(n4360), .ZN(n4334)
         );
  OAI21_X1 U5368 ( .B1(n4377), .B2(n4335), .A(n4334), .ZN(U2940) );
  INV_X1 U5369 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n4337) );
  INV_X1 U5370 ( .A(DATAI_3_), .ZN(n4615) );
  NOR2_X1 U5371 ( .A1(n4570), .A2(n4615), .ZN(n4357) );
  AOI21_X1 U5372 ( .B1(n5902), .B2(EAX_REG_3__SCAN_IN), .A(n4357), .ZN(n4336)
         );
  OAI21_X1 U5373 ( .B1(n4377), .B2(n4337), .A(n4336), .ZN(U2942) );
  INV_X1 U5374 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n4339) );
  INV_X1 U5375 ( .A(DATAI_5_), .ZN(n4577) );
  NOR2_X1 U5376 ( .A1(n4570), .A2(n4577), .ZN(n4371) );
  AOI21_X1 U5377 ( .B1(n5902), .B2(EAX_REG_5__SCAN_IN), .A(n4371), .ZN(n4338)
         );
  OAI21_X1 U5378 ( .B1(n4377), .B2(n4339), .A(n4338), .ZN(U2944) );
  INV_X1 U5379 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n4341) );
  INV_X1 U5380 ( .A(DATAI_11_), .ZN(n4934) );
  NOR2_X1 U5381 ( .A1(n4570), .A2(n4934), .ZN(n4351) );
  AOI21_X1 U5382 ( .B1(n5902), .B2(EAX_REG_11__SCAN_IN), .A(n4351), .ZN(n4340)
         );
  OAI21_X1 U5383 ( .B1(n4377), .B2(n4341), .A(n4340), .ZN(U2950) );
  INV_X1 U5384 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n4344) );
  AOI21_X1 U5385 ( .B1(n5902), .B2(EAX_REG_7__SCAN_IN), .A(n4342), .ZN(n4343)
         );
  OAI21_X1 U5386 ( .B1(n4377), .B2(n4344), .A(n4343), .ZN(U2946) );
  INV_X1 U5387 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n4346) );
  INV_X1 U5388 ( .A(DATAI_13_), .ZN(n5038) );
  NOR2_X1 U5389 ( .A1(n4570), .A2(n5038), .ZN(n4354) );
  AOI21_X1 U5390 ( .B1(n5902), .B2(EAX_REG_13__SCAN_IN), .A(n4354), .ZN(n4345)
         );
  OAI21_X1 U5391 ( .B1(n4377), .B2(n4346), .A(n4345), .ZN(U2952) );
  INV_X1 U5392 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n4348) );
  INV_X1 U5393 ( .A(DATAI_8_), .ZN(n4664) );
  NOR2_X1 U5394 ( .A1(n4570), .A2(n4664), .ZN(n4365) );
  AOI21_X1 U5395 ( .B1(n5902), .B2(EAX_REG_8__SCAN_IN), .A(n4365), .ZN(n4347)
         );
  OAI21_X1 U5396 ( .B1(n4377), .B2(n4348), .A(n4347), .ZN(U2947) );
  INV_X1 U5397 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n4350) );
  INV_X1 U5398 ( .A(DATAI_4_), .ZN(n4613) );
  NOR2_X1 U5399 ( .A1(n4570), .A2(n4613), .ZN(n4368) );
  AOI21_X1 U5400 ( .B1(n5902), .B2(EAX_REG_4__SCAN_IN), .A(n4368), .ZN(n4349)
         );
  OAI21_X1 U5401 ( .B1(n4377), .B2(n4350), .A(n4349), .ZN(U2943) );
  INV_X1 U5402 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n4353) );
  AOI21_X1 U5403 ( .B1(n5902), .B2(EAX_REG_27__SCAN_IN), .A(n4351), .ZN(n4352)
         );
  OAI21_X1 U5404 ( .B1(n4377), .B2(n4353), .A(n4352), .ZN(U2935) );
  INV_X1 U5405 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n4356) );
  AOI21_X1 U5406 ( .B1(n5902), .B2(EAX_REG_29__SCAN_IN), .A(n4354), .ZN(n4355)
         );
  OAI21_X1 U5407 ( .B1(n4377), .B2(n4356), .A(n4355), .ZN(U2937) );
  INV_X1 U5408 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4359) );
  AOI21_X1 U5409 ( .B1(n5902), .B2(EAX_REG_19__SCAN_IN), .A(n4357), .ZN(n4358)
         );
  OAI21_X1 U5410 ( .B1(n4377), .B2(n4359), .A(n4358), .ZN(U2927) );
  INV_X1 U5411 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4362) );
  AOI21_X1 U5412 ( .B1(n5902), .B2(EAX_REG_17__SCAN_IN), .A(n4360), .ZN(n4361)
         );
  OAI21_X1 U5413 ( .B1(n4377), .B2(n4362), .A(n4361), .ZN(U2925) );
  INV_X1 U5414 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n4364) );
  INV_X1 U5415 ( .A(DATAI_6_), .ZN(n4617) );
  NOR2_X1 U5416 ( .A1(n4570), .A2(n4617), .ZN(n4374) );
  AOI21_X1 U5417 ( .B1(n5902), .B2(EAX_REG_6__SCAN_IN), .A(n4374), .ZN(n4363)
         );
  OAI21_X1 U5418 ( .B1(n4377), .B2(n4364), .A(n4363), .ZN(U2945) );
  INV_X1 U5419 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n4367) );
  AOI21_X1 U5420 ( .B1(n5902), .B2(EAX_REG_24__SCAN_IN), .A(n4365), .ZN(n4366)
         );
  OAI21_X1 U5421 ( .B1(n4377), .B2(n4367), .A(n4366), .ZN(U2932) );
  INV_X1 U5422 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n4370) );
  AOI21_X1 U5423 ( .B1(n5902), .B2(EAX_REG_20__SCAN_IN), .A(n4368), .ZN(n4369)
         );
  OAI21_X1 U5424 ( .B1(n4377), .B2(n4370), .A(n4369), .ZN(U2928) );
  INV_X1 U5425 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n4373) );
  AOI21_X1 U5426 ( .B1(n5902), .B2(EAX_REG_21__SCAN_IN), .A(n4371), .ZN(n4372)
         );
  OAI21_X1 U5427 ( .B1(n4377), .B2(n4373), .A(n4372), .ZN(U2929) );
  INV_X1 U5428 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n4376) );
  AOI21_X1 U5429 ( .B1(n5902), .B2(EAX_REG_22__SCAN_IN), .A(n4374), .ZN(n4375)
         );
  OAI21_X1 U5430 ( .B1(n4377), .B2(n4376), .A(n4375), .ZN(U2930) );
  INV_X1 U5431 ( .A(n4379), .ZN(n4565) );
  NAND2_X1 U5432 ( .A1(n4565), .A2(n4250), .ZN(n4380) );
  NOR2_X1 U5433 ( .A1(n4232), .A2(n4380), .ZN(n4381) );
  AND2_X1 U5434 ( .A1(n3013), .A2(n4381), .ZN(n4382) );
  INV_X1 U5435 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4384) );
  AND2_X1 U5436 ( .A1(n6373), .A2(n4384), .ZN(n4527) );
  INV_X1 U5437 ( .A(n4527), .ZN(n4389) );
  INV_X1 U5438 ( .A(n4385), .ZN(n6371) );
  INV_X1 U5439 ( .A(n3102), .ZN(n4387) );
  INV_X1 U5440 ( .A(n4386), .ZN(n5048) );
  NAND3_X1 U5441 ( .A1(n6371), .A2(n4387), .A3(n5048), .ZN(n4388) );
  OAI211_X1 U5442 ( .C1(n6120), .C2(n4532), .A(n4389), .B(n4388), .ZN(n6374)
         );
  NOR2_X1 U5443 ( .A1(n4826), .A2(n6504), .ZN(n5040) );
  AOI22_X1 U5444 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4390), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6012), .ZN(n5041) );
  AOI222_X1 U5445 ( .A1(n6374), .A2(n5045), .B1(n5040), .B2(n5041), .C1(n4391), 
        .C2(n5047), .ZN(n4393) );
  INV_X1 U5446 ( .A(n6508), .ZN(n6503) );
  INV_X1 U5447 ( .A(n5047), .ZN(n6412) );
  NOR2_X1 U5448 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6412), .ZN(n6502)
         );
  OAI21_X1 U5449 ( .B1(n6502), .B2(n6503), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n4392) );
  OAI21_X1 U5450 ( .B1(n4393), .B2(n6503), .A(n4392), .ZN(U3460) );
  XNOR2_X1 U5451 ( .A(n4394), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4473)
         );
  NOR2_X1 U5452 ( .A1(n6016), .A2(n5719), .ZN(n5727) );
  INV_X1 U5453 ( .A(n5727), .ZN(n4397) );
  INV_X1 U5454 ( .A(n5726), .ZN(n4395) );
  AOI21_X1 U5455 ( .B1(n4395), .B2(n4431), .A(n6504), .ZN(n4396) );
  AOI21_X1 U5456 ( .B1(n4397), .B2(n6504), .A(n4396), .ZN(n4402) );
  INV_X1 U5457 ( .A(n4398), .ZN(n4399) );
  AOI21_X1 U5458 ( .B1(n6504), .B2(n4400), .A(n4399), .ZN(n5250) );
  INV_X1 U5459 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6513) );
  NOR2_X1 U5460 ( .A1(n5819), .A2(n6513), .ZN(n4471) );
  AOI21_X1 U5461 ( .B1(n6010), .B2(n5250), .A(n4471), .ZN(n4401) );
  OAI211_X1 U5462 ( .C1(n4473), .C2(n5623), .A(n4402), .B(n4401), .ZN(U3018)
         );
  INV_X1 U5463 ( .A(n5250), .ZN(n4408) );
  INV_X1 U5464 ( .A(n4403), .ZN(n4404) );
  AOI21_X1 U5465 ( .B1(n4406), .B2(n4405), .A(n4404), .ZN(n5249) );
  INV_X1 U5466 ( .A(n5249), .ZN(n4612) );
  OAI222_X1 U5467 ( .A1(n4408), .A2(n5309), .B1(n4407), .B2(n5311), .C1(n4612), 
        .C2(n5312), .ZN(U2859) );
  INV_X1 U5468 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4413) );
  NAND2_X1 U5469 ( .A1(n4409), .A2(n6373), .ZN(n4410) );
  NAND2_X1 U5470 ( .A1(n5908), .A2(n4410), .ZN(n4411) );
  INV_X1 U5471 ( .A(n6434), .ZN(n4838) );
  NOR2_X4 U5472 ( .A1(n5871), .A2(n6529), .ZN(n5887) );
  AOI22_X1 U5473 ( .A1(n6529), .A2(UWORD_REG_7__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4412) );
  OAI21_X1 U5474 ( .B1(n4413), .B2(n5859), .A(n4412), .ZN(U2900) );
  INV_X1 U5475 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5892) );
  AOI22_X1 U5476 ( .A1(n6529), .A2(UWORD_REG_9__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4414) );
  OAI21_X1 U5477 ( .B1(n5892), .B2(n5859), .A(n4414), .ZN(U2898) );
  INV_X1 U5478 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4416) );
  AOI22_X1 U5479 ( .A1(n6529), .A2(UWORD_REG_8__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4415) );
  OAI21_X1 U5480 ( .B1(n4416), .B2(n5859), .A(n4415), .ZN(U2899) );
  AOI22_X1 U5481 ( .A1(n6529), .A2(UWORD_REG_0__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4417) );
  OAI21_X1 U5482 ( .B1(n4301), .B2(n5859), .A(n4417), .ZN(U2907) );
  INV_X1 U5483 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4419) );
  AOI22_X1 U5484 ( .A1(n6529), .A2(UWORD_REG_6__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4418) );
  OAI21_X1 U5485 ( .B1(n4419), .B2(n5859), .A(n4418), .ZN(U2901) );
  INV_X1 U5486 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4421) );
  AOI22_X1 U5487 ( .A1(n6529), .A2(UWORD_REG_5__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4420) );
  OAI21_X1 U5488 ( .B1(n4421), .B2(n5859), .A(n4420), .ZN(U2902) );
  INV_X1 U5489 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4423) );
  AOI22_X1 U5490 ( .A1(n6529), .A2(UWORD_REG_4__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4422) );
  OAI21_X1 U5491 ( .B1(n4423), .B2(n5859), .A(n4422), .ZN(U2903) );
  INV_X1 U5492 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4425) );
  AOI22_X1 U5493 ( .A1(n6529), .A2(UWORD_REG_3__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4424) );
  OAI21_X1 U5494 ( .B1(n4425), .B2(n5859), .A(n4424), .ZN(U2904) );
  AOI22_X1 U5495 ( .A1(n6529), .A2(UWORD_REG_2__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4426) );
  OAI21_X1 U5496 ( .B1(n4323), .B2(n5859), .A(n4426), .ZN(U2905) );
  INV_X1 U5497 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4428) );
  AOI22_X1 U5498 ( .A1(n6529), .A2(UWORD_REG_1__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4427) );
  OAI21_X1 U5499 ( .B1(n4428), .B2(n5859), .A(n4427), .ZN(U2906) );
  INV_X1 U5500 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4430) );
  AOI22_X1 U5501 ( .A1(n6529), .A2(UWORD_REG_10__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4429) );
  OAI21_X1 U5502 ( .B1(n4430), .B2(n5859), .A(n4429), .ZN(U2897) );
  OAI21_X1 U5503 ( .B1(n5727), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4431), 
        .ZN(n4439) );
  XNOR2_X1 U5504 ( .A(n4433), .B(n4432), .ZN(n4863) );
  NAND3_X1 U5505 ( .A1(n4605), .A2(n6012), .A3(n4434), .ZN(n4437) );
  AND2_X1 U5506 ( .A1(n6000), .A2(REIP_REG_1__SCAN_IN), .ZN(n4860) );
  AOI21_X1 U5507 ( .B1(n6010), .B2(n4435), .A(n4860), .ZN(n4436) );
  OAI211_X1 U5508 ( .C1(n4863), .C2(n5623), .A(n4437), .B(n4436), .ZN(n4438)
         );
  AOI21_X1 U5509 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n4439), .A(n4438), 
        .ZN(n4440) );
  INV_X1 U5510 ( .A(n4440), .ZN(U3017) );
  NOR2_X1 U5511 ( .A1(n4443), .A2(n4442), .ZN(n4444) );
  NOR2_X1 U5512 ( .A1(n4441), .A2(n4444), .ZN(n5942) );
  INV_X1 U5513 ( .A(n5942), .ZN(n4616) );
  XNOR2_X1 U5514 ( .A(n4445), .B(n4454), .ZN(n6009) );
  AOI22_X1 U5515 ( .A1(n5306), .A2(n6009), .B1(EBX_REG_2__SCAN_IN), .B2(n5305), 
        .ZN(n4446) );
  OAI21_X1 U5516 ( .B1(n4616), .B2(n5312), .A(n4446), .ZN(U2857) );
  AOI21_X1 U5517 ( .B1(n4441), .B2(n4457), .A(n4447), .ZN(n4448) );
  NOR2_X1 U5518 ( .A1(n4553), .A2(n4448), .ZN(n4896) );
  INV_X1 U5519 ( .A(n4896), .ZN(n5824) );
  OAI21_X1 U5520 ( .B1(n4449), .B2(n4450), .A(n4549), .ZN(n4451) );
  INV_X1 U5521 ( .A(n4451), .ZN(n5992) );
  AOI22_X1 U5522 ( .A1(n5306), .A2(n5992), .B1(EBX_REG_4__SCAN_IN), .B2(n5305), 
        .ZN(n4452) );
  OAI21_X1 U5523 ( .B1(n5824), .B2(n5312), .A(n4452), .ZN(U2855) );
  INV_X1 U5524 ( .A(n4445), .ZN(n4455) );
  AOI21_X1 U5525 ( .B1(n4455), .B2(n4454), .A(n4453), .ZN(n4456) );
  OR2_X1 U5526 ( .A1(n4456), .A2(n4449), .ZN(n4883) );
  INV_X1 U5527 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4458) );
  XNOR2_X1 U5528 ( .A(n4441), .B(n4457), .ZN(n5927) );
  OAI222_X1 U5529 ( .A1(n4883), .A2(n5309), .B1(n4458), .B2(n5311), .C1(n5927), 
        .C2(n5312), .ZN(U2856) );
  INV_X1 U5530 ( .A(n4459), .ZN(n4461) );
  NAND2_X1 U5531 ( .A1(n4553), .A2(n4552), .ZN(n4460) );
  NAND2_X1 U5532 ( .A1(n4461), .A2(n4460), .ZN(n4463) );
  AND2_X1 U5533 ( .A1(n4463), .A2(n4462), .ZN(n4877) );
  INV_X1 U5534 ( .A(n4877), .ZN(n4948) );
  INV_X1 U5535 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U5536 ( .A1(n4551), .A2(n4464), .ZN(n4465) );
  AND2_X1 U5537 ( .A1(n4561), .A2(n4465), .ZN(n4940) );
  INV_X1 U5538 ( .A(n4940), .ZN(n4466) );
  OAI222_X1 U5539 ( .A1(n4948), .A2(n5312), .B1(n5311), .B2(n4467), .C1(n4466), 
        .C2(n5309), .ZN(U2853) );
  OAI21_X1 U5540 ( .B1(n4468), .B2(n5936), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4469) );
  INV_X1 U5541 ( .A(n4469), .ZN(n4470) );
  AOI211_X1 U5542 ( .C1(n5249), .C2(n5941), .A(n4471), .B(n4470), .ZN(n4472)
         );
  OAI21_X1 U5543 ( .B1(n5753), .B2(n4473), .A(n4472), .ZN(U2986) );
  NAND3_X1 U5544 ( .A1(n6265), .A2(n6381), .A3(n4976), .ZN(n4672) );
  NOR2_X1 U5545 ( .A1(n4485), .A2(n6303), .ZN(n4623) );
  INV_X1 U5546 ( .A(n4618), .ZN(n4474) );
  NOR2_X1 U5547 ( .A1(n4474), .A2(n4974), .ZN(n4486) );
  OAI21_X1 U5548 ( .B1(n4486), .B2(n6303), .A(n4743), .ZN(n6065) );
  AOI211_X1 U5549 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4792), .A(n4623), .B(
        n6065), .ZN(n4484) );
  INV_X1 U5550 ( .A(n3033), .ZN(n4579) );
  NAND3_X1 U5551 ( .A1(n3590), .A2(n6028), .A3(n4579), .ZN(n4665) );
  NAND2_X1 U5552 ( .A1(n4476), .A2(n4478), .ZN(n6228) );
  OR2_X1 U5553 ( .A1(n6309), .A2(n4970), .ZN(n6358) );
  OAI21_X1 U5554 ( .B1(n4762), .B2(n6364), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4482) );
  NAND2_X1 U5555 ( .A1(n4481), .A2(n6120), .ZN(n4704) );
  NAND3_X1 U5556 ( .A1(n4482), .A2(n6317), .A3(n4666), .ZN(n4483) );
  NAND2_X1 U5557 ( .A1(n4786), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4491) );
  NAND2_X1 U5558 ( .A1(DATAI_5_), .A2(n4743), .ZN(n6248) );
  AND2_X1 U5559 ( .A1(n4485), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6264) );
  INV_X1 U5560 ( .A(n6264), .ZN(n6062) );
  INV_X1 U5561 ( .A(n4486), .ZN(n6057) );
  OAI22_X1 U5562 ( .A1(n4666), .A2(n6305), .B1(n6062), .B2(n6057), .ZN(n4789)
         );
  INV_X1 U5563 ( .A(n4762), .ZN(n4787) );
  INV_X1 U5564 ( .A(DATAI_21_), .ZN(n4487) );
  NOR2_X1 U5565 ( .A1(n5499), .A2(n4487), .ZN(n6245) );
  INV_X1 U5566 ( .A(DATAI_29_), .ZN(n4488) );
  INV_X1 U5567 ( .A(n6348), .ZN(n6080) );
  OAI22_X1 U5568 ( .A1(n4787), .A2(n6351), .B1(n6080), .B2(n6358), .ZN(n4489)
         );
  AOI21_X1 U5569 ( .B1(n6347), .B2(n4789), .A(n4489), .ZN(n4490) );
  OAI211_X1 U5570 ( .C1(n4792), .C2(n4718), .A(n4491), .B(n4490), .ZN(U3025)
         );
  INV_X1 U5571 ( .A(n6322), .ZN(n4730) );
  NAND2_X1 U5572 ( .A1(n4786), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U5573 ( .A1(DATAI_1_), .A2(n4743), .ZN(n6235) );
  INV_X1 U5574 ( .A(DATAI_17_), .ZN(n4492) );
  NOR2_X1 U5575 ( .A1(n5499), .A2(n4492), .ZN(n6232) );
  INV_X1 U5576 ( .A(n6232), .ZN(n6327) );
  INV_X1 U5577 ( .A(DATAI_25_), .ZN(n4493) );
  INV_X1 U5578 ( .A(n6324), .ZN(n6071) );
  OAI22_X1 U5579 ( .A1(n4787), .A2(n6327), .B1(n6071), .B2(n6358), .ZN(n4494)
         );
  AOI21_X1 U5580 ( .B1(n6323), .B2(n4789), .A(n4494), .ZN(n4495) );
  OAI211_X1 U5581 ( .C1(n4792), .C2(n4730), .A(n4496), .B(n4495), .ZN(U3021)
         );
  NAND2_X1 U5582 ( .A1(n4786), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4501) );
  NAND2_X1 U5583 ( .A1(DATAI_0_), .A2(n4743), .ZN(n6231) );
  INV_X1 U5584 ( .A(DATAI_16_), .ZN(n4497) );
  NOR2_X1 U5585 ( .A1(n5499), .A2(n4497), .ZN(n6318) );
  INV_X1 U5586 ( .A(n6318), .ZN(n6273) );
  INV_X1 U5587 ( .A(DATAI_24_), .ZN(n4498) );
  INV_X1 U5588 ( .A(n6270), .ZN(n6321) );
  OAI22_X1 U5589 ( .A1(n4787), .A2(n6273), .B1(n6321), .B2(n6358), .ZN(n4499)
         );
  AOI21_X1 U5590 ( .B1(n6308), .B2(n4789), .A(n4499), .ZN(n4500) );
  OAI211_X1 U5591 ( .C1(n4726), .C2(n4792), .A(n4501), .B(n4500), .ZN(U3020)
         );
  INV_X1 U5592 ( .A(n6334), .ZN(n4722) );
  NAND2_X1 U5593 ( .A1(n4786), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U5594 ( .A1(DATAI_3_), .A2(n4743), .ZN(n6241) );
  INV_X1 U5595 ( .A(DATAI_19_), .ZN(n4502) );
  NOR2_X1 U5596 ( .A1(n5499), .A2(n4502), .ZN(n6336) );
  INV_X1 U5597 ( .A(n6336), .ZN(n6283) );
  NAND2_X1 U5598 ( .A1(n5941), .A2(DATAI_27_), .ZN(n6339) );
  OAI22_X1 U5599 ( .A1(n4787), .A2(n6283), .B1(n6339), .B2(n6358), .ZN(n4503)
         );
  AOI21_X1 U5600 ( .B1(n6335), .B2(n4789), .A(n4503), .ZN(n4504) );
  OAI211_X1 U5601 ( .C1(n4792), .C2(n4722), .A(n4505), .B(n4504), .ZN(U3023)
         );
  INV_X1 U5602 ( .A(n6360), .ZN(n4714) );
  NAND2_X1 U5603 ( .A1(n4786), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4509) );
  NAND2_X1 U5604 ( .A1(DATAI_7_), .A2(n4743), .ZN(n6258) );
  INV_X1 U5605 ( .A(DATAI_23_), .ZN(n4506) );
  NOR2_X1 U5606 ( .A1(n5499), .A2(n4506), .ZN(n6365) );
  NAND2_X1 U5607 ( .A1(n5941), .A2(DATAI_31_), .ZN(n6370) );
  OAI22_X1 U5608 ( .A1(n4787), .A2(n6299), .B1(n6370), .B2(n6358), .ZN(n4507)
         );
  AOI21_X1 U5609 ( .B1(n6363), .B2(n4789), .A(n4507), .ZN(n4508) );
  OAI211_X1 U5610 ( .C1(n4792), .C2(n4714), .A(n4509), .B(n4508), .ZN(U3027)
         );
  INV_X1 U5611 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5754) );
  AND2_X1 U5612 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5754), .ZN(n4539) );
  INV_X1 U5613 ( .A(n4532), .ZN(n6372) );
  NAND2_X1 U5614 ( .A1(n4510), .A2(n6388), .ZN(n4525) );
  INV_X1 U5615 ( .A(n4525), .ZN(n4521) );
  NOR2_X1 U5616 ( .A1(n4386), .A2(n6645), .ZN(n4511) );
  XNOR2_X1 U5617 ( .A(n4511), .B(n4523), .ZN(n4520) );
  NAND2_X1 U5618 ( .A1(n6645), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4512) );
  INV_X1 U5619 ( .A(n4512), .ZN(n4513) );
  MUX2_X1 U5620 ( .A(n4513), .B(n4512), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4518) );
  INV_X1 U5621 ( .A(n4514), .ZN(n4526) );
  INV_X1 U5622 ( .A(n4515), .ZN(n4516) );
  OAI211_X1 U5623 ( .C1(n4386), .C2(n4523), .A(n4517), .B(n4516), .ZN(n5625)
         );
  AOI22_X1 U5624 ( .A1(n6373), .A2(n4518), .B1(n4526), .B2(n5625), .ZN(n4519)
         );
  OAI21_X1 U5625 ( .B1(n4521), .B2(n4520), .A(n4519), .ZN(n4522) );
  AOI21_X1 U5626 ( .B1(n3031), .B2(n6372), .A(n4522), .ZN(n5627) );
  MUX2_X1 U5627 ( .A(n4523), .B(n5627), .S(n6375), .Z(n6383) );
  MUX2_X1 U5628 ( .A(n4525), .B(n4526), .S(n4386), .Z(n4524) );
  AOI21_X1 U5629 ( .B1(n6373), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4524), 
        .ZN(n4530) );
  MUX2_X1 U5630 ( .A(n4526), .B(n4525), .S(n4386), .Z(n4528) );
  NOR2_X1 U5631 ( .A1(n4528), .A2(n4527), .ZN(n4529) );
  MUX2_X1 U5632 ( .A(n4530), .B(n4529), .S(n6645), .Z(n4531) );
  OAI21_X1 U5633 ( .B1(n4481), .B2(n4532), .A(n4531), .ZN(n5046) );
  INV_X1 U5634 ( .A(n5046), .ZN(n4533) );
  NAND2_X1 U5635 ( .A1(n6375), .A2(n4533), .ZN(n4534) );
  OAI21_X1 U5636 ( .B1(n6375), .B2(n6645), .A(n4534), .ZN(n6378) );
  NOR3_X1 U5637 ( .A1(n6383), .A2(STATE2_REG_1__SCAN_IN), .A3(n6378), .ZN(
        n4535) );
  AOI21_X1 U5638 ( .B1(n4536), .B2(n4539), .A(n4535), .ZN(n6403) );
  NOR2_X1 U5639 ( .A1(n6403), .A2(n3102), .ZN(n4545) );
  OAI22_X1 U5640 ( .A1(n6375), .A2(n4538), .B1(n4537), .B2(n3013), .ZN(n4540)
         );
  AOI22_X1 U5641 ( .A1(n4540), .A2(n4826), .B1(n4539), .B2(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6401) );
  INV_X1 U5642 ( .A(n6401), .ZN(n4543) );
  NOR3_X1 U5643 ( .A1(n4545), .A2(n4543), .A3(FLUSH_REG_SCAN_IN), .ZN(n4542)
         );
  INV_X1 U5644 ( .A(n4541), .ZN(n6499) );
  INV_X1 U5645 ( .A(n4743), .ZN(n4669) );
  NOR3_X1 U5646 ( .A1(n4545), .A2(n4544), .A3(n4543), .ZN(n6409) );
  INV_X1 U5647 ( .A(n3029), .ZN(n6149) );
  NAND2_X1 U5648 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6501), .ZN(n4636) );
  INV_X1 U5649 ( .A(n4636), .ZN(n4546) );
  OAI22_X1 U5650 ( .A1(n4970), .A2(n6305), .B1(n6149), .B2(n4546), .ZN(n4547)
         );
  OAI21_X1 U5651 ( .B1(n6409), .B2(n4547), .A(n6024), .ZN(n4548) );
  OAI21_X1 U5652 ( .B1(n6024), .B2(n6216), .A(n4548), .ZN(U3465) );
  OAI21_X1 U5653 ( .B1(n4138), .B2(n4137), .A(n4551), .ZN(n5981) );
  XOR2_X1 U5654 ( .A(n4553), .B(n4552), .Z(n5923) );
  INV_X1 U5655 ( .A(n5923), .ZN(n4578) );
  INV_X1 U5656 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4554) );
  OAI222_X1 U5657 ( .A1(n5981), .A2(n5309), .B1(n5312), .B2(n4578), .C1(n4554), 
        .C2(n5311), .ZN(U2854) );
  NAND2_X1 U5658 ( .A1(n4557), .A2(n4462), .ZN(n4558) );
  AND2_X1 U5659 ( .A1(n4556), .A2(n4558), .ZN(n5915) );
  INV_X1 U5660 ( .A(n5915), .ZN(n4576) );
  INV_X1 U5661 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4562) );
  INV_X1 U5662 ( .A(n4559), .ZN(n4560) );
  XNOR2_X1 U5663 ( .A(n4561), .B(n4560), .ZN(n5975) );
  INV_X1 U5664 ( .A(n5975), .ZN(n5795) );
  OAI222_X1 U5665 ( .A1(n4576), .A2(n5312), .B1(n4562), .B2(n5311), .C1(n5795), 
        .C2(n5309), .ZN(U2852) );
  NAND2_X1 U5666 ( .A1(n4563), .A2(n3205), .ZN(n4564) );
  NOR2_X1 U5667 ( .A1(n4565), .A2(n4564), .ZN(n4567) );
  AND2_X1 U5668 ( .A1(n3176), .A2(n3280), .ZN(n4574) );
  INV_X1 U5669 ( .A(n4574), .ZN(n4572) );
  OAI222_X1 U5670 ( .A1(n4576), .A2(n5361), .B1(n5359), .B2(n4575), .C1(n5357), 
        .C2(n3646), .ZN(U2884) );
  INV_X1 U5671 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5880) );
  OAI222_X1 U5672 ( .A1(n5361), .A2(n4578), .B1(n5357), .B2(n5880), .C1(n4577), 
        .C2(n5359), .ZN(U2886) );
  NAND3_X1 U5673 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6265), .A3(n6381), .ZN(n6034) );
  NOR2_X1 U5674 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6034), .ZN(n4583)
         );
  NOR2_X1 U5675 ( .A1(n4665), .A2(n4970), .ZN(n4763) );
  NOR2_X1 U5676 ( .A1(n4638), .A2(n4579), .ZN(n4580) );
  NAND2_X1 U5677 ( .A1(n6317), .A2(n5750), .ZN(n6310) );
  OAI21_X1 U5678 ( .B1(n4763), .B2(n6051), .A(n6310), .ZN(n4581) );
  NAND2_X1 U5679 ( .A1(n4481), .A2(n4378), .ZN(n4972) );
  AOI21_X1 U5680 ( .B1(n4581), .B2(n6030), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4582) );
  OAI21_X1 U5681 ( .B1(n4974), .B2(n6303), .A(n4743), .ZN(n6266) );
  NOR2_X1 U5682 ( .A1(n4623), .A2(n6266), .ZN(n4981) );
  NAND2_X1 U5683 ( .A1(n4796), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4586) );
  NAND2_X1 U5684 ( .A1(n4974), .A2(n6265), .ZN(n6122) );
  OAI22_X1 U5685 ( .A1(n6030), .A2(n6305), .B1(n6062), .B2(n6122), .ZN(n4800)
         );
  INV_X1 U5686 ( .A(n4763), .ZN(n4798) );
  OAI22_X1 U5687 ( .A1(n6370), .A2(n4798), .B1(n4797), .B2(n6299), .ZN(n4584)
         );
  AOI21_X1 U5688 ( .B1(n6363), .B2(n4800), .A(n4584), .ZN(n4585) );
  OAI211_X1 U5689 ( .C1(n4803), .C2(n4714), .A(n4586), .B(n4585), .ZN(U3043)
         );
  NAND2_X1 U5690 ( .A1(n4796), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4589) );
  OAI22_X1 U5691 ( .A1(n6080), .A2(n4798), .B1(n4797), .B2(n6351), .ZN(n4587)
         );
  AOI21_X1 U5692 ( .B1(n6347), .B2(n4800), .A(n4587), .ZN(n4588) );
  OAI211_X1 U5693 ( .C1(n4803), .C2(n4718), .A(n4589), .B(n4588), .ZN(U3041)
         );
  NAND2_X1 U5694 ( .A1(n4796), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4592) );
  OAI22_X1 U5695 ( .A1(n6339), .A2(n4798), .B1(n4797), .B2(n6283), .ZN(n4590)
         );
  AOI21_X1 U5696 ( .B1(n6335), .B2(n4800), .A(n4590), .ZN(n4591) );
  OAI211_X1 U5697 ( .C1(n4803), .C2(n4722), .A(n4592), .B(n4591), .ZN(U3039)
         );
  NAND2_X1 U5698 ( .A1(n4796), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4595) );
  OAI22_X1 U5699 ( .A1(n6071), .A2(n4798), .B1(n4797), .B2(n6327), .ZN(n4593)
         );
  AOI21_X1 U5700 ( .B1(n6323), .B2(n4800), .A(n4593), .ZN(n4594) );
  OAI211_X1 U5701 ( .C1(n4803), .C2(n4730), .A(n4595), .B(n4594), .ZN(U3037)
         );
  NAND2_X1 U5702 ( .A1(n4796), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4598) );
  OAI22_X1 U5703 ( .A1(n4798), .A2(n6321), .B1(n6273), .B2(n4797), .ZN(n4596)
         );
  AOI21_X1 U5704 ( .B1(n6308), .B2(n4800), .A(n4596), .ZN(n4597) );
  OAI211_X1 U5705 ( .C1(n4726), .C2(n4803), .A(n4598), .B(n4597), .ZN(U3036)
         );
  OAI21_X1 U5706 ( .B1(n4600), .B2(n4601), .A(n4603), .ZN(n4879) );
  AND2_X1 U5707 ( .A1(n6000), .A2(REIP_REG_6__SCAN_IN), .ZN(n4874) );
  AOI21_X1 U5709 ( .B1(n5586), .B2(n5983), .A(n5582), .ZN(n4604) );
  INV_X1 U5710 ( .A(n4604), .ZN(n6014) );
  AOI21_X1 U5711 ( .B1(n4606), .B2(n4605), .A(n6014), .ZN(n5989) );
  OAI21_X1 U5712 ( .B1(n5983), .B2(n6013), .A(n5721), .ZN(n4925) );
  INV_X1 U5713 ( .A(n4925), .ZN(n6002) );
  OAI33_X1 U5714 ( .A1(1'b0), .A2(n5989), .A3(n4607), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6002), .B3(n4606), .ZN(n4609) );
  AOI211_X1 U5715 ( .C1(n6010), .C2(n4940), .A(n4874), .B(n4609), .ZN(n4610)
         );
  OAI21_X1 U5716 ( .B1(n5623), .B2(n4879), .A(n4610), .ZN(U3012) );
  OAI222_X1 U5717 ( .A1(n4612), .A2(n5361), .B1(n5359), .B2(n4611), .C1(n5357), 
        .C2(n4304), .ZN(U2891) );
  INV_X1 U5718 ( .A(EAX_REG_4__SCAN_IN), .ZN(n5882) );
  OAI222_X1 U5719 ( .A1(n5824), .A2(n5361), .B1(n5359), .B2(n4613), .C1(n5357), 
        .C2(n5882), .ZN(U2887) );
  INV_X1 U5720 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5886) );
  OAI222_X1 U5721 ( .A1(n5846), .A2(n5361), .B1(n5359), .B2(n4614), .C1(n5357), 
        .C2(n5886), .ZN(U2890) );
  INV_X1 U5722 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6699) );
  OAI222_X1 U5723 ( .A1(n5927), .A2(n5361), .B1(n5359), .B2(n4615), .C1(n5357), 
        .C2(n6699), .ZN(U2888) );
  INV_X1 U5724 ( .A(DATAI_2_), .ZN(n6686) );
  OAI222_X1 U5725 ( .A1(n4616), .A2(n5361), .B1(n5359), .B2(n6686), .C1(n5357), 
        .C2(n4320), .ZN(U2889) );
  OAI222_X1 U5726 ( .A1(n4948), .A2(n5361), .B1(n5359), .B2(n4617), .C1(n5357), 
        .C2(n3639), .ZN(U2885) );
  OR2_X1 U5727 ( .A1(n4481), .A2(n4378), .ZN(n6218) );
  INV_X1 U5728 ( .A(n6218), .ZN(n4622) );
  AOI21_X1 U5729 ( .B1(n4622), .B2(n3031), .A(n6305), .ZN(n4621) );
  NAND2_X1 U5730 ( .A1(n3033), .A2(n6260), .ZN(n4703) );
  OAI21_X1 U5731 ( .B1(n6210), .B2(n6253), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4620) );
  NOR2_X1 U5732 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6381), .ZN(n6221)
         );
  NAND2_X1 U5733 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6221), .ZN(n6223) );
  NOR2_X1 U5734 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6223), .ZN(n4751)
         );
  OR2_X1 U5735 ( .A1(n4974), .A2(n4618), .ZN(n4709) );
  AOI21_X1 U5736 ( .B1(n4709), .B2(STATE2_REG_2__SCAN_IN), .A(n4669), .ZN(
        n4701) );
  OAI211_X1 U5737 ( .C1(n6501), .C2(n4751), .A(n6062), .B(n4701), .ZN(n4619)
         );
  INV_X1 U5738 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5739 ( .A1(n4622), .A2(n6317), .ZN(n6058) );
  INV_X1 U5740 ( .A(n4623), .ZN(n6262) );
  OAI22_X1 U5741 ( .A1(n6058), .A2(n6261), .B1(n6262), .B2(n4709), .ZN(n4749)
         );
  INV_X1 U5742 ( .A(n6210), .ZN(n4747) );
  OAI22_X1 U5743 ( .A1(n4747), .A2(n6080), .B1(n6351), .B2(n4746), .ZN(n4624)
         );
  AOI21_X1 U5744 ( .B1(n6347), .B2(n4749), .A(n4624), .ZN(n4626) );
  NAND2_X1 U5745 ( .A1(n6346), .A2(n4751), .ZN(n4625) );
  OAI211_X1 U5746 ( .C1(n4755), .C2(n4627), .A(n4626), .B(n4625), .ZN(U3121)
         );
  INV_X1 U5747 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4631) );
  OAI22_X1 U5748 ( .A1(n4747), .A2(n6071), .B1(n6327), .B2(n4746), .ZN(n4628)
         );
  AOI21_X1 U5749 ( .B1(n6323), .B2(n4749), .A(n4628), .ZN(n4630) );
  NAND2_X1 U5750 ( .A1(n6322), .A2(n4751), .ZN(n4629) );
  OAI211_X1 U5751 ( .C1(n4755), .C2(n4631), .A(n4630), .B(n4629), .ZN(U3117)
         );
  INV_X1 U5752 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4635) );
  OAI22_X1 U5753 ( .A1(n4747), .A2(n6321), .B1(n6273), .B2(n4746), .ZN(n4632)
         );
  AOI21_X1 U5754 ( .B1(n6308), .B2(n4749), .A(n4632), .ZN(n4634) );
  NAND2_X1 U5755 ( .A1(n6307), .A2(n4751), .ZN(n4633) );
  OAI211_X1 U5756 ( .C1(n4755), .C2(n4635), .A(n4634), .B(n4633), .ZN(U3116)
         );
  NAND2_X1 U5757 ( .A1(n6024), .A2(n4636), .ZN(n4663) );
  NAND2_X1 U5758 ( .A1(n6024), .A2(n6317), .ZN(n4662) );
  INV_X1 U5759 ( .A(n4662), .ZN(n4650) );
  OR2_X1 U5760 ( .A1(n3033), .A2(n5750), .ZN(n6060) );
  OR2_X1 U5761 ( .A1(n6228), .A2(n6060), .ZN(n6215) );
  NAND2_X1 U5762 ( .A1(n3033), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6027) );
  OR2_X1 U5763 ( .A1(n6119), .A2(n6027), .ZN(n6148) );
  NAND2_X1 U5764 ( .A1(n4638), .A2(n5750), .ZN(n4639) );
  NAND4_X1 U5765 ( .A1(n6181), .A2(n6215), .A3(n6148), .A4(n4639), .ZN(n4640)
         );
  INV_X1 U5766 ( .A(n6024), .ZN(n4651) );
  AOI22_X1 U5767 ( .A1(n4650), .A2(n4640), .B1(n4651), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4641) );
  OAI21_X1 U5768 ( .B1(n6261), .B2(n4663), .A(n4641), .ZN(U3462) );
  INV_X1 U5769 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4645) );
  OAI22_X1 U5770 ( .A1(n4747), .A2(n6339), .B1(n6283), .B2(n4746), .ZN(n4642)
         );
  AOI21_X1 U5771 ( .B1(n6335), .B2(n4749), .A(n4642), .ZN(n4644) );
  NAND2_X1 U5772 ( .A1(n6334), .A2(n4751), .ZN(n4643) );
  OAI211_X1 U5773 ( .C1(n4755), .C2(n4645), .A(n4644), .B(n4643), .ZN(U3119)
         );
  INV_X1 U5774 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4649) );
  OAI22_X1 U5775 ( .A1(n4747), .A2(n6370), .B1(n6299), .B2(n4746), .ZN(n4646)
         );
  AOI21_X1 U5776 ( .B1(n6363), .B2(n4749), .A(n4646), .ZN(n4648) );
  NAND2_X1 U5777 ( .A1(n6360), .A2(n4751), .ZN(n4647) );
  OAI211_X1 U5778 ( .C1(n4755), .C2(n4649), .A(n4648), .B(n4647), .ZN(U3123)
         );
  OAI211_X1 U5779 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3033), .A(n4650), .B(
        n6027), .ZN(n4653) );
  NAND2_X1 U5780 ( .A1(n4651), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4652) );
  OAI211_X1 U5781 ( .C1(n4663), .C2(n6120), .A(n4653), .B(n4652), .ZN(U3464)
         );
  AOI21_X1 U5782 ( .B1(n4655), .B2(n4556), .A(n4654), .ZN(n4872) );
  INV_X1 U5783 ( .A(n4872), .ZN(n4913) );
  OR2_X1 U5784 ( .A1(n4657), .A2(n4656), .ZN(n4658) );
  NAND2_X1 U5785 ( .A1(n4834), .A2(n4658), .ZN(n5966) );
  INV_X1 U5786 ( .A(n5966), .ZN(n4659) );
  AOI22_X1 U5787 ( .A1(n5306), .A2(n4659), .B1(EBX_REG_8__SCAN_IN), .B2(n5305), 
        .ZN(n4660) );
  OAI21_X1 U5788 ( .B1(n4913), .B2(n5312), .A(n4660), .ZN(U2851) );
  XNOR2_X1 U5789 ( .A(n6028), .B(n6027), .ZN(n4661) );
  OAI222_X1 U5790 ( .A1(n6024), .A2(n6381), .B1(n4663), .B2(n4481), .C1(n4662), 
        .C2(n4661), .ZN(U3463) );
  INV_X1 U5791 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5876) );
  OAI222_X1 U5792 ( .A1(n4913), .A2(n5361), .B1(n5359), .B2(n4664), .C1(n5357), 
        .C2(n5876), .ZN(U2883) );
  NOR2_X1 U5793 ( .A1(n6216), .A2(n4672), .ZN(n4667) );
  OAI21_X1 U5794 ( .B1(n4665), .B2(n5750), .A(n6317), .ZN(n4673) );
  INV_X1 U5795 ( .A(n4666), .ZN(n4668) );
  AOI21_X1 U5796 ( .B1(n4668), .B2(n3029), .A(n4667), .ZN(n4674) );
  INV_X1 U5797 ( .A(n4674), .ZN(n4671) );
  AOI21_X1 U5798 ( .B1(n6216), .B2(STATE2_REG_3__SCAN_IN), .A(n4669), .ZN(
        n6314) );
  AOI21_X1 U5799 ( .B1(n6305), .B2(n4672), .A(n6222), .ZN(n4670) );
  OAI22_X1 U5800 ( .A1(n4674), .A2(n4673), .B1(n6303), .B2(n4672), .ZN(n4760)
         );
  AOI22_X1 U5801 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4761), .B1(n6323), 
        .B2(n4760), .ZN(n4676) );
  AOI22_X1 U5802 ( .A1(n6232), .A2(n4763), .B1(n4762), .B2(n6324), .ZN(n4675)
         );
  OAI211_X1 U5803 ( .C1(n4730), .C2(n4766), .A(n4676), .B(n4675), .ZN(U3029)
         );
  AOI22_X1 U5804 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4761), .B1(n6308), 
        .B2(n4760), .ZN(n4678) );
  AOI22_X1 U5805 ( .A1(n6318), .A2(n4763), .B1(n4762), .B2(n6270), .ZN(n4677)
         );
  OAI211_X1 U5806 ( .C1(n4726), .C2(n4766), .A(n4678), .B(n4677), .ZN(U3028)
         );
  AOI22_X1 U5807 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4761), .B1(n6363), 
        .B2(n4760), .ZN(n4680) );
  INV_X1 U5808 ( .A(n6370), .ZN(n6295) );
  AOI22_X1 U5809 ( .A1(n6365), .A2(n4763), .B1(n4762), .B2(n6295), .ZN(n4679)
         );
  OAI211_X1 U5810 ( .C1(n4714), .C2(n4766), .A(n4680), .B(n4679), .ZN(U3035)
         );
  AOI22_X1 U5811 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4761), .B1(n6347), 
        .B2(n4760), .ZN(n4682) );
  AOI22_X1 U5812 ( .A1(n6245), .A2(n4763), .B1(n4762), .B2(n6348), .ZN(n4681)
         );
  OAI211_X1 U5813 ( .C1(n4718), .C2(n4766), .A(n4682), .B(n4681), .ZN(U3033)
         );
  AOI22_X1 U5814 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4761), .B1(n6335), 
        .B2(n4760), .ZN(n4684) );
  INV_X1 U5815 ( .A(n6339), .ZN(n6280) );
  AOI22_X1 U5816 ( .A1(n6336), .A2(n4763), .B1(n4762), .B2(n6280), .ZN(n4683)
         );
  OAI211_X1 U5817 ( .C1(n4722), .C2(n4766), .A(n4684), .B(n4683), .ZN(U3031)
         );
  NAND3_X1 U5818 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6381), .A3(n4976), .ZN(n4700) );
  OR2_X1 U5819 ( .A1(n6216), .A2(n4700), .ZN(n4823) );
  NAND2_X1 U5820 ( .A1(n3031), .A2(n3029), .ZN(n6300) );
  OR2_X1 U5821 ( .A1(n6300), .A2(n4704), .ZN(n4685) );
  AND2_X1 U5822 ( .A1(n4685), .A2(n4823), .ZN(n4689) );
  INV_X1 U5823 ( .A(n4689), .ZN(n4687) );
  OAI21_X1 U5824 ( .B1(n6181), .B2(n6060), .A(n6317), .ZN(n4688) );
  AOI21_X1 U5825 ( .B1(n6305), .B2(n4700), .A(n6222), .ZN(n4686) );
  OAI21_X1 U5826 ( .B1(n4687), .B2(n4688), .A(n4686), .ZN(n4818) );
  OAI22_X1 U5827 ( .A1(n4689), .A2(n4688), .B1(n6303), .B2(n4700), .ZN(n4817)
         );
  AOI22_X1 U5828 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4818), .B1(n6347), 
        .B2(n4817), .ZN(n4691) );
  AOI22_X1 U5829 ( .A1(n5004), .A2(n6245), .B1(n4819), .B2(n6348), .ZN(n4690)
         );
  OAI211_X1 U5830 ( .C1(n4823), .C2(n4718), .A(n4691), .B(n4690), .ZN(U3097)
         );
  AOI22_X1 U5831 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4818), .B1(n6308), 
        .B2(n4817), .ZN(n4693) );
  AOI22_X1 U5832 ( .A1(n5004), .A2(n6318), .B1(n4819), .B2(n6270), .ZN(n4692)
         );
  OAI211_X1 U5833 ( .C1(n4823), .C2(n4726), .A(n4693), .B(n4692), .ZN(U3092)
         );
  AOI22_X1 U5834 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4818), .B1(n6323), 
        .B2(n4817), .ZN(n4695) );
  AOI22_X1 U5835 ( .A1(n5004), .A2(n6232), .B1(n4819), .B2(n6324), .ZN(n4694)
         );
  OAI211_X1 U5836 ( .C1(n4823), .C2(n4730), .A(n4695), .B(n4694), .ZN(U3093)
         );
  AOI22_X1 U5837 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4818), .B1(n6335), 
        .B2(n4817), .ZN(n4697) );
  AOI22_X1 U5838 ( .A1(n5004), .A2(n6336), .B1(n4819), .B2(n6280), .ZN(n4696)
         );
  OAI211_X1 U5839 ( .C1(n4823), .C2(n4722), .A(n4697), .B(n4696), .ZN(U3095)
         );
  AOI22_X1 U5840 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4818), .B1(n6363), 
        .B2(n4817), .ZN(n4699) );
  AOI22_X1 U5841 ( .A1(n5004), .A2(n6365), .B1(n4819), .B2(n6295), .ZN(n4698)
         );
  OAI211_X1 U5842 ( .C1(n4823), .C2(n4714), .A(n4699), .B(n4698), .ZN(U3099)
         );
  NOR2_X1 U5843 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4700), .ZN(n4702)
         );
  OAI211_X1 U5844 ( .C1(n6501), .C2(n4702), .A(n6262), .B(n4701), .ZN(n4707)
         );
  AOI21_X1 U5845 ( .B1(n4810), .B2(n6154), .A(n5750), .ZN(n4705) );
  NOR2_X1 U5846 ( .A1(n6261), .A2(n4704), .ZN(n4708) );
  NOR3_X1 U5847 ( .A1(n4705), .A2(n4708), .A3(n6305), .ZN(n4706) );
  NAND2_X1 U5848 ( .A1(n4809), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4713) );
  INV_X1 U5849 ( .A(n4708), .ZN(n4710) );
  OAI22_X1 U5850 ( .A1(n4710), .A2(n6305), .B1(n6062), .B2(n4709), .ZN(n4812)
         );
  OAI22_X1 U5851 ( .A1(n4810), .A2(n6299), .B1(n6370), .B2(n6154), .ZN(n4711)
         );
  AOI21_X1 U5852 ( .B1(n6363), .B2(n4812), .A(n4711), .ZN(n4712) );
  OAI211_X1 U5853 ( .C1(n4816), .C2(n4714), .A(n4713), .B(n4712), .ZN(U3091)
         );
  NAND2_X1 U5854 ( .A1(n4809), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4717) );
  OAI22_X1 U5855 ( .A1(n4810), .A2(n6351), .B1(n6080), .B2(n6154), .ZN(n4715)
         );
  AOI21_X1 U5856 ( .B1(n6347), .B2(n4812), .A(n4715), .ZN(n4716) );
  OAI211_X1 U5857 ( .C1(n4816), .C2(n4718), .A(n4717), .B(n4716), .ZN(U3089)
         );
  NAND2_X1 U5858 ( .A1(n4809), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4721) );
  OAI22_X1 U5859 ( .A1(n4810), .A2(n6283), .B1(n6339), .B2(n6154), .ZN(n4719)
         );
  AOI21_X1 U5860 ( .B1(n6335), .B2(n4812), .A(n4719), .ZN(n4720) );
  OAI211_X1 U5861 ( .C1(n4816), .C2(n4722), .A(n4721), .B(n4720), .ZN(U3087)
         );
  NAND2_X1 U5862 ( .A1(n4809), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4725) );
  OAI22_X1 U5863 ( .A1(n4810), .A2(n6273), .B1(n6321), .B2(n6154), .ZN(n4723)
         );
  AOI21_X1 U5864 ( .B1(n6308), .B2(n4812), .A(n4723), .ZN(n4724) );
  OAI211_X1 U5865 ( .C1(n4726), .C2(n4816), .A(n4725), .B(n4724), .ZN(U3084)
         );
  NAND2_X1 U5866 ( .A1(n4809), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4729) );
  OAI22_X1 U5867 ( .A1(n4810), .A2(n6327), .B1(n6071), .B2(n6154), .ZN(n4727)
         );
  AOI21_X1 U5868 ( .B1(n6323), .B2(n4812), .A(n4727), .ZN(n4728) );
  OAI211_X1 U5869 ( .C1(n4816), .C2(n4730), .A(n4729), .B(n4728), .ZN(U3085)
         );
  INV_X1 U5870 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4736) );
  NAND2_X1 U5871 ( .A1(DATAI_4_), .A2(n4743), .ZN(n6244) );
  INV_X1 U5872 ( .A(DATAI_28_), .ZN(n4731) );
  INV_X1 U5873 ( .A(n6284), .ZN(n6345) );
  INV_X1 U5874 ( .A(DATAI_20_), .ZN(n4732) );
  INV_X1 U5875 ( .A(n6342), .ZN(n6287) );
  OAI22_X1 U5876 ( .A1(n4747), .A2(n6345), .B1(n6287), .B2(n4746), .ZN(n4733)
         );
  AOI21_X1 U5877 ( .B1(n6341), .B2(n4749), .A(n4733), .ZN(n4735) );
  NAND2_X1 U5878 ( .A1(n6340), .A2(n4751), .ZN(n4734) );
  OAI211_X1 U5879 ( .C1(n4755), .C2(n4736), .A(n4735), .B(n4734), .ZN(U3120)
         );
  INV_X1 U5880 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4742) );
  NAND2_X1 U5881 ( .A1(DATAI_2_), .A2(n4743), .ZN(n6238) );
  INV_X1 U5882 ( .A(DATAI_26_), .ZN(n4737) );
  NOR2_X1 U5883 ( .A1(n5499), .A2(n4737), .ZN(n6276) );
  INV_X1 U5884 ( .A(n6276), .ZN(n6333) );
  INV_X1 U5885 ( .A(DATAI_18_), .ZN(n4738) );
  NOR2_X1 U5886 ( .A1(n5499), .A2(n4738), .ZN(n6330) );
  OAI22_X1 U5887 ( .A1(n4747), .A2(n6333), .B1(n6279), .B2(n4746), .ZN(n4739)
         );
  AOI21_X1 U5888 ( .B1(n6329), .B2(n4749), .A(n4739), .ZN(n4741) );
  NAND2_X1 U5889 ( .A1(n6328), .A2(n4751), .ZN(n4740) );
  OAI211_X1 U5890 ( .C1(n4755), .C2(n4742), .A(n4741), .B(n4740), .ZN(U3118)
         );
  INV_X1 U5891 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4754) );
  NAND2_X1 U5892 ( .A1(DATAI_6_), .A2(n4743), .ZN(n6252) );
  INV_X1 U5893 ( .A(DATAI_30_), .ZN(n4744) );
  INV_X1 U5894 ( .A(n6355), .ZN(n6083) );
  INV_X1 U5895 ( .A(DATAI_22_), .ZN(n4745) );
  NOR2_X1 U5896 ( .A1(n5499), .A2(n4745), .ZN(n6249) );
  INV_X1 U5897 ( .A(n6249), .ZN(n6359) );
  OAI22_X1 U5898 ( .A1(n4747), .A2(n6083), .B1(n6359), .B2(n4746), .ZN(n4748)
         );
  AOI21_X1 U5899 ( .B1(n6353), .B2(n4749), .A(n4748), .ZN(n4753) );
  NAND2_X1 U5900 ( .A1(n6352), .A2(n4751), .ZN(n4752) );
  OAI211_X1 U5901 ( .C1(n4755), .C2(n4754), .A(n4753), .B(n4752), .ZN(U3122)
         );
  INV_X1 U5902 ( .A(n6340), .ZN(n4815) );
  AOI22_X1 U5903 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4761), .B1(n6341), 
        .B2(n4760), .ZN(n4757) );
  AOI22_X1 U5904 ( .A1(n6342), .A2(n4763), .B1(n4762), .B2(n6284), .ZN(n4756)
         );
  OAI211_X1 U5905 ( .C1(n4815), .C2(n4766), .A(n4757), .B(n4756), .ZN(U3032)
         );
  INV_X1 U5906 ( .A(n6352), .ZN(n4822) );
  AOI22_X1 U5907 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4761), .B1(n6353), 
        .B2(n4760), .ZN(n4759) );
  AOI22_X1 U5908 ( .A1(n6249), .A2(n4763), .B1(n4762), .B2(n6355), .ZN(n4758)
         );
  OAI211_X1 U5909 ( .C1(n4822), .C2(n4766), .A(n4759), .B(n4758), .ZN(U3034)
         );
  INV_X1 U5910 ( .A(n6328), .ZN(n4806) );
  AOI22_X1 U5911 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4761), .B1(n6329), 
        .B2(n4760), .ZN(n4765) );
  AOI22_X1 U5912 ( .A1(n6330), .A2(n4763), .B1(n4762), .B2(n6276), .ZN(n4764)
         );
  OAI211_X1 U5913 ( .C1(n4806), .C2(n4766), .A(n4765), .B(n4764), .ZN(U3030)
         );
  INV_X1 U5914 ( .A(n4767), .ZN(n4768) );
  OAI21_X1 U5915 ( .B1(n4654), .B2(n4769), .A(n4767), .ZN(n4921) );
  AOI22_X1 U5916 ( .A1(n5072), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n5352), .ZN(n4770) );
  OAI21_X1 U5917 ( .B1(n4921), .B2(n5361), .A(n4770), .ZN(U2882) );
  NAND2_X1 U5918 ( .A1(n4786), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4773) );
  OAI22_X1 U5919 ( .A1(n4787), .A2(n6359), .B1(n6083), .B2(n6358), .ZN(n4771)
         );
  AOI21_X1 U5920 ( .B1(n6353), .B2(n4789), .A(n4771), .ZN(n4772) );
  OAI211_X1 U5921 ( .C1(n4792), .C2(n4822), .A(n4773), .B(n4772), .ZN(U3026)
         );
  NAND2_X1 U5922 ( .A1(n4796), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4776) );
  OAI22_X1 U5923 ( .A1(n6345), .A2(n4798), .B1(n4797), .B2(n6287), .ZN(n4774)
         );
  AOI21_X1 U5924 ( .B1(n6341), .B2(n4800), .A(n4774), .ZN(n4775) );
  OAI211_X1 U5925 ( .C1(n4803), .C2(n4815), .A(n4776), .B(n4775), .ZN(U3040)
         );
  NAND2_X1 U5926 ( .A1(n4786), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4779) );
  OAI22_X1 U5927 ( .A1(n4787), .A2(n6279), .B1(n6333), .B2(n6358), .ZN(n4777)
         );
  AOI21_X1 U5928 ( .B1(n6329), .B2(n4789), .A(n4777), .ZN(n4778) );
  OAI211_X1 U5929 ( .C1(n4792), .C2(n4806), .A(n4779), .B(n4778), .ZN(U3022)
         );
  NAND2_X1 U5930 ( .A1(n4796), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4782) );
  OAI22_X1 U5931 ( .A1(n6083), .A2(n4798), .B1(n4797), .B2(n6359), .ZN(n4780)
         );
  AOI21_X1 U5932 ( .B1(n6353), .B2(n4800), .A(n4780), .ZN(n4781) );
  OAI211_X1 U5933 ( .C1(n4803), .C2(n4822), .A(n4782), .B(n4781), .ZN(U3042)
         );
  NAND2_X1 U5934 ( .A1(n4809), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4785) );
  OAI22_X1 U5935 ( .A1(n4810), .A2(n6359), .B1(n6083), .B2(n6154), .ZN(n4783)
         );
  AOI21_X1 U5936 ( .B1(n6353), .B2(n4812), .A(n4783), .ZN(n4784) );
  OAI211_X1 U5937 ( .C1(n4816), .C2(n4822), .A(n4785), .B(n4784), .ZN(U3090)
         );
  NAND2_X1 U5938 ( .A1(n4786), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4791) );
  OAI22_X1 U5939 ( .A1(n4787), .A2(n6287), .B1(n6345), .B2(n6358), .ZN(n4788)
         );
  AOI21_X1 U5940 ( .B1(n6341), .B2(n4789), .A(n4788), .ZN(n4790) );
  OAI211_X1 U5941 ( .C1(n4792), .C2(n4815), .A(n4791), .B(n4790), .ZN(U3024)
         );
  NAND2_X1 U5942 ( .A1(n4809), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4795) );
  OAI22_X1 U5943 ( .A1(n4810), .A2(n6279), .B1(n6333), .B2(n6154), .ZN(n4793)
         );
  AOI21_X1 U5944 ( .B1(n6329), .B2(n4812), .A(n4793), .ZN(n4794) );
  OAI211_X1 U5945 ( .C1(n4816), .C2(n4806), .A(n4795), .B(n4794), .ZN(U3086)
         );
  NAND2_X1 U5946 ( .A1(n4796), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4802) );
  OAI22_X1 U5947 ( .A1(n6333), .A2(n4798), .B1(n4797), .B2(n6279), .ZN(n4799)
         );
  AOI21_X1 U5948 ( .B1(n6329), .B2(n4800), .A(n4799), .ZN(n4801) );
  OAI211_X1 U5949 ( .C1(n4803), .C2(n4806), .A(n4802), .B(n4801), .ZN(U3038)
         );
  AOI22_X1 U5950 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4818), .B1(n6329), 
        .B2(n4817), .ZN(n4805) );
  AOI22_X1 U5951 ( .A1(n5004), .A2(n6330), .B1(n4819), .B2(n6276), .ZN(n4804)
         );
  OAI211_X1 U5952 ( .C1(n4823), .C2(n4806), .A(n4805), .B(n4804), .ZN(U3094)
         );
  AOI22_X1 U5953 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4818), .B1(n6341), 
        .B2(n4817), .ZN(n4808) );
  AOI22_X1 U5954 ( .A1(n5004), .A2(n6342), .B1(n4819), .B2(n6284), .ZN(n4807)
         );
  OAI211_X1 U5955 ( .C1(n4823), .C2(n4815), .A(n4808), .B(n4807), .ZN(U3096)
         );
  NAND2_X1 U5956 ( .A1(n4809), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4814) );
  OAI22_X1 U5957 ( .A1(n4810), .A2(n6287), .B1(n6345), .B2(n6154), .ZN(n4811)
         );
  AOI21_X1 U5958 ( .B1(n6341), .B2(n4812), .A(n4811), .ZN(n4813) );
  OAI211_X1 U5959 ( .C1(n4816), .C2(n4815), .A(n4814), .B(n4813), .ZN(U3088)
         );
  AOI22_X1 U5960 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4818), .B1(n6353), 
        .B2(n4817), .ZN(n4821) );
  AOI22_X1 U5961 ( .A1(n5004), .A2(n6249), .B1(n4819), .B2(n6355), .ZN(n4820)
         );
  OAI211_X1 U5962 ( .C1(n4823), .C2(n4822), .A(n4821), .B(n4820), .ZN(U3098)
         );
  INV_X1 U5963 ( .A(n6424), .ZN(n6532) );
  AOI21_X1 U5964 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6532), .A(n6414), .ZN(
        n6415) );
  AOI21_X1 U5965 ( .B1(n6414), .B2(n5091), .A(n6415), .ZN(n4825) );
  AND2_X1 U5966 ( .A1(n4824), .A2(n4077), .ZN(n6420) );
  INV_X1 U5967 ( .A(n4917), .ZN(n4849) );
  NOR2_X1 U5968 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4842) );
  INV_X1 U5969 ( .A(n4842), .ZN(n4830) );
  NAND2_X1 U5970 ( .A1(n3208), .A2(n4830), .ZN(n4840) );
  NAND2_X1 U5971 ( .A1(n4831), .A2(EBX_REG_31__SCAN_IN), .ZN(n4832) );
  NOR2_X1 U5972 ( .A1(n4840), .A2(n4832), .ZN(n4833) );
  INV_X1 U5973 ( .A(n4834), .ZN(n4837) );
  INV_X1 U5974 ( .A(n4836), .ZN(n4865) );
  OAI21_X1 U5975 ( .B1(n4837), .B2(n2999), .A(n4865), .ZN(n5956) );
  NOR2_X1 U5976 ( .A1(n5849), .A2(n5956), .ZN(n4848) );
  NAND2_X1 U5977 ( .A1(n4838), .A2(n4842), .ZN(n6408) );
  NAND2_X1 U5978 ( .A1(n3092), .A2(n6408), .ZN(n4839) );
  OAI21_X1 U5979 ( .B1(EBX_REG_31__SCAN_IN), .B2(n4840), .A(n4839), .ZN(n4841)
         );
  AND2_X2 U5980 ( .A1(n6526), .A2(n4841), .ZN(n5831) );
  AND3_X1 U5981 ( .A1(n4843), .A2(n4842), .A3(n3208), .ZN(n4844) );
  INV_X1 U5982 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6453) );
  INV_X1 U5983 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6515) );
  INV_X1 U5984 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6451) );
  INV_X1 U5985 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6448) );
  NOR3_X1 U5986 ( .A1(n6515), .A2(n6451), .A3(n6448), .ZN(n5816) );
  NAND2_X1 U5987 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5816), .ZN(n5809) );
  NOR2_X1 U5988 ( .A1(n6453), .A2(n5809), .ZN(n4939) );
  NAND2_X1 U5989 ( .A1(REIP_REG_6__SCAN_IN), .A2(n4939), .ZN(n5796) );
  NOR2_X1 U5990 ( .A1(n6456), .A2(n5796), .ZN(n4907) );
  OAI21_X1 U5991 ( .B1(n5833), .B2(n4952), .A(n5858), .ZN(n5788) );
  AOI22_X1 U5992 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5831), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5788), .ZN(n4845) );
  INV_X1 U5993 ( .A(n6000), .ZN(n5819) );
  OAI211_X1 U5994 ( .C1(n5821), .C2(n4846), .A(n4845), .B(n5819), .ZN(n4847)
         );
  AOI211_X1 U5995 ( .C1(n5776), .C2(n4849), .A(n4848), .B(n4847), .ZN(n4852)
         );
  INV_X1 U5996 ( .A(n4952), .ZN(n4906) );
  INV_X1 U5997 ( .A(n5790), .ZN(n4850) );
  NOR2_X1 U5998 ( .A1(n4850), .A2(REIP_REG_9__SCAN_IN), .ZN(n5789) );
  INV_X1 U5999 ( .A(n5789), .ZN(n4851) );
  OAI211_X1 U6000 ( .C1(n4921), .C2(n5785), .A(n4852), .B(n4851), .ZN(U2818)
         );
  INV_X1 U6001 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4853) );
  OAI222_X1 U6002 ( .A1(n4921), .A2(n5312), .B1(n4853), .B2(n5311), .C1(n5309), 
        .C2(n5956), .ZN(U2850) );
  NOR2_X1 U6003 ( .A1(n4768), .A2(n4855), .ZN(n4856) );
  AOI22_X1 U6004 ( .A1(n5072), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n5352), .ZN(n4857) );
  OAI21_X1 U6005 ( .B1(n5786), .B2(n5361), .A(n4857), .ZN(U2881) );
  INV_X1 U6006 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U6007 ( .A1(n5494), .A2(n4858), .ZN(n4862) );
  NOR2_X1 U6008 ( .A1(n5846), .A2(n5499), .ZN(n4859) );
  AOI211_X1 U6009 ( .C1(n5936), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4860), 
        .B(n4859), .ZN(n4861) );
  OAI211_X1 U6010 ( .C1(n4863), .C2(n5753), .A(n4862), .B(n4861), .ZN(U2985)
         );
  INV_X1 U6011 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6543) );
  AND2_X1 U6012 ( .A1(n4865), .A2(n4864), .ZN(n4866) );
  OR2_X1 U6013 ( .A1(n3038), .A2(n4866), .ZN(n5781) );
  OAI222_X1 U6014 ( .A1(n5786), .A2(n5312), .B1(n5311), .B2(n6543), .C1(n5781), 
        .C2(n5309), .ZN(U2849) );
  OAI21_X1 U6015 ( .B1(n4867), .B2(n4869), .A(n4868), .ZN(n5965) );
  AOI22_X1 U6016 ( .A1(n5936), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6000), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4870) );
  OAI21_X1 U6017 ( .B1(n5946), .B2(n4908), .A(n4870), .ZN(n4871) );
  AOI21_X1 U6018 ( .B1(n4872), .B2(n5941), .A(n4871), .ZN(n4873) );
  OAI21_X1 U6019 ( .B1(n5965), .B2(n5753), .A(n4873), .ZN(U2978) );
  AOI21_X1 U6020 ( .B1(n5936), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4874), 
        .ZN(n4875) );
  OAI21_X1 U6021 ( .B1(n5946), .B2(n4943), .A(n4875), .ZN(n4876) );
  AOI21_X1 U6022 ( .B1(n4877), .B2(n5941), .A(n4876), .ZN(n4878) );
  OAI21_X1 U6023 ( .B1(n4879), .B2(n5753), .A(n4878), .ZN(U2980) );
  NAND2_X1 U6024 ( .A1(n6526), .A2(n5745), .ZN(n4880) );
  NAND2_X1 U6025 ( .A1(n4880), .A2(n5785), .ZN(n5854) );
  INV_X1 U6026 ( .A(n5854), .ZN(n5823) );
  OAI21_X1 U6027 ( .B1(n5833), .B2(n5816), .A(n5858), .ZN(n5827) );
  OR2_X1 U6028 ( .A1(n5833), .A2(REIP_REG_1__SCAN_IN), .ZN(n5845) );
  AND2_X1 U6029 ( .A1(n5858), .A2(REIP_REG_2__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U6030 ( .A1(n5845), .A2(n4881), .ZN(n5835) );
  NAND2_X1 U6031 ( .A1(n5835), .A2(n6451), .ZN(n4888) );
  NAND2_X1 U6032 ( .A1(n6526), .A2(n4882), .ZN(n5847) );
  INV_X1 U6033 ( .A(n4883), .ZN(n6001) );
  AOI22_X1 U6034 ( .A1(n5832), .A2(n6001), .B1(n5831), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4886) );
  INV_X1 U6035 ( .A(n5935), .ZN(n4884) );
  AOI22_X1 U6036 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n5843), .B1(n5776), 
        .B2(n4884), .ZN(n4885) );
  OAI211_X1 U6037 ( .C1(n6261), .C2(n5847), .A(n4886), .B(n4885), .ZN(n4887)
         );
  AOI21_X1 U6038 ( .B1(n5827), .B2(n4888), .A(n4887), .ZN(n4889) );
  OAI21_X1 U6039 ( .B1(n5823), .B2(n5927), .A(n4889), .ZN(U2824) );
  OAI21_X1 U6040 ( .B1(n4890), .B2(n4893), .A(n4892), .ZN(n5993) );
  NAND2_X1 U6041 ( .A1(n6000), .A2(REIP_REG_4__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U6042 ( .A1(n5936), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4894)
         );
  OAI211_X1 U6043 ( .C1(n5946), .C2(n5822), .A(n5990), .B(n4894), .ZN(n4895)
         );
  AOI21_X1 U6044 ( .B1(n4896), .B2(n5941), .A(n4895), .ZN(n4897) );
  OAI21_X1 U6045 ( .B1(n5993), .B2(n5753), .A(n4897), .ZN(U2982) );
  NOR2_X1 U6046 ( .A1(n4854), .A2(n4900), .ZN(n4901) );
  OR2_X1 U6047 ( .A1(n4899), .A2(n4901), .ZN(n4966) );
  OAI21_X1 U6048 ( .B1(n3038), .B2(n4902), .A(n5028), .ZN(n4949) );
  INV_X1 U6049 ( .A(n4949), .ZN(n5948) );
  AOI22_X1 U6050 ( .A1(n5306), .A2(n5948), .B1(EBX_REG_11__SCAN_IN), .B2(n5305), .ZN(n4903) );
  OAI21_X1 U6051 ( .B1(n4966), .B2(n5312), .A(n4903), .ZN(U2848) );
  AOI22_X1 U6052 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n5843), .B1(
        REIP_REG_8__SCAN_IN), .B2(n5788), .ZN(n4904) );
  OAI211_X1 U6053 ( .C1(n5851), .C2(n4905), .A(n4904), .B(n5819), .ZN(n4911)
         );
  INV_X1 U6054 ( .A(n5833), .ZN(n5817) );
  AND3_X1 U6055 ( .A1(n5817), .A2(n4907), .A3(n4906), .ZN(n4910) );
  OAI22_X1 U6056 ( .A1(n5848), .A2(n4908), .B1(n5849), .B2(n5966), .ZN(n4909)
         );
  NOR3_X1 U6057 ( .A1(n4911), .A2(n4910), .A3(n4909), .ZN(n4912) );
  OAI21_X1 U6058 ( .B1(n5785), .B2(n4913), .A(n4912), .ZN(U2819) );
  XNOR2_X1 U6059 ( .A(n5436), .B(n5963), .ZN(n4915) );
  XNOR2_X1 U6060 ( .A(n4914), .B(n4915), .ZN(n5960) );
  NAND2_X1 U6061 ( .A1(n5960), .A2(n5940), .ZN(n4920) );
  INV_X1 U6062 ( .A(REIP_REG_9__SCAN_IN), .ZN(n4916) );
  NOR2_X1 U6063 ( .A1(n5819), .A2(n4916), .ZN(n5957) );
  NOR2_X1 U6064 ( .A1(n5946), .A2(n4917), .ZN(n4918) );
  AOI211_X1 U6065 ( .C1(n5936), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n5957), 
        .B(n4918), .ZN(n4919) );
  OAI211_X1 U6066 ( .C1(n5499), .C2(n4921), .A(n4920), .B(n4919), .ZN(U2977)
         );
  NAND2_X1 U6067 ( .A1(n4959), .A2(n4922), .ZN(n4924) );
  XOR2_X1 U6068 ( .A(n4924), .B(n4923), .Z(n5014) );
  NAND2_X1 U6069 ( .A1(n4929), .A2(n4925), .ZN(n5979) );
  NOR2_X1 U6070 ( .A1(n4926), .A2(n5979), .ZN(n5959) );
  OAI211_X1 U6071 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5959), .B(n4927), .ZN(n4933) );
  INV_X1 U6072 ( .A(n5586), .ZN(n5057) );
  OAI22_X1 U6073 ( .A1(n4929), .A2(n5721), .B1(n5057), .B2(n4928), .ZN(n4930)
         );
  NOR2_X1 U6074 ( .A1(n5582), .A2(n4930), .ZN(n5977) );
  OAI21_X1 U6075 ( .B1(n5968), .B2(n5615), .A(n5977), .ZN(n5955) );
  INV_X1 U6076 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6460) );
  OAI22_X1 U6077 ( .A1(n5967), .A2(n5781), .B1(n6460), .B2(n5819), .ZN(n4931)
         );
  AOI21_X1 U6078 ( .B1(n5955), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n4931), 
        .ZN(n4932) );
  OAI211_X1 U6079 ( .C1(n5014), .C2(n5623), .A(n4933), .B(n4932), .ZN(U3008)
         );
  INV_X1 U6080 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6564) );
  OAI222_X1 U6081 ( .A1(n4966), .A2(n5361), .B1(n5359), .B2(n4934), .C1(n5357), 
        .C2(n6564), .ZN(U2880) );
  OAI21_X1 U6082 ( .B1(n4899), .B2(n4936), .A(n4935), .ZN(n5774) );
  XNOR2_X1 U6083 ( .A(n5028), .B(n4937), .ZN(n5769) );
  AOI22_X1 U6084 ( .A1(n5306), .A2(n5769), .B1(EBX_REG_12__SCAN_IN), .B2(n5305), .ZN(n4938) );
  OAI21_X1 U6085 ( .B1(n5774), .B2(n5312), .A(n4938), .ZN(U2847) );
  AND2_X1 U6086 ( .A1(n5817), .A2(n4939), .ZN(n4944) );
  NAND2_X1 U6087 ( .A1(n5833), .A2(n5858), .ZN(n5193) );
  NOR2_X1 U6088 ( .A1(n4944), .A2(n5253), .ZN(n5811) );
  AOI22_X1 U6089 ( .A1(n5832), .A2(n4940), .B1(n5831), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4942) );
  AOI21_X1 U6090 ( .B1(n5843), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6000), 
        .ZN(n4941) );
  OAI211_X1 U6091 ( .C1(n4943), .C2(n5848), .A(n4942), .B(n4941), .ZN(n4946)
         );
  INV_X1 U6092 ( .A(n4944), .ZN(n4945) );
  NOR2_X1 U6093 ( .A1(n4945), .A2(REIP_REG_6__SCAN_IN), .ZN(n5804) );
  AOI211_X1 U6094 ( .C1(n5811), .C2(REIP_REG_6__SCAN_IN), .A(n4946), .B(n5804), 
        .ZN(n4947) );
  OAI21_X1 U6095 ( .B1(n5785), .B2(n4948), .A(n4947), .ZN(U2821) );
  NAND2_X1 U6096 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n4950) );
  NOR2_X1 U6097 ( .A1(REIP_REG_11__SCAN_IN), .A2(n4950), .ZN(n4956) );
  OAI22_X1 U6098 ( .A1(n4962), .A2(n5848), .B1(n5849), .B2(n4949), .ZN(n4955)
         );
  INV_X1 U6099 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6670) );
  NOR2_X1 U6100 ( .A1(n6670), .A2(n4950), .ZN(n4951) );
  NAND3_X1 U6101 ( .A1(n4952), .A2(n4951), .A3(n5858), .ZN(n5077) );
  NAND2_X1 U6102 ( .A1(n5193), .A2(n5077), .ZN(n5779) );
  AOI22_X1 U6103 ( .A1(EBX_REG_11__SCAN_IN), .A2(n5831), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n5843), .ZN(n4953) );
  OAI211_X1 U6104 ( .C1(n6670), .C2(n5779), .A(n4953), .B(n5819), .ZN(n4954)
         );
  AOI211_X1 U6105 ( .C1(n5790), .C2(n4956), .A(n4955), .B(n4954), .ZN(n4957)
         );
  OAI21_X1 U6106 ( .B1(n5785), .B2(n4966), .A(n4957), .ZN(U2816) );
  NAND2_X1 U6107 ( .A1(n4958), .A2(n4959), .ZN(n4961) );
  XNOR2_X1 U6108 ( .A(n5436), .B(n5953), .ZN(n4960) );
  XNOR2_X1 U6109 ( .A(n4961), .B(n4960), .ZN(n5950) );
  NAND2_X1 U6110 ( .A1(n5950), .A2(n5940), .ZN(n4965) );
  NOR2_X1 U6111 ( .A1(n5819), .A2(n6670), .ZN(n5947) );
  NOR2_X1 U6112 ( .A1(n5946), .A2(n4962), .ZN(n4963) );
  AOI211_X1 U6113 ( .C1(n5936), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5947), 
        .B(n4963), .ZN(n4964) );
  OAI211_X1 U6114 ( .C1(n5499), .C2(n4966), .A(n4965), .B(n4964), .ZN(U2975)
         );
  INV_X1 U6115 ( .A(DATAI_12_), .ZN(n4968) );
  OAI222_X1 U6116 ( .A1(n5774), .A2(n5361), .B1(n4968), .B2(n5359), .C1(n4967), 
        .C2(n5357), .ZN(U2879) );
  INV_X1 U6117 ( .A(n5004), .ZN(n4969) );
  NAND2_X1 U6118 ( .A1(n4969), .A2(n6317), .ZN(n4971) );
  NAND2_X1 U6119 ( .A1(n3033), .A2(n4970), .ZN(n6118) );
  OAI21_X1 U6120 ( .B1(n4971), .B2(n6208), .A(n6310), .ZN(n4978) );
  INV_X1 U6121 ( .A(n4972), .ZN(n4973) );
  INV_X1 U6122 ( .A(n4974), .ZN(n6263) );
  NOR2_X1 U6123 ( .A1(n6263), .A2(n6265), .ZN(n4975) );
  NOR3_X1 U6124 ( .A1(n6265), .A2(n4976), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n6189) );
  NAND2_X1 U6125 ( .A1(n6216), .A2(n6189), .ZN(n4979) );
  INV_X1 U6126 ( .A(n6184), .ZN(n4977) );
  AOI22_X1 U6127 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4979), .B1(n4978), .B2(
        n4977), .ZN(n4980) );
  OAI211_X1 U6128 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6303), .A(n4981), .B(n4980), .ZN(n5003) );
  AOI22_X1 U6129 ( .A1(n5004), .A2(n6270), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5003), .ZN(n4982) );
  OAI21_X1 U6130 ( .B1(n5006), .B2(n6273), .A(n4982), .ZN(n4983) );
  AOI21_X1 U6131 ( .B1(n6307), .B2(n5008), .A(n4983), .ZN(n4984) );
  OAI21_X1 U6132 ( .B1(n5010), .B2(n6231), .A(n4984), .ZN(U3100) );
  AOI22_X1 U6133 ( .A1(n5004), .A2(n6295), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5003), .ZN(n4985) );
  OAI21_X1 U6134 ( .B1(n5006), .B2(n6299), .A(n4985), .ZN(n4986) );
  AOI21_X1 U6135 ( .B1(n6360), .B2(n5008), .A(n4986), .ZN(n4987) );
  OAI21_X1 U6136 ( .B1(n5010), .B2(n6258), .A(n4987), .ZN(U3107) );
  AOI22_X1 U6137 ( .A1(n5004), .A2(n6280), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5003), .ZN(n4988) );
  OAI21_X1 U6138 ( .B1(n5006), .B2(n6283), .A(n4988), .ZN(n4989) );
  AOI21_X1 U6139 ( .B1(n6334), .B2(n5008), .A(n4989), .ZN(n4990) );
  OAI21_X1 U6140 ( .B1(n5010), .B2(n6241), .A(n4990), .ZN(U3103) );
  AOI22_X1 U6141 ( .A1(n5004), .A2(n6284), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5003), .ZN(n4991) );
  OAI21_X1 U6142 ( .B1(n5006), .B2(n6287), .A(n4991), .ZN(n4992) );
  AOI21_X1 U6143 ( .B1(n6340), .B2(n5008), .A(n4992), .ZN(n4993) );
  OAI21_X1 U6144 ( .B1(n5010), .B2(n6244), .A(n4993), .ZN(U3104) );
  AOI22_X1 U6145 ( .A1(n5004), .A2(n6276), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5003), .ZN(n4994) );
  OAI21_X1 U6146 ( .B1(n5006), .B2(n6279), .A(n4994), .ZN(n4995) );
  AOI21_X1 U6147 ( .B1(n6328), .B2(n5008), .A(n4995), .ZN(n4996) );
  OAI21_X1 U6148 ( .B1(n5010), .B2(n6238), .A(n4996), .ZN(U3102) );
  AOI22_X1 U6149 ( .A1(n5004), .A2(n6348), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5003), .ZN(n4997) );
  OAI21_X1 U6150 ( .B1(n5006), .B2(n6351), .A(n4997), .ZN(n4998) );
  AOI21_X1 U6151 ( .B1(n6346), .B2(n5008), .A(n4998), .ZN(n4999) );
  OAI21_X1 U6152 ( .B1(n5010), .B2(n6248), .A(n4999), .ZN(U3105) );
  AOI22_X1 U6153 ( .A1(n5004), .A2(n6324), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5003), .ZN(n5000) );
  OAI21_X1 U6154 ( .B1(n5006), .B2(n6327), .A(n5000), .ZN(n5001) );
  AOI21_X1 U6155 ( .B1(n6322), .B2(n5008), .A(n5001), .ZN(n5002) );
  OAI21_X1 U6156 ( .B1(n5010), .B2(n6235), .A(n5002), .ZN(U3101) );
  AOI22_X1 U6157 ( .A1(n5004), .A2(n6355), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5003), .ZN(n5005) );
  OAI21_X1 U6158 ( .B1(n5006), .B2(n6359), .A(n5005), .ZN(n5007) );
  AOI21_X1 U6159 ( .B1(n6352), .B2(n5008), .A(n5007), .ZN(n5009) );
  OAI21_X1 U6160 ( .B1(n5010), .B2(n6252), .A(n5009), .ZN(U3106) );
  OAI22_X1 U6161 ( .A1(n5492), .A2(n6711), .B1(n5819), .B2(n6460), .ZN(n5012)
         );
  NOR2_X1 U6162 ( .A1(n5786), .A2(n5499), .ZN(n5011) );
  AOI211_X1 U6163 ( .C1(n5494), .C2(n5783), .A(n5012), .B(n5011), .ZN(n5013)
         );
  OAI21_X1 U6164 ( .B1(n5014), .B2(n5753), .A(n5013), .ZN(U2976) );
  XNOR2_X1 U6165 ( .A(n5015), .B(n5016), .ZN(n5737) );
  INV_X1 U6166 ( .A(n5737), .ZN(n5024) );
  INV_X1 U6167 ( .A(n5018), .ZN(n5019) );
  AOI21_X1 U6168 ( .B1(n5017), .B2(n5020), .A(n5019), .ZN(n5025) );
  AOI22_X1 U6169 ( .A1(n5936), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n6000), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n5021) );
  OAI21_X1 U6170 ( .B1(n5946), .B2(n5032), .A(n5021), .ZN(n5022) );
  AOI21_X1 U6171 ( .B1(n5025), .B2(n5941), .A(n5022), .ZN(n5023) );
  OAI21_X1 U6172 ( .B1(n5024), .B2(n5753), .A(n5023), .ZN(U2973) );
  INV_X1 U6173 ( .A(n5025), .ZN(n5039) );
  OAI21_X1 U6174 ( .B1(n5028), .B2(n5027), .A(n5026), .ZN(n5029) );
  NAND2_X1 U6175 ( .A1(n5029), .A2(n5237), .ZN(n5031) );
  INV_X1 U6176 ( .A(n5031), .ZN(n5738) );
  AOI22_X1 U6177 ( .A1(n5306), .A2(n5738), .B1(EBX_REG_13__SCAN_IN), .B2(n5305), .ZN(n5030) );
  OAI21_X1 U6178 ( .B1(n5039), .B2(n5312), .A(n5030), .ZN(U2846) );
  NAND2_X1 U6179 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5243) );
  INV_X1 U6180 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6463) );
  INV_X1 U6181 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6465) );
  NAND4_X1 U6182 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(n5790), .ZN(n5780) );
  AOI21_X1 U6183 ( .B1(n6463), .B2(n6465), .A(n5780), .ZN(n5036) );
  OAI22_X1 U6184 ( .A1(n5032), .A2(n5848), .B1(n5849), .B2(n5031), .ZN(n5035)
         );
  AOI22_X1 U6185 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5831), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n5843), .ZN(n5033) );
  OAI211_X1 U6186 ( .C1(n6463), .C2(n5779), .A(n5033), .B(n5819), .ZN(n5034)
         );
  AOI211_X1 U6187 ( .C1(n5243), .C2(n5036), .A(n5035), .B(n5034), .ZN(n5037)
         );
  OAI21_X1 U6188 ( .B1(n5039), .B2(n5785), .A(n5037), .ZN(U2814) );
  OAI222_X1 U6189 ( .A1(n5039), .A2(n5361), .B1(n5359), .B2(n5038), .C1(n5357), 
        .C2(n3732), .ZN(U2878) );
  INV_X1 U6190 ( .A(n5040), .ZN(n5042) );
  NOR2_X1 U6191 ( .A1(n5042), .A2(n5041), .ZN(n5044) );
  NOR3_X1 U6192 ( .A1(n5048), .A2(n6645), .A3(n6412), .ZN(n5043) );
  AOI211_X1 U6193 ( .C1(n5046), .C2(n5045), .A(n5044), .B(n5043), .ZN(n5050)
         );
  AOI21_X1 U6194 ( .B1(n5048), .B2(n5047), .A(n6503), .ZN(n5049) );
  OAI22_X1 U6195 ( .A1(n5050), .A2(n6503), .B1(n5049), .B2(n3612), .ZN(U3459)
         );
  NOR2_X1 U6196 ( .A1(n5053), .A2(n3056), .ZN(n5054) );
  XNOR2_X1 U6197 ( .A(n5051), .B(n5054), .ZN(n5068) );
  OAI22_X1 U6198 ( .A1(n6013), .A2(n5055), .B1(n5720), .B2(n5721), .ZN(n5949)
         );
  NAND3_X1 U6199 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5060), .A3(n5949), .ZN(n5056) );
  OAI21_X1 U6200 ( .B1(n5819), .B2(n6465), .A(n5056), .ZN(n5063) );
  NOR2_X1 U6201 ( .A1(n5057), .A2(n5725), .ZN(n5058) );
  AOI211_X1 U6202 ( .C1(n6016), .C2(n5720), .A(n5058), .B(n5582), .ZN(n5954)
         );
  INV_X1 U6203 ( .A(n6013), .ZN(n5059) );
  OAI21_X1 U6204 ( .B1(n6016), .B2(n5059), .A(n5953), .ZN(n5061) );
  AOI21_X1 U6205 ( .B1(n5954), .B2(n5061), .A(n5060), .ZN(n5062) );
  AOI211_X1 U6206 ( .C1(n6010), .C2(n5769), .A(n5063), .B(n5062), .ZN(n5064)
         );
  OAI21_X1 U6207 ( .B1(n5068), .B2(n5623), .A(n5064), .ZN(U3006) );
  INV_X1 U6208 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5771) );
  OAI22_X1 U6209 ( .A1(n5492), .A2(n5771), .B1(n5819), .B2(n6465), .ZN(n5066)
         );
  NOR2_X1 U6210 ( .A1(n5774), .A2(n5499), .ZN(n5065) );
  AOI211_X1 U6211 ( .C1(n5494), .C2(n5777), .A(n5066), .B(n5065), .ZN(n5067)
         );
  OAI21_X1 U6212 ( .B1(n5068), .B2(n5753), .A(n5067), .ZN(U2974) );
  INV_X1 U6213 ( .A(n5218), .ZN(n5070) );
  OAI21_X1 U6214 ( .B1(n3007), .B2(n5071), .A(n5070), .ZN(n5479) );
  AOI22_X1 U6215 ( .A1(n5072), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n5352), .ZN(n5073) );
  OAI21_X1 U6216 ( .B1(n5479), .B2(n5361), .A(n5073), .ZN(U2876) );
  INV_X1 U6217 ( .A(n5482), .ZN(n5076) );
  NOR2_X1 U6218 ( .A1(n5239), .A2(n5074), .ZN(n5075) );
  OR2_X1 U6219 ( .A1(n5221), .A2(n5075), .ZN(n5620) );
  OAI22_X1 U6220 ( .A1(n5848), .A2(n5076), .B1(n5849), .B2(n5620), .ZN(n5082)
         );
  NAND3_X1 U6221 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .ZN(n5078) );
  NOR2_X1 U6222 ( .A1(n5077), .A2(n5078), .ZN(n5094) );
  NOR2_X1 U6223 ( .A1(n5253), .A2(n5094), .ZN(n5235) );
  INV_X1 U6224 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6469) );
  AOI22_X1 U6225 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5235), .B1(n5225), .B2(
        n6469), .ZN(n5079) );
  OAI211_X1 U6226 ( .C1(n5821), .C2(n5080), .A(n5079), .B(n5819), .ZN(n5081)
         );
  AOI211_X1 U6227 ( .C1(EBX_REG_15__SCAN_IN), .C2(n5831), .A(n5082), .B(n5081), 
        .ZN(n5083) );
  OAI21_X1 U6228 ( .B1(n5479), .B2(n5785), .A(n5083), .ZN(U2812) );
  INV_X1 U6229 ( .A(n5084), .ZN(n5116) );
  AOI21_X1 U6230 ( .B1(n5936), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5085), 
        .ZN(n5086) );
  OAI21_X1 U6231 ( .B1(n5946), .B2(n5116), .A(n5086), .ZN(n5087) );
  AOI21_X1 U6232 ( .B1(n5115), .B2(n5941), .A(n5087), .ZN(n5088) );
  OAI21_X1 U6233 ( .B1(n5089), .B2(n5753), .A(n5088), .ZN(U2956) );
  NAND2_X1 U6234 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(n5090), .ZN(n5092) );
  NAND3_X1 U6235 ( .A1(n5093), .A2(n5092), .A3(n5091), .ZN(U2788) );
  INV_X1 U6236 ( .A(n5314), .ZN(n5114) );
  INV_X1 U6237 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6476) );
  NAND3_X1 U6238 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        n5225), .ZN(n5212) );
  NAND3_X1 U6239 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        n5202), .ZN(n5682) );
  NAND4_X1 U6240 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5666), .ZN(n5630) );
  NAND3_X1 U6241 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5150) );
  NOR2_X1 U6242 ( .A1(n5630), .A2(n5150), .ZN(n5163) );
  NAND3_X1 U6243 ( .A1(n5163), .A2(REIP_REG_27__SCAN_IN), .A3(
        REIP_REG_28__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U6244 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n5110) );
  INV_X1 U6245 ( .A(n5110), .ZN(n5099) );
  NAND2_X1 U6246 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5098) );
  INV_X1 U6247 ( .A(n5150), .ZN(n5097) );
  NAND3_X1 U6248 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5096) );
  NAND4_X1 U6249 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5094), .A3(
        REIP_REG_16__SCAN_IN), .A4(REIP_REG_15__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6250 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5179) );
  NOR2_X1 U6251 ( .A1(n5192), .A2(n5179), .ZN(n5095) );
  AOI21_X1 U6252 ( .B1(n5095), .B2(REIP_REG_20__SCAN_IN), .A(n5253), .ZN(n5687) );
  AOI21_X1 U6253 ( .B1(n5193), .B2(n5096), .A(n5687), .ZN(n5661) );
  OAI21_X1 U6254 ( .B1(n5253), .B2(n5097), .A(n5661), .ZN(n5636) );
  AOI21_X1 U6255 ( .B1(n5817), .B2(n5098), .A(n5636), .ZN(n5128) );
  OAI21_X1 U6256 ( .B1(n5137), .B2(n5099), .A(n5128), .ZN(n5121) );
  OAI22_X1 U6257 ( .A1(n5101), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5100), .ZN(n5107) );
  INV_X1 U6258 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6259 ( .A1(n5296), .A2(n5255), .ZN(n5130) );
  OAI21_X2 U6260 ( .B1(n5103), .B2(n5296), .A(n3093), .ZN(n5129) );
  AOI21_X2 U6261 ( .B1(n5129), .B2(n5105), .A(n5104), .ZN(n5106) );
  NAND2_X1 U6262 ( .A1(n5843), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5109)
         );
  NAND4_X1 U6263 ( .A1(n6526), .A2(n3092), .A3(EBX_REG_31__SCAN_IN), .A4(n6408), .ZN(n5108) );
  OAI211_X1 U6264 ( .C1(n5505), .C2(n5849), .A(n5109), .B(n5108), .ZN(n5112)
         );
  NOR3_X1 U6265 ( .A1(n5137), .A2(REIP_REG_31__SCAN_IN), .A3(n5110), .ZN(n5111) );
  OAI21_X1 U6266 ( .B1(n5114), .B2(n5785), .A(n5113), .ZN(U2796) );
  OAI22_X1 U6267 ( .A1(n5117), .A2(n5821), .B1(n5848), .B2(n5116), .ZN(n5120)
         );
  NOR2_X1 U6268 ( .A1(n5118), .A2(n5849), .ZN(n5119) );
  AOI211_X1 U6269 ( .C1(EBX_REG_30__SCAN_IN), .C2(n5831), .A(n5120), .B(n5119), 
        .ZN(n5124) );
  INV_X1 U6270 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6492) );
  NOR2_X1 U6271 ( .A1(n5137), .A2(n6492), .ZN(n5122) );
  OAI21_X1 U6272 ( .B1(n5122), .B2(REIP_REG_30__SCAN_IN), .A(n5121), .ZN(n5123) );
  OAI211_X1 U6273 ( .C1(n5319), .C2(n5785), .A(n5124), .B(n5123), .ZN(U2797)
         );
  AOI21_X1 U6274 ( .B1(n5127), .B2(n5125), .A(n5126), .ZN(n5367) );
  INV_X1 U6275 ( .A(n5367), .ZN(n5322) );
  INV_X1 U6276 ( .A(n5128), .ZN(n5153) );
  INV_X1 U6277 ( .A(n5129), .ZN(n5133) );
  OAI211_X1 U6278 ( .C1(n5296), .C2(n5131), .A(n5102), .B(n5130), .ZN(n5132)
         );
  NAND2_X1 U6279 ( .A1(n5133), .A2(n5132), .ZN(n5511) );
  OAI22_X1 U6280 ( .A1(n5134), .A2(n5821), .B1(n5848), .B2(n5365), .ZN(n5135)
         );
  AOI21_X1 U6281 ( .B1(n5831), .B2(EBX_REG_29__SCAN_IN), .A(n5135), .ZN(n5136)
         );
  OAI21_X1 U6282 ( .B1(n5511), .B2(n5849), .A(n5136), .ZN(n5139) );
  NOR2_X1 U6283 ( .A1(n5137), .A2(REIP_REG_29__SCAN_IN), .ZN(n5138) );
  AOI211_X1 U6284 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5153), .A(n5139), .B(n5138), .ZN(n5140) );
  OAI21_X1 U6285 ( .B1(n5322), .B2(n5785), .A(n5140), .ZN(U2798) );
  BUF_X1 U6286 ( .A(n5141), .Z(n5142) );
  OR2_X1 U6287 ( .A1(n5160), .A2(n5144), .ZN(n5145) );
  NAND2_X1 U6288 ( .A1(n5102), .A2(n5145), .ZN(n5518) );
  INV_X1 U6289 ( .A(n5146), .ZN(n5378) );
  OAI22_X1 U6290 ( .A1(n5147), .A2(n5821), .B1(n5848), .B2(n5378), .ZN(n5148)
         );
  AOI21_X1 U6291 ( .B1(n5831), .B2(EBX_REG_28__SCAN_IN), .A(n5148), .ZN(n5149)
         );
  OAI21_X1 U6292 ( .B1(n5518), .B2(n5849), .A(n5149), .ZN(n5152) );
  INV_X1 U6293 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6488) );
  NOR4_X1 U6294 ( .A1(n5630), .A2(n5150), .A3(REIP_REG_28__SCAN_IN), .A4(n6488), .ZN(n5151) );
  AOI211_X1 U6295 ( .C1(REIP_REG_28__SCAN_IN), .C2(n5153), .A(n5152), .B(n5151), .ZN(n5154) );
  OAI21_X1 U6296 ( .B1(n5376), .B2(n5785), .A(n5154), .ZN(U2799) );
  AOI21_X1 U6297 ( .B1(n5156), .B2(n5155), .A(n5142), .ZN(n5389) );
  INV_X1 U6298 ( .A(n5389), .ZN(n5327) );
  AOI22_X1 U6299 ( .A1(EBX_REG_27__SCAN_IN), .A2(n5831), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5843), .ZN(n5157) );
  OAI21_X1 U6300 ( .B1(n5387), .B2(n5848), .A(n5157), .ZN(n5162) );
  NOR2_X1 U6301 ( .A1(n5264), .A2(n5158), .ZN(n5159) );
  OR2_X1 U6302 ( .A1(n5160), .A2(n5159), .ZN(n5531) );
  NOR2_X1 U6303 ( .A1(n5531), .A2(n5849), .ZN(n5161) );
  AOI211_X1 U6304 ( .C1(n5636), .C2(REIP_REG_27__SCAN_IN), .A(n5162), .B(n5161), .ZN(n5165) );
  NAND2_X1 U6305 ( .A1(n5163), .A2(n6488), .ZN(n5164) );
  OAI211_X1 U6306 ( .C1(n5327), .C2(n5785), .A(n5165), .B(n5164), .ZN(U2800)
         );
  INV_X1 U6307 ( .A(n5166), .ZN(n5168) );
  AOI21_X1 U6308 ( .B1(n5168), .B2(n3035), .A(n5167), .ZN(n5416) );
  INV_X1 U6309 ( .A(n5416), .ZN(n5334) );
  INV_X1 U6310 ( .A(n5661), .ZN(n5641) );
  INV_X1 U6311 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6482) );
  INV_X1 U6312 ( .A(n5630), .ZN(n5647) );
  AOI22_X1 U6313 ( .A1(n5843), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .B1(n6482), 
        .B2(n5647), .ZN(n5169) );
  OAI21_X1 U6314 ( .B1(n5848), .B2(n5414), .A(n5169), .ZN(n5175) );
  OR2_X1 U6315 ( .A1(n5276), .A2(n5171), .ZN(n5172) );
  NAND2_X1 U6316 ( .A1(n5170), .A2(n5172), .ZN(n5552) );
  INV_X1 U6317 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5173) );
  OAI22_X1 U6318 ( .A1(n5552), .A2(n5849), .B1(n5173), .B2(n5851), .ZN(n5174)
         );
  AOI211_X1 U6319 ( .C1(n5641), .C2(REIP_REG_24__SCAN_IN), .A(n5175), .B(n5174), .ZN(n5176) );
  OAI21_X1 U6320 ( .B1(n5334), .B2(n5785), .A(n5176), .ZN(U2803) );
  INV_X1 U6321 ( .A(n3062), .ZN(n5190) );
  AOI21_X1 U6322 ( .B1(n3042), .B2(n5190), .A(n5178), .ZN(n5449) );
  INV_X1 U6323 ( .A(n5449), .ZN(n5346) );
  OAI211_X1 U6324 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5202), .B(n5179), .ZN(n5188) );
  NAND3_X1 U6325 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5193), .A3(n5192), .ZN(
        n5186) );
  AOI21_X1 U6326 ( .B1(n5843), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6000), 
        .ZN(n5185) );
  MUX2_X1 U6327 ( .A(n5293), .B(n5180), .S(n5296), .Z(n5195) );
  OR2_X1 U6328 ( .A1(n5208), .A2(n5195), .ZN(n5196) );
  XNOR2_X1 U6329 ( .A(n5196), .B(n5181), .ZN(n5600) );
  INV_X1 U6330 ( .A(n5600), .ZN(n5301) );
  AOI22_X1 U6331 ( .A1(n5832), .A2(n5301), .B1(n5831), .B2(EBX_REG_19__SCAN_IN), .ZN(n5184) );
  INV_X1 U6332 ( .A(n5447), .ZN(n5182) );
  NAND2_X1 U6333 ( .A1(n5776), .A2(n5182), .ZN(n5183) );
  AND4_X1 U6334 ( .A1(n5186), .A2(n5185), .A3(n5184), .A4(n5183), .ZN(n5187)
         );
  OAI211_X1 U6335 ( .C1(n5346), .C2(n5785), .A(n5188), .B(n5187), .ZN(U2808)
         );
  INV_X1 U6336 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U6337 ( .A1(n5193), .A2(n5192), .ZN(n5211) );
  AOI22_X1 U6338 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5831), .B1(n5451), .B2(n5776), .ZN(n5194) );
  OAI21_X1 U6339 ( .B1(n6473), .B2(n5211), .A(n5194), .ZN(n5201) );
  INV_X1 U6340 ( .A(n5208), .ZN(n5198) );
  INV_X1 U6341 ( .A(n5195), .ZN(n5197) );
  OAI21_X1 U6342 ( .B1(n5198), .B2(n5197), .A(n5196), .ZN(n5605) );
  AOI21_X1 U6343 ( .B1(n5843), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6000), 
        .ZN(n5199) );
  OAI21_X1 U6344 ( .B1(n5849), .B2(n5605), .A(n5199), .ZN(n5200) );
  AOI211_X1 U6345 ( .C1(n5202), .C2(n6473), .A(n5201), .B(n5200), .ZN(n5203)
         );
  OAI21_X1 U6346 ( .B1(n5452), .B2(n5785), .A(n5203), .ZN(U2809) );
  NAND2_X1 U6347 ( .A1(n5218), .A2(n5217), .ZN(n5216) );
  AOI21_X1 U6348 ( .B1(n5204), .B2(n5216), .A(n3088), .ZN(n5697) );
  INV_X1 U6349 ( .A(n5697), .ZN(n5351) );
  NAND2_X1 U6350 ( .A1(n5221), .A2(n5219), .ZN(n5207) );
  INV_X1 U6351 ( .A(n5205), .ZN(n5206) );
  NAND2_X1 U6352 ( .A1(n5207), .A2(n5206), .ZN(n5209) );
  AND2_X1 U6353 ( .A1(n5209), .A2(n5208), .ZN(n5703) );
  AOI22_X1 U6354 ( .A1(EBX_REG_17__SCAN_IN), .A2(n5831), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n5843), .ZN(n5210) );
  OAI211_X1 U6355 ( .C1(n5848), .C2(n5700), .A(n5210), .B(n5819), .ZN(n5214)
         );
  AOI21_X1 U6356 ( .B1(n6551), .B2(n5212), .A(n5211), .ZN(n5213) );
  AOI211_X1 U6357 ( .C1(n5703), .C2(n5832), .A(n5214), .B(n5213), .ZN(n5215)
         );
  OAI21_X1 U6358 ( .B1(n5351), .B2(n5785), .A(n5215), .ZN(U2810) );
  OAI21_X1 U6359 ( .B1(n5218), .B2(n5217), .A(n5216), .ZN(n5475) );
  INV_X1 U6360 ( .A(n5219), .ZN(n5220) );
  XNOR2_X1 U6361 ( .A(n5221), .B(n5220), .ZN(n5708) );
  INV_X1 U6362 ( .A(n5222), .ZN(n5472) );
  AOI21_X1 U6363 ( .B1(n5776), .B2(n5472), .A(n6000), .ZN(n5223) );
  OAI21_X1 U6364 ( .B1(n5821), .B2(n5470), .A(n5223), .ZN(n5229) );
  AOI22_X1 U6365 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5831), .B1(
        REIP_REG_16__SCAN_IN), .B2(n5235), .ZN(n5227) );
  NAND2_X1 U6366 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5224) );
  OAI211_X1 U6367 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n5225), .B(n5224), .ZN(n5226) );
  NAND2_X1 U6368 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  AOI211_X1 U6369 ( .C1(n5832), .C2(n5708), .A(n5229), .B(n5228), .ZN(n5230)
         );
  OAI21_X1 U6370 ( .B1(n5475), .B2(n5785), .A(n5230), .ZN(U2811) );
  INV_X1 U6371 ( .A(n3006), .ZN(n5234) );
  NAND3_X1 U6372 ( .A1(n5018), .A2(n5232), .A3(n5231), .ZN(n5233) );
  NAND2_X1 U6373 ( .A1(n5234), .A2(n5233), .ZN(n5498) );
  INV_X1 U6374 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6679) );
  AOI22_X1 U6375 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n5843), .B1(
        REIP_REG_14__SCAN_IN), .B2(n5235), .ZN(n5242) );
  AND2_X1 U6376 ( .A1(n5237), .A2(n5236), .ZN(n5238) );
  NOR2_X1 U6377 ( .A1(n5239), .A2(n5238), .ZN(n5717) );
  OAI21_X1 U6378 ( .B1(n5848), .B2(n5489), .A(n5819), .ZN(n5240) );
  AOI21_X1 U6379 ( .B1(n5832), .B2(n5717), .A(n5240), .ZN(n5241) );
  OAI211_X1 U6380 ( .C1(n6679), .C2(n5851), .A(n5242), .B(n5241), .ZN(n5245)
         );
  NOR3_X1 U6381 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5243), .A3(n5780), .ZN(n5244) );
  NOR2_X1 U6382 ( .A1(n5245), .A2(n5244), .ZN(n5246) );
  OAI21_X1 U6383 ( .B1(n5498), .B2(n5785), .A(n5246), .ZN(U2813) );
  OAI21_X1 U6384 ( .B1(n5843), .B2(n5776), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5247) );
  OAI21_X1 U6385 ( .B1(n5847), .B2(n6149), .A(n5247), .ZN(n5248) );
  AOI21_X1 U6386 ( .B1(n5249), .B2(n5854), .A(n5248), .ZN(n5252) );
  AOI22_X1 U6387 ( .A1(n5250), .A2(n5832), .B1(n5831), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5251) );
  OAI211_X1 U6388 ( .C1(n5253), .C2(n6513), .A(n5252), .B(n5251), .ZN(U2827)
         );
  INV_X1 U6389 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5254) );
  OAI22_X1 U6390 ( .A1(n5505), .A2(n5309), .B1(n5311), .B2(n5254), .ZN(U2828)
         );
  OAI222_X1 U6391 ( .A1(n5312), .A2(n5322), .B1(n5255), .B2(n5311), .C1(n5511), 
        .C2(n5309), .ZN(U2830) );
  OAI22_X1 U6392 ( .A1(n5518), .A2(n5309), .B1(n5256), .B2(n5311), .ZN(n5257)
         );
  INV_X1 U6393 ( .A(n5257), .ZN(n5258) );
  OAI21_X1 U6394 ( .B1(n5376), .B2(n5312), .A(n5258), .ZN(U2831) );
  INV_X1 U6395 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5259) );
  OAI222_X1 U6396 ( .A1(n5312), .A2(n5327), .B1(n5259), .B2(n5311), .C1(n5531), 
        .C2(n5309), .ZN(U2832) );
  OAI21_X1 U6397 ( .B1(n5260), .B2(n5261), .A(n5155), .ZN(n5633) );
  AND2_X1 U6398 ( .A1(n5270), .A2(n5262), .ZN(n5263) );
  NOR2_X1 U6399 ( .A1(n5264), .A2(n5263), .ZN(n5631) );
  AOI22_X1 U6400 ( .A1(n5631), .A2(n5306), .B1(EBX_REG_26__SCAN_IN), .B2(n5305), .ZN(n5265) );
  OAI21_X1 U6401 ( .B1(n5633), .B2(n5312), .A(n5265), .ZN(U2833) );
  NOR2_X1 U6402 ( .A1(n5167), .A2(n5266), .ZN(n5267) );
  INV_X1 U6403 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6404 ( .A1(n5170), .A2(n5268), .ZN(n5269) );
  NAND2_X1 U6405 ( .A1(n5270), .A2(n5269), .ZN(n5643) );
  OAI222_X1 U6406 ( .A1(n5644), .A2(n5312), .B1(n5271), .B2(n5311), .C1(n5309), 
        .C2(n5643), .ZN(U2834) );
  OAI222_X1 U6407 ( .A1(n5312), .A2(n5334), .B1(n5311), .B2(n5173), .C1(n5552), 
        .C2(n5309), .ZN(U2835) );
  INV_X1 U6408 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5277) );
  INV_X1 U6409 ( .A(n5272), .ZN(n5273) );
  AOI21_X1 U6410 ( .B1(n5289), .B2(n5274), .A(n5273), .ZN(n5275) );
  OR2_X1 U6411 ( .A1(n5276), .A2(n5275), .ZN(n5655) );
  OAI222_X1 U6412 ( .A1(n5312), .A2(n5654), .B1(n5277), .B2(n5311), .C1(n5655), 
        .C2(n5309), .ZN(U2836) );
  AOI21_X1 U6413 ( .B1(n5280), .B2(n5278), .A(n5279), .ZN(n5665) );
  INV_X1 U6414 ( .A(n5665), .ZN(n5339) );
  XNOR2_X1 U6415 ( .A(n5289), .B(n5281), .ZN(n5664) );
  AOI22_X1 U6416 ( .A1(n5664), .A2(n5306), .B1(EBX_REG_22__SCAN_IN), .B2(n5305), .ZN(n5282) );
  OAI21_X1 U6417 ( .B1(n5339), .B2(n5312), .A(n5282), .ZN(U2837) );
  NAND2_X1 U6418 ( .A1(n5283), .A2(n5284), .ZN(n5285) );
  NAND2_X1 U6419 ( .A1(n5278), .A2(n5285), .ZN(n5675) );
  INV_X1 U6420 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5290) );
  AND2_X1 U6421 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  NOR2_X1 U6422 ( .A1(n5289), .A2(n5288), .ZN(n5577) );
  INV_X1 U6423 ( .A(n5577), .ZN(n5674) );
  OAI222_X1 U6424 ( .A1(n5675), .A2(n5312), .B1(n5290), .B2(n5311), .C1(n5309), 
        .C2(n5674), .ZN(U2838) );
  OR2_X1 U6425 ( .A1(n5178), .A2(n5291), .ZN(n5292) );
  NAND2_X1 U6426 ( .A1(n5283), .A2(n5292), .ZN(n5684) );
  INV_X1 U6427 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5300) );
  INV_X1 U6428 ( .A(n5293), .ZN(n5297) );
  MUX2_X1 U6429 ( .A(n5297), .B(n5296), .S(n5295), .Z(n5299) );
  XNOR2_X1 U6430 ( .A(n5299), .B(n5298), .ZN(n5683) );
  OAI222_X1 U6431 ( .A1(n5684), .A2(n5312), .B1(n5311), .B2(n5300), .C1(n5683), 
        .C2(n5309), .ZN(U2839) );
  AOI22_X1 U6432 ( .A1(n5301), .A2(n5306), .B1(EBX_REG_19__SCAN_IN), .B2(n5305), .ZN(n5302) );
  OAI21_X1 U6433 ( .B1(n5346), .B2(n5312), .A(n5302), .ZN(U2840) );
  OAI222_X1 U6434 ( .A1(n5605), .A2(n5309), .B1(n5311), .B2(n4179), .C1(n5452), 
        .C2(n5312), .ZN(U2841) );
  INV_X1 U6435 ( .A(n5703), .ZN(n5303) );
  OAI222_X1 U6436 ( .A1(n5351), .A2(n5312), .B1(n5304), .B2(n5311), .C1(n5309), 
        .C2(n5303), .ZN(U2842) );
  AOI22_X1 U6437 ( .A1(n5708), .A2(n5306), .B1(EBX_REG_16__SCAN_IN), .B2(n5305), .ZN(n5307) );
  OAI21_X1 U6438 ( .B1(n5475), .B2(n5312), .A(n5307), .ZN(U2843) );
  OAI222_X1 U6439 ( .A1(n5620), .A2(n5309), .B1(n5308), .B2(n5311), .C1(n5479), 
        .C2(n5312), .ZN(U2844) );
  INV_X1 U6440 ( .A(n5717), .ZN(n5310) );
  OAI222_X1 U6441 ( .A1(n5498), .A2(n5312), .B1(n5311), .B2(n6679), .C1(n5310), 
        .C2(n5309), .ZN(U2845) );
  NAND3_X1 U6442 ( .A1(n5314), .A2(n5313), .A3(n5357), .ZN(n5316) );
  AOI22_X1 U6443 ( .A1(n5353), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5352), .ZN(n5315) );
  NAND2_X1 U6444 ( .A1(n5316), .A2(n5315), .ZN(U2860) );
  AOI22_X1 U6445 ( .A1(n5353), .A2(DATAI_30_), .B1(n5352), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6446 ( .A1(n5354), .A2(DATAI_14_), .ZN(n5317) );
  OAI211_X1 U6447 ( .C1(n5319), .C2(n5361), .A(n5318), .B(n5317), .ZN(U2861)
         );
  AOI22_X1 U6448 ( .A1(n5353), .A2(DATAI_29_), .B1(n5352), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6449 ( .A1(n5354), .A2(DATAI_13_), .ZN(n5320) );
  OAI211_X1 U6450 ( .C1(n5322), .C2(n5361), .A(n5321), .B(n5320), .ZN(U2862)
         );
  AOI22_X1 U6451 ( .A1(n5353), .A2(DATAI_28_), .B1(n5352), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6452 ( .A1(n5354), .A2(DATAI_12_), .ZN(n5323) );
  OAI211_X1 U6453 ( .C1(n5376), .C2(n5361), .A(n5324), .B(n5323), .ZN(U2863)
         );
  AOI22_X1 U6454 ( .A1(n5353), .A2(DATAI_27_), .B1(n5352), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6455 ( .A1(n5354), .A2(DATAI_11_), .ZN(n5325) );
  OAI211_X1 U6456 ( .C1(n5327), .C2(n5361), .A(n5326), .B(n5325), .ZN(U2864)
         );
  AOI22_X1 U6457 ( .A1(n5353), .A2(DATAI_26_), .B1(n5352), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6458 ( .A1(n5354), .A2(DATAI_10_), .ZN(n5328) );
  OAI211_X1 U6459 ( .C1(n5633), .C2(n5361), .A(n5329), .B(n5328), .ZN(U2865)
         );
  AOI22_X1 U6460 ( .A1(n5353), .A2(DATAI_25_), .B1(n5352), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6461 ( .A1(n5354), .A2(DATAI_9_), .ZN(n5330) );
  OAI211_X1 U6462 ( .C1(n5644), .C2(n5361), .A(n5331), .B(n5330), .ZN(U2866)
         );
  AOI22_X1 U6463 ( .A1(n5353), .A2(DATAI_24_), .B1(n5352), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6464 ( .A1(n5354), .A2(DATAI_8_), .ZN(n5332) );
  OAI211_X1 U6465 ( .C1(n5334), .C2(n5361), .A(n5333), .B(n5332), .ZN(U2867)
         );
  AOI22_X1 U6466 ( .A1(n5353), .A2(DATAI_23_), .B1(n5352), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6467 ( .A1(n5354), .A2(DATAI_7_), .ZN(n5335) );
  OAI211_X1 U6468 ( .C1(n5654), .C2(n5361), .A(n5336), .B(n5335), .ZN(U2868)
         );
  AOI22_X1 U6469 ( .A1(n5353), .A2(DATAI_22_), .B1(n5352), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6470 ( .A1(n5354), .A2(DATAI_6_), .ZN(n5337) );
  OAI211_X1 U6471 ( .C1(n5339), .C2(n5361), .A(n5338), .B(n5337), .ZN(U2869)
         );
  AOI22_X1 U6472 ( .A1(n5353), .A2(DATAI_21_), .B1(n5352), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6473 ( .A1(n5354), .A2(DATAI_5_), .ZN(n5340) );
  OAI211_X1 U6474 ( .C1(n5675), .C2(n5361), .A(n5341), .B(n5340), .ZN(U2870)
         );
  AOI22_X1 U6475 ( .A1(n5353), .A2(DATAI_20_), .B1(n5352), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6476 ( .A1(n5354), .A2(DATAI_4_), .ZN(n5342) );
  OAI211_X1 U6477 ( .C1(n5684), .C2(n5361), .A(n5343), .B(n5342), .ZN(U2871)
         );
  AOI22_X1 U6478 ( .A1(n5353), .A2(DATAI_19_), .B1(n5352), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U6479 ( .A1(n5354), .A2(DATAI_3_), .ZN(n5344) );
  OAI211_X1 U6480 ( .C1(n5346), .C2(n5361), .A(n5345), .B(n5344), .ZN(U2872)
         );
  AOI22_X1 U6481 ( .A1(n5353), .A2(DATAI_18_), .B1(n5352), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6482 ( .A1(n5354), .A2(DATAI_2_), .ZN(n5347) );
  OAI211_X1 U6483 ( .C1(n5452), .C2(n5361), .A(n5348), .B(n5347), .ZN(U2873)
         );
  AOI22_X1 U6484 ( .A1(n5353), .A2(DATAI_17_), .B1(n5352), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6485 ( .A1(n5354), .A2(DATAI_1_), .ZN(n5349) );
  OAI211_X1 U6486 ( .C1(n5351), .C2(n5361), .A(n5350), .B(n5349), .ZN(U2874)
         );
  AOI22_X1 U6487 ( .A1(n5353), .A2(DATAI_16_), .B1(n5352), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6488 ( .A1(n5354), .A2(DATAI_0_), .ZN(n5355) );
  OAI211_X1 U6489 ( .C1(n5475), .C2(n5361), .A(n5356), .B(n5355), .ZN(U2875)
         );
  INV_X1 U6490 ( .A(DATAI_14_), .ZN(n5360) );
  OAI222_X1 U6491 ( .A1(n5498), .A2(n5361), .B1(n5360), .B2(n5359), .C1(n5358), 
        .C2(n5357), .ZN(U2877) );
  NAND2_X1 U6492 ( .A1(n5362), .A2(n5371), .ZN(n5363) );
  XNOR2_X1 U6493 ( .A(n5363), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5517)
         );
  AND2_X1 U6494 ( .A1(n6000), .A2(REIP_REG_29__SCAN_IN), .ZN(n5513) );
  AOI21_X1 U6495 ( .B1(n5936), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5513), 
        .ZN(n5364) );
  OAI21_X1 U6496 ( .B1(n5946), .B2(n5365), .A(n5364), .ZN(n5366) );
  AOI21_X1 U6497 ( .B1(n5367), .B2(n5941), .A(n5366), .ZN(n5368) );
  OAI21_X1 U6498 ( .B1(n5517), .B2(n5753), .A(n5368), .ZN(U2957) );
  INV_X1 U6499 ( .A(n5383), .ZN(n5375) );
  NOR2_X1 U6500 ( .A1(n5369), .A2(n5392), .ZN(n5382) );
  INV_X1 U6501 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U6502 ( .A1(n6539), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5373) );
  NAND3_X1 U6503 ( .A1(n5383), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5370), .ZN(n5372) );
  OAI211_X1 U6504 ( .C1(n5382), .C2(n5373), .A(n5372), .B(n5371), .ZN(n5374)
         );
  INV_X1 U6505 ( .A(n5376), .ZN(n5380) );
  AND2_X1 U6506 ( .A1(n6000), .A2(REIP_REG_28__SCAN_IN), .ZN(n5522) );
  AOI21_X1 U6507 ( .B1(n5936), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5522), 
        .ZN(n5377) );
  OAI21_X1 U6508 ( .B1(n5946), .B2(n5378), .A(n5377), .ZN(n5379) );
  AOI21_X1 U6509 ( .B1(n5380), .B2(n5941), .A(n5379), .ZN(n5381) );
  OAI21_X1 U6510 ( .B1(n5527), .B2(n5753), .A(n5381), .ZN(U2958) );
  NOR2_X1 U6511 ( .A1(n5383), .A2(n5382), .ZN(n5384) );
  XNOR2_X1 U6512 ( .A(n5384), .B(n6539), .ZN(n5536) );
  NAND2_X1 U6513 ( .A1(n6000), .A2(REIP_REG_27__SCAN_IN), .ZN(n5530) );
  INV_X1 U6514 ( .A(n5530), .ZN(n5385) );
  AOI21_X1 U6515 ( .B1(n5936), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5385), 
        .ZN(n5386) );
  OAI21_X1 U6516 ( .B1(n5946), .B2(n5387), .A(n5386), .ZN(n5388) );
  AOI21_X1 U6517 ( .B1(n5389), .B2(n5941), .A(n5388), .ZN(n5390) );
  OAI21_X1 U6518 ( .B1(n5536), .B2(n5753), .A(n5390), .ZN(U2959) );
  NAND2_X1 U6519 ( .A1(n5392), .A2(n5391), .ZN(n5394) );
  XOR2_X1 U6520 ( .A(n5394), .B(n5393), .Z(n5544) );
  INV_X1 U6521 ( .A(n5633), .ZN(n5398) );
  INV_X1 U6522 ( .A(n5629), .ZN(n5396) );
  AND2_X1 U6523 ( .A1(n6000), .A2(REIP_REG_26__SCAN_IN), .ZN(n5541) );
  AOI21_X1 U6524 ( .B1(n5936), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5541), 
        .ZN(n5395) );
  OAI21_X1 U6525 ( .B1(n5946), .B2(n5396), .A(n5395), .ZN(n5397) );
  AOI21_X1 U6526 ( .B1(n5398), .B2(n5941), .A(n5397), .ZN(n5399) );
  OAI21_X1 U6527 ( .B1(n5544), .B2(n5753), .A(n5399), .ZN(U2960) );
  OAI21_X1 U6528 ( .B1(n5401), .B2(n5400), .A(n5369), .ZN(n5402) );
  INV_X1 U6529 ( .A(n5402), .ZN(n5550) );
  INV_X1 U6530 ( .A(n5644), .ZN(n5405) );
  AND2_X1 U6531 ( .A1(n6000), .A2(REIP_REG_25__SCAN_IN), .ZN(n5546) );
  AOI21_X1 U6532 ( .B1(n5936), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5546), 
        .ZN(n5403) );
  OAI21_X1 U6533 ( .B1(n5946), .B2(n5640), .A(n5403), .ZN(n5404) );
  AOI21_X1 U6534 ( .B1(n5405), .B2(n5941), .A(n5404), .ZN(n5406) );
  OAI21_X1 U6535 ( .B1(n5550), .B2(n5753), .A(n5406), .ZN(U2961) );
  NAND2_X2 U6536 ( .A1(n5428), .A2(n3081), .ZN(n5418) );
  OR2_X2 U6537 ( .A1(n5418), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5410)
         );
  INV_X1 U6538 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6698) );
  MUX2_X1 U6539 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .B(n6698), .S(n5467), 
        .Z(n5407) );
  NAND3_X1 U6540 ( .A1(n5410), .A2(n5409), .A3(n5408), .ZN(n5412) );
  XNOR2_X1 U6541 ( .A(n5412), .B(n5411), .ZN(n5557) );
  NAND2_X1 U6542 ( .A1(n6000), .A2(REIP_REG_24__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U6543 ( .A1(n5936), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5413)
         );
  OAI211_X1 U6544 ( .C1(n5946), .C2(n5414), .A(n5551), .B(n5413), .ZN(n5415)
         );
  AOI21_X1 U6545 ( .B1(n5416), .B2(n5941), .A(n5415), .ZN(n5417) );
  OAI21_X1 U6546 ( .B1(n5557), .B2(n5753), .A(n5417), .ZN(U2962) );
  INV_X1 U6547 ( .A(n5419), .ZN(n5420) );
  NOR2_X1 U6548 ( .A1(n5421), .A2(n5420), .ZN(n5422) );
  XNOR2_X1 U6549 ( .A(n5418), .B(n5422), .ZN(n5570) );
  INV_X1 U6550 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5423) );
  NOR2_X1 U6551 ( .A1(n5819), .A2(n5423), .ZN(n5568) );
  NOR2_X1 U6552 ( .A1(n5492), .A2(n5424), .ZN(n5425) );
  AOI211_X1 U6553 ( .C1(n5494), .C2(n5663), .A(n5568), .B(n5425), .ZN(n5427)
         );
  NAND2_X1 U6554 ( .A1(n5665), .A2(n5941), .ZN(n5426) );
  OAI211_X1 U6555 ( .C1(n5570), .C2(n5753), .A(n5427), .B(n5426), .ZN(U2964)
         );
  OAI21_X1 U6556 ( .B1(n5430), .B2(n5429), .A(n5428), .ZN(n5572) );
  NAND2_X1 U6557 ( .A1(n5572), .A2(n5940), .ZN(n5433) );
  INV_X1 U6558 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6478) );
  NOR2_X1 U6559 ( .A1(n5819), .A2(n6478), .ZN(n5576) );
  NOR2_X1 U6560 ( .A1(n5946), .A2(n5672), .ZN(n5431) );
  AOI211_X1 U6561 ( .C1(n5936), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5576), 
        .B(n5431), .ZN(n5432) );
  OAI211_X1 U6562 ( .C1(n5499), .C2(n5675), .A(n5433), .B(n5432), .ZN(U2965)
         );
  XNOR2_X1 U6563 ( .A(n5436), .B(n5435), .ZN(n5437) );
  XNOR2_X1 U6564 ( .A(n5445), .B(n5437), .ZN(n5595) );
  NAND2_X1 U6565 ( .A1(n6000), .A2(REIP_REG_20__SCAN_IN), .ZN(n5591) );
  OAI21_X1 U6566 ( .B1(n5492), .B2(n5690), .A(n5591), .ZN(n5439) );
  NOR2_X1 U6567 ( .A1(n5684), .A2(n5499), .ZN(n5438) );
  AOI211_X1 U6568 ( .C1(n5494), .C2(n5681), .A(n5439), .B(n5438), .ZN(n5440)
         );
  OAI21_X1 U6569 ( .B1(n5595), .B2(n5753), .A(n5440), .ZN(U2966) );
  OR2_X1 U6570 ( .A1(n4086), .A2(n5442), .ZN(n5443) );
  AOI22_X1 U6571 ( .A1(n5445), .A2(n5444), .B1(n5441), .B2(n5443), .ZN(n5604)
         );
  NAND2_X1 U6572 ( .A1(n6000), .A2(REIP_REG_19__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U6573 ( .A1(n5936), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5446)
         );
  OAI211_X1 U6574 ( .C1(n5946), .C2(n5447), .A(n5598), .B(n5446), .ZN(n5448)
         );
  AOI21_X1 U6575 ( .B1(n5449), .B2(n5941), .A(n5448), .ZN(n5450) );
  OAI21_X1 U6576 ( .B1(n5604), .B2(n5753), .A(n5450), .ZN(U2967) );
  INV_X1 U6577 ( .A(n5451), .ZN(n5465) );
  INV_X1 U6578 ( .A(n5452), .ZN(n5453) );
  NAND2_X1 U6579 ( .A1(n5453), .A2(n5941), .ZN(n5464) );
  INV_X1 U6580 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5613) );
  AND2_X1 U6581 ( .A1(n5436), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5455)
         );
  INV_X1 U6582 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U6583 ( .A1(n5587), .A2(n5457), .ZN(n5458) );
  OR3_X1 U6584 ( .A1(n5456), .A2(n5436), .A3(n5458), .ZN(n5694) );
  INV_X1 U6585 ( .A(n5694), .ZN(n5459) );
  NOR2_X1 U6586 ( .A1(n5695), .A2(n5459), .ZN(n5460) );
  XOR2_X1 U6587 ( .A(n5613), .B(n5460), .Z(n5610) );
  INV_X1 U6588 ( .A(n5610), .ZN(n5461) );
  NAND2_X1 U6589 ( .A1(n6000), .A2(REIP_REG_18__SCAN_IN), .ZN(n5606) );
  OAI21_X1 U6590 ( .B1(n5753), .B2(n5461), .A(n5606), .ZN(n5462) );
  AOI21_X1 U6591 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n5936), .A(n5462), 
        .ZN(n5463) );
  OAI211_X1 U6592 ( .C1(n5465), .C2(n5946), .A(n5464), .B(n5463), .ZN(U2968)
         );
  MUX2_X1 U6593 ( .A(n5457), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .S(n5467), 
        .Z(n5468) );
  XNOR2_X1 U6594 ( .A(n5466), .B(n5468), .ZN(n5709) );
  NAND2_X1 U6595 ( .A1(n5709), .A2(n5940), .ZN(n5474) );
  INV_X1 U6596 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5469) );
  OAI22_X1 U6597 ( .A1(n5492), .A2(n5470), .B1(n5819), .B2(n5469), .ZN(n5471)
         );
  AOI21_X1 U6598 ( .B1(n5472), .B2(n5494), .A(n5471), .ZN(n5473) );
  OAI211_X1 U6599 ( .C1(n5499), .C2(n5475), .A(n5474), .B(n5473), .ZN(U2970)
         );
  INV_X1 U6600 ( .A(n5456), .ZN(n5477) );
  AOI21_X1 U6601 ( .B1(n5478), .B2(n3014), .A(n5477), .ZN(n5624) );
  NAND2_X1 U6602 ( .A1(n6000), .A2(REIP_REG_15__SCAN_IN), .ZN(n5619) );
  OAI21_X1 U6603 ( .B1(n5492), .B2(n5080), .A(n5619), .ZN(n5481) );
  NOR2_X1 U6604 ( .A1(n5479), .A2(n5499), .ZN(n5480) );
  AOI211_X1 U6605 ( .C1(n5494), .C2(n5482), .A(n5481), .B(n5480), .ZN(n5483)
         );
  OAI21_X1 U6606 ( .B1(n5624), .B2(n5753), .A(n5483), .ZN(U2971) );
  INV_X1 U6607 ( .A(n5485), .ZN(n5487) );
  NOR2_X1 U6608 ( .A1(n5487), .A2(n5486), .ZN(n5488) );
  XNOR2_X1 U6609 ( .A(n5484), .B(n5488), .ZN(n5718) );
  NAND2_X1 U6610 ( .A1(n5718), .A2(n5940), .ZN(n5497) );
  INV_X1 U6611 ( .A(n5489), .ZN(n5495) );
  INV_X1 U6612 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5490) );
  OAI22_X1 U6613 ( .A1(n5492), .A2(n5491), .B1(n5819), .B2(n5490), .ZN(n5493)
         );
  AOI21_X1 U6614 ( .B1(n5495), .B2(n5494), .A(n5493), .ZN(n5496) );
  OAI211_X1 U6615 ( .C1(n5499), .C2(n5498), .A(n5497), .B(n5496), .ZN(U2972)
         );
  OAI21_X1 U6616 ( .B1(n5615), .B2(n5500), .A(n5529), .ZN(n5504) );
  INV_X1 U6617 ( .A(n5500), .ZN(n5501) );
  NOR3_X1 U6618 ( .A1(n5528), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5501), 
        .ZN(n5502) );
  AOI211_X1 U6619 ( .C1(INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n5504), .A(n5503), .B(n5502), .ZN(n5508) );
  INV_X1 U6620 ( .A(n5505), .ZN(n5506) );
  NAND2_X1 U6621 ( .A1(n5506), .A2(n6010), .ZN(n5507) );
  OAI211_X1 U6622 ( .C1(n5509), .C2(n5623), .A(n5508), .B(n5507), .ZN(U2987)
         );
  OAI21_X1 U6623 ( .B1(n5528), .B2(n5510), .A(n3515), .ZN(n5514) );
  NOR2_X1 U6624 ( .A1(n5511), .A2(n5967), .ZN(n5512) );
  AOI211_X1 U6625 ( .C1(n5515), .C2(n5514), .A(n5513), .B(n5512), .ZN(n5516)
         );
  OAI21_X1 U6626 ( .B1(n5517), .B2(n5623), .A(n5516), .ZN(U2989) );
  INV_X1 U6627 ( .A(n5518), .ZN(n5523) );
  NOR3_X1 U6628 ( .A1(n5528), .A2(n5520), .A3(n5519), .ZN(n5521) );
  AOI211_X1 U6629 ( .C1(n5523), .C2(n6010), .A(n5522), .B(n5521), .ZN(n5526)
         );
  INV_X1 U6630 ( .A(n5529), .ZN(n5524) );
  NAND2_X1 U6631 ( .A1(n5524), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5525) );
  OAI211_X1 U6632 ( .C1(n5527), .C2(n5623), .A(n5526), .B(n5525), .ZN(U2990)
         );
  INV_X1 U6633 ( .A(n5528), .ZN(n5534) );
  NOR2_X1 U6634 ( .A1(n5529), .A2(n6539), .ZN(n5533) );
  OAI21_X1 U6635 ( .B1(n5531), .B2(n5967), .A(n5530), .ZN(n5532) );
  AOI211_X1 U6636 ( .C1(n5534), .C2(n6539), .A(n5533), .B(n5532), .ZN(n5535)
         );
  OAI21_X1 U6637 ( .B1(n5536), .B2(n5623), .A(n5535), .ZN(U2991) );
  INV_X1 U6638 ( .A(n5547), .ZN(n5537) );
  AOI211_X1 U6639 ( .C1(n3517), .C2(n5539), .A(n5538), .B(n5537), .ZN(n5540)
         );
  AOI211_X1 U6640 ( .C1(n6010), .C2(n5631), .A(n5541), .B(n5540), .ZN(n5543)
         );
  NAND2_X1 U6641 ( .A1(n5555), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5542) );
  OAI211_X1 U6642 ( .C1(n5544), .C2(n5623), .A(n5543), .B(n5542), .ZN(U2992)
         );
  NOR2_X1 U6643 ( .A1(n5643), .A2(n5967), .ZN(n5545) );
  AOI211_X1 U6644 ( .C1(n5547), .C2(n3517), .A(n5546), .B(n5545), .ZN(n5549)
         );
  NAND2_X1 U6645 ( .A1(n5555), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5548) );
  OAI211_X1 U6646 ( .C1(n5550), .C2(n5623), .A(n5549), .B(n5548), .ZN(U2993)
         );
  OAI21_X1 U6647 ( .B1(n5559), .B2(n6698), .A(n5411), .ZN(n5554) );
  OAI21_X1 U6648 ( .B1(n5552), .B2(n5967), .A(n5551), .ZN(n5553) );
  AOI21_X1 U6649 ( .B1(n5555), .B2(n5554), .A(n5553), .ZN(n5556) );
  OAI21_X1 U6650 ( .B1(n5557), .B2(n5623), .A(n5556), .ZN(U2994) );
  NAND2_X1 U6651 ( .A1(n5558), .A2(n6021), .ZN(n5564) );
  NOR2_X1 U6652 ( .A1(n5559), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5562)
         );
  OAI21_X1 U6653 ( .B1(n5655), .B2(n5967), .A(n5560), .ZN(n5561) );
  NOR2_X1 U6654 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  OAI211_X1 U6655 ( .C1(n5566), .C2(n6698), .A(n5564), .B(n5563), .ZN(U2995)
         );
  AOI21_X1 U6656 ( .B1(n5571), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5565) );
  NOR2_X1 U6657 ( .A1(n5566), .A2(n5565), .ZN(n5567) );
  AOI211_X1 U6658 ( .C1(n6010), .C2(n5664), .A(n5568), .B(n5567), .ZN(n5569)
         );
  OAI21_X1 U6659 ( .B1(n5570), .B2(n5623), .A(n5569), .ZN(U2996) );
  INV_X1 U6660 ( .A(n5571), .ZN(n5580) );
  NAND2_X1 U6661 ( .A1(n5572), .A2(n6021), .ZN(n5579) );
  NOR2_X1 U6662 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  AOI211_X1 U6663 ( .C1(n6010), .C2(n5577), .A(n5576), .B(n5575), .ZN(n5578)
         );
  OAI211_X1 U6664 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5580), .A(n5579), .B(n5578), .ZN(U2997) );
  AOI21_X1 U6665 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5581), .A(n5721), 
        .ZN(n5583) );
  AOI211_X1 U6666 ( .C1(n5586), .C2(n5584), .A(n5583), .B(n5582), .ZN(n5701)
         );
  INV_X1 U6667 ( .A(n5701), .ZN(n5585) );
  AOI21_X1 U6668 ( .B1(n5587), .B2(n5586), .A(n5585), .ZN(n5614) );
  OAI21_X1 U6669 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5615), .A(n5614), 
        .ZN(n5602) );
  NAND2_X1 U6670 ( .A1(n5949), .A2(n5588), .ZN(n5707) );
  NOR2_X1 U6671 ( .A1(n5707), .A2(n5589), .ZN(n5597) );
  XNOR2_X1 U6672 ( .A(n5596), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5590)
         );
  NAND2_X1 U6673 ( .A1(n5597), .A2(n5590), .ZN(n5592) );
  OAI211_X1 U6674 ( .C1(n5967), .C2(n5683), .A(n5592), .B(n5591), .ZN(n5593)
         );
  AOI21_X1 U6675 ( .B1(n5602), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5593), 
        .ZN(n5594) );
  OAI21_X1 U6676 ( .B1(n5595), .B2(n5623), .A(n5594), .ZN(U2998) );
  NAND2_X1 U6677 ( .A1(n5597), .A2(n5596), .ZN(n5599) );
  OAI211_X1 U6678 ( .C1(n5600), .C2(n5967), .A(n5599), .B(n5598), .ZN(n5601)
         );
  AOI21_X1 U6679 ( .B1(n5602), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5601), 
        .ZN(n5603) );
  OAI21_X1 U6680 ( .B1(n5604), .B2(n5623), .A(n5603), .ZN(U2999) );
  INV_X1 U6681 ( .A(n5605), .ZN(n5609) );
  INV_X1 U6682 ( .A(n5606), .ZN(n5608) );
  NOR3_X1 U6683 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5587), .A3(n5707), 
        .ZN(n5607) );
  AOI211_X1 U6684 ( .C1(n5609), .C2(n6010), .A(n5608), .B(n5607), .ZN(n5612)
         );
  NAND2_X1 U6685 ( .A1(n6021), .A2(n5610), .ZN(n5611) );
  OAI211_X1 U6686 ( .C1(n5614), .C2(n5613), .A(n5612), .B(n5611), .ZN(U3000)
         );
  OAI21_X1 U6687 ( .B1(n5615), .B2(n5616), .A(n5954), .ZN(n5710) );
  AND3_X1 U6688 ( .A1(n5617), .A2(n5949), .A3(n5616), .ZN(n5711) );
  INV_X1 U6689 ( .A(n5711), .ZN(n5618) );
  OAI211_X1 U6690 ( .C1(n5967), .C2(n5620), .A(n5619), .B(n5618), .ZN(n5621)
         );
  AOI21_X1 U6691 ( .B1(n5710), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5621), 
        .ZN(n5622) );
  OAI21_X1 U6692 ( .B1(n5624), .B2(n5623), .A(n5622), .ZN(U3003) );
  INV_X1 U6693 ( .A(n5625), .ZN(n5626) );
  OAI22_X1 U6694 ( .A1(n5627), .A2(n6510), .B1(n5626), .B2(n6412), .ZN(n5628)
         );
  MUX2_X1 U6695 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5628), .S(n6508), 
        .Z(U3456) );
  AND2_X1 U6696 ( .A1(n5887), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6697 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n5843), .B1(n5629), 
        .B2(n5776), .ZN(n5638) );
  NAND2_X1 U6698 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5646) );
  INV_X1 U6699 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6486) );
  OAI21_X1 U6700 ( .B1(n5646), .B2(n5630), .A(n6486), .ZN(n5635) );
  INV_X1 U6701 ( .A(n5631), .ZN(n5632) );
  OAI22_X1 U6702 ( .A1(n5633), .A2(n5785), .B1(n5632), .B2(n5849), .ZN(n5634)
         );
  AOI21_X1 U6703 ( .B1(n5636), .B2(n5635), .A(n5634), .ZN(n5637) );
  OAI211_X1 U6704 ( .C1(n5639), .C2(n5851), .A(n5638), .B(n5637), .ZN(U2801)
         );
  AOI22_X1 U6705 ( .A1(EBX_REG_25__SCAN_IN), .A2(n5831), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5843), .ZN(n5651) );
  INV_X1 U6706 ( .A(n5640), .ZN(n5642) );
  AOI22_X1 U6707 ( .A1(n5642), .A2(n5776), .B1(REIP_REG_25__SCAN_IN), .B2(
        n5641), .ZN(n5650) );
  OAI22_X1 U6708 ( .A1(n5644), .A2(n5785), .B1(n5849), .B2(n5643), .ZN(n5645)
         );
  INV_X1 U6709 ( .A(n5645), .ZN(n5649) );
  OAI211_X1 U6710 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5647), .B(n5646), .ZN(n5648) );
  NAND4_X1 U6711 ( .A1(n5651), .A2(n5650), .A3(n5649), .A4(n5648), .ZN(U2802)
         );
  AND2_X1 U6712 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5666), .ZN(n5662) );
  AOI21_X1 U6713 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5662), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5660) );
  OAI22_X1 U6714 ( .A1(n4095), .A2(n5821), .B1(n5652), .B2(n5848), .ZN(n5653)
         );
  AOI21_X1 U6715 ( .B1(EBX_REG_23__SCAN_IN), .B2(n5831), .A(n5653), .ZN(n5659)
         );
  INV_X1 U6716 ( .A(n5654), .ZN(n5657) );
  INV_X1 U6717 ( .A(n5785), .ZN(n5803) );
  INV_X1 U6718 ( .A(n5655), .ZN(n5656) );
  AOI22_X1 U6719 ( .A1(n5657), .A2(n5803), .B1(n5656), .B2(n5832), .ZN(n5658)
         );
  OAI211_X1 U6720 ( .C1(n5661), .C2(n5660), .A(n5659), .B(n5658), .ZN(U2804)
         );
  AOI22_X1 U6721 ( .A1(EBX_REG_22__SCAN_IN), .A2(n5831), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n5843), .ZN(n5671) );
  AOI22_X1 U6722 ( .A1(n5663), .A2(n5776), .B1(n5662), .B2(n5423), .ZN(n5670)
         );
  AOI22_X1 U6723 ( .A1(n5665), .A2(n5803), .B1(n5832), .B2(n5664), .ZN(n5669)
         );
  NAND2_X1 U6724 ( .A1(n6478), .A2(n5666), .ZN(n5677) );
  INV_X1 U6725 ( .A(n5677), .ZN(n5667) );
  OAI21_X1 U6726 ( .B1(n5687), .B2(n5667), .A(REIP_REG_22__SCAN_IN), .ZN(n5668) );
  NAND4_X1 U6727 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), .ZN(U2805)
         );
  AOI22_X1 U6728 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5831), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5843), .ZN(n5680) );
  INV_X1 U6729 ( .A(n5672), .ZN(n5673) );
  AOI22_X1 U6730 ( .A1(n5673), .A2(n5776), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5687), .ZN(n5679) );
  OAI22_X1 U6731 ( .A1(n5675), .A2(n5785), .B1(n5849), .B2(n5674), .ZN(n5676)
         );
  INV_X1 U6732 ( .A(n5676), .ZN(n5678) );
  NAND4_X1 U6733 ( .A1(n5680), .A2(n5679), .A3(n5678), .A4(n5677), .ZN(U2806)
         );
  AOI22_X1 U6734 ( .A1(EBX_REG_20__SCAN_IN), .A2(n5831), .B1(n5681), .B2(n5776), .ZN(n5689) );
  NAND2_X1 U6735 ( .A1(n5682), .A2(n6476), .ZN(n5686) );
  OAI22_X1 U6736 ( .A1(n5684), .A2(n5785), .B1(n5849), .B2(n5683), .ZN(n5685)
         );
  AOI21_X1 U6737 ( .B1(n5687), .B2(n5686), .A(n5685), .ZN(n5688) );
  OAI211_X1 U6738 ( .C1(n5690), .C2(n5821), .A(n5689), .B(n5688), .ZN(U2807)
         );
  AOI22_X1 U6739 ( .A1(n6000), .A2(REIP_REG_17__SCAN_IN), .B1(n5936), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U6740 ( .A1(n5691), .A2(n5587), .ZN(n5693) );
  NAND2_X1 U6741 ( .A1(n5691), .A2(n5457), .ZN(n5692) );
  AOI22_X1 U6742 ( .A1(n5454), .A2(n5693), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5692), .ZN(n5696) );
  OAI21_X1 U6743 ( .B1(n5696), .B2(n5695), .A(n5694), .ZN(n5704) );
  AOI22_X1 U6744 ( .A1(n5704), .A2(n5940), .B1(n5941), .B2(n5697), .ZN(n5698)
         );
  OAI211_X1 U6745 ( .C1(n5946), .C2(n5700), .A(n5699), .B(n5698), .ZN(U2969)
         );
  OAI22_X1 U6746 ( .A1(n5587), .A2(n5701), .B1(n5819), .B2(n6551), .ZN(n5702)
         );
  INV_X1 U6747 ( .A(n5702), .ZN(n5706) );
  AOI22_X1 U6748 ( .A1(n5704), .A2(n6021), .B1(n6010), .B2(n5703), .ZN(n5705)
         );
  OAI211_X1 U6749 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5707), .A(n5706), .B(n5705), .ZN(U3001) );
  AOI22_X1 U6750 ( .A1(n5709), .A2(n6021), .B1(n6010), .B2(n5708), .ZN(n5716)
         );
  NAND2_X1 U6751 ( .A1(n6000), .A2(REIP_REG_16__SCAN_IN), .ZN(n5715) );
  OAI21_X1 U6752 ( .B1(n5711), .B2(n5710), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n5714) );
  NAND3_X1 U6753 ( .A1(n5712), .A2(n5457), .A3(n5949), .ZN(n5713) );
  NAND4_X1 U6754 ( .A1(n5716), .A2(n5715), .A3(n5714), .A4(n5713), .ZN(U3002)
         );
  AOI22_X1 U6755 ( .A1(n5718), .A2(n6021), .B1(n6010), .B2(n5717), .ZN(n5732)
         );
  NAND2_X1 U6756 ( .A1(n6000), .A2(REIP_REG_14__SCAN_IN), .ZN(n5731) );
  NAND3_X1 U6757 ( .A1(n5719), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n5725), 
        .ZN(n5723) );
  OR2_X1 U6758 ( .A1(n5721), .A2(n5720), .ZN(n5722) );
  AOI211_X1 U6759 ( .C1(n5723), .C2(n5722), .A(INSTADDRPOINTER_REG_13__SCAN_IN), .B(n5724), .ZN(n5736) );
  INV_X1 U6760 ( .A(n5724), .ZN(n5728) );
  NAND2_X1 U6761 ( .A1(n5728), .A2(n5725), .ZN(n5734) );
  OAI21_X1 U6762 ( .B1(n3499), .B2(n5734), .A(n5726), .ZN(n5733) );
  OAI211_X1 U6763 ( .C1(n5728), .C2(n5727), .A(n5954), .B(n5733), .ZN(n5739)
         );
  OAI21_X1 U6764 ( .B1(n5736), .B2(n5739), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5730) );
  NAND4_X1 U6765 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5728), .A3(n6577), .A4(n5949), .ZN(n5729) );
  NAND4_X1 U6766 ( .A1(n5732), .A2(n5731), .A3(n5730), .A4(n5729), .ZN(U3004)
         );
  OAI22_X1 U6767 ( .A1(n5819), .A2(n6463), .B1(n5734), .B2(n5733), .ZN(n5735)
         );
  AOI211_X1 U6768 ( .C1(n5737), .C2(n6021), .A(n5736), .B(n5735), .ZN(n5741)
         );
  AOI22_X1 U6769 ( .A1(n5739), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .B1(n6010), .B2(n5738), .ZN(n5740) );
  NAND2_X1 U6770 ( .A1(n5741), .A2(n5740), .ZN(U3005) );
  AOI21_X1 U6771 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6446), .A(n6437), .ZN(n5748) );
  INV_X1 U6772 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5742) );
  AOI21_X1 U6773 ( .B1(n5748), .B2(n5742), .A(n6464), .ZN(U2789) );
  INV_X1 U6774 ( .A(n5743), .ZN(n6397) );
  OAI22_X1 U6775 ( .A1(n6397), .A2(n5745), .B1(n4238), .B2(n5744), .ZN(n5752)
         );
  OAI21_X1 U6776 ( .B1(n5752), .B2(n6418), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5746) );
  OAI21_X1 U6777 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6419), .A(n5746), .ZN(
        U2790) );
  INV_X2 U6778 ( .A(n6464), .ZN(n6537) );
  NOR2_X1 U6779 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5749) );
  OAI21_X1 U6780 ( .B1(n5749), .B2(D_C_N_REG_SCAN_IN), .A(n6537), .ZN(n5747)
         );
  OAI21_X1 U6781 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6537), .A(n5747), .ZN(
        U2791) );
  NOR2_X1 U6782 ( .A1(n6464), .A2(n5748), .ZN(n6498) );
  OAI21_X1 U6783 ( .B1(BS16_N), .B2(n5749), .A(n6498), .ZN(n6497) );
  OAI21_X1 U6784 ( .B1(n6498), .B2(n5750), .A(n6497), .ZN(U2792) );
  AOI21_X1 U6785 ( .B1(n5751), .B2(n6434), .A(READY_N), .ZN(n6530) );
  NOR2_X1 U6786 ( .A1(n5752), .A2(n6530), .ZN(n6398) );
  NOR2_X1 U6787 ( .A1(n6398), .A2(n6418), .ZN(n6525) );
  OAI21_X1 U6788 ( .B1(n6525), .B2(n5754), .A(n5753), .ZN(U2793) );
  NOR4_X1 U6789 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5758) );
  NOR4_X1 U6790 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n5757) );
  NOR4_X1 U6791 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5756) );
  NOR4_X1 U6792 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5755) );
  NAND4_X1 U6793 ( .A1(n5758), .A2(n5757), .A3(n5756), .A4(n5755), .ZN(n5764)
         );
  NOR4_X1 U6794 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n5762) );
  AOI211_X1 U6795 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_17__SCAN_IN), .B(
        DATAWIDTH_REG_12__SCAN_IN), .ZN(n5761) );
  NOR4_X1 U6796 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n5760)
         );
  NOR4_X1 U6797 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n5759) );
  NAND4_X1 U6798 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n5763)
         );
  NOR2_X1 U6799 ( .A1(n5764), .A2(n5763), .ZN(n6518) );
  INV_X1 U6800 ( .A(n6518), .ZN(n5767) );
  NAND2_X1 U6801 ( .A1(n6518), .A2(n6513), .ZN(n6514) );
  NOR3_X1 U6802 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(n6514), .ZN(n5766) );
  AOI21_X1 U6803 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n5767), .A(n5766), .ZN(
        n5765) );
  OAI21_X1 U6804 ( .B1(n6515), .B2(n5767), .A(n5765), .ZN(U2794) );
  NAND2_X1 U6805 ( .A1(n6518), .A2(n6515), .ZN(n6519) );
  AOI21_X1 U6806 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(n5767), .A(n5766), .ZN(
        n5768) );
  OAI21_X1 U6807 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(n6519), .A(n5768), .ZN(
        U2795) );
  NAND2_X1 U6808 ( .A1(n5832), .A2(n5769), .ZN(n5770) );
  OAI211_X1 U6809 ( .C1(n5821), .C2(n5771), .A(n5770), .B(n5819), .ZN(n5772)
         );
  AOI21_X1 U6810 ( .B1(n5831), .B2(EBX_REG_12__SCAN_IN), .A(n5772), .ZN(n5773)
         );
  OAI21_X1 U6811 ( .B1(n5774), .B2(n5785), .A(n5773), .ZN(n5775) );
  AOI21_X1 U6812 ( .B1(n5777), .B2(n5776), .A(n5775), .ZN(n5778) );
  OAI221_X1 U6813 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5780), .C1(n6465), .C2(
        n5779), .A(n5778), .ZN(U2815) );
  OAI22_X1 U6814 ( .A1(n5851), .A2(n6543), .B1(n5849), .B2(n5781), .ZN(n5782)
         );
  AOI211_X1 U6815 ( .C1(n5843), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6000), 
        .B(n5782), .ZN(n5794) );
  INV_X1 U6816 ( .A(n5783), .ZN(n5784) );
  OAI22_X1 U6817 ( .A1(n5786), .A2(n5785), .B1(n5848), .B2(n5784), .ZN(n5787)
         );
  INV_X1 U6818 ( .A(n5787), .ZN(n5793) );
  OAI21_X1 U6819 ( .B1(n5789), .B2(n5788), .A(REIP_REG_10__SCAN_IN), .ZN(n5792) );
  NAND3_X1 U6820 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5790), .A3(n6460), .ZN(n5791) );
  NAND4_X1 U6821 ( .A1(n5794), .A2(n5793), .A3(n5792), .A4(n5791), .ZN(U2817)
         );
  OR2_X1 U6822 ( .A1(n5849), .A2(n5795), .ZN(n5801) );
  NOR2_X1 U6823 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5796), .ZN(n5797) );
  NAND2_X1 U6824 ( .A1(n5817), .A2(n5797), .ZN(n5800) );
  AOI21_X1 U6825 ( .B1(n5843), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6000), 
        .ZN(n5799) );
  NAND2_X1 U6826 ( .A1(n5831), .A2(EBX_REG_7__SCAN_IN), .ZN(n5798) );
  NAND4_X1 U6827 ( .A1(n5801), .A2(n5800), .A3(n5799), .A4(n5798), .ZN(n5802)
         );
  AOI21_X1 U6828 ( .B1(n5915), .B2(n5803), .A(n5802), .ZN(n5806) );
  OAI21_X1 U6829 ( .B1(n5811), .B2(n5804), .A(REIP_REG_7__SCAN_IN), .ZN(n5805)
         );
  OAI211_X1 U6830 ( .C1(n5848), .C2(n5918), .A(n5806), .B(n5805), .ZN(U2820)
         );
  OAI22_X1 U6831 ( .A1(n5807), .A2(n5821), .B1(n5849), .B2(n5981), .ZN(n5808)
         );
  AOI211_X1 U6832 ( .C1(n5831), .C2(EBX_REG_5__SCAN_IN), .A(n6000), .B(n5808), 
        .ZN(n5813) );
  OAI21_X1 U6833 ( .B1(n5833), .B2(n5809), .A(n6453), .ZN(n5810) );
  AOI22_X1 U6834 ( .A1(n5811), .A2(n5810), .B1(n5923), .B2(n5854), .ZN(n5812)
         );
  OAI211_X1 U6835 ( .C1(n5926), .C2(n5848), .A(n5813), .B(n5812), .ZN(U2822)
         );
  INV_X1 U6836 ( .A(n5847), .ZN(n5815) );
  AOI22_X1 U6837 ( .A1(n5832), .A2(n5992), .B1(n5815), .B2(n5814), .ZN(n5829)
         );
  INV_X1 U6838 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5820) );
  INV_X1 U6839 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6450) );
  NAND3_X1 U6840 ( .A1(n5817), .A2(n5816), .A3(n6450), .ZN(n5818) );
  OAI211_X1 U6841 ( .C1(n5821), .C2(n5820), .A(n5819), .B(n5818), .ZN(n5826)
         );
  OAI22_X1 U6842 ( .A1(n5824), .A2(n5823), .B1(n5822), .B2(n5848), .ZN(n5825)
         );
  AOI211_X1 U6843 ( .C1(REIP_REG_4__SCAN_IN), .C2(n5827), .A(n5826), .B(n5825), 
        .ZN(n5828) );
  OAI211_X1 U6844 ( .C1(n5830), .C2(n5851), .A(n5829), .B(n5828), .ZN(U2823)
         );
  AOI22_X1 U6845 ( .A1(n5832), .A2(n6009), .B1(n5831), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5842) );
  OAI21_X1 U6846 ( .B1(n5833), .B2(n6515), .A(n6448), .ZN(n5834) );
  NAND2_X1 U6847 ( .A1(n5835), .A2(n5834), .ZN(n5840) );
  NAND2_X1 U6848 ( .A1(n5843), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5836)
         );
  OAI21_X1 U6849 ( .B1(n5847), .B2(n4481), .A(n5836), .ZN(n5837) );
  INV_X1 U6850 ( .A(n5837), .ZN(n5839) );
  NAND2_X1 U6851 ( .A1(n5854), .A2(n5942), .ZN(n5838) );
  AND3_X1 U6852 ( .A1(n5840), .A2(n5839), .A3(n5838), .ZN(n5841) );
  OAI211_X1 U6853 ( .C1(n5945), .C2(n5848), .A(n5842), .B(n5841), .ZN(U2825)
         );
  NAND2_X1 U6854 ( .A1(n5843), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5844)
         );
  AND2_X1 U6855 ( .A1(n5845), .A2(n5844), .ZN(n5857) );
  INV_X1 U6856 ( .A(n5846), .ZN(n5855) );
  OAI22_X1 U6857 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n5848), .B1(n5847), 
        .B2(n6120), .ZN(n5853) );
  INV_X1 U6858 ( .A(n4327), .ZN(n5850) );
  OAI22_X1 U6859 ( .A1(n5851), .A2(n4117), .B1(n5850), .B2(n5849), .ZN(n5852)
         );
  AOI211_X1 U6860 ( .C1(n5855), .C2(n5854), .A(n5853), .B(n5852), .ZN(n5856)
         );
  OAI211_X1 U6861 ( .C1(n5858), .C2(n6515), .A(n5857), .B(n5856), .ZN(U2826)
         );
  INV_X1 U6862 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n5861) );
  INV_X1 U6863 ( .A(n5859), .ZN(n5864) );
  AOI22_X1 U6864 ( .A1(n5887), .A2(DATAO_REG_30__SCAN_IN), .B1(n5864), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5860) );
  OAI21_X1 U6865 ( .B1(n6405), .B2(n5861), .A(n5860), .ZN(U2893) );
  AOI22_X1 U6866 ( .A1(n5887), .A2(DATAO_REG_29__SCAN_IN), .B1(n5864), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5862) );
  OAI21_X1 U6867 ( .B1(n6405), .B2(n4356), .A(n5862), .ZN(U2894) );
  INV_X1 U6868 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6696) );
  AOI22_X1 U6869 ( .A1(n5887), .A2(DATAO_REG_28__SCAN_IN), .B1(n5864), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5863) );
  OAI21_X1 U6870 ( .B1(n6405), .B2(n6696), .A(n5863), .ZN(U2895) );
  AOI22_X1 U6871 ( .A1(n5887), .A2(DATAO_REG_27__SCAN_IN), .B1(n5864), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5865) );
  OAI21_X1 U6872 ( .B1(n6405), .B2(n4353), .A(n5865), .ZN(U2896) );
  INV_X1 U6873 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5909) );
  INV_X2 U6874 ( .A(n6405), .ZN(n6529) );
  AOI22_X1 U6875 ( .A1(n6529), .A2(LWORD_REG_15__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5866) );
  OAI21_X1 U6876 ( .B1(n5909), .B2(n5889), .A(n5866), .ZN(U2908) );
  AOI22_X1 U6877 ( .A1(n6529), .A2(LWORD_REG_14__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5867) );
  OAI21_X1 U6878 ( .B1(n5358), .B2(n5889), .A(n5867), .ZN(U2909) );
  AOI22_X1 U6879 ( .A1(n6529), .A2(LWORD_REG_13__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5868) );
  OAI21_X1 U6880 ( .B1(n3732), .B2(n5889), .A(n5868), .ZN(U2910) );
  AOI22_X1 U6881 ( .A1(n6529), .A2(LWORD_REG_12__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5869) );
  OAI21_X1 U6882 ( .B1(n4967), .B2(n5889), .A(n5869), .ZN(U2911) );
  AOI22_X1 U6883 ( .A1(n6529), .A2(LWORD_REG_11__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n5870) );
  OAI21_X1 U6884 ( .B1(n6564), .B2(n5889), .A(n5870), .ZN(U2912) );
  INV_X1 U6885 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6663) );
  AOI22_X1 U6886 ( .A1(EAX_REG_10__SCAN_IN), .A2(n5871), .B1(n5887), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5872) );
  OAI21_X1 U6887 ( .B1(n6405), .B2(n6663), .A(n5872), .ZN(U2913) );
  INV_X1 U6888 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5874) );
  AOI22_X1 U6889 ( .A1(n6529), .A2(LWORD_REG_9__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5873) );
  OAI21_X1 U6890 ( .B1(n5874), .B2(n5889), .A(n5873), .ZN(U2914) );
  AOI22_X1 U6891 ( .A1(n6529), .A2(LWORD_REG_8__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5875) );
  OAI21_X1 U6892 ( .B1(n5876), .B2(n5889), .A(n5875), .ZN(U2915) );
  AOI22_X1 U6893 ( .A1(n6529), .A2(LWORD_REG_7__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5877) );
  OAI21_X1 U6894 ( .B1(n3646), .B2(n5889), .A(n5877), .ZN(U2916) );
  AOI22_X1 U6895 ( .A1(n6529), .A2(LWORD_REG_6__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5878) );
  OAI21_X1 U6896 ( .B1(n3639), .B2(n5889), .A(n5878), .ZN(U2917) );
  AOI22_X1 U6897 ( .A1(n6529), .A2(LWORD_REG_5__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5879) );
  OAI21_X1 U6898 ( .B1(n5880), .B2(n5889), .A(n5879), .ZN(U2918) );
  AOI22_X1 U6899 ( .A1(n6529), .A2(LWORD_REG_4__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n5881) );
  OAI21_X1 U6900 ( .B1(n5882), .B2(n5889), .A(n5881), .ZN(U2919) );
  AOI22_X1 U6901 ( .A1(n6529), .A2(LWORD_REG_3__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5883) );
  OAI21_X1 U6902 ( .B1(n6699), .B2(n5889), .A(n5883), .ZN(U2920) );
  AOI22_X1 U6903 ( .A1(n6529), .A2(LWORD_REG_2__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5884) );
  OAI21_X1 U6904 ( .B1(n4320), .B2(n5889), .A(n5884), .ZN(U2921) );
  AOI22_X1 U6905 ( .A1(n6529), .A2(LWORD_REG_1__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5885) );
  OAI21_X1 U6906 ( .B1(n5886), .B2(n5889), .A(n5885), .ZN(U2922) );
  AOI22_X1 U6907 ( .A1(n6529), .A2(LWORD_REG_0__SCAN_IN), .B1(n5887), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5888) );
  OAI21_X1 U6908 ( .B1(n4304), .B2(n5889), .A(n5888), .ZN(U2923) );
  NAND2_X1 U6909 ( .A1(n5906), .A2(DATAI_9_), .ZN(n5896) );
  INV_X1 U6910 ( .A(n5896), .ZN(n5890) );
  AOI21_X1 U6911 ( .B1(n5905), .B2(UWORD_REG_9__SCAN_IN), .A(n5890), .ZN(n5891) );
  OAI21_X1 U6912 ( .B1(n5892), .B2(n5908), .A(n5891), .ZN(U2933) );
  AOI22_X1 U6913 ( .A1(EAX_REG_26__SCAN_IN), .A2(n5902), .B1(n5905), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U6914 ( .A1(n5906), .A2(DATAI_10_), .ZN(n5898) );
  NAND2_X1 U6915 ( .A1(n5893), .A2(n5898), .ZN(U2934) );
  AOI22_X1 U6916 ( .A1(EAX_REG_28__SCAN_IN), .A2(n5902), .B1(n5905), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U6917 ( .A1(n5906), .A2(DATAI_12_), .ZN(n5900) );
  NAND2_X1 U6918 ( .A1(n5894), .A2(n5900), .ZN(U2936) );
  AOI22_X1 U6919 ( .A1(EAX_REG_30__SCAN_IN), .A2(n5902), .B1(n5905), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U6920 ( .A1(n5906), .A2(DATAI_14_), .ZN(n5903) );
  NAND2_X1 U6921 ( .A1(n5895), .A2(n5903), .ZN(U2938) );
  AOI22_X1 U6922 ( .A1(EAX_REG_9__SCAN_IN), .A2(n5902), .B1(n5905), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U6923 ( .A1(n5897), .A2(n5896), .ZN(U2948) );
  AOI22_X1 U6924 ( .A1(EAX_REG_10__SCAN_IN), .A2(n5902), .B1(n5905), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U6925 ( .A1(n5899), .A2(n5898), .ZN(U2949) );
  AOI22_X1 U6926 ( .A1(EAX_REG_12__SCAN_IN), .A2(n5902), .B1(n5905), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U6927 ( .A1(n5901), .A2(n5900), .ZN(U2951) );
  AOI22_X1 U6928 ( .A1(EAX_REG_14__SCAN_IN), .A2(n5902), .B1(n5905), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U6929 ( .A1(n5904), .A2(n5903), .ZN(U2953) );
  AOI22_X1 U6930 ( .A1(n5906), .A2(DATAI_15_), .B1(n5905), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n5907) );
  OAI21_X1 U6931 ( .B1(n5909), .B2(n5908), .A(n5907), .ZN(U2954) );
  AOI22_X1 U6932 ( .A1(n6000), .A2(REIP_REG_7__SCAN_IN), .B1(n5936), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5917) );
  OAI21_X1 U6933 ( .B1(n3019), .B2(n5913), .A(n5912), .ZN(n5914) );
  INV_X1 U6934 ( .A(n5914), .ZN(n5974) );
  AOI22_X1 U6935 ( .A1(n5974), .A2(n5940), .B1(n5941), .B2(n5915), .ZN(n5916)
         );
  OAI211_X1 U6936 ( .C1(n5946), .C2(n5918), .A(n5917), .B(n5916), .ZN(U2979)
         );
  AOI22_X1 U6937 ( .A1(n6000), .A2(REIP_REG_5__SCAN_IN), .B1(n5936), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5925) );
  OAI21_X1 U6938 ( .B1(n3011), .B2(n5921), .A(n3010), .ZN(n5922) );
  INV_X1 U6939 ( .A(n5922), .ZN(n5985) );
  AOI22_X1 U6940 ( .A1(n5985), .A2(n5940), .B1(n5941), .B2(n5923), .ZN(n5924)
         );
  OAI211_X1 U6941 ( .C1(n5946), .C2(n5926), .A(n5925), .B(n5924), .ZN(U2981)
         );
  AOI22_X1 U6942 ( .A1(n6000), .A2(REIP_REG_3__SCAN_IN), .B1(n5936), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5934) );
  INV_X1 U6943 ( .A(n5927), .ZN(n5932) );
  OR2_X1 U6944 ( .A1(n5929), .A2(n5928), .ZN(n5930) );
  AND2_X1 U6945 ( .A1(n5931), .A2(n5930), .ZN(n6004) );
  AOI22_X1 U6946 ( .A1(n5941), .A2(n5932), .B1(n6004), .B2(n5940), .ZN(n5933)
         );
  OAI211_X1 U6947 ( .C1(n5946), .C2(n5935), .A(n5934), .B(n5933), .ZN(U2983)
         );
  AOI22_X1 U6948 ( .A1(n6000), .A2(REIP_REG_2__SCAN_IN), .B1(n5936), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5944) );
  INV_X1 U6949 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6669) );
  XNOR2_X1 U6950 ( .A(n5938), .B(n6669), .ZN(n5939) );
  XNOR2_X1 U6951 ( .A(n5937), .B(n5939), .ZN(n6020) );
  AOI22_X1 U6952 ( .A1(n5942), .A2(n5941), .B1(n5940), .B2(n6020), .ZN(n5943)
         );
  OAI211_X1 U6953 ( .C1(n5946), .C2(n5945), .A(n5944), .B(n5943), .ZN(U2984)
         );
  AOI21_X1 U6954 ( .B1(n6010), .B2(n5948), .A(n5947), .ZN(n5952) );
  AOI22_X1 U6955 ( .A1(n6021), .A2(n5950), .B1(n5953), .B2(n5949), .ZN(n5951)
         );
  OAI211_X1 U6956 ( .C1(n5954), .C2(n5953), .A(n5952), .B(n5951), .ZN(U3007)
         );
  INV_X1 U6957 ( .A(n5955), .ZN(n5964) );
  INV_X1 U6958 ( .A(n5956), .ZN(n5958) );
  AOI21_X1 U6959 ( .B1(n6010), .B2(n5958), .A(n5957), .ZN(n5962) );
  AOI22_X1 U6960 ( .A1(n5960), .A2(n6021), .B1(n5959), .B2(n5963), .ZN(n5961)
         );
  OAI211_X1 U6961 ( .C1(n5964), .C2(n5963), .A(n5962), .B(n5961), .ZN(U3009)
         );
  INV_X1 U6962 ( .A(n5965), .ZN(n5971) );
  INV_X1 U6963 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6458) );
  OAI22_X1 U6964 ( .A1(n5967), .A2(n5966), .B1(n6458), .B2(n5819), .ZN(n5970)
         );
  AOI211_X1 U6965 ( .C1(n5978), .C2(n5973), .A(n5968), .B(n5979), .ZN(n5969)
         );
  AOI211_X1 U6966 ( .C1(n5971), .C2(n6021), .A(n5970), .B(n5969), .ZN(n5972)
         );
  OAI21_X1 U6967 ( .B1(n5977), .B2(n5973), .A(n5972), .ZN(U3010) );
  AOI222_X1 U6968 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6000), .B1(n6010), .B2(
        n5975), .C1(n6021), .C2(n5974), .ZN(n5976) );
  OAI221_X1 U6969 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5979), .C1(n5978), .C2(n5977), .A(n5976), .ZN(U3011) );
  AOI21_X1 U6970 ( .B1(n6016), .B2(n5980), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n5988) );
  INV_X1 U6971 ( .A(n5981), .ZN(n5982) );
  AOI22_X1 U6972 ( .A1(n6010), .A2(n5982), .B1(n6000), .B2(REIP_REG_5__SCAN_IN), .ZN(n5987) );
  NOR4_X1 U6973 ( .A1(n6013), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n5983), 
        .A4(n5995), .ZN(n5984) );
  AOI21_X1 U6974 ( .B1(n5985), .B2(n6021), .A(n5984), .ZN(n5986) );
  OAI211_X1 U6975 ( .C1(n5989), .C2(n5988), .A(n5987), .B(n5986), .ZN(U3013)
         );
  AOI21_X1 U6976 ( .B1(n6016), .B2(n6011), .A(n6014), .ZN(n6008) );
  INV_X1 U6977 ( .A(n5990), .ZN(n5991) );
  AOI21_X1 U6978 ( .B1(n6010), .B2(n5992), .A(n5991), .ZN(n5998) );
  INV_X1 U6979 ( .A(n5993), .ZN(n5996) );
  AOI211_X1 U6980 ( .C1(n6007), .C2(n5999), .A(n6002), .B(n6011), .ZN(n5994)
         );
  AOI22_X1 U6981 ( .A1(n5996), .A2(n6021), .B1(n5995), .B2(n5994), .ZN(n5997)
         );
  OAI211_X1 U6982 ( .C1(n6008), .C2(n5999), .A(n5998), .B(n5997), .ZN(U3014)
         );
  AOI22_X1 U6983 ( .A1(n6010), .A2(n6001), .B1(n6000), .B2(REIP_REG_3__SCAN_IN), .ZN(n6006) );
  NOR2_X1 U6984 ( .A1(n6011), .A2(n6002), .ZN(n6003) );
  AOI22_X1 U6985 ( .A1(n6004), .A2(n6021), .B1(n6003), .B2(n6007), .ZN(n6005)
         );
  OAI211_X1 U6986 ( .C1(n6008), .C2(n6007), .A(n6006), .B(n6005), .ZN(U3015)
         );
  AOI22_X1 U6987 ( .A1(n6016), .A2(n6011), .B1(n6010), .B2(n6009), .ZN(n6023)
         );
  NOR3_X1 U6988 ( .A1(n6013), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n6012), 
        .ZN(n6019) );
  AOI21_X1 U6989 ( .B1(n6016), .B2(n6015), .A(n6014), .ZN(n6017) );
  NOR2_X1 U6990 ( .A1(n6017), .A2(n6669), .ZN(n6018) );
  AOI211_X1 U6991 ( .C1(n6021), .C2(n6020), .A(n6019), .B(n6018), .ZN(n6022)
         );
  OAI211_X1 U6992 ( .C1(n5819), .C2(n6448), .A(n6023), .B(n6022), .ZN(U3016)
         );
  NOR2_X1 U6993 ( .A1(n6025), .A2(n6024), .ZN(U3019) );
  NOR2_X1 U6994 ( .A1(n6185), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6052)
         );
  AOI22_X1 U6995 ( .A1(n6307), .A2(n6052), .B1(n6270), .B2(n6051), .ZN(n6038)
         );
  INV_X1 U6996 ( .A(n6027), .ZN(n6182) );
  NAND3_X1 U6997 ( .A1(n6181), .A2(n6028), .A3(n6182), .ZN(n6029) );
  NAND2_X1 U6998 ( .A1(n6029), .A2(n6317), .ZN(n6036) );
  INV_X1 U6999 ( .A(n6030), .ZN(n6031) );
  AOI21_X1 U7000 ( .B1(n6031), .B2(n3029), .A(n6052), .ZN(n6035) );
  INV_X1 U7001 ( .A(n6035), .ZN(n6033) );
  AOI21_X1 U7002 ( .B1(n6305), .B2(n6034), .A(n6222), .ZN(n6032) );
  OAI22_X1 U7003 ( .A1(n6036), .A2(n6035), .B1(n6034), .B2(n6303), .ZN(n6053)
         );
  AOI22_X1 U7004 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6054), .B1(n6308), 
        .B2(n6053), .ZN(n6037) );
  OAI211_X1 U7005 ( .C1(n6273), .C2(n6089), .A(n6038), .B(n6037), .ZN(U3044)
         );
  AOI22_X1 U7006 ( .A1(n6322), .A2(n6052), .B1(n6324), .B2(n6051), .ZN(n6040)
         );
  AOI22_X1 U7007 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6054), .B1(n6323), 
        .B2(n6053), .ZN(n6039) );
  OAI211_X1 U7008 ( .C1(n6327), .C2(n6089), .A(n6040), .B(n6039), .ZN(U3045)
         );
  AOI22_X1 U7009 ( .A1(n6328), .A2(n6052), .B1(n6276), .B2(n6051), .ZN(n6042)
         );
  AOI22_X1 U7010 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6054), .B1(n6329), 
        .B2(n6053), .ZN(n6041) );
  OAI211_X1 U7011 ( .C1(n6279), .C2(n6089), .A(n6042), .B(n6041), .ZN(U3046)
         );
  AOI22_X1 U7012 ( .A1(n6334), .A2(n6052), .B1(n6280), .B2(n6051), .ZN(n6044)
         );
  AOI22_X1 U7013 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6054), .B1(n6335), 
        .B2(n6053), .ZN(n6043) );
  OAI211_X1 U7014 ( .C1(n6283), .C2(n6089), .A(n6044), .B(n6043), .ZN(U3047)
         );
  AOI22_X1 U7015 ( .A1(n6340), .A2(n6052), .B1(n6284), .B2(n6051), .ZN(n6046)
         );
  AOI22_X1 U7016 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6054), .B1(n6341), 
        .B2(n6053), .ZN(n6045) );
  OAI211_X1 U7017 ( .C1(n6287), .C2(n6089), .A(n6046), .B(n6045), .ZN(U3048)
         );
  AOI22_X1 U7018 ( .A1(n6346), .A2(n6052), .B1(n6348), .B2(n6051), .ZN(n6048)
         );
  AOI22_X1 U7019 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6054), .B1(n6347), 
        .B2(n6053), .ZN(n6047) );
  OAI211_X1 U7020 ( .C1(n6351), .C2(n6089), .A(n6048), .B(n6047), .ZN(U3049)
         );
  AOI22_X1 U7021 ( .A1(n6352), .A2(n6052), .B1(n6355), .B2(n6051), .ZN(n6050)
         );
  AOI22_X1 U7022 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6054), .B1(n6353), 
        .B2(n6053), .ZN(n6049) );
  OAI211_X1 U7023 ( .C1(n6359), .C2(n6089), .A(n6050), .B(n6049), .ZN(U3050)
         );
  AOI22_X1 U7024 ( .A1(n6360), .A2(n6052), .B1(n6295), .B2(n6051), .ZN(n6056)
         );
  AOI22_X1 U7025 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6054), .B1(n6363), 
        .B2(n6053), .ZN(n6055) );
  OAI211_X1 U7026 ( .C1(n6299), .C2(n6089), .A(n6056), .B(n6055), .ZN(U3051)
         );
  OAI22_X1 U7027 ( .A1(n6058), .A2(n3031), .B1(n6057), .B2(n6262), .ZN(n6085)
         );
  NAND2_X1 U7028 ( .A1(n6221), .A2(n6265), .ZN(n6092) );
  NOR2_X1 U7029 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6092), .ZN(n6084)
         );
  AOI22_X1 U7030 ( .A1(n6308), .A2(n6085), .B1(n6307), .B2(n6084), .ZN(n6068)
         );
  INV_X1 U7031 ( .A(n6089), .ZN(n6061) );
  NOR2_X1 U7032 ( .A1(n6218), .A2(n6059), .ZN(n6091) );
  OAI21_X1 U7033 ( .B1(n6119), .B2(n6060), .A(n6317), .ZN(n6090) );
  AOI211_X1 U7034 ( .C1(n6061), .C2(n6310), .A(n6091), .B(n6090), .ZN(n6064)
         );
  OAI21_X1 U7035 ( .B1(n6084), .B2(n6501), .A(n6062), .ZN(n6063) );
  NOR2_X2 U7036 ( .A1(n6119), .A2(n6066), .ZN(n6113) );
  AOI22_X1 U7037 ( .A1(n6086), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6318), 
        .B2(n6113), .ZN(n6067) );
  OAI211_X1 U7038 ( .C1(n6321), .C2(n6089), .A(n6068), .B(n6067), .ZN(U3052)
         );
  AOI22_X1 U7039 ( .A1(n6323), .A2(n6085), .B1(n6322), .B2(n6084), .ZN(n6070)
         );
  AOI22_X1 U7040 ( .A1(n6086), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6232), 
        .B2(n6113), .ZN(n6069) );
  OAI211_X1 U7041 ( .C1(n6071), .C2(n6089), .A(n6070), .B(n6069), .ZN(U3053)
         );
  AOI22_X1 U7042 ( .A1(n6329), .A2(n6085), .B1(n6328), .B2(n6084), .ZN(n6073)
         );
  AOI22_X1 U7043 ( .A1(n6086), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6330), 
        .B2(n6113), .ZN(n6072) );
  OAI211_X1 U7044 ( .C1(n6333), .C2(n6089), .A(n6073), .B(n6072), .ZN(U3054)
         );
  AOI22_X1 U7045 ( .A1(n6335), .A2(n6085), .B1(n6334), .B2(n6084), .ZN(n6075)
         );
  AOI22_X1 U7046 ( .A1(n6086), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6336), 
        .B2(n6113), .ZN(n6074) );
  OAI211_X1 U7047 ( .C1(n6339), .C2(n6089), .A(n6075), .B(n6074), .ZN(U3055)
         );
  AOI22_X1 U7048 ( .A1(n6341), .A2(n6085), .B1(n6340), .B2(n6084), .ZN(n6077)
         );
  AOI22_X1 U7049 ( .A1(n6086), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6342), 
        .B2(n6113), .ZN(n6076) );
  OAI211_X1 U7050 ( .C1(n6345), .C2(n6089), .A(n6077), .B(n6076), .ZN(U3056)
         );
  AOI22_X1 U7051 ( .A1(n6347), .A2(n6085), .B1(n6346), .B2(n6084), .ZN(n6079)
         );
  AOI22_X1 U7052 ( .A1(n6086), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6245), 
        .B2(n6113), .ZN(n6078) );
  OAI211_X1 U7053 ( .C1(n6080), .C2(n6089), .A(n6079), .B(n6078), .ZN(U3057)
         );
  AOI22_X1 U7054 ( .A1(n6353), .A2(n6085), .B1(n6352), .B2(n6084), .ZN(n6082)
         );
  AOI22_X1 U7055 ( .A1(n6086), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6249), 
        .B2(n6113), .ZN(n6081) );
  OAI211_X1 U7056 ( .C1(n6083), .C2(n6089), .A(n6082), .B(n6081), .ZN(U3058)
         );
  AOI22_X1 U7057 ( .A1(n6363), .A2(n6085), .B1(n6360), .B2(n6084), .ZN(n6088)
         );
  AOI22_X1 U7058 ( .A1(n6086), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6365), 
        .B2(n6113), .ZN(n6087) );
  OAI211_X1 U7059 ( .C1(n6370), .C2(n6089), .A(n6088), .B(n6087), .ZN(U3059)
         );
  INV_X1 U7060 ( .A(n6090), .ZN(n6095) );
  NOR2_X1 U7061 ( .A1(n6216), .A2(n6092), .ZN(n6112) );
  AOI21_X1 U7062 ( .B1(n6091), .B2(n3029), .A(n6112), .ZN(n6094) );
  INV_X1 U7063 ( .A(n6094), .ZN(n6093) );
  INV_X1 U7064 ( .A(n6092), .ZN(n6097) );
  NOR2_X2 U7065 ( .A1(n6119), .A2(n6227), .ZN(n6143) );
  AOI22_X1 U7066 ( .A1(n6307), .A2(n6112), .B1(n6318), .B2(n6143), .ZN(n6099)
         );
  NAND2_X1 U7067 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  OAI211_X1 U7068 ( .C1(n6317), .C2(n6097), .A(n6096), .B(n6314), .ZN(n6114)
         );
  AOI22_X1 U7069 ( .A1(n6114), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n6270), 
        .B2(n6113), .ZN(n6098) );
  OAI211_X1 U7070 ( .C1(n6117), .C2(n6231), .A(n6099), .B(n6098), .ZN(U3060)
         );
  AOI22_X1 U7071 ( .A1(n6322), .A2(n6112), .B1(n6232), .B2(n6143), .ZN(n6101)
         );
  AOI22_X1 U7072 ( .A1(n6114), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n6324), 
        .B2(n6113), .ZN(n6100) );
  OAI211_X1 U7073 ( .C1(n6117), .C2(n6235), .A(n6101), .B(n6100), .ZN(U3061)
         );
  AOI22_X1 U7074 ( .A1(n6328), .A2(n6112), .B1(n6330), .B2(n6143), .ZN(n6103)
         );
  AOI22_X1 U7075 ( .A1(n6114), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n6276), 
        .B2(n6113), .ZN(n6102) );
  OAI211_X1 U7076 ( .C1(n6117), .C2(n6238), .A(n6103), .B(n6102), .ZN(U3062)
         );
  AOI22_X1 U7077 ( .A1(n6334), .A2(n6112), .B1(n6336), .B2(n6143), .ZN(n6105)
         );
  AOI22_X1 U7078 ( .A1(n6114), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n6280), 
        .B2(n6113), .ZN(n6104) );
  OAI211_X1 U7079 ( .C1(n6117), .C2(n6241), .A(n6105), .B(n6104), .ZN(U3063)
         );
  AOI22_X1 U7080 ( .A1(n6340), .A2(n6112), .B1(n6342), .B2(n6143), .ZN(n6107)
         );
  AOI22_X1 U7081 ( .A1(n6114), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n6284), 
        .B2(n6113), .ZN(n6106) );
  OAI211_X1 U7082 ( .C1(n6117), .C2(n6244), .A(n6107), .B(n6106), .ZN(U3064)
         );
  AOI22_X1 U7083 ( .A1(n6346), .A2(n6112), .B1(n6245), .B2(n6143), .ZN(n6109)
         );
  AOI22_X1 U7084 ( .A1(n6114), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n6348), 
        .B2(n6113), .ZN(n6108) );
  OAI211_X1 U7085 ( .C1(n6117), .C2(n6248), .A(n6109), .B(n6108), .ZN(U3065)
         );
  AOI22_X1 U7086 ( .A1(n6352), .A2(n6112), .B1(n6249), .B2(n6143), .ZN(n6111)
         );
  AOI22_X1 U7087 ( .A1(n6114), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n6355), 
        .B2(n6113), .ZN(n6110) );
  OAI211_X1 U7088 ( .C1(n6117), .C2(n6252), .A(n6111), .B(n6110), .ZN(U3066)
         );
  AOI22_X1 U7089 ( .A1(n6360), .A2(n6112), .B1(n6365), .B2(n6143), .ZN(n6116)
         );
  AOI22_X1 U7090 ( .A1(n6114), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n6295), 
        .B2(n6113), .ZN(n6115) );
  OAI211_X1 U7091 ( .C1(n6117), .C2(n6258), .A(n6116), .B(n6115), .ZN(U3067)
         );
  INV_X1 U7092 ( .A(n6301), .ZN(n6121) );
  NAND2_X1 U7093 ( .A1(n6261), .A2(n6121), .ZN(n6150) );
  OAI22_X1 U7094 ( .A1(n6150), .A2(n6305), .B1(n6122), .B2(n6262), .ZN(n6142)
         );
  NOR2_X1 U7095 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6156), .ZN(n6141)
         );
  AOI22_X1 U7096 ( .A1(n6308), .A2(n6142), .B1(n6307), .B2(n6141), .ZN(n6128)
         );
  OAI21_X1 U7097 ( .B1(n6174), .B2(n6143), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6123) );
  NAND3_X1 U7098 ( .A1(n6123), .A2(n6317), .A3(n6150), .ZN(n6126) );
  INV_X1 U7099 ( .A(n6141), .ZN(n6124) );
  AOI211_X1 U7100 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6124), .A(n6264), .B(
        n6266), .ZN(n6125) );
  NAND3_X1 U7101 ( .A1(n6265), .A2(n6126), .A3(n6125), .ZN(n6144) );
  AOI22_X1 U7102 ( .A1(n6144), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6270), 
        .B2(n6143), .ZN(n6127) );
  OAI211_X1 U7103 ( .C1(n6273), .C2(n6147), .A(n6128), .B(n6127), .ZN(U3068)
         );
  AOI22_X1 U7104 ( .A1(n6323), .A2(n6142), .B1(n6322), .B2(n6141), .ZN(n6130)
         );
  AOI22_X1 U7105 ( .A1(n6144), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6324), 
        .B2(n6143), .ZN(n6129) );
  OAI211_X1 U7106 ( .C1(n6327), .C2(n6147), .A(n6130), .B(n6129), .ZN(U3069)
         );
  AOI22_X1 U7107 ( .A1(n6329), .A2(n6142), .B1(n6328), .B2(n6141), .ZN(n6132)
         );
  AOI22_X1 U7108 ( .A1(n6144), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6276), 
        .B2(n6143), .ZN(n6131) );
  OAI211_X1 U7109 ( .C1(n6279), .C2(n6147), .A(n6132), .B(n6131), .ZN(U3070)
         );
  AOI22_X1 U7110 ( .A1(n6335), .A2(n6142), .B1(n6334), .B2(n6141), .ZN(n6134)
         );
  AOI22_X1 U7111 ( .A1(n6144), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6280), 
        .B2(n6143), .ZN(n6133) );
  OAI211_X1 U7112 ( .C1(n6283), .C2(n6147), .A(n6134), .B(n6133), .ZN(U3071)
         );
  AOI22_X1 U7113 ( .A1(n6341), .A2(n6142), .B1(n6340), .B2(n6141), .ZN(n6136)
         );
  AOI22_X1 U7114 ( .A1(n6144), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6284), 
        .B2(n6143), .ZN(n6135) );
  OAI211_X1 U7115 ( .C1(n6287), .C2(n6147), .A(n6136), .B(n6135), .ZN(U3072)
         );
  AOI22_X1 U7116 ( .A1(n6347), .A2(n6142), .B1(n6346), .B2(n6141), .ZN(n6138)
         );
  AOI22_X1 U7117 ( .A1(n6144), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6348), 
        .B2(n6143), .ZN(n6137) );
  OAI211_X1 U7118 ( .C1(n6351), .C2(n6147), .A(n6138), .B(n6137), .ZN(U3073)
         );
  AOI22_X1 U7119 ( .A1(n6353), .A2(n6142), .B1(n6352), .B2(n6141), .ZN(n6140)
         );
  AOI22_X1 U7120 ( .A1(n6144), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6355), 
        .B2(n6143), .ZN(n6139) );
  OAI211_X1 U7121 ( .C1(n6359), .C2(n6147), .A(n6140), .B(n6139), .ZN(U3074)
         );
  AOI22_X1 U7122 ( .A1(n6363), .A2(n6142), .B1(n6360), .B2(n6141), .ZN(n6146)
         );
  AOI22_X1 U7123 ( .A1(n6144), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6295), 
        .B2(n6143), .ZN(n6145) );
  OAI211_X1 U7124 ( .C1(n6299), .C2(n6147), .A(n6146), .B(n6145), .ZN(U3075)
         );
  NAND2_X1 U7125 ( .A1(n6317), .A2(n6148), .ZN(n6158) );
  OR2_X1 U7126 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  OAI22_X1 U7127 ( .A1(n6303), .A2(n6156), .B1(n6158), .B2(n6155), .ZN(n6152)
         );
  INV_X1 U7128 ( .A(n6153), .ZN(n6175) );
  AOI22_X1 U7129 ( .A1(n6307), .A2(n6175), .B1(n6318), .B2(n6176), .ZN(n6161)
         );
  INV_X1 U7130 ( .A(n6155), .ZN(n6159) );
  AOI21_X1 U7131 ( .B1(n6156), .B2(n6305), .A(n6222), .ZN(n6157) );
  AOI22_X1 U7132 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6177), .B1(n6270), 
        .B2(n6174), .ZN(n6160) );
  OAI211_X1 U7133 ( .C1(n6180), .C2(n6231), .A(n6161), .B(n6160), .ZN(U3076)
         );
  AOI22_X1 U7134 ( .A1(n6322), .A2(n6175), .B1(n6232), .B2(n6176), .ZN(n6163)
         );
  AOI22_X1 U7135 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6177), .B1(n6324), 
        .B2(n6174), .ZN(n6162) );
  OAI211_X1 U7136 ( .C1(n6180), .C2(n6235), .A(n6163), .B(n6162), .ZN(U3077)
         );
  AOI22_X1 U7137 ( .A1(n6328), .A2(n6175), .B1(n6330), .B2(n6176), .ZN(n6165)
         );
  AOI22_X1 U7138 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6177), .B1(n6276), 
        .B2(n6174), .ZN(n6164) );
  OAI211_X1 U7139 ( .C1(n6180), .C2(n6238), .A(n6165), .B(n6164), .ZN(U3078)
         );
  AOI22_X1 U7140 ( .A1(n6334), .A2(n6175), .B1(n6280), .B2(n6174), .ZN(n6167)
         );
  AOI22_X1 U7141 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6177), .B1(n6336), 
        .B2(n6176), .ZN(n6166) );
  OAI211_X1 U7142 ( .C1(n6180), .C2(n6241), .A(n6167), .B(n6166), .ZN(U3079)
         );
  AOI22_X1 U7143 ( .A1(n6340), .A2(n6175), .B1(n6342), .B2(n6176), .ZN(n6169)
         );
  AOI22_X1 U7144 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6177), .B1(n6284), 
        .B2(n6174), .ZN(n6168) );
  OAI211_X1 U7145 ( .C1(n6180), .C2(n6244), .A(n6169), .B(n6168), .ZN(U3080)
         );
  AOI22_X1 U7146 ( .A1(n6346), .A2(n6175), .B1(n6348), .B2(n6174), .ZN(n6171)
         );
  AOI22_X1 U7147 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6177), .B1(n6245), 
        .B2(n6176), .ZN(n6170) );
  OAI211_X1 U7148 ( .C1(n6180), .C2(n6248), .A(n6171), .B(n6170), .ZN(U3081)
         );
  AOI22_X1 U7149 ( .A1(n6352), .A2(n6175), .B1(n6249), .B2(n6176), .ZN(n6173)
         );
  AOI22_X1 U7150 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6177), .B1(n6355), 
        .B2(n6174), .ZN(n6172) );
  OAI211_X1 U7151 ( .C1(n6180), .C2(n6252), .A(n6173), .B(n6172), .ZN(U3082)
         );
  AOI22_X1 U7152 ( .A1(n6360), .A2(n6175), .B1(n6295), .B2(n6174), .ZN(n6179)
         );
  AOI22_X1 U7153 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6177), .B1(n6365), 
        .B2(n6176), .ZN(n6178) );
  OAI211_X1 U7154 ( .C1(n6180), .C2(n6258), .A(n6179), .B(n6178), .ZN(U3083)
         );
  INV_X1 U7155 ( .A(n6181), .ZN(n6183) );
  AOI21_X1 U7156 ( .B1(n6183), .B2(n6182), .A(n6305), .ZN(n6188) );
  NAND2_X1 U7157 ( .A1(n6184), .A2(n3029), .ZN(n6187) );
  NOR2_X1 U7158 ( .A1(n6185), .A2(n6265), .ZN(n6209) );
  INV_X1 U7159 ( .A(n6209), .ZN(n6186) );
  NAND2_X1 U7160 ( .A1(n6187), .A2(n6186), .ZN(n6192) );
  AOI22_X1 U7161 ( .A1(n6307), .A2(n6209), .B1(n6318), .B2(n6210), .ZN(n6195)
         );
  INV_X1 U7162 ( .A(n6188), .ZN(n6193) );
  INV_X1 U7163 ( .A(n6189), .ZN(n6190) );
  AOI21_X1 U7164 ( .B1(n6305), .B2(n6190), .A(n6222), .ZN(n6191) );
  AOI22_X1 U7165 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6211), .B1(n6270), 
        .B2(n6208), .ZN(n6194) );
  OAI211_X1 U7166 ( .C1(n6214), .C2(n6231), .A(n6195), .B(n6194), .ZN(U3108)
         );
  AOI22_X1 U7167 ( .A1(n6322), .A2(n6209), .B1(n6324), .B2(n6208), .ZN(n6197)
         );
  AOI22_X1 U7168 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6211), .B1(n6232), 
        .B2(n6210), .ZN(n6196) );
  OAI211_X1 U7169 ( .C1(n6214), .C2(n6235), .A(n6197), .B(n6196), .ZN(U3109)
         );
  AOI22_X1 U7170 ( .A1(n6328), .A2(n6209), .B1(n6330), .B2(n6210), .ZN(n6199)
         );
  AOI22_X1 U7171 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6211), .B1(n6276), 
        .B2(n6208), .ZN(n6198) );
  OAI211_X1 U7172 ( .C1(n6214), .C2(n6238), .A(n6199), .B(n6198), .ZN(U3110)
         );
  AOI22_X1 U7173 ( .A1(n6334), .A2(n6209), .B1(n6280), .B2(n6208), .ZN(n6201)
         );
  AOI22_X1 U7174 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6211), .B1(n6336), 
        .B2(n6210), .ZN(n6200) );
  OAI211_X1 U7175 ( .C1(n6214), .C2(n6241), .A(n6201), .B(n6200), .ZN(U3111)
         );
  AOI22_X1 U7176 ( .A1(n6340), .A2(n6209), .B1(n6284), .B2(n6208), .ZN(n6203)
         );
  AOI22_X1 U7177 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6211), .B1(n6342), 
        .B2(n6210), .ZN(n6202) );
  OAI211_X1 U7178 ( .C1(n6214), .C2(n6244), .A(n6203), .B(n6202), .ZN(U3112)
         );
  AOI22_X1 U7179 ( .A1(n6346), .A2(n6209), .B1(n6245), .B2(n6210), .ZN(n6205)
         );
  AOI22_X1 U7180 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6211), .B1(n6348), 
        .B2(n6208), .ZN(n6204) );
  OAI211_X1 U7181 ( .C1(n6214), .C2(n6248), .A(n6205), .B(n6204), .ZN(U3113)
         );
  AOI22_X1 U7182 ( .A1(n6352), .A2(n6209), .B1(n6355), .B2(n6208), .ZN(n6207)
         );
  AOI22_X1 U7183 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6211), .B1(n6249), 
        .B2(n6210), .ZN(n6206) );
  OAI211_X1 U7184 ( .C1(n6214), .C2(n6252), .A(n6207), .B(n6206), .ZN(U3114)
         );
  AOI22_X1 U7185 ( .A1(n6360), .A2(n6209), .B1(n6295), .B2(n6208), .ZN(n6213)
         );
  AOI22_X1 U7186 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6211), .B1(n6365), 
        .B2(n6210), .ZN(n6212) );
  OAI211_X1 U7187 ( .C1(n6214), .C2(n6258), .A(n6213), .B(n6212), .ZN(U3115)
         );
  NOR2_X1 U7188 ( .A1(n6303), .A2(n6265), .ZN(n6220) );
  NAND2_X1 U7189 ( .A1(n6317), .A2(n6215), .ZN(n6226) );
  INV_X1 U7190 ( .A(n6226), .ZN(n6219) );
  NOR2_X1 U7191 ( .A1(n6216), .A2(n6223), .ZN(n6254) );
  INV_X1 U7192 ( .A(n6254), .ZN(n6217) );
  OAI21_X1 U7193 ( .B1(n6300), .B2(n6218), .A(n6217), .ZN(n6225) );
  AOI22_X1 U7194 ( .A1(n6307), .A2(n6254), .B1(n6270), .B2(n6253), .ZN(n6230)
         );
  AOI21_X1 U7195 ( .B1(n6305), .B2(n6223), .A(n6222), .ZN(n6224) );
  OAI21_X1 U7196 ( .B1(n6226), .B2(n6225), .A(n6224), .ZN(n6255) );
  NOR2_X2 U7197 ( .A1(n6228), .A2(n6227), .ZN(n6294) );
  AOI22_X1 U7198 ( .A1(n6255), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n6318), 
        .B2(n6294), .ZN(n6229) );
  OAI211_X1 U7199 ( .C1(n6259), .C2(n6231), .A(n6230), .B(n6229), .ZN(U3124)
         );
  AOI22_X1 U7200 ( .A1(n6322), .A2(n6254), .B1(n6324), .B2(n6253), .ZN(n6234)
         );
  AOI22_X1 U7201 ( .A1(n6255), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n6232), 
        .B2(n6294), .ZN(n6233) );
  OAI211_X1 U7202 ( .C1(n6259), .C2(n6235), .A(n6234), .B(n6233), .ZN(U3125)
         );
  AOI22_X1 U7203 ( .A1(n6328), .A2(n6254), .B1(n6330), .B2(n6294), .ZN(n6237)
         );
  AOI22_X1 U7204 ( .A1(n6255), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n6276), 
        .B2(n6253), .ZN(n6236) );
  OAI211_X1 U7205 ( .C1(n6259), .C2(n6238), .A(n6237), .B(n6236), .ZN(U3126)
         );
  AOI22_X1 U7206 ( .A1(n6334), .A2(n6254), .B1(n6280), .B2(n6253), .ZN(n6240)
         );
  AOI22_X1 U7207 ( .A1(n6255), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n6336), 
        .B2(n6294), .ZN(n6239) );
  OAI211_X1 U7208 ( .C1(n6259), .C2(n6241), .A(n6240), .B(n6239), .ZN(U3127)
         );
  AOI22_X1 U7209 ( .A1(n6340), .A2(n6254), .B1(n6284), .B2(n6253), .ZN(n6243)
         );
  AOI22_X1 U7210 ( .A1(n6255), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n6342), 
        .B2(n6294), .ZN(n6242) );
  OAI211_X1 U7211 ( .C1(n6259), .C2(n6244), .A(n6243), .B(n6242), .ZN(U3128)
         );
  AOI22_X1 U7212 ( .A1(n6346), .A2(n6254), .B1(n6348), .B2(n6253), .ZN(n6247)
         );
  AOI22_X1 U7213 ( .A1(n6255), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n6245), 
        .B2(n6294), .ZN(n6246) );
  OAI211_X1 U7214 ( .C1(n6259), .C2(n6248), .A(n6247), .B(n6246), .ZN(U3129)
         );
  AOI22_X1 U7215 ( .A1(n6352), .A2(n6254), .B1(n6355), .B2(n6253), .ZN(n6251)
         );
  AOI22_X1 U7216 ( .A1(n6255), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n6249), 
        .B2(n6294), .ZN(n6250) );
  OAI211_X1 U7217 ( .C1(n6259), .C2(n6252), .A(n6251), .B(n6250), .ZN(U3130)
         );
  AOI22_X1 U7218 ( .A1(n6360), .A2(n6254), .B1(n6295), .B2(n6253), .ZN(n6257)
         );
  AOI22_X1 U7219 ( .A1(n6255), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n6365), 
        .B2(n6294), .ZN(n6256) );
  OAI211_X1 U7220 ( .C1(n6259), .C2(n6258), .A(n6257), .B(n6256), .ZN(U3131)
         );
  OAI33_X1 U7221 ( .A1(n6263), .A2(n6265), .A3(n6262), .B1(n6301), .B2(n6305), 
        .B3(n6261), .ZN(n6293) );
  NOR2_X1 U7222 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6304), .ZN(n6292)
         );
  AOI22_X1 U7223 ( .A1(n6308), .A2(n6293), .B1(n6307), .B2(n6292), .ZN(n6272)
         );
  NOR3_X1 U7224 ( .A1(n6266), .A2(n6265), .A3(n6264), .ZN(n6269) );
  INV_X1 U7225 ( .A(n6369), .ZN(n6354) );
  OAI21_X1 U7226 ( .B1(n6354), .B2(n6294), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6267) );
  NAND3_X1 U7227 ( .A1(n6301), .A2(n6317), .A3(n6267), .ZN(n6268) );
  OAI211_X1 U7228 ( .C1(n6292), .C2(n6501), .A(n6269), .B(n6268), .ZN(n6296)
         );
  AOI22_X1 U7229 ( .A1(n6296), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n6270), 
        .B2(n6294), .ZN(n6271) );
  OAI211_X1 U7230 ( .C1(n6273), .C2(n6369), .A(n6272), .B(n6271), .ZN(U3132)
         );
  AOI22_X1 U7231 ( .A1(n6323), .A2(n6293), .B1(n6322), .B2(n6292), .ZN(n6275)
         );
  AOI22_X1 U7232 ( .A1(n6296), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n6324), 
        .B2(n6294), .ZN(n6274) );
  OAI211_X1 U7233 ( .C1(n6327), .C2(n6369), .A(n6275), .B(n6274), .ZN(U3133)
         );
  AOI22_X1 U7234 ( .A1(n6329), .A2(n6293), .B1(n6328), .B2(n6292), .ZN(n6278)
         );
  AOI22_X1 U7235 ( .A1(n6296), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n6276), 
        .B2(n6294), .ZN(n6277) );
  OAI211_X1 U7236 ( .C1(n6279), .C2(n6369), .A(n6278), .B(n6277), .ZN(U3134)
         );
  AOI22_X1 U7237 ( .A1(n6335), .A2(n6293), .B1(n6334), .B2(n6292), .ZN(n6282)
         );
  AOI22_X1 U7238 ( .A1(n6296), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n6280), 
        .B2(n6294), .ZN(n6281) );
  OAI211_X1 U7239 ( .C1(n6283), .C2(n6369), .A(n6282), .B(n6281), .ZN(U3135)
         );
  AOI22_X1 U7240 ( .A1(n6341), .A2(n3043), .B1(n6340), .B2(n6292), .ZN(n6286)
         );
  AOI22_X1 U7241 ( .A1(n6296), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n6284), 
        .B2(n6294), .ZN(n6285) );
  OAI211_X1 U7242 ( .C1(n6287), .C2(n6369), .A(n6286), .B(n6285), .ZN(U3136)
         );
  AOI22_X1 U7243 ( .A1(n6347), .A2(n3043), .B1(n6346), .B2(n6292), .ZN(n6289)
         );
  AOI22_X1 U7244 ( .A1(n6296), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n6348), 
        .B2(n6294), .ZN(n6288) );
  OAI211_X1 U7245 ( .C1(n6351), .C2(n6369), .A(n6289), .B(n6288), .ZN(U3137)
         );
  AOI22_X1 U7246 ( .A1(n6353), .A2(n3043), .B1(n6352), .B2(n6292), .ZN(n6291)
         );
  AOI22_X1 U7247 ( .A1(n6296), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n6355), 
        .B2(n6294), .ZN(n6290) );
  OAI211_X1 U7248 ( .C1(n6359), .C2(n6369), .A(n6291), .B(n6290), .ZN(U3138)
         );
  AOI22_X1 U7249 ( .A1(n6363), .A2(n3043), .B1(n6360), .B2(n6292), .ZN(n6298)
         );
  AOI22_X1 U7250 ( .A1(n6296), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n6295), 
        .B2(n6294), .ZN(n6297) );
  OAI211_X1 U7251 ( .C1(n6299), .C2(n6369), .A(n6298), .B(n6297), .ZN(U3139)
         );
  OR2_X1 U7252 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  AND2_X1 U7253 ( .A1(n6302), .A2(n6306), .ZN(n6312) );
  OAI22_X1 U7254 ( .A1(n6312), .A2(n6305), .B1(n6304), .B2(n6303), .ZN(n6362)
         );
  INV_X1 U7255 ( .A(n6306), .ZN(n6361) );
  AOI22_X1 U7256 ( .A1(n6308), .A2(n6362), .B1(n6361), .B2(n6307), .ZN(n6320)
         );
  INV_X1 U7257 ( .A(n6309), .ZN(n6311) );
  OAI21_X1 U7258 ( .B1(n6311), .B2(n5499), .A(n6310), .ZN(n6313) );
  NAND2_X1 U7259 ( .A1(n6313), .A2(n6312), .ZN(n6315) );
  OAI211_X1 U7260 ( .C1(n6317), .C2(n6316), .A(n6315), .B(n6314), .ZN(n6366)
         );
  AOI22_X1 U7261 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6366), .B1(n6318), 
        .B2(n6364), .ZN(n6319) );
  OAI211_X1 U7262 ( .C1(n6321), .C2(n6369), .A(n6320), .B(n6319), .ZN(U3140)
         );
  AOI22_X1 U7263 ( .A1(n6323), .A2(n6362), .B1(n6361), .B2(n6322), .ZN(n6326)
         );
  AOI22_X1 U7264 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6366), .B1(n6324), 
        .B2(n6354), .ZN(n6325) );
  OAI211_X1 U7265 ( .C1(n6327), .C2(n6358), .A(n6326), .B(n6325), .ZN(U3141)
         );
  AOI22_X1 U7266 ( .A1(n6329), .A2(n6362), .B1(n6361), .B2(n6328), .ZN(n6332)
         );
  AOI22_X1 U7267 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6366), .B1(n6330), 
        .B2(n6364), .ZN(n6331) );
  OAI211_X1 U7268 ( .C1(n6333), .C2(n6369), .A(n6332), .B(n6331), .ZN(U3142)
         );
  AOI22_X1 U7269 ( .A1(n6335), .A2(n6362), .B1(n6361), .B2(n6334), .ZN(n6338)
         );
  AOI22_X1 U7270 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6366), .B1(n6336), 
        .B2(n6364), .ZN(n6337) );
  OAI211_X1 U7271 ( .C1(n6339), .C2(n6369), .A(n6338), .B(n6337), .ZN(U3143)
         );
  AOI22_X1 U7272 ( .A1(n6341), .A2(n6362), .B1(n6361), .B2(n6340), .ZN(n6344)
         );
  AOI22_X1 U7273 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6366), .B1(n6342), 
        .B2(n6364), .ZN(n6343) );
  OAI211_X1 U7274 ( .C1(n6345), .C2(n6369), .A(n6344), .B(n6343), .ZN(U3144)
         );
  AOI22_X1 U7275 ( .A1(n6347), .A2(n6362), .B1(n6361), .B2(n6346), .ZN(n6350)
         );
  AOI22_X1 U7276 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6366), .B1(n6348), 
        .B2(n6354), .ZN(n6349) );
  OAI211_X1 U7277 ( .C1(n6351), .C2(n6358), .A(n6350), .B(n6349), .ZN(U3145)
         );
  AOI22_X1 U7278 ( .A1(n6353), .A2(n6362), .B1(n6361), .B2(n6352), .ZN(n6357)
         );
  AOI22_X1 U7279 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6366), .B1(n6355), 
        .B2(n6354), .ZN(n6356) );
  OAI211_X1 U7280 ( .C1(n6359), .C2(n6358), .A(n6357), .B(n6356), .ZN(U3146)
         );
  AOI22_X1 U7281 ( .A1(n6363), .A2(n6362), .B1(n6361), .B2(n6360), .ZN(n6368)
         );
  AOI22_X1 U7282 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6366), .B1(n6365), 
        .B2(n6364), .ZN(n6367) );
  OAI211_X1 U7283 ( .C1(n6370), .C2(n6369), .A(n6368), .B(n6367), .ZN(U3147)
         );
  AOI22_X1 U7284 ( .A1(n3029), .A2(n6372), .B1(n6371), .B2(n3095), .ZN(n6506)
         );
  NAND2_X1 U7285 ( .A1(n6373), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6511) );
  AND3_X1 U7286 ( .A1(n6506), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6511), 
        .ZN(n6377) );
  NAND2_X1 U7287 ( .A1(n6375), .A2(n6374), .ZN(n6376) );
  AOI222_X1 U7288 ( .A1(n6377), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n6377), .B2(n6376), .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6376), 
        .ZN(n6382) );
  INV_X1 U7289 ( .A(n6382), .ZN(n6379) );
  OAI21_X1 U7290 ( .B1(n6379), .B2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n6378), 
        .ZN(n6380) );
  OAI21_X1 U7291 ( .B1(n6382), .B2(n6381), .A(n6380), .ZN(n6384) );
  INV_X1 U7292 ( .A(n6384), .ZN(n6387) );
  INV_X1 U7293 ( .A(n6383), .ZN(n6386) );
  AOI21_X1 U7294 ( .B1(n6384), .B2(n6383), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n6385) );
  AOI21_X1 U7295 ( .B1(n6387), .B2(n6386), .A(n6385), .ZN(n6404) );
  INV_X1 U7296 ( .A(n6388), .ZN(n6390) );
  NOR3_X1 U7297 ( .A1(n6390), .A2(n6389), .A3(n4238), .ZN(n6394) );
  INV_X1 U7298 ( .A(n6391), .ZN(n6392) );
  OAI22_X1 U7299 ( .A1(n6397), .A2(n6394), .B1(n6393), .B2(n6392), .ZN(n6395)
         );
  AOI21_X1 U7300 ( .B1(n6397), .B2(n6396), .A(n6395), .ZN(n6524) );
  OAI21_X1 U7301 ( .B1(MORE_REG_SCAN_IN), .B2(FLUSH_REG_SCAN_IN), .A(n6398), 
        .ZN(n6399) );
  AND4_X1 U7302 ( .A1(n6401), .A2(n6524), .A3(n6400), .A4(n6399), .ZN(n6402)
         );
  OAI211_X1 U7303 ( .C1(n6404), .C2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n6403), .B(n6402), .ZN(n6410) );
  OAI22_X1 U7304 ( .A1(n6410), .A2(n6418), .B1(n6405), .B2(n6528), .ZN(n6406)
         );
  OAI21_X1 U7305 ( .B1(n6408), .B2(n6407), .A(n6406), .ZN(n6500) );
  OAI21_X1 U7306 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6528), .A(n6500), .ZN(
        n6417) );
  AOI211_X1 U7307 ( .C1(n6411), .C2(n6410), .A(n6409), .B(n6417), .ZN(n6416)
         );
  OAI21_X1 U7308 ( .B1(n6412), .B2(n6424), .A(n6500), .ZN(n6413) );
  AOI22_X1 U7309 ( .A1(n6416), .A2(n6415), .B1(n6414), .B2(n6413), .ZN(U3148)
         );
  NOR2_X1 U7310 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6427) );
  NAND2_X1 U7311 ( .A1(n6417), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6423) );
  OAI21_X1 U7312 ( .B1(READY_N), .B2(n6419), .A(n6418), .ZN(n6421) );
  AOI21_X1 U7313 ( .B1(n6500), .B2(n6421), .A(n6420), .ZN(n6422) );
  OAI21_X1 U7314 ( .B1(n6427), .B2(n6423), .A(n6422), .ZN(U3149) );
  OAI211_X1 U7315 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6528), .A(n6499), .B(
        n6424), .ZN(n6426) );
  OAI21_X1 U7316 ( .B1(n6427), .B2(n6426), .A(n6425), .ZN(U3150) );
  AND2_X1 U7317 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6428), .ZN(U3151) );
  AND2_X1 U7318 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6428), .ZN(U3152) );
  AND2_X1 U7319 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6428), .ZN(U3153) );
  AND2_X1 U7320 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6428), .ZN(U3154) );
  AND2_X1 U7321 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6428), .ZN(U3155) );
  AND2_X1 U7322 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6428), .ZN(U3156) );
  AND2_X1 U7323 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6428), .ZN(U3157) );
  AND2_X1 U7324 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6428), .ZN(U3158) );
  AND2_X1 U7325 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6428), .ZN(U3159) );
  AND2_X1 U7326 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6428), .ZN(U3160) );
  AND2_X1 U7327 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6428), .ZN(U3161) );
  AND2_X1 U7328 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6428), .ZN(U3162) );
  INV_X1 U7329 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6712) );
  NOR2_X1 U7330 ( .A1(n6498), .A2(n6712), .ZN(U3163) );
  AND2_X1 U7331 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6428), .ZN(U3164) );
  INV_X1 U7332 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6553) );
  NOR2_X1 U7333 ( .A1(n6498), .A2(n6553), .ZN(U3165) );
  AND2_X1 U7334 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6428), .ZN(U3166) );
  AND2_X1 U7335 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6428), .ZN(U3167) );
  AND2_X1 U7336 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6428), .ZN(U3168) );
  AND2_X1 U7337 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6428), .ZN(U3169) );
  INV_X1 U7338 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6575) );
  NOR2_X1 U7339 ( .A1(n6498), .A2(n6575), .ZN(U3170) );
  AND2_X1 U7340 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6428), .ZN(U3171) );
  AND2_X1 U7341 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6428), .ZN(U3172) );
  AND2_X1 U7342 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6428), .ZN(U3173) );
  AND2_X1 U7343 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6428), .ZN(U3174) );
  AND2_X1 U7344 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6428), .ZN(U3175) );
  AND2_X1 U7345 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6428), .ZN(U3176) );
  AND2_X1 U7346 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6428), .ZN(U3177) );
  AND2_X1 U7347 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6428), .ZN(U3178) );
  AND2_X1 U7348 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6428), .ZN(U3179) );
  INV_X1 U7349 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6563) );
  NOR2_X1 U7350 ( .A1(n6498), .A2(n6563), .ZN(U3180) );
  NOR2_X1 U7351 ( .A1(n6446), .A2(n6429), .ZN(n6439) );
  INV_X1 U7352 ( .A(HOLD), .ZN(n6681) );
  NOR2_X1 U7353 ( .A1(n6446), .A2(n6681), .ZN(n6436) );
  AOI21_X1 U7354 ( .B1(STATE_REG_1__SCAN_IN), .B2(READY_N), .A(n6436), .ZN(
        n6443) );
  NOR2_X1 U7355 ( .A1(n6429), .A2(n6681), .ZN(n6432) );
  INV_X1 U7356 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6431) );
  INV_X1 U7357 ( .A(NA_N), .ZN(n6440) );
  AOI211_X1 U7358 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6440), .A(
        STATE_REG_0__SCAN_IN), .B(n6439), .ZN(n6445) );
  AOI221_X1 U7359 ( .B1(n6432), .B2(n6537), .C1(n6431), .C2(n6537), .A(n6445), 
        .ZN(n6430) );
  OAI21_X1 U7360 ( .B1(n6439), .B2(n6443), .A(n6430), .ZN(U3181) );
  NOR2_X1 U7361 ( .A1(n6437), .A2(n6431), .ZN(n6441) );
  NOR2_X1 U7362 ( .A1(n6441), .A2(n6432), .ZN(n6435) );
  NAND2_X1 U7363 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6433) );
  OAI211_X1 U7364 ( .C1(n6436), .C2(n6435), .A(n6434), .B(n6433), .ZN(U3182)
         );
  AOI221_X1 U7365 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6528), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6438) );
  AOI221_X1 U7366 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6438), .C2(HOLD), .A(n6437), .ZN(n6444) );
  AOI21_X1 U7367 ( .B1(n6441), .B2(n6440), .A(n6439), .ZN(n6442) );
  OAI22_X1 U7368 ( .A1(n6445), .A2(n6444), .B1(n6443), .B2(n6442), .ZN(U3183)
         );
  NAND2_X1 U7369 ( .A1(n6446), .A2(n6464), .ZN(n6484) );
  AOI22_X1 U7370 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6734), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6537), .ZN(n6447) );
  OAI21_X1 U7371 ( .B1(n6448), .B2(n6484), .A(n6447), .ZN(U3184) );
  AOI22_X1 U7372 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6734), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6537), .ZN(n6449) );
  OAI21_X1 U7373 ( .B1(n6451), .B2(n6484), .A(n6449), .ZN(U3185) );
  INV_X1 U7374 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6666) );
  OAI222_X1 U7375 ( .A1(n6494), .A2(n6451), .B1(n6666), .B2(n6464), .C1(n6450), 
        .C2(n6484), .ZN(U3186) );
  INV_X1 U7376 ( .A(n6484), .ZN(n6733) );
  AOI22_X1 U7377 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6537), .ZN(n6452) );
  OAI21_X1 U7378 ( .B1(n6453), .B2(n6494), .A(n6452), .ZN(U3188) );
  AOI22_X1 U7379 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6734), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6537), .ZN(n6454) );
  OAI21_X1 U7380 ( .B1(n6456), .B2(n6484), .A(n6454), .ZN(U3189) );
  AOI22_X1 U7381 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6537), .ZN(n6455) );
  OAI21_X1 U7382 ( .B1(n6456), .B2(n6494), .A(n6455), .ZN(U3190) );
  AOI22_X1 U7383 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6537), .ZN(n6457) );
  OAI21_X1 U7384 ( .B1(n6458), .B2(n6494), .A(n6457), .ZN(U3191) );
  AOI22_X1 U7385 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6734), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6537), .ZN(n6459) );
  OAI21_X1 U7386 ( .B1(n6460), .B2(n6484), .A(n6459), .ZN(U3192) );
  AOI22_X1 U7387 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6734), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6537), .ZN(n6461) );
  OAI21_X1 U7388 ( .B1(n6670), .B2(n6484), .A(n6461), .ZN(U3193) );
  AOI22_X1 U7389 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6734), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6537), .ZN(n6462) );
  OAI21_X1 U7390 ( .B1(n6465), .B2(n6484), .A(n6462), .ZN(U3194) );
  INV_X1 U7391 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6721) );
  OAI222_X1 U7392 ( .A1(n6494), .A2(n6465), .B1(n6721), .B2(n6464), .C1(n6463), 
        .C2(n6484), .ZN(U3195) );
  AOI222_X1 U7393 ( .A1(n6734), .A2(REIP_REG_13__SCAN_IN), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6537), .C1(REIP_REG_14__SCAN_IN), .C2(
        n6733), .ZN(n6466) );
  INV_X1 U7394 ( .A(n6466), .ZN(U3196) );
  AOI22_X1 U7395 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6734), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6537), .ZN(n6467) );
  OAI21_X1 U7396 ( .B1(n6469), .B2(n6484), .A(n6467), .ZN(U3197) );
  AOI22_X1 U7397 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6537), .ZN(n6468) );
  OAI21_X1 U7398 ( .B1(n6469), .B2(n6494), .A(n6468), .ZN(U3198) );
  AOI22_X1 U7399 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6537), .ZN(n6470) );
  OAI21_X1 U7400 ( .B1(n5469), .B2(n6494), .A(n6470), .ZN(U3199) );
  AOI222_X1 U7401 ( .A1(n6733), .A2(REIP_REG_18__SCAN_IN), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6537), .C1(REIP_REG_17__SCAN_IN), .C2(
        n6734), .ZN(n6471) );
  INV_X1 U7402 ( .A(n6471), .ZN(U3200) );
  AOI22_X1 U7403 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6537), .ZN(n6472) );
  OAI21_X1 U7404 ( .B1(n6473), .B2(n6494), .A(n6472), .ZN(U3201) );
  AOI22_X1 U7405 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6734), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6537), .ZN(n6474) );
  OAI21_X1 U7406 ( .B1(n6476), .B2(n6484), .A(n6474), .ZN(U3202) );
  AOI22_X1 U7407 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6537), .ZN(n6475) );
  OAI21_X1 U7408 ( .B1(n6476), .B2(n6494), .A(n6475), .ZN(U3203) );
  AOI22_X1 U7409 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6537), .ZN(n6477) );
  OAI21_X1 U7410 ( .B1(n6478), .B2(n6494), .A(n6477), .ZN(U3204) );
  AOI22_X1 U7411 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6537), .ZN(n6479) );
  OAI21_X1 U7412 ( .B1(n5423), .B2(n6494), .A(n6479), .ZN(U3205) );
  AOI22_X1 U7413 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6734), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6537), .ZN(n6480) );
  OAI21_X1 U7414 ( .B1(n6482), .B2(n6484), .A(n6480), .ZN(U3206) );
  AOI22_X1 U7415 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6537), .ZN(n6481) );
  OAI21_X1 U7416 ( .B1(n6482), .B2(n6494), .A(n6481), .ZN(U3207) );
  AOI22_X1 U7417 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6734), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6537), .ZN(n6483) );
  OAI21_X1 U7418 ( .B1(n6486), .B2(n6484), .A(n6483), .ZN(U3208) );
  AOI22_X1 U7419 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6537), .ZN(n6485) );
  OAI21_X1 U7420 ( .B1(n6486), .B2(n6494), .A(n6485), .ZN(U3209) );
  AOI22_X1 U7421 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6537), .ZN(n6487) );
  OAI21_X1 U7422 ( .B1(n6488), .B2(n6494), .A(n6487), .ZN(U3210) );
  INV_X1 U7423 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6490) );
  AOI22_X1 U7424 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6537), .ZN(n6489) );
  OAI21_X1 U7425 ( .B1(n6490), .B2(n6494), .A(n6489), .ZN(U3211) );
  AOI22_X1 U7426 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6537), .ZN(n6491) );
  OAI21_X1 U7427 ( .B1(n6492), .B2(n6494), .A(n6491), .ZN(U3212) );
  INV_X1 U7428 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6495) );
  AOI22_X1 U7429 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6537), .ZN(n6493) );
  OAI21_X1 U7430 ( .B1(n6495), .B2(n6494), .A(n6493), .ZN(U3213) );
  MUX2_X1 U7431 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6537), .Z(U3445) );
  MUX2_X1 U7432 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6537), .Z(U3446) );
  MUX2_X1 U7433 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6537), .Z(U3447) );
  MUX2_X1 U7434 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6537), .Z(U3448) );
  OAI21_X1 U7435 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6498), .A(n6497), .ZN(
        n6496) );
  INV_X1 U7436 ( .A(n6496), .ZN(U3451) );
  INV_X1 U7437 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6512) );
  OAI21_X1 U7438 ( .B1(n6498), .B2(n6512), .A(n6497), .ZN(U3452) );
  OAI221_X1 U7439 ( .B1(n6501), .B2(STATE2_REG_0__SCAN_IN), .C1(n6501), .C2(
        n6500), .A(n6499), .ZN(U3453) );
  AOI211_X1 U7440 ( .C1(STATE2_REG_1__SCAN_IN), .C2(n6504), .A(n6503), .B(
        n6502), .ZN(n6505) );
  OAI21_X1 U7441 ( .B1(n6506), .B2(n6510), .A(n6505), .ZN(n6507) );
  OAI21_X1 U7442 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6508), .A(n6507), 
        .ZN(n6509) );
  OAI21_X1 U7443 ( .B1(n6511), .B2(n6510), .A(n6509), .ZN(U3461) );
  INV_X1 U7444 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6695) );
  AOI221_X1 U7445 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6513), .C1(n6695), 
        .C2(n6512), .A(n6519), .ZN(n6517) );
  OAI22_X1 U7446 ( .A1(n6518), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(n6515), 
        .B2(n6514), .ZN(n6516) );
  NOR2_X1 U7447 ( .A1(n6517), .A2(n6516), .ZN(U3468) );
  OAI22_X1 U7448 ( .A1(n6519), .A2(REIP_REG_0__SCAN_IN), .B1(n6518), .B2(
        BYTEENABLE_REG_0__SCAN_IN), .ZN(n6520) );
  INV_X1 U7449 ( .A(n6520), .ZN(U3469) );
  NAND2_X1 U7450 ( .A1(n6537), .A2(W_R_N_REG_SCAN_IN), .ZN(n6521) );
  OAI21_X1 U7451 ( .B1(n6537), .B2(READREQUEST_REG_SCAN_IN), .A(n6521), .ZN(
        U3470) );
  INV_X1 U7452 ( .A(MORE_REG_SCAN_IN), .ZN(n6523) );
  INV_X1 U7453 ( .A(n6525), .ZN(n6522) );
  AOI22_X1 U7454 ( .A1(n6525), .A2(n6524), .B1(n6523), .B2(n6522), .ZN(U3471)
         );
  AOI211_X1 U7455 ( .C1(n6529), .C2(n6528), .A(n6527), .B(n6526), .ZN(n6536)
         );
  OAI211_X1 U7456 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6531), .A(n6530), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6533) );
  AOI21_X1 U7457 ( .B1(n6533), .B2(STATE2_REG_0__SCAN_IN), .A(n6532), .ZN(
        n6535) );
  NAND2_X1 U7458 ( .A1(n6536), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6534) );
  OAI21_X1 U7459 ( .B1(n6536), .B2(n6535), .A(n6534), .ZN(U3472) );
  MUX2_X1 U7460 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6537), .Z(U3473) );
  AOI22_X1 U7461 ( .A1(n6539), .A2(keyinput101), .B1(keyinput96), .B2(n6699), 
        .ZN(n6538) );
  OAI221_X1 U7462 ( .B1(n6539), .B2(keyinput101), .C1(n6699), .C2(keyinput96), 
        .A(n6538), .ZN(n6549) );
  INV_X1 U7463 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6718) );
  AOI22_X1 U7464 ( .A1(n6670), .A2(keyinput73), .B1(n6718), .B2(keyinput125), 
        .ZN(n6540) );
  OAI221_X1 U7465 ( .B1(n6670), .B2(keyinput73), .C1(n6718), .C2(keyinput125), 
        .A(n6540), .ZN(n6548) );
  INV_X1 U7466 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6542) );
  AOI22_X1 U7467 ( .A1(n6543), .A2(keyinput80), .B1(n6542), .B2(keyinput106), 
        .ZN(n6541) );
  OAI221_X1 U7468 ( .B1(n6543), .B2(keyinput80), .C1(n6542), .C2(keyinput106), 
        .A(n6541), .ZN(n6547) );
  XOR2_X1 U7469 ( .A(n4353), .B(keyinput95), .Z(n6545) );
  XNOR2_X1 U7470 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .B(keyinput109), .ZN(n6544) );
  NAND2_X1 U7471 ( .A1(n6545), .A2(n6544), .ZN(n6546) );
  NOR4_X1 U7472 ( .A1(n6549), .A2(n6548), .A3(n6547), .A4(n6546), .ZN(n6588)
         );
  AOI22_X1 U7473 ( .A1(n6695), .A2(keyinput70), .B1(n6551), .B2(keyinput79), 
        .ZN(n6550) );
  OAI221_X1 U7474 ( .B1(n6695), .B2(keyinput70), .C1(n6551), .C2(keyinput79), 
        .A(n6550), .ZN(n6561) );
  AOI22_X1 U7475 ( .A1(n6686), .A2(keyinput78), .B1(keyinput71), .B2(n6553), 
        .ZN(n6552) );
  OAI221_X1 U7476 ( .B1(n6686), .B2(keyinput78), .C1(n6553), .C2(keyinput71), 
        .A(n6552), .ZN(n6560) );
  INV_X1 U7477 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6720) );
  INV_X1 U7478 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6555) );
  AOI22_X1 U7479 ( .A1(n6720), .A2(keyinput115), .B1(n6555), .B2(keyinput104), 
        .ZN(n6554) );
  OAI221_X1 U7480 ( .B1(n6720), .B2(keyinput115), .C1(n6555), .C2(keyinput104), 
        .A(n6554), .ZN(n6559) );
  INV_X1 U7481 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6680) );
  XOR2_X1 U7482 ( .A(n6680), .B(keyinput87), .Z(n6557) );
  XNOR2_X1 U7483 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .B(keyinput108), .ZN(n6556) );
  NAND2_X1 U7484 ( .A1(n6557), .A2(n6556), .ZN(n6558) );
  NOR4_X1 U7485 ( .A1(n6561), .A2(n6560), .A3(n6559), .A4(n6558), .ZN(n6587)
         );
  AOI22_X1 U7486 ( .A1(n6564), .A2(keyinput121), .B1(keyinput123), .B2(n6563), 
        .ZN(n6562) );
  OAI221_X1 U7487 ( .B1(n6564), .B2(keyinput121), .C1(n6563), .C2(keyinput123), 
        .A(n6562), .ZN(n6573) );
  INV_X1 U7488 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n6566) );
  AOI22_X1 U7489 ( .A1(n6566), .A2(keyinput110), .B1(n4356), .B2(keyinput118), 
        .ZN(n6565) );
  OAI221_X1 U7490 ( .B1(n6566), .B2(keyinput110), .C1(n4356), .C2(keyinput118), 
        .A(n6565), .ZN(n6572) );
  INV_X1 U7491 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6568) );
  AOI22_X1 U7492 ( .A1(n6568), .A2(keyinput65), .B1(keyinput124), .B2(n6721), 
        .ZN(n6567) );
  OAI221_X1 U7493 ( .B1(n6568), .B2(keyinput65), .C1(n6721), .C2(keyinput124), 
        .A(n6567), .ZN(n6571) );
  INV_X1 U7494 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6664) );
  INV_X1 U7495 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n6667) );
  AOI22_X1 U7496 ( .A1(n6664), .A2(keyinput116), .B1(n6667), .B2(keyinput89), 
        .ZN(n6569) );
  OAI221_X1 U7497 ( .B1(n6664), .B2(keyinput116), .C1(n6667), .C2(keyinput89), 
        .A(n6569), .ZN(n6570) );
  NOR4_X1 U7498 ( .A1(n6573), .A2(n6572), .A3(n6571), .A4(n6570), .ZN(n6586)
         );
  AOI22_X1 U7499 ( .A1(n6712), .A2(keyinput72), .B1(keyinput127), .B2(n6575), 
        .ZN(n6574) );
  OAI221_X1 U7500 ( .B1(n6712), .B2(keyinput72), .C1(n6575), .C2(keyinput127), 
        .A(n6574), .ZN(n6584) );
  AOI22_X1 U7501 ( .A1(n6696), .A2(keyinput112), .B1(n6577), .B2(keyinput94), 
        .ZN(n6576) );
  OAI221_X1 U7502 ( .B1(n6696), .B2(keyinput112), .C1(n6577), .C2(keyinput94), 
        .A(n6576), .ZN(n6583) );
  INV_X1 U7503 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6687) );
  XOR2_X1 U7504 ( .A(n6687), .B(keyinput86), .Z(n6581) );
  INV_X1 U7505 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6704) );
  XOR2_X1 U7506 ( .A(n6704), .B(keyinput98), .Z(n6580) );
  XNOR2_X1 U7507 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput83), .ZN(
        n6579) );
  XNOR2_X1 U7508 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .B(keyinput90), .ZN(n6578) );
  NAND4_X1 U7509 ( .A1(n6581), .A2(n6580), .A3(n6579), .A4(n6578), .ZN(n6582)
         );
  NOR3_X1 U7510 ( .A1(n6584), .A2(n6583), .A3(n6582), .ZN(n6585) );
  AND4_X1 U7511 ( .A1(n6588), .A2(n6587), .A3(n6586), .A4(n6585), .ZN(n6732)
         );
  OAI22_X1 U7512 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(keyinput122), .B1(
        INSTQUEUE_REG_14__1__SCAN_IN), .B2(keyinput120), .ZN(n6589) );
  AOI221_X1 U7513 ( .B1(INSTQUEUE_REG_9__5__SCAN_IN), .B2(keyinput122), .C1(
        keyinput120), .C2(INSTQUEUE_REG_14__1__SCAN_IN), .A(n6589), .ZN(n6596)
         );
  OAI22_X1 U7514 ( .A1(STATE2_REG_2__SCAN_IN), .A2(keyinput114), .B1(
        keyinput84), .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6590) );
  AOI221_X1 U7515 ( .B1(STATE2_REG_2__SCAN_IN), .B2(keyinput114), .C1(
        INSTQUEUE_REG_6__2__SCAN_IN), .C2(keyinput84), .A(n6590), .ZN(n6595)
         );
  OAI22_X1 U7516 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(keyinput93), .B1(
        BS16_N), .B2(keyinput68), .ZN(n6591) );
  AOI221_X1 U7517 ( .B1(INSTQUEUE_REG_2__6__SCAN_IN), .B2(keyinput93), .C1(
        keyinput68), .C2(BS16_N), .A(n6591), .ZN(n6594) );
  OAI22_X1 U7518 ( .A1(DATAO_REG_1__SCAN_IN), .A2(keyinput119), .B1(
        keyinput111), .B2(ADDRESS_REG_16__SCAN_IN), .ZN(n6592) );
  AOI221_X1 U7519 ( .B1(DATAO_REG_1__SCAN_IN), .B2(keyinput119), .C1(
        ADDRESS_REG_16__SCAN_IN), .C2(keyinput111), .A(n6592), .ZN(n6593) );
  NAND4_X1 U7520 ( .A1(n6596), .A2(n6595), .A3(n6594), .A4(n6593), .ZN(n6624)
         );
  OAI22_X1 U7521 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(keyinput92), .B1(
        DATAO_REG_25__SCAN_IN), .B2(keyinput74), .ZN(n6597) );
  AOI221_X1 U7522 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput92), 
        .C1(keyinput74), .C2(DATAO_REG_25__SCAN_IN), .A(n6597), .ZN(n6604) );
  OAI22_X1 U7523 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(keyinput107), .B1(
        keyinput81), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6598) );
  AOI221_X1 U7524 ( .B1(INSTQUEUE_REG_5__2__SCAN_IN), .B2(keyinput107), .C1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .C2(keyinput81), .A(n6598), .ZN(n6603)
         );
  OAI22_X1 U7525 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(keyinput69), .B1(
        keyinput102), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6599) );
  AOI221_X1 U7526 ( .B1(INSTQUEUE_REG_9__2__SCAN_IN), .B2(keyinput69), .C1(
        INSTADDRPOINTER_REG_2__SCAN_IN), .C2(keyinput102), .A(n6599), .ZN(
        n6602) );
  OAI22_X1 U7527 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(keyinput91), .B1(
        INSTQUEUE_REG_7__2__SCAN_IN), .B2(keyinput76), .ZN(n6600) );
  AOI221_X1 U7528 ( .B1(INSTQUEUE_REG_11__5__SCAN_IN), .B2(keyinput91), .C1(
        keyinput76), .C2(INSTQUEUE_REG_7__2__SCAN_IN), .A(n6600), .ZN(n6601)
         );
  NAND4_X1 U7529 ( .A1(n6604), .A2(n6603), .A3(n6602), .A4(n6601), .ZN(n6623)
         );
  OAI22_X1 U7530 ( .A1(EBX_REG_14__SCAN_IN), .A2(keyinput64), .B1(
        EAX_REG_25__SCAN_IN), .B2(keyinput100), .ZN(n6605) );
  AOI221_X1 U7531 ( .B1(EBX_REG_14__SCAN_IN), .B2(keyinput64), .C1(keyinput100), .C2(EAX_REG_25__SCAN_IN), .A(n6605), .ZN(n6612) );
  OAI22_X1 U7532 ( .A1(REIP_REG_16__SCAN_IN), .A2(keyinput88), .B1(keyinput105), .B2(DATAO_REG_24__SCAN_IN), .ZN(n6606) );
  AOI221_X1 U7533 ( .B1(REIP_REG_16__SCAN_IN), .B2(keyinput88), .C1(
        DATAO_REG_24__SCAN_IN), .C2(keyinput105), .A(n6606), .ZN(n6611) );
  OAI22_X1 U7534 ( .A1(n6701), .A2(keyinput75), .B1(keyinput99), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6607) );
  AOI221_X1 U7535 ( .B1(n6701), .B2(keyinput75), .C1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .C2(keyinput99), .A(n6607), .ZN(n6610) );
  OAI22_X1 U7536 ( .A1(EAX_REG_24__SCAN_IN), .A2(keyinput117), .B1(keyinput85), 
        .B2(DATAI_8_), .ZN(n6608) );
  AOI221_X1 U7537 ( .B1(EAX_REG_24__SCAN_IN), .B2(keyinput117), .C1(DATAI_8_), 
        .C2(keyinput85), .A(n6608), .ZN(n6609) );
  NAND4_X1 U7538 ( .A1(n6612), .A2(n6611), .A3(n6610), .A4(n6609), .ZN(n6622)
         );
  OAI22_X1 U7539 ( .A1(n6645), .A2(keyinput113), .B1(
        INSTADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput103), .ZN(n6613) );
  AOI221_X1 U7540 ( .B1(n6645), .B2(keyinput113), .C1(keyinput103), .C2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A(n6613), .ZN(n6620) );
  OAI22_X1 U7541 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput82), .B1(
        LWORD_REG_10__SCAN_IN), .B2(keyinput66), .ZN(n6614) );
  AOI221_X1 U7542 ( .B1(PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput82), .C1(
        keyinput66), .C2(LWORD_REG_10__SCAN_IN), .A(n6614), .ZN(n6619) );
  OAI22_X1 U7543 ( .A1(ADDRESS_REG_2__SCAN_IN), .A2(keyinput67), .B1(HOLD), 
        .B2(keyinput126), .ZN(n6615) );
  AOI221_X1 U7544 ( .B1(ADDRESS_REG_2__SCAN_IN), .B2(keyinput67), .C1(
        keyinput126), .C2(HOLD), .A(n6615), .ZN(n6618) );
  OAI22_X1 U7545 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(keyinput97), .B1(
        UWORD_REG_14__SCAN_IN), .B2(keyinput77), .ZN(n6616) );
  AOI221_X1 U7546 ( .B1(INSTQUEUE_REG_12__6__SCAN_IN), .B2(keyinput97), .C1(
        keyinput77), .C2(UWORD_REG_14__SCAN_IN), .A(n6616), .ZN(n6617) );
  NAND4_X1 U7547 ( .A1(n6620), .A2(n6619), .A3(n6618), .A4(n6617), .ZN(n6621)
         );
  NOR4_X1 U7548 ( .A1(n6624), .A2(n6623), .A3(n6622), .A4(n6621), .ZN(n6731)
         );
  AOI22_X1 U7549 ( .A1(DATAI_8_), .A2(keyinput21), .B1(EAX_REG_25__SCAN_IN), 
        .B2(keyinput36), .ZN(n6625) );
  OAI221_X1 U7550 ( .B1(DATAI_8_), .B2(keyinput21), .C1(EAX_REG_25__SCAN_IN), 
        .C2(keyinput36), .A(n6625), .ZN(n6632) );
  AOI22_X1 U7551 ( .A1(REIP_REG_17__SCAN_IN), .A2(keyinput15), .B1(
        EAX_REG_11__SCAN_IN), .B2(keyinput57), .ZN(n6626) );
  OAI221_X1 U7552 ( .B1(REIP_REG_17__SCAN_IN), .B2(keyinput15), .C1(
        EAX_REG_11__SCAN_IN), .C2(keyinput57), .A(n6626), .ZN(n6631) );
  AOI22_X1 U7553 ( .A1(EAX_REG_24__SCAN_IN), .A2(keyinput53), .B1(
        INSTADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput30), .ZN(n6627) );
  OAI221_X1 U7554 ( .B1(EAX_REG_24__SCAN_IN), .B2(keyinput53), .C1(
        INSTADDRPOINTER_REG_14__SCAN_IN), .C2(keyinput30), .A(n6627), .ZN(
        n6630) );
  AOI22_X1 U7555 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(keyinput56), .B1(
        INSTQUEUE_REG_1__5__SCAN_IN), .B2(keyinput42), .ZN(n6628) );
  OAI221_X1 U7556 ( .B1(INSTQUEUE_REG_14__1__SCAN_IN), .B2(keyinput56), .C1(
        INSTQUEUE_REG_1__5__SCAN_IN), .C2(keyinput42), .A(n6628), .ZN(n6629)
         );
  NOR4_X1 U7557 ( .A1(n6632), .A2(n6631), .A3(n6630), .A4(n6629), .ZN(n6661)
         );
  AOI22_X1 U7558 ( .A1(UWORD_REG_11__SCAN_IN), .A2(keyinput31), .B1(
        INSTQUEUE_REG_11__5__SCAN_IN), .B2(keyinput27), .ZN(n6633) );
  OAI221_X1 U7559 ( .B1(UWORD_REG_11__SCAN_IN), .B2(keyinput31), .C1(
        INSTQUEUE_REG_11__5__SCAN_IN), .C2(keyinput27), .A(n6633), .ZN(n6640)
         );
  AOI22_X1 U7560 ( .A1(EBX_REG_10__SCAN_IN), .A2(keyinput16), .B1(
        INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput37), .ZN(n6634) );
  OAI221_X1 U7561 ( .B1(EBX_REG_10__SCAN_IN), .B2(keyinput16), .C1(
        INSTADDRPOINTER_REG_27__SCAN_IN), .C2(keyinput37), .A(n6634), .ZN(
        n6639) );
  AOI22_X1 U7562 ( .A1(ADDRESS_REG_16__SCAN_IN), .A2(keyinput47), .B1(
        INSTQUEUE_REG_7__7__SCAN_IN), .B2(keyinput45), .ZN(n6635) );
  OAI221_X1 U7563 ( .B1(ADDRESS_REG_16__SCAN_IN), .B2(keyinput47), .C1(
        INSTQUEUE_REG_7__7__SCAN_IN), .C2(keyinput45), .A(n6635), .ZN(n6638)
         );
  AOI22_X1 U7564 ( .A1(DATAO_REG_1__SCAN_IN), .A2(keyinput55), .B1(
        INSTQUEUE_REG_9__5__SCAN_IN), .B2(keyinput58), .ZN(n6636) );
  OAI221_X1 U7565 ( .B1(DATAO_REG_1__SCAN_IN), .B2(keyinput55), .C1(
        INSTQUEUE_REG_9__5__SCAN_IN), .C2(keyinput58), .A(n6636), .ZN(n6637)
         );
  NOR4_X1 U7566 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .ZN(n6660)
         );
  AOI22_X1 U7567 ( .A1(UWORD_REG_14__SCAN_IN), .A2(keyinput13), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput1), .ZN(n6641) );
  OAI221_X1 U7568 ( .B1(UWORD_REG_14__SCAN_IN), .B2(keyinput13), .C1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .C2(keyinput1), .A(n6641), .ZN(n6649)
         );
  AOI22_X1 U7569 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(keyinput33), .B1(
        STATE2_REG_2__SCAN_IN), .B2(keyinput50), .ZN(n6642) );
  OAI221_X1 U7570 ( .B1(INSTQUEUE_REG_12__6__SCAN_IN), .B2(keyinput33), .C1(
        STATE2_REG_2__SCAN_IN), .C2(keyinput50), .A(n6642), .ZN(n6648) );
  AOI22_X1 U7571 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(keyinput63), .B1(
        DATAO_REG_10__SCAN_IN), .B2(keyinput46), .ZN(n6643) );
  OAI221_X1 U7572 ( .B1(DATAWIDTH_REG_12__SCAN_IN), .B2(keyinput63), .C1(
        DATAO_REG_10__SCAN_IN), .C2(keyinput46), .A(n6643), .ZN(n6647) );
  AOI22_X1 U7573 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(keyinput19), .B1(
        n6645), .B2(keyinput49), .ZN(n6644) );
  OAI221_X1 U7574 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(keyinput19), 
        .C1(n6645), .C2(keyinput49), .A(n6644), .ZN(n6646) );
  NOR4_X1 U7575 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .ZN(n6659)
         );
  AOI22_X1 U7576 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(keyinput59), .B1(
        DATAWIDTH_REG_17__SCAN_IN), .B2(keyinput7), .ZN(n6650) );
  OAI221_X1 U7577 ( .B1(DATAWIDTH_REG_2__SCAN_IN), .B2(keyinput59), .C1(
        DATAWIDTH_REG_17__SCAN_IN), .C2(keyinput7), .A(n6650), .ZN(n6657) );
  AOI22_X1 U7578 ( .A1(UWORD_REG_13__SCAN_IN), .A2(keyinput54), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput18), .ZN(n6651) );
  OAI221_X1 U7579 ( .B1(UWORD_REG_13__SCAN_IN), .B2(keyinput54), .C1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .C2(keyinput18), .A(n6651), .ZN(n6656) );
  AOI22_X1 U7580 ( .A1(DATAO_REG_25__SCAN_IN), .A2(keyinput10), .B1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput28), .ZN(n6652) );
  OAI221_X1 U7581 ( .B1(DATAO_REG_25__SCAN_IN), .B2(keyinput10), .C1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput28), .A(n6652), .ZN(
        n6655) );
  AOI22_X1 U7582 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(keyinput12), .B1(
        INSTQUEUE_REG_11__4__SCAN_IN), .B2(keyinput40), .ZN(n6653) );
  OAI221_X1 U7583 ( .B1(INSTQUEUE_REG_7__2__SCAN_IN), .B2(keyinput12), .C1(
        INSTQUEUE_REG_11__4__SCAN_IN), .C2(keyinput40), .A(n6653), .ZN(n6654)
         );
  NOR4_X1 U7584 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6658)
         );
  NAND4_X1 U7585 ( .A1(n6661), .A2(n6660), .A3(n6659), .A4(n6658), .ZN(n6730)
         );
  AOI22_X1 U7586 ( .A1(n6664), .A2(keyinput52), .B1(n6663), .B2(keyinput2), 
        .ZN(n6662) );
  OAI221_X1 U7587 ( .B1(n6664), .B2(keyinput52), .C1(n6663), .C2(keyinput2), 
        .A(n6662), .ZN(n6677) );
  AOI22_X1 U7588 ( .A1(n6667), .A2(keyinput25), .B1(keyinput3), .B2(n6666), 
        .ZN(n6665) );
  OAI221_X1 U7589 ( .B1(n6667), .B2(keyinput25), .C1(n6666), .C2(keyinput3), 
        .A(n6665), .ZN(n6676) );
  AOI22_X1 U7590 ( .A1(n6670), .A2(keyinput9), .B1(n6669), .B2(keyinput38), 
        .ZN(n6668) );
  OAI221_X1 U7591 ( .B1(n6670), .B2(keyinput9), .C1(n6669), .C2(keyinput38), 
        .A(n6668), .ZN(n6675) );
  INV_X1 U7592 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n6671) );
  XOR2_X1 U7593 ( .A(keyinput41), .B(n6671), .Z(n6673) );
  XNOR2_X1 U7594 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .B(keyinput44), .ZN(n6672)
         );
  NAND2_X1 U7595 ( .A1(n6673), .A2(n6672), .ZN(n6674) );
  NOR4_X1 U7596 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n6728)
         );
  AOI22_X1 U7597 ( .A1(n6680), .A2(keyinput23), .B1(keyinput0), .B2(n6679), 
        .ZN(n6678) );
  OAI221_X1 U7598 ( .B1(n6680), .B2(keyinput23), .C1(n6679), .C2(keyinput0), 
        .A(n6678), .ZN(n6684) );
  XOR2_X1 U7599 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .B(keyinput29), .Z(n6683)
         );
  XNOR2_X1 U7600 ( .A(n6681), .B(keyinput62), .ZN(n6682) );
  OR3_X1 U7601 ( .A1(n6684), .A2(n6683), .A3(n6682), .ZN(n6693) );
  AOI22_X1 U7602 ( .A1(n6687), .A2(keyinput22), .B1(keyinput14), .B2(n6686), 
        .ZN(n6685) );
  OAI221_X1 U7603 ( .B1(n6687), .B2(keyinput22), .C1(n6686), .C2(keyinput14), 
        .A(n6685), .ZN(n6692) );
  INV_X1 U7604 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6690) );
  AOI22_X1 U7605 ( .A1(n6690), .A2(keyinput43), .B1(keyinput5), .B2(n6689), 
        .ZN(n6688) );
  OAI221_X1 U7606 ( .B1(n6690), .B2(keyinput43), .C1(n6689), .C2(keyinput5), 
        .A(n6688), .ZN(n6691) );
  NOR3_X1 U7607 ( .A1(n6693), .A2(n6692), .A3(n6691), .ZN(n6727) );
  AOI22_X1 U7608 ( .A1(n6696), .A2(keyinput48), .B1(keyinput6), .B2(n6695), 
        .ZN(n6694) );
  OAI221_X1 U7609 ( .B1(n6696), .B2(keyinput48), .C1(n6695), .C2(keyinput6), 
        .A(n6694), .ZN(n6708) );
  AOI22_X1 U7610 ( .A1(n6699), .A2(keyinput32), .B1(n6698), .B2(keyinput39), 
        .ZN(n6697) );
  OAI221_X1 U7611 ( .B1(n6699), .B2(keyinput32), .C1(n6698), .C2(keyinput39), 
        .A(n6697), .ZN(n6707) );
  AOI22_X1 U7612 ( .A1(n6702), .A2(keyinput17), .B1(n6701), .B2(keyinput11), 
        .ZN(n6700) );
  OAI221_X1 U7613 ( .B1(n6702), .B2(keyinput17), .C1(n6701), .C2(keyinput11), 
        .A(n6700), .ZN(n6706) );
  AOI22_X1 U7614 ( .A1(n5469), .A2(keyinput24), .B1(n6704), .B2(keyinput34), 
        .ZN(n6703) );
  OAI221_X1 U7615 ( .B1(n5469), .B2(keyinput24), .C1(n6704), .C2(keyinput34), 
        .A(n6703), .ZN(n6705) );
  NOR4_X1 U7616 ( .A1(n6708), .A2(n6707), .A3(n6706), .A4(n6705), .ZN(n6726)
         );
  INV_X1 U7617 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6710) );
  AOI22_X1 U7618 ( .A1(n6711), .A2(keyinput35), .B1(n6710), .B2(keyinput20), 
        .ZN(n6709) );
  OAI221_X1 U7619 ( .B1(n6711), .B2(keyinput35), .C1(n6710), .C2(keyinput20), 
        .A(n6709), .ZN(n6715) );
  XOR2_X1 U7620 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .B(keyinput26), .Z(n6714)
         );
  XNOR2_X1 U7621 ( .A(n6712), .B(keyinput8), .ZN(n6713) );
  OR3_X1 U7622 ( .A1(n6715), .A2(n6714), .A3(n6713), .ZN(n6724) );
  INV_X1 U7623 ( .A(BS16_N), .ZN(n6717) );
  AOI22_X1 U7624 ( .A1(n6718), .A2(keyinput61), .B1(keyinput4), .B2(n6717), 
        .ZN(n6716) );
  OAI221_X1 U7625 ( .B1(n6718), .B2(keyinput61), .C1(n6717), .C2(keyinput4), 
        .A(n6716), .ZN(n6723) );
  AOI22_X1 U7626 ( .A1(n6721), .A2(keyinput60), .B1(n6720), .B2(keyinput51), 
        .ZN(n6719) );
  OAI221_X1 U7627 ( .B1(n6721), .B2(keyinput60), .C1(n6720), .C2(keyinput51), 
        .A(n6719), .ZN(n6722) );
  NOR3_X1 U7628 ( .A1(n6724), .A2(n6723), .A3(n6722), .ZN(n6725) );
  NAND4_X1 U7629 ( .A1(n6728), .A2(n6727), .A3(n6726), .A4(n6725), .ZN(n6729)
         );
  AOI211_X1 U7630 ( .C1(n6732), .C2(n6731), .A(n6730), .B(n6729), .ZN(n6736)
         );
  AOI222_X1 U7631 ( .A1(n6537), .A2(ADDRESS_REG_3__SCAN_IN), .B1(
        REIP_REG_4__SCAN_IN), .B2(n6734), .C1(REIP_REG_5__SCAN_IN), .C2(n6733), 
        .ZN(n6735) );
  XNOR2_X1 U7632 ( .A(n6736), .B(n6735), .ZN(U3187) );
  CLKBUF_X1 U34460 ( .A(n3220), .Z(n4831) );
  CLKBUF_X1 U3457 ( .A(n3318), .Z(n3005) );
  INV_X1 U3534 ( .A(n4077), .ZN(n4074) );
endmodule

