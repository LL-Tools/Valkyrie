

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4925;

  CLKBUF_X1 U2383 ( .A(n2715), .Z(n3980) );
  XNOR2_X1 U2384 ( .A(n2210), .B(IR_REG_2__SCAN_IN), .ZN(n4437) );
  NAND2_X1 U2385 ( .A1(n2715), .A2(n4430), .ZN(n3045) );
  INV_X1 U2386 ( .A(n3516), .ZN(n3659) );
  INV_X2 U2387 ( .A(n2150), .ZN(n3656) );
  INV_X1 U2388 ( .A(n4580), .ZN(n3055) );
  AND2_X1 U2389 ( .A1(n3918), .A2(n3915), .ZN(n3879) );
  OAI21_X1 U2390 ( .B1(n3188), .B2(n3932), .A(n3930), .ZN(n3197) );
  NAND2_X1 U2391 ( .A1(n2451), .A2(IR_REG_31__SCAN_IN), .ZN(n2210) );
  AND3_X1 U2392 ( .A1(n2426), .A2(n2160), .A3(n2409), .ZN(n2141) );
  INV_X4 U2393 ( .A(n2142), .ZN(n2698) );
  NOR2_X2 U2395 ( .A1(n2159), .A2(n2867), .ZN(n2866) );
  XNOR2_X2 U2396 ( .A(n2763), .B(n2762), .ZN(n2828) );
  OR2_X1 U2397 ( .A1(n3342), .A2(n3872), .ZN(n3343) );
  OR2_X1 U2398 ( .A1(n4088), .A2(n4423), .ZN(n2813) );
  NAND2_X1 U2399 ( .A1(n2327), .A2(n3924), .ZN(n3172) );
  NAND2_X1 U2400 ( .A1(n2348), .A2(n2347), .ZN(n3011) );
  NAND2_X2 U2401 ( .A1(n2919), .A2(n4531), .ZN(n3801) );
  OR2_X1 U2402 ( .A1(n2861), .A2(n4797), .ZN(n2348) );
  INV_X2 U2403 ( .A(n4661), .ZN(n2143) );
  AND3_X1 U2404 ( .A1(n2467), .A2(n2466), .A3(n2465), .ZN(n2964) );
  INV_X2 U2405 ( .A(n4002), .ZN(U4043) );
  INV_X1 U2406 ( .A(n2981), .ZN(n3056) );
  NAND2_X1 U2407 ( .A1(n3980), .A2(n2937), .ZN(n4375) );
  CLKBUF_X3 U2408 ( .A(n2462), .Z(n2944) );
  NAND2_X1 U2409 ( .A1(n2822), .A2(n2819), .ZN(n2468) );
  XNOR2_X1 U2410 ( .A(n2707), .B(n2706), .ZN(n2715) );
  CLKBUF_X3 U2411 ( .A(n2458), .Z(n2636) );
  INV_X1 U2412 ( .A(n2752), .ZN(n4430) );
  NAND2_X1 U2413 ( .A1(n2705), .A2(IR_REG_31__SCAN_IN), .ZN(n2707) );
  OR2_X1 U2414 ( .A1(n2761), .A2(n2760), .ZN(n2772) );
  OR2_X1 U2415 ( .A1(n2434), .A2(n2431), .ZN(n2432) );
  NAND2_X1 U2416 ( .A1(n2768), .A2(IR_REG_31__SCAN_IN), .ZN(n2763) );
  OR2_X1 U2417 ( .A1(n2760), .A2(n2431), .ZN(n2764) );
  AND2_X1 U2418 ( .A1(n2565), .A2(n2427), .ZN(n2308) );
  AND4_X1 U2419 ( .A1(n2618), .A2(n2425), .A3(n2424), .A4(n2423), .ZN(n2426)
         );
  NOR2_X1 U2420 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2618)
         );
  NOR2_X1 U2422 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2365)
         );
  NOR2_X1 U2423 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2232)
         );
  NOR2_X1 U2424 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2231)
         );
  NOR2_X1 U2425 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2425)
         );
  NOR2_X1 U2426 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2424)
         );
  NOR2_X1 U2427 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2423)
         );
  INV_X1 U2428 ( .A(IR_REG_20__SCAN_IN), .ZN(n2706) );
  NAND2_X1 U2429 ( .A1(n4162), .A2(n3701), .ZN(n2281) );
  INV_X1 U2430 ( .A(n3875), .ZN(n2272) );
  INV_X1 U2431 ( .A(n3675), .ZN(n3027) );
  AND2_X1 U2432 ( .A1(n2892), .A2(n2891), .ZN(n3514) );
  NOR2_X1 U2433 ( .A1(n3777), .A2(n2399), .ZN(n2398) );
  NOR2_X1 U2434 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2234)
         );
  NOR2_X1 U2435 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2233)
         );
  INV_X1 U2436 ( .A(n3890), .ZN(n2291) );
  AOI21_X1 U2437 ( .B1(n3925), .B2(n2516), .A(n2176), .ZN(n2305) );
  NAND2_X1 U2438 ( .A1(n4001), .A2(n4572), .ZN(n3922) );
  NAND2_X1 U2439 ( .A1(n2262), .A2(n3063), .ZN(n4589) );
  AND2_X1 U2440 ( .A1(n2478), .A2(n3062), .ZN(n2262) );
  AND2_X1 U2441 ( .A1(n2819), .A2(n2436), .ZN(n2462) );
  AND2_X1 U2442 ( .A1(n3922), .A2(n3919), .ZN(n4590) );
  AND2_X1 U2443 ( .A1(n2330), .A2(n2404), .ZN(n2329) );
  AND2_X1 U2444 ( .A1(n2620), .A2(n2567), .ZN(n2209) );
  INV_X1 U2445 ( .A(n2390), .ZN(n2386) );
  NAND2_X1 U2446 ( .A1(n3654), .A2(n2369), .ZN(n2195) );
  INV_X1 U2447 ( .A(n3767), .ZN(n2206) );
  XNOR2_X1 U2448 ( .A(n2346), .B(n2932), .ZN(n2929) );
  AOI21_X1 U2449 ( .B1(n2319), .B2(n2323), .A(n2317), .ZN(n2316) );
  INV_X1 U2450 ( .A(n2319), .ZN(n2318) );
  AND2_X1 U2451 ( .A1(n2321), .A2(n3848), .ZN(n2319) );
  AND2_X1 U2452 ( .A1(n2291), .A2(n2690), .ZN(n2287) );
  AND2_X1 U2453 ( .A1(n4165), .A2(n4319), .ZN(n2689) );
  NAND2_X1 U2454 ( .A1(n4151), .A2(n4170), .ZN(n2681) );
  AOI21_X1 U2455 ( .B1(n2277), .B2(n2278), .A(n2161), .ZN(n2276) );
  INV_X1 U2457 ( .A(n2292), .ZN(n4219) );
  AND2_X1 U2458 ( .A1(n2297), .A2(n2301), .ZN(n2296) );
  NAND2_X1 U2459 ( .A1(n2294), .A2(n3898), .ZN(n2293) );
  AOI21_X1 U2460 ( .B1(n2313), .B2(n2315), .A(n2311), .ZN(n2310) );
  INV_X1 U2461 ( .A(n3824), .ZN(n2311) );
  INV_X1 U2462 ( .A(n2267), .ZN(n2266) );
  AOI21_X1 U2463 ( .B1(n2268), .B2(n2547), .A(n2148), .ZN(n2267) );
  OAI21_X1 U2464 ( .B1(n3190), .B2(n2536), .A(n2535), .ZN(n3198) );
  NAND2_X1 U2465 ( .A1(n2724), .A2(n3927), .ZN(n3188) );
  OAI22_X1 U2466 ( .A1(n3137), .A2(n2506), .B1(n3163), .B2(n4000), .ZN(n3184)
         );
  OAI21_X1 U2467 ( .B1(n2794), .B2(n2179), .A(n2250), .ZN(n2247) );
  NOR2_X1 U2468 ( .A1(n4090), .A2(n4598), .ZN(n2250) );
  NAND2_X1 U2469 ( .A1(n2705), .A2(n2648), .ZN(n4081) );
  NOR2_X1 U2470 ( .A1(n4075), .A2(n4076), .ZN(n4526) );
  NAND2_X1 U2471 ( .A1(n4526), .A2(n4527), .ZN(n4524) );
  NAND2_X1 U2472 ( .A1(n2969), .A2(n2236), .ZN(n3909) );
  INV_X1 U2473 ( .A(IR_REG_27__SCAN_IN), .ZN(n2430) );
  INV_X1 U2474 ( .A(IR_REG_28__SCAN_IN), .ZN(n2429) );
  NOR2_X1 U2475 ( .A1(n2675), .A2(n4702), .ZN(n2683) );
  NAND2_X1 U2476 ( .A1(n4471), .A2(n3263), .ZN(n3265) );
  NOR2_X1 U2477 ( .A1(n4499), .A2(n2221), .ZN(n4058) );
  AND2_X1 U2478 ( .A1(n4056), .A2(REG2_REG_15__SCAN_IN), .ZN(n2221) );
  OR2_X1 U2479 ( .A1(n2571), .A2(n4623), .ZN(n2584) );
  AND3_X1 U2480 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2499) );
  NAND2_X1 U2481 ( .A1(n2964), .A2(n2981), .ZN(n3913) );
  AND2_X1 U2482 ( .A1(n2936), .A2(n2985), .ZN(n2991) );
  INV_X1 U2483 ( .A(n2825), .ZN(n2785) );
  NAND2_X1 U2484 ( .A1(n2170), .A2(n2299), .ZN(n2298) );
  NAND2_X1 U2485 ( .A1(n2300), .A2(n2649), .ZN(n2299) );
  INV_X1 U2486 ( .A(n2638), .ZN(n2300) );
  AND2_X1 U2487 ( .A1(n4278), .A2(n2649), .ZN(n2301) );
  AND2_X1 U2488 ( .A1(n2334), .A2(n3557), .ZN(n2333) );
  NOR2_X1 U2489 ( .A1(n3501), .A2(n3523), .ZN(n2334) );
  NAND2_X1 U2490 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2756) );
  AND2_X1 U2491 ( .A1(n2426), .A2(n2160), .ZN(n2405) );
  INV_X1 U2492 ( .A(IR_REG_21__SCAN_IN), .ZN(n4731) );
  AND2_X1 U2493 ( .A1(n2209), .A2(n2208), .ZN(n2207) );
  INV_X1 U2494 ( .A(IR_REG_17__SCAN_IN), .ZN(n2208) );
  OR2_X1 U2495 ( .A1(n2555), .A2(IR_REG_10__SCAN_IN), .ZN(n2556) );
  INV_X1 U2496 ( .A(IR_REG_2__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U2497 ( .A1(n2368), .A2(n3796), .ZN(n2367) );
  INV_X1 U2498 ( .A(n2370), .ZN(n2368) );
  NOR2_X1 U2499 ( .A1(n2388), .A2(n2383), .ZN(n2382) );
  INV_X1 U2500 ( .A(n3737), .ZN(n2383) );
  AND2_X1 U2501 ( .A1(n2369), .A2(n3651), .ZN(n2188) );
  NOR2_X1 U2502 ( .A1(n2153), .A2(n3691), .ZN(n2192) );
  AOI21_X1 U2503 ( .B1(n2969), .B2(n3670), .A(n2968), .ZN(n2975) );
  AOI21_X1 U2504 ( .B1(n2896), .B2(n3514), .A(n2154), .ZN(n2970) );
  NAND2_X1 U2505 ( .A1(n2654), .A2(REG3_REG_21__SCAN_IN), .ZN(n2659) );
  OAI21_X1 U2506 ( .B1(n3716), .B2(n2180), .A(n2394), .ZN(n3758) );
  AOI21_X1 U2507 ( .B1(n3645), .B2(n2395), .A(n2181), .ZN(n2394) );
  INV_X1 U2508 ( .A(n2398), .ZN(n2395) );
  OAI21_X1 U2509 ( .B1(n3115), .B2(n3516), .A(n3076), .ZN(n3077) );
  AND2_X1 U2510 ( .A1(n3498), .A2(n3497), .ZN(n3552) );
  NOR2_X1 U2511 ( .A1(n3576), .A2(n2391), .ZN(n2390) );
  INV_X1 U2512 ( .A(n3570), .ZN(n2391) );
  NAND2_X1 U2513 ( .A1(n2371), .A2(n2171), .ZN(n2370) );
  INV_X1 U2514 ( .A(n3725), .ZN(n2371) );
  AND2_X1 U2515 ( .A1(n4430), .A2(n4429), .ZN(n2905) );
  AOI21_X1 U2516 ( .B1(n4034), .B2(REG2_REG_3__SCAN_IN), .A(n2219), .ZN(n2851)
         );
  NOR2_X1 U2517 ( .A1(n2220), .A2(n2858), .ZN(n2219) );
  OR2_X1 U2518 ( .A1(n2870), .A2(n2869), .ZN(n2354) );
  NAND2_X1 U2519 ( .A1(n4031), .A2(n2860), .ZN(n2346) );
  XNOR2_X1 U2520 ( .A(n2876), .B(n2349), .ZN(n2861) );
  INV_X1 U2521 ( .A(n3011), .ZN(n3013) );
  OAI21_X1 U2522 ( .B1(n3259), .B2(n2224), .A(n2222), .ZN(n3261) );
  AOI21_X1 U2523 ( .B1(n2225), .B2(n2223), .A(n2169), .ZN(n2222) );
  INV_X1 U2524 ( .A(n2225), .ZN(n2224) );
  NAND2_X1 U2525 ( .A1(n4459), .A2(REG2_REG_10__SCAN_IN), .ZN(n4458) );
  NAND2_X1 U2526 ( .A1(n4504), .A2(n4045), .ZN(n4046) );
  NAND2_X1 U2527 ( .A1(n4071), .A2(n2360), .ZN(n2359) );
  NAND2_X1 U2528 ( .A1(n4063), .A2(n2361), .ZN(n2360) );
  INV_X1 U2529 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2361) );
  NOR2_X1 U2530 ( .A1(n3904), .A2(n3893), .ZN(n2256) );
  INV_X1 U2531 ( .A(n2258), .ZN(n2252) );
  OR2_X1 U2532 ( .A1(n2324), .A2(n3852), .ZN(n2321) );
  AND2_X1 U2533 ( .A1(n2326), .A2(n4110), .ZN(n2324) );
  NAND2_X1 U2534 ( .A1(n3799), .A2(n4145), .ZN(n2690) );
  NAND2_X1 U2535 ( .A1(n2279), .A2(n2281), .ZN(n2277) );
  NAND2_X1 U2536 ( .A1(n2666), .A2(n2281), .ZN(n2278) );
  AOI22_X1 U2537 ( .A1(n4219), .A2(n2658), .B1(n4238), .B2(n4221), .ZN(n4211)
         );
  AND2_X1 U2538 ( .A1(n2650), .A2(REG3_REG_20__SCAN_IN), .ZN(n2654) );
  AND2_X1 U2539 ( .A1(n2297), .A2(n3898), .ZN(n4239) );
  AOI21_X1 U2540 ( .B1(n3477), .B2(n2627), .A(n2626), .ZN(n4275) );
  NAND2_X1 U2541 ( .A1(n4275), .A2(n4278), .ZN(n4274) );
  INV_X1 U2542 ( .A(n2265), .ZN(n2264) );
  OAI21_X1 U2543 ( .B1(n2144), .B2(n2151), .A(n3331), .ZN(n2265) );
  NAND2_X1 U2544 ( .A1(n2271), .A2(n2270), .ZN(n2269) );
  INV_X1 U2545 ( .A(n3198), .ZN(n2271) );
  NAND2_X1 U2546 ( .A1(n2269), .A2(n2268), .ZN(n3356) );
  NAND2_X1 U2547 ( .A1(n3197), .A2(n3945), .ZN(n2725) );
  AND2_X1 U2548 ( .A1(n3364), .A2(n3366), .ZN(n3875) );
  AOI21_X1 U2549 ( .B1(n2305), .B2(n2303), .A(n2177), .ZN(n2302) );
  INV_X1 U2550 ( .A(n2305), .ZN(n2304) );
  OAI21_X1 U2551 ( .B1(n3172), .B2(n2723), .A(n3928), .ZN(n3208) );
  AND2_X1 U2552 ( .A1(n2722), .A2(n3928), .ZN(n3925) );
  NAND2_X1 U2553 ( .A1(n2498), .A2(n2497), .ZN(n3137) );
  OAI21_X1 U2554 ( .B1(n4575), .B2(n2721), .A(n3922), .ZN(n3102) );
  AND2_X1 U2555 ( .A1(n2239), .A2(n2238), .ZN(n2241) );
  NOR2_X1 U2556 ( .A1(n2237), .A2(n2236), .ZN(n2235) );
  INV_X1 U2557 ( .A(n2452), .ZN(n2237) );
  NAND2_X1 U2558 ( .A1(n3984), .A2(n2744), .ZN(n4282) );
  NOR2_X1 U2559 ( .A1(n4300), .A2(n4303), .ZN(n4301) );
  OAI21_X1 U2560 ( .B1(n2254), .B2(n2256), .A(n4593), .ZN(n2243) );
  NAND2_X1 U2561 ( .A1(n2704), .A2(n2168), .ZN(n2794) );
  NAND2_X1 U2562 ( .A1(n2282), .A2(n2284), .ZN(n2704) );
  AOI21_X1 U2563 ( .B1(n2285), .B2(n2286), .A(n2178), .ZN(n2284) );
  NAND2_X1 U2564 ( .A1(n2255), .A2(n2257), .ZN(n2254) );
  NAND2_X1 U2565 ( .A1(n2261), .A2(n2167), .ZN(n2257) );
  NAND2_X1 U2566 ( .A1(n3893), .A2(n2258), .ZN(n2255) );
  OR2_X1 U2567 ( .A1(n2807), .A2(n3840), .ZN(n4300) );
  NAND2_X1 U2568 ( .A1(n4115), .A2(n3674), .ZN(n2807) );
  NOR2_X1 U2569 ( .A1(n4132), .A2(n4307), .ZN(n4115) );
  NAND2_X1 U2570 ( .A1(n4211), .A2(n4210), .ZN(n4337) );
  INV_X1 U2571 ( .A(n3997), .ZN(n3372) );
  INV_X1 U2572 ( .A(n3996), .ZN(n3437) );
  NAND2_X1 U2573 ( .A1(n2435), .A2(n3689), .ZN(n2437) );
  MUX2_X1 U2574 ( .A(IR_REG_31__SCAN_IN), .B(n2433), .S(IR_REG_29__SCAN_IN), 
        .Z(n2435) );
  INV_X1 U2575 ( .A(IR_REG_8__SCAN_IN), .ZN(n4713) );
  INV_X1 U2576 ( .A(IR_REG_1__SCAN_IN), .ZN(n2363) );
  NAND2_X1 U2577 ( .A1(n2376), .A2(n2379), .ZN(n3286) );
  OR2_X1 U2578 ( .A1(n3158), .A2(n2377), .ZN(n2376) );
  NAND2_X1 U2579 ( .A1(n3025), .A2(n3026), .ZN(n2196) );
  AOI21_X1 U2580 ( .B1(n2374), .B2(n2377), .A(n2373), .ZN(n2372) );
  NAND2_X1 U2581 ( .A1(n3158), .A2(n2374), .ZN(n2199) );
  NOR2_X1 U2582 ( .A1(n3283), .A2(n3284), .ZN(n2373) );
  NAND2_X1 U2583 ( .A1(n2978), .A2(n2977), .ZN(n2198) );
  AND2_X1 U2584 ( .A1(n2980), .A2(n2979), .ZN(n3812) );
  OAI21_X1 U2585 ( .B1(n3728), .B2(n2142), .A(n2688), .ZN(n4165) );
  INV_X1 U2586 ( .A(n3115), .ZN(n4001) );
  NAND2_X1 U2587 ( .A1(n2474), .A2(n2473), .ZN(n4580) );
  XNOR2_X1 U2588 ( .A(n2851), .B(n2932), .ZN(n2928) );
  NOR2_X1 U2589 ( .A1(n4515), .A2(REG1_REG_16__SCAN_IN), .ZN(n4516) );
  XNOR2_X1 U2590 ( .A(n4046), .B(n4057), .ZN(n4515) );
  NAND2_X1 U2591 ( .A1(n2358), .A2(n4480), .ZN(n2357) );
  NAND2_X1 U2592 ( .A1(n2359), .A2(n4521), .ZN(n2358) );
  AOI21_X1 U2593 ( .B1(n4523), .B2(ADDR_REG_18__SCAN_IN), .A(n4522), .ZN(n2356) );
  NOR2_X1 U2594 ( .A1(n2359), .A2(n4521), .ZN(n4520) );
  XNOR2_X1 U2595 ( .A(n2343), .B(n4078), .ZN(n4083) );
  NAND2_X1 U2596 ( .A1(n4524), .A2(n2185), .ZN(n2343) );
  AND2_X1 U2597 ( .A1(n2853), .A2(n2922), .ZN(n4525) );
  NOR2_X1 U2598 ( .A1(n4520), .A2(n2230), .ZN(n2229) );
  AND2_X1 U2599 ( .A1(n4074), .A2(REG2_REG_18__SCAN_IN), .ZN(n2230) );
  AOI21_X1 U2600 ( .B1(n2794), .B2(n2256), .A(n2254), .ZN(n2253) );
  OR2_X1 U2601 ( .A1(n2794), .A2(n2252), .ZN(n2251) );
  XOR2_X1 U2602 ( .A(n3860), .B(n2794), .Z(n4094) );
  NAND2_X1 U2603 ( .A1(n3183), .A2(n2516), .ZN(n3207) );
  AND2_X1 U2604 ( .A1(n2143), .A2(n4658), .ZN(n4220) );
  NAND2_X1 U2605 ( .A1(n2918), .A2(n2917), .ZN(n4531) );
  INV_X1 U2606 ( .A(n3548), .ZN(n3549) );
  INV_X1 U2607 ( .A(n2718), .ZN(n3878) );
  INV_X1 U2608 ( .A(IR_REG_22__SCAN_IN), .ZN(n2406) );
  INV_X1 U2609 ( .A(n3645), .ZN(n2396) );
  INV_X1 U2610 ( .A(n2174), .ZN(n2393) );
  INV_X1 U2612 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2880) );
  OR2_X1 U2613 ( .A1(n3258), .A2(n4533), .ZN(n2227) );
  INV_X1 U2614 ( .A(n2227), .ZN(n2223) );
  AOI21_X1 U2615 ( .B1(n3266), .B2(n2214), .A(n2213), .ZN(n2212) );
  AND2_X1 U2616 ( .A1(n3894), .A2(n4157), .ZN(n3965) );
  OR2_X1 U2617 ( .A1(n2295), .A2(n3897), .ZN(n2294) );
  INV_X1 U2618 ( .A(n2298), .ZN(n2295) );
  NAND2_X1 U2619 ( .A1(n2612), .A2(n2415), .ZN(n2629) );
  AOI21_X1 U2620 ( .B1(n2314), .B2(n3954), .A(n3331), .ZN(n2313) );
  INV_X1 U2621 ( .A(n2727), .ZN(n2314) );
  INV_X1 U2622 ( .A(n3954), .ZN(n2315) );
  INV_X1 U2623 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2583) );
  NOR2_X1 U2624 ( .A1(n2549), .A2(n2548), .ZN(n2570) );
  INV_X1 U2625 ( .A(n2516), .ZN(n2303) );
  NOR2_X1 U2626 ( .A1(n2507), .A2(n2880), .ZN(n2517) );
  NAND2_X1 U2627 ( .A1(n2698), .A2(REG3_REG_1__SCAN_IN), .ZN(n2239) );
  NAND2_X1 U2628 ( .A1(n2462), .A2(REG1_REG_1__SCAN_IN), .ZN(n2240) );
  INV_X1 U2629 ( .A(n2287), .ZN(n2285) );
  NOR2_X1 U2630 ( .A1(n2261), .A2(n2167), .ZN(n2258) );
  NAND2_X1 U2631 ( .A1(n2787), .A2(n2637), .ZN(n2337) );
  NAND2_X1 U2632 ( .A1(n3066), .A2(n3918), .ZN(n4575) );
  AND2_X1 U2633 ( .A1(n2428), .A2(n2427), .ZN(n2330) );
  INV_X1 U2634 ( .A(IR_REG_19__SCAN_IN), .ZN(n4730) );
  AND3_X1 U2635 ( .A1(n4720), .A2(n4713), .A3(n2531), .ZN(n2532) );
  INV_X1 U2636 ( .A(IR_REG_6__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U2637 ( .A1(n3225), .A2(n3226), .ZN(n2379) );
  OR2_X1 U2638 ( .A1(n2659), .A2(n4868), .ZN(n2667) );
  INV_X1 U2639 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2537) );
  INV_X1 U2640 ( .A(n3998), .ZN(n3607) );
  AND2_X1 U2641 ( .A1(n2375), .A2(n2379), .ZN(n2374) );
  INV_X1 U2642 ( .A(n3285), .ZN(n2375) );
  NAND2_X1 U2643 ( .A1(n2163), .A2(n2378), .ZN(n2377) );
  INV_X1 U2644 ( .A(n2412), .ZN(n2378) );
  AND2_X1 U2645 ( .A1(n2204), .A2(n3769), .ZN(n2203) );
  NAND2_X1 U2646 ( .A1(n3767), .A2(n2205), .ZN(n2204) );
  INV_X1 U2647 ( .A(n3618), .ZN(n2205) );
  NAND2_X1 U2648 ( .A1(n3569), .A2(n3568), .ZN(n3570) );
  INV_X1 U2649 ( .A(n3567), .ZN(n3568) );
  INV_X1 U2650 ( .A(n3566), .ZN(n3569) );
  NAND2_X1 U2651 ( .A1(n2446), .A2(n2445), .ZN(n2458) );
  OR2_X1 U2652 ( .A1(n2802), .A2(n2410), .ZN(n2446) );
  AND2_X1 U2653 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2410)
         );
  INV_X1 U2654 ( .A(n2893), .ZN(n2894) );
  NAND2_X1 U2655 ( .A1(n3619), .A2(n3618), .ZN(n3766) );
  NOR2_X1 U2656 ( .A1(n3636), .A2(n3717), .ZN(n2399) );
  INV_X1 U2657 ( .A(n4133), .ZN(n3802) );
  OR2_X1 U2658 ( .A1(n3665), .A2(n3664), .ZN(n3796) );
  AND2_X1 U2659 ( .A1(n2592), .A2(REG3_REG_15__SCAN_IN), .ZN(n2612) );
  OR2_X1 U2660 ( .A1(n2691), .A2(n2684), .ZN(n3728) );
  NAND4_X1 U2661 ( .A1(n2457), .A2(n2456), .A3(n2455), .A4(n2454), .ZN(n2896)
         );
  NAND2_X1 U2662 ( .A1(n2462), .A2(REG1_REG_0__SCAN_IN), .ZN(n2454) );
  INV_X1 U2663 ( .A(IR_REG_4__SCAN_IN), .ZN(n2421) );
  NAND2_X1 U2664 ( .A1(n2354), .A2(n2353), .ZN(n2352) );
  NAND2_X1 U2665 ( .A1(n4434), .A2(REG2_REG_5__SCAN_IN), .ZN(n2353) );
  AOI21_X1 U2666 ( .B1(n2884), .B2(REG2_REG_6__SCAN_IN), .A(n2351), .ZN(n2886)
         );
  AND2_X1 U2667 ( .A1(n2352), .A2(n4433), .ZN(n2351) );
  AND2_X1 U2668 ( .A1(n2172), .A2(n4452), .ZN(n2225) );
  NAND2_X1 U2669 ( .A1(n3259), .A2(n2227), .ZN(n2226) );
  NAND2_X1 U2670 ( .A1(n4481), .A2(REG2_REG_12__SCAN_IN), .ZN(n4479) );
  XNOR2_X1 U2671 ( .A(n4053), .B(n4498), .ZN(n4491) );
  OAI21_X1 U2672 ( .B1(REG2_REG_13__SCAN_IN), .B2(n4051), .A(n2350), .ZN(n4053) );
  NAND2_X1 U2673 ( .A1(n2211), .A2(n3255), .ZN(n2350) );
  OAI21_X1 U2674 ( .B1(n2215), .B2(n4481), .A(n2212), .ZN(n2211) );
  INV_X1 U2675 ( .A(n3266), .ZN(n2215) );
  XNOR2_X1 U2676 ( .A(n4058), .B(n4057), .ZN(n4512) );
  NAND2_X1 U2677 ( .A1(n4512), .A2(n4510), .ZN(n4511) );
  AND2_X1 U2678 ( .A1(n3839), .A2(n3862), .ZN(n2325) );
  AND2_X1 U2679 ( .A1(n2743), .A2(n3862), .ZN(n4125) );
  AND2_X1 U2680 ( .A1(n2636), .A2(DATAI_20_), .ZN(n4245) );
  NAND2_X1 U2681 ( .A1(n2312), .A2(n3954), .ZN(n3828) );
  NAND2_X1 U2682 ( .A1(n3367), .A2(n2727), .ZN(n2312) );
  NAND2_X1 U2683 ( .A1(n3138), .A2(n3936), .ZN(n2327) );
  AND2_X1 U2684 ( .A1(n2491), .A2(n2490), .ZN(n4574) );
  AOI22_X1 U2685 ( .A1(n4589), .A2(n2487), .B1(n2488), .B2(n4590), .ZN(n3101)
         );
  INV_X1 U2686 ( .A(IR_REG_23__SCAN_IN), .ZN(n4607) );
  NAND2_X1 U2687 ( .A1(n3067), .A2(n3879), .ZN(n3066) );
  NAND2_X1 U2688 ( .A1(n2146), .A2(n2719), .ZN(n3063) );
  NAND2_X1 U2689 ( .A1(n2718), .A2(n3908), .ZN(n2986) );
  OR2_X1 U2690 ( .A1(n2718), .A2(n2991), .ZN(n2992) );
  AND2_X1 U2691 ( .A1(n2753), .A2(n2752), .ZN(n2937) );
  NOR3_X1 U2692 ( .A1(n4207), .A2(n2340), .A3(n3701), .ZN(n4168) );
  NOR2_X1 U2693 ( .A1(n4207), .A2(n3701), .ZN(n4187) );
  OR2_X1 U2694 ( .A1(n2145), .A2(n4205), .ZN(n4207) );
  AOI21_X1 U2695 ( .B1(n4275), .B2(n2301), .A(n2298), .ZN(n4240) );
  NOR3_X1 U2696 ( .A1(n4285), .A2(n4266), .A3(n4284), .ZN(n4267) );
  AND2_X1 U2697 ( .A1(n3419), .A2(n2149), .ZN(n3478) );
  NAND2_X1 U2698 ( .A1(n3478), .A2(n3572), .ZN(n4285) );
  AND4_X1 U2699 ( .A1(n2607), .A2(n2606), .A3(n2605), .A4(n2604), .ZN(n4368)
         );
  AND4_X1 U2700 ( .A1(n2589), .A2(n2588), .A3(n2587), .A4(n2586), .ZN(n3518)
         );
  NAND2_X1 U2701 ( .A1(n3419), .A2(n2334), .ZN(n3346) );
  INV_X1 U2702 ( .A(n4379), .ZN(n3558) );
  INV_X1 U2703 ( .A(n3523), .ZN(n3517) );
  NAND2_X1 U2704 ( .A1(n3419), .A2(n3418), .ZN(n3421) );
  INV_X1 U2705 ( .A(n3593), .ZN(n3357) );
  AND2_X1 U2706 ( .A1(n3358), .A2(n3357), .ZN(n3419) );
  NOR2_X1 U2707 ( .A1(n3322), .A2(n3398), .ZN(n3358) );
  OR2_X1 U2708 ( .A1(n3199), .A2(n3389), .ZN(n3322) );
  INV_X1 U2709 ( .A(n3296), .ZN(n3292) );
  NAND2_X1 U2710 ( .A1(n3217), .A2(n3292), .ZN(n3199) );
  AND2_X1 U2711 ( .A1(n2520), .A2(n2519), .ZN(n3289) );
  NAND2_X1 U2712 ( .A1(n2331), .A2(n3229), .ZN(n3215) );
  NOR2_X1 U2713 ( .A1(n3215), .A2(n3536), .ZN(n3217) );
  INV_X1 U2714 ( .A(n4282), .ZN(n4576) );
  NOR2_X1 U2715 ( .A1(n4583), .A2(n4582), .ZN(n4586) );
  AND2_X1 U2716 ( .A1(n2911), .A2(n2905), .ZN(n4363) );
  INV_X1 U2717 ( .A(n4362), .ZN(n4571) );
  INV_X1 U2718 ( .A(n4367), .ZN(n4581) );
  AND2_X1 U2719 ( .A1(n2236), .A2(n2939), .ZN(n3007) );
  NAND2_X1 U2720 ( .A1(n3056), .A2(n3007), .ZN(n2342) );
  AND3_X1 U2721 ( .A1(n2782), .A2(n2901), .A3(n3041), .ZN(n2790) );
  NOR2_X1 U2722 ( .A1(n2402), .A2(IR_REG_26__SCAN_IN), .ZN(n2401) );
  NAND2_X1 U2723 ( .A1(n2404), .A2(n2403), .ZN(n2402) );
  INV_X1 U2724 ( .A(IR_REG_29__SCAN_IN), .ZN(n2403) );
  NAND2_X1 U2725 ( .A1(n2443), .A2(IR_REG_31__SCAN_IN), .ZN(n2802) );
  NAND2_X1 U2726 ( .A1(n2757), .A2(n2330), .ZN(n2443) );
  NAND2_X1 U2727 ( .A1(n2759), .A2(n2758), .ZN(n2761) );
  NAND2_X1 U2728 ( .A1(n2431), .A2(n2427), .ZN(n2758) );
  INV_X1 U2729 ( .A(IR_REG_24__SCAN_IN), .ZN(n2762) );
  NAND2_X1 U2730 ( .A1(n2568), .A2(n2209), .ZN(n2623) );
  AND2_X1 U2731 ( .A1(n2608), .A2(n2601), .ZN(n4056) );
  AND2_X1 U2732 ( .A1(n2568), .A2(n2567), .ZN(n2621) );
  AND2_X1 U2733 ( .A1(n2559), .A2(n2577), .ZN(n3256) );
  INV_X1 U2734 ( .A(IR_REG_7__SCAN_IN), .ZN(n2531) );
  NOR2_X1 U2735 ( .A1(n2492), .A2(IR_REG_5__SCAN_IN), .ZN(n2533) );
  INV_X1 U2736 ( .A(IR_REG_3__SCAN_IN), .ZN(n4721) );
  NAND2_X1 U2737 ( .A1(n2194), .A2(n2190), .ZN(n3690) );
  NOR2_X1 U2738 ( .A1(n2191), .A2(n2153), .ZN(n2190) );
  INV_X1 U2739 ( .A(n2193), .ZN(n2191) );
  NAND2_X1 U2740 ( .A1(n3696), .A2(n3645), .ZN(n3699) );
  OR2_X1 U2741 ( .A1(n2447), .A2(n2461), .ZN(n2466) );
  AND2_X1 U2742 ( .A1(n2464), .A2(n2463), .ZN(n2465) );
  AOI21_X1 U2743 ( .B1(n2386), .B2(n2387), .A(n2385), .ZN(n2384) );
  INV_X1 U2744 ( .A(n3785), .ZN(n2385) );
  NAND2_X1 U2745 ( .A1(n2189), .A2(n3673), .ZN(n3681) );
  NAND2_X1 U2746 ( .A1(n2187), .A2(n2186), .ZN(n3592) );
  NAND2_X1 U2747 ( .A1(n3654), .A2(n3757), .ZN(n3727) );
  INV_X1 U2748 ( .A(n2201), .ZN(n3129) );
  OR2_X1 U2749 ( .A1(n3079), .A2(n3078), .ZN(n3080) );
  NAND2_X1 U2750 ( .A1(n2400), .A2(n2397), .ZN(n3776) );
  INV_X1 U2751 ( .A(n2399), .ZN(n2397) );
  NAND2_X1 U2752 ( .A1(n2389), .A2(n3575), .ZN(n3787) );
  NAND2_X1 U2753 ( .A1(n2392), .A2(n2390), .ZN(n2389) );
  NAND2_X1 U2754 ( .A1(n2366), .A2(n2370), .ZN(n3794) );
  INV_X1 U2755 ( .A(n3806), .ZN(n3819) );
  OAI21_X1 U2756 ( .B1(n4134), .B2(n2142), .A(n2696), .ZN(n4308) );
  NAND2_X1 U2757 ( .A1(n2673), .A2(n2672), .ZN(n4162) );
  OAI211_X1 U2758 ( .C1(n4224), .C2(n2142), .A(n2657), .B(n2656), .ZN(n4201)
         );
  OAI211_X1 U2759 ( .C1(n4247), .C2(n2142), .A(n2653), .B(n2652), .ZN(n4341)
         );
  NAND2_X1 U2760 ( .A1(n2645), .A2(n2644), .ZN(n4279) );
  INV_X1 U2761 ( .A(n4374), .ZN(n3994) );
  INV_X1 U2762 ( .A(n4368), .ZN(n3995) );
  NAND4_X1 U2763 ( .A1(n2564), .A2(n2563), .A3(n2562), .A4(n2561), .ZN(n3594)
         );
  INV_X1 U2764 ( .A(n3289), .ZN(n3999) );
  INV_X1 U2765 ( .A(n2964), .ZN(n3711) );
  CLKBUF_X1 U2766 ( .A(n2896), .Z(n2936) );
  AND2_X1 U2767 ( .A1(n2839), .A2(n2838), .ZN(n2853) );
  NAND2_X1 U2768 ( .A1(n2847), .A2(n2846), .ZN(n4020) );
  XNOR2_X1 U2769 ( .A(n4437), .B(n2856), .ZN(n4025) );
  OAI21_X1 U2770 ( .B1(n2928), .B2(n2218), .A(n2217), .ZN(n2216) );
  INV_X1 U2771 ( .A(n2354), .ZN(n2868) );
  NAND2_X1 U2772 ( .A1(n2346), .A2(n4435), .ZN(n2344) );
  XNOR2_X1 U2773 ( .A(n2352), .B(n2349), .ZN(n2884) );
  INV_X1 U2774 ( .A(n2348), .ZN(n2877) );
  NAND2_X1 U2775 ( .A1(n2878), .A2(n4433), .ZN(n2347) );
  XNOR2_X1 U2776 ( .A(n3259), .B(n3258), .ZN(n3260) );
  AND2_X1 U2777 ( .A1(n2226), .A2(n2172), .ZN(n4451) );
  NAND2_X1 U2778 ( .A1(n2226), .A2(n2225), .ZN(n4450) );
  NAND2_X1 U2779 ( .A1(n4458), .A2(n3262), .ZN(n4472) );
  NAND2_X1 U2780 ( .A1(n4472), .A2(n4473), .ZN(n4471) );
  NAND2_X1 U2781 ( .A1(n4479), .A2(n3266), .ZN(n4051) );
  NOR2_X1 U2782 ( .A1(n4501), .A2(n4500), .ZN(n4499) );
  NOR2_X1 U2783 ( .A1(n4516), .A2(n4047), .ZN(n4050) );
  NAND2_X1 U2784 ( .A1(n2320), .A2(n2321), .ZN(n2795) );
  NAND2_X1 U2785 ( .A1(n2743), .A2(n2322), .ZN(n2320) );
  NAND2_X1 U2786 ( .A1(n2283), .A2(n2286), .ZN(n4111) );
  NAND2_X1 U2787 ( .A1(n2290), .A2(n2287), .ZN(n2283) );
  NAND2_X1 U2788 ( .A1(n2442), .A2(n2441), .ZN(n4120) );
  INV_X1 U2789 ( .A(n2689), .ZN(n2288) );
  NAND2_X1 U2790 ( .A1(n2290), .A2(n2690), .ZN(n2289) );
  NAND2_X1 U2791 ( .A1(n2275), .A2(n2277), .ZN(n4156) );
  OR2_X1 U2792 ( .A1(n4211), .A2(n2278), .ZN(n2275) );
  NAND2_X1 U2793 ( .A1(n4337), .A2(n2666), .ZN(n4176) );
  NAND2_X1 U2794 ( .A1(n4274), .A2(n2638), .ZN(n4253) );
  INV_X1 U2795 ( .A(n4364), .ZN(n4265) );
  INV_X1 U2796 ( .A(n2263), .ZN(n3332) );
  AOI21_X1 U2797 ( .B1(n3198), .B2(n2144), .A(n2151), .ZN(n2263) );
  NAND2_X1 U2798 ( .A1(n2269), .A2(n2273), .ZN(n3316) );
  NAND4_X1 U2799 ( .A1(n2543), .A2(n2542), .A3(n2541), .A4(n2540), .ZN(n3997)
         );
  INV_X1 U2800 ( .A(n3925), .ZN(n2306) );
  INV_X1 U2801 ( .A(n3184), .ZN(n2307) );
  AND2_X1 U2802 ( .A1(n2143), .A2(n4362), .ZN(n4222) );
  AND2_X1 U2803 ( .A1(n2143), .A2(n4363), .ZN(n4146) );
  AND3_X1 U2804 ( .A1(n2484), .A2(n2411), .A3(n2483), .ZN(n3115) );
  OR2_X1 U2805 ( .A1(n2447), .A2(n2482), .ZN(n2483) );
  NAND2_X1 U2806 ( .A1(n2249), .A2(n2248), .ZN(n2811) );
  OR2_X1 U2807 ( .A1(n4090), .A2(n4593), .ZN(n2248) );
  INV_X1 U2808 ( .A(n4604), .ZN(n4602) );
  XNOR2_X1 U2809 ( .A(n4301), .B(n2332), .ZN(n4440) );
  INV_X1 U2810 ( .A(n4296), .ZN(n2332) );
  OR2_X1 U2811 ( .A1(n4302), .A2(n4301), .ZN(n4444) );
  NAND2_X1 U2812 ( .A1(n2246), .A2(n2245), .ZN(n2244) );
  INV_X1 U2813 ( .A(n2247), .ZN(n2246) );
  INV_X1 U2814 ( .A(n2243), .ZN(n2242) );
  NAND2_X1 U2815 ( .A1(n2917), .A2(n2825), .ZN(n4549) );
  INV_X1 U2816 ( .A(n2437), .ZN(n2819) );
  INV_X1 U2817 ( .A(n2911), .ZN(n2979) );
  NAND2_X1 U2818 ( .A1(n3032), .A2(STATE_REG_SCAN_IN), .ZN(n4551) );
  XNOR2_X1 U2819 ( .A(n2713), .B(IR_REG_22__SCAN_IN), .ZN(n4429) );
  INV_X1 U2820 ( .A(n4081), .ZN(n4667) );
  INV_X1 U2821 ( .A(n3128), .ZN(n2200) );
  AND2_X1 U2822 ( .A1(n2198), .A2(n2197), .ZN(n2984) );
  INV_X1 U2823 ( .A(n2355), .ZN(n4529) );
  OAI21_X1 U2824 ( .B1(n4520), .B2(n2357), .A(n2356), .ZN(n2355) );
  XNOR2_X1 U2825 ( .A(n2229), .B(n2228), .ZN(n4085) );
  INV_X1 U2826 ( .A(n4073), .ZN(n2228) );
  NAND2_X1 U2827 ( .A1(n2253), .A2(n2251), .ZN(n4086) );
  OR2_X1 U2828 ( .A1(n4095), .A2(n4372), .ZN(n2788) );
  OR2_X1 U2829 ( .A1(n4095), .A2(n4423), .ZN(n2792) );
  AND2_X1 U2830 ( .A1(n2147), .A2(n2268), .ZN(n2144) );
  OR3_X1 U2831 ( .A1(n4285), .A2(n2337), .A3(n2184), .ZN(n2145) );
  AND2_X1 U2832 ( .A1(n2993), .A2(n2459), .ZN(n2146) );
  NAND2_X1 U2833 ( .A1(n2202), .A2(n2175), .ZN(n2400) );
  NOR2_X1 U2834 ( .A1(n2582), .A2(n2581), .ZN(n2147) );
  INV_X1 U2835 ( .A(n3851), .ZN(n2317) );
  NAND2_X1 U2836 ( .A1(n3355), .A2(n2579), .ZN(n2148) );
  AND2_X1 U2837 ( .A1(n2333), .A2(n4373), .ZN(n2149) );
  INV_X1 U2838 ( .A(n4170), .ZN(n2340) );
  AND2_X1 U2839 ( .A1(n3045), .A2(n2962), .ZN(n2150) );
  INV_X1 U2840 ( .A(n2948), .ZN(n2746) );
  AND3_X1 U2841 ( .A1(n2308), .A2(n2141), .A3(n2401), .ZN(n2434) );
  AND2_X1 U2842 ( .A1(n2147), .A2(n2266), .ZN(n2151) );
  OR2_X1 U2843 ( .A1(n3561), .A2(n3560), .ZN(n2152) );
  AND2_X1 U2844 ( .A1(n2308), .A2(n2141), .ZN(n2760) );
  NAND2_X1 U2845 ( .A1(n2708), .A2(n4731), .ZN(n2711) );
  NAND2_X1 U2846 ( .A1(n2367), .A2(n3795), .ZN(n2153) );
  AND2_X1 U2847 ( .A1(n2985), .A2(n3027), .ZN(n2154) );
  NOR2_X1 U2848 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2450)
         );
  INV_X1 U2849 ( .A(n2448), .ZN(n2945) );
  INV_X1 U2850 ( .A(n2448), .ZN(n2798) );
  NAND2_X1 U2851 ( .A1(n2202), .A2(n2203), .ZN(n3716) );
  NAND2_X1 U2852 ( .A1(n2392), .A2(n3570), .ZN(n3746) );
  NAND2_X1 U2853 ( .A1(n2436), .A2(n2437), .ZN(n2447) );
  INV_X1 U2854 ( .A(n3712), .ZN(n2236) );
  AND2_X1 U2855 ( .A1(n4308), .A2(n3802), .ZN(n2155) );
  AND2_X1 U2856 ( .A1(n2197), .A2(n2196), .ZN(n2156) );
  AND2_X1 U2857 ( .A1(n2698), .A2(n4606), .ZN(n2157) );
  NAND2_X1 U2858 ( .A1(n2765), .A2(n4427), .ZN(n2891) );
  AND2_X1 U2859 ( .A1(n3766), .A2(n3767), .ZN(n2158) );
  AND2_X1 U2860 ( .A1(n2345), .A2(n2344), .ZN(n2159) );
  AND2_X1 U2861 ( .A1(n4731), .A2(n2406), .ZN(n2160) );
  NAND2_X1 U2862 ( .A1(n2450), .A2(n2420), .ZN(n2475) );
  INV_X1 U2863 ( .A(n2323), .ZN(n2322) );
  NAND2_X1 U2864 ( .A1(n3842), .A2(n2325), .ZN(n2323) );
  AND2_X1 U2865 ( .A1(n2485), .A2(n2477), .ZN(n4436) );
  INV_X1 U2866 ( .A(IR_REG_25__SCAN_IN), .ZN(n2427) );
  AND2_X1 U2867 ( .A1(n2272), .A2(n2273), .ZN(n2268) );
  INV_X1 U2868 ( .A(n3225), .ZN(n2380) );
  NOR2_X1 U2869 ( .A1(n4151), .A2(n4170), .ZN(n2161) );
  AND2_X1 U2870 ( .A1(n3796), .A2(n2371), .ZN(n2369) );
  NAND2_X1 U2871 ( .A1(n2405), .A2(n2565), .ZN(n2162) );
  INV_X1 U2872 ( .A(IR_REG_26__SCAN_IN), .ZN(n2428) );
  NAND2_X1 U2873 ( .A1(n2380), .A2(n3227), .ZN(n2163) );
  OR2_X1 U2874 ( .A1(n2155), .A2(n2689), .ZN(n2164) );
  INV_X1 U2875 ( .A(n2444), .ZN(n2404) );
  AND2_X1 U2876 ( .A1(n2289), .A2(n2288), .ZN(n2165) );
  AND2_X1 U2877 ( .A1(n2193), .A2(n2192), .ZN(n2166) );
  NAND2_X1 U2878 ( .A1(n2164), .A2(n2291), .ZN(n2286) );
  INV_X1 U2879 ( .A(n4433), .ZN(n2349) );
  INV_X1 U2880 ( .A(IR_REG_0__SCAN_IN), .ZN(n2364) );
  AND2_X1 U2881 ( .A1(n4120), .A2(n4096), .ZN(n2167) );
  OR2_X1 U2882 ( .A1(n4102), .A2(n4117), .ZN(n2168) );
  NAND2_X1 U2883 ( .A1(n3601), .A2(n3394), .ZN(n3487) );
  AND2_X1 U2884 ( .A1(n3257), .A2(REG2_REG_9__SCAN_IN), .ZN(n2169) );
  OR2_X1 U2885 ( .A1(n4279), .A2(n4266), .ZN(n2170) );
  AND2_X1 U2886 ( .A1(n3658), .A2(n3657), .ZN(n2171) );
  INV_X1 U2887 ( .A(n3904), .ZN(n2261) );
  INV_X1 U2888 ( .A(n3501), .ZN(n3418) );
  NAND2_X1 U2889 ( .A1(n3258), .A2(n4533), .ZN(n2172) );
  OR2_X1 U2890 ( .A1(n4285), .A2(n4284), .ZN(n2173) );
  NOR3_X1 U2891 ( .A1(n4207), .A2(n2339), .A3(n3802), .ZN(n2341) );
  INV_X1 U2892 ( .A(n2547), .ZN(n2270) );
  OR2_X1 U2893 ( .A1(n3718), .A2(n3635), .ZN(n2174) );
  INV_X1 U2894 ( .A(n2338), .ZN(n4144) );
  NOR2_X1 U2895 ( .A1(n4207), .A2(n2339), .ZN(n2338) );
  AND2_X1 U2896 ( .A1(n2203), .A2(n2174), .ZN(n2175) );
  AND2_X1 U2897 ( .A1(n3289), .A2(n3288), .ZN(n2176) );
  INV_X1 U2898 ( .A(n2388), .ZN(n2387) );
  NAND2_X1 U2899 ( .A1(n3575), .A2(n2183), .ZN(n2388) );
  AND2_X1 U2900 ( .A1(n3999), .A2(n3536), .ZN(n2177) );
  NOR2_X1 U2901 ( .A1(n4129), .A2(n4307), .ZN(n2178) );
  OR2_X1 U2902 ( .A1(n2252), .A2(n4382), .ZN(n2179) );
  INV_X1 U2903 ( .A(n2666), .ZN(n2280) );
  OR2_X1 U2904 ( .A1(n2396), .A2(n2393), .ZN(n2180) );
  NAND2_X1 U2905 ( .A1(n3650), .A2(n3651), .ZN(n2181) );
  OAI21_X1 U2906 ( .B1(n4210), .B2(n2280), .A(n2674), .ZN(n2279) );
  INV_X1 U2907 ( .A(n3897), .ZN(n2297) );
  NAND2_X1 U2908 ( .A1(n3909), .A2(n3912), .ZN(n2718) );
  AND2_X2 U2909 ( .A1(n3044), .A2(n4531), .ZN(n4661) );
  NOR2_X1 U2910 ( .A1(n3158), .A2(n2412), .ZN(n2182) );
  NAND2_X1 U2911 ( .A1(n2307), .A2(n2306), .ZN(n3183) );
  OAI21_X1 U2912 ( .B1(n3184), .B2(n2304), .A(n2302), .ZN(n3190) );
  NAND2_X1 U2913 ( .A1(n2199), .A2(n2372), .ZN(n3531) );
  OR2_X1 U2914 ( .A1(n3582), .A2(n3581), .ZN(n2183) );
  OR2_X1 U2915 ( .A1(n4266), .A2(n4340), .ZN(n2184) );
  OAI21_X1 U2916 ( .B1(n3198), .B2(n2151), .A(n2264), .ZN(n3330) );
  INV_X1 U2917 ( .A(n2336), .ZN(n4349) );
  NOR3_X1 U2918 ( .A1(n4285), .A2(n2337), .A3(n4266), .ZN(n2336) );
  NAND2_X1 U2919 ( .A1(n3419), .A2(n2333), .ZN(n2335) );
  INV_X1 U2920 ( .A(n3738), .ZN(n4373) );
  AND2_X1 U2921 ( .A1(n3959), .A2(n3955), .ZN(n3873) );
  INV_X1 U2922 ( .A(n4189), .ZN(n3701) );
  INV_X1 U2923 ( .A(n2969), .ZN(n2965) );
  AND2_X2 U2924 ( .A1(n2790), .A2(n3043), .ZN(n4600) );
  INV_X1 U2925 ( .A(n2719), .ZN(n3880) );
  AND2_X1 U2926 ( .A1(n2853), .A2(n3987), .ZN(n4480) );
  NAND2_X1 U2927 ( .A1(n4241), .A2(n4353), .ZN(n4593) );
  INV_X1 U2928 ( .A(n2331), .ZN(n3176) );
  NOR2_X1 U2929 ( .A1(n3142), .A2(n3163), .ZN(n2331) );
  NAND2_X1 U2930 ( .A1(n2929), .A2(REG1_REG_4__SCAN_IN), .ZN(n2345) );
  OAI21_X1 U2931 ( .B1(n2895), .B2(n2967), .A(n2894), .ZN(n2899) );
  INV_X1 U2932 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2213) );
  INV_X1 U2933 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2214) );
  XNOR2_X1 U2934 ( .A(n2432), .B(IR_REG_30__SCAN_IN), .ZN(n2822) );
  OR2_X1 U2935 ( .A1(n4554), .A2(n4077), .ZN(n2185) );
  OAI21_X1 U2936 ( .B1(n3592), .B2(n3590), .A(n3588), .ZN(n3550) );
  NAND2_X1 U2937 ( .A1(n3487), .A2(n3486), .ZN(n2186) );
  OAI21_X1 U2938 ( .B1(n3487), .B2(n3486), .A(n3485), .ZN(n2187) );
  INV_X1 U2939 ( .A(n4375), .ZN(n4584) );
  INV_X2 U2940 ( .A(n2967), .ZN(n3670) );
  NAND2_X2 U2941 ( .A1(n4375), .A2(n3027), .ZN(n2967) );
  NAND2_X4 U2942 ( .A1(n3045), .A2(n2891), .ZN(n3675) );
  OR2_X2 U2943 ( .A1(n3653), .A2(n2195), .ZN(n2194) );
  NAND2_X1 U2944 ( .A1(n3654), .A2(n2188), .ZN(n2193) );
  NAND2_X1 U2945 ( .A1(n3653), .A2(n3652), .ZN(n3757) );
  NAND2_X1 U2946 ( .A1(n2166), .A2(n2194), .ZN(n2189) );
  OR2_X1 U2947 ( .A1(n2978), .A2(n2977), .ZN(n2197) );
  AND2_X2 U2948 ( .A1(n2201), .A2(n2200), .ZN(n3158) );
  OR2_X2 U2949 ( .A1(n3125), .A2(n2407), .ZN(n2201) );
  OR2_X2 U2950 ( .A1(n3619), .A2(n2206), .ZN(n2202) );
  NAND2_X1 U2951 ( .A1(n2568), .A2(n2207), .ZN(n2646) );
  INV_X1 U2952 ( .A(n2216), .ZN(n2870) );
  NAND2_X1 U2953 ( .A1(n2852), .A2(n4435), .ZN(n2217) );
  INV_X1 U2954 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2218) );
  INV_X1 U2955 ( .A(n2850), .ZN(n2220) );
  NAND4_X1 U2956 ( .A1(n2234), .A2(n2233), .A3(n2232), .A4(n2231), .ZN(n2422)
         );
  NAND4_X1 U2957 ( .A1(n2239), .A2(n2240), .A3(n2238), .A4(n2452), .ZN(n2969)
         );
  NAND3_X1 U2958 ( .A1(n2241), .A2(n2240), .A3(n2235), .ZN(n3912) );
  NAND2_X1 U2959 ( .A1(n2469), .A2(REG0_REG_1__SCAN_IN), .ZN(n2238) );
  OAI21_X1 U2960 ( .B1(n2794), .B2(n2254), .A(n2242), .ZN(n2245) );
  NAND2_X1 U2961 ( .A1(n2244), .A2(n2259), .ZN(n2814) );
  NAND3_X1 U2962 ( .A1(n2253), .A2(n2251), .A3(n2260), .ZN(n2249) );
  NAND2_X1 U2963 ( .A1(n4598), .A2(n2812), .ZN(n2259) );
  INV_X1 U2964 ( .A(n4090), .ZN(n2260) );
  OR2_X1 U2965 ( .A1(n3372), .A2(n3605), .ZN(n2273) );
  NAND2_X1 U2966 ( .A1(n4211), .A2(n2277), .ZN(n2274) );
  NAND2_X1 U2967 ( .A1(n2274), .A2(n2276), .ZN(n2682) );
  INV_X1 U2968 ( .A(n4142), .ZN(n2290) );
  NAND2_X1 U2969 ( .A1(n4142), .A2(n2286), .ZN(n2282) );
  AOI21_X1 U2970 ( .B1(n4275), .B2(n2296), .A(n2293), .ZN(n2292) );
  AND2_X1 U2971 ( .A1(n2141), .A2(n2565), .ZN(n2757) );
  NOR2_X1 U2972 ( .A1(n4054), .A2(n4490), .ZN(n4501) );
  NAND2_X1 U2973 ( .A1(n2431), .A2(n2363), .ZN(n2362) );
  AOI21_X1 U2974 ( .B1(n3345), .B2(n2602), .A(n2408), .ZN(n3463) );
  NAND2_X1 U2975 ( .A1(n3330), .A2(n2591), .ZN(n3345) );
  NAND2_X1 U2976 ( .A1(n2471), .A2(n2470), .ZN(n2472) );
  NAND2_X1 U2977 ( .A1(n3464), .A2(n2611), .ZN(n3477) );
  NAND2_X1 U2978 ( .A1(n3367), .A2(n2313), .ZN(n2309) );
  NAND2_X1 U2979 ( .A1(n2309), .A2(n2310), .ZN(n3342) );
  OAI21_X1 U2980 ( .B1(n2743), .B2(n2318), .A(n2316), .ZN(n2796) );
  AOI21_X1 U2981 ( .B1(n2743), .B2(n2325), .A(n3850), .ZN(n4108) );
  INV_X1 U2982 ( .A(n3850), .ZN(n2326) );
  NAND2_X1 U2983 ( .A1(n2757), .A2(n2329), .ZN(n2328) );
  NAND2_X1 U2984 ( .A1(n2328), .A2(IR_REG_31__SCAN_IN), .ZN(n2433) );
  OR2_X1 U2985 ( .A1(n2718), .A2(n3908), .ZN(n2999) );
  INV_X1 U2986 ( .A(n2335), .ZN(n3467) );
  NAND3_X1 U2987 ( .A1(n4170), .A2(n4145), .A3(n4189), .ZN(n2339) );
  INV_X1 U2988 ( .A(n2341), .ZN(n4132) );
  NAND3_X1 U2989 ( .A1(n3056), .A2(n3007), .A3(n3065), .ZN(n4583) );
  NAND2_X1 U2990 ( .A1(n2342), .A2(n3092), .ZN(n3071) );
  AND2_X1 U2991 ( .A1(n3008), .A2(n2342), .ZN(n4567) );
  MUX2_X1 U2992 ( .A(n2845), .B(REG2_REG_1__SCAN_IN), .S(n4006), .Z(n2847) );
  NAND4_X1 U2994 ( .A1(n2365), .A2(n2421), .A3(n2420), .A4(n2364), .ZN(n2492)
         );
  NAND3_X1 U2995 ( .A1(n3654), .A2(n3757), .A3(n2371), .ZN(n2366) );
  NAND2_X1 U2996 ( .A1(n2381), .A2(n2384), .ZN(n3614) );
  NAND3_X1 U2997 ( .A1(n3565), .A2(n2382), .A3(n2152), .ZN(n2381) );
  NAND3_X1 U2998 ( .A1(n3565), .A2(n2152), .A3(n3737), .ZN(n2392) );
  NAND2_X1 U2999 ( .A1(n2400), .A2(n2398), .ZN(n3696) );
  AND2_X1 U3000 ( .A1(n2565), .A2(n2426), .ZN(n2708) );
  OAI21_X2 U3001 ( .B1(n3102), .B2(n3100), .A(n3934), .ZN(n3138) );
  OR2_X1 U3002 ( .A1(n2142), .A2(n2460), .ZN(n2467) );
  OR2_X1 U3003 ( .A1(n2142), .A2(n2453), .ZN(n2457) );
  CLKBUF_X1 U3004 ( .A(n3550), .Z(n3510) );
  INV_X1 U3005 ( .A(n4372), .ZN(n3310) );
  AND2_X1 U3006 ( .A1(n3124), .A2(n3123), .ZN(n2407) );
  AND2_X1 U3007 ( .A1(n3558), .A2(n3557), .ZN(n2408) );
  AND2_X1 U3008 ( .A1(n4607), .A2(n2762), .ZN(n2409) );
  INV_X1 U3009 ( .A(n4205), .ZN(n3638) );
  AND2_X1 U3010 ( .A1(n2636), .A2(DATAI_22_), .ZN(n4205) );
  AND2_X1 U3011 ( .A1(n2665), .A2(n2664), .ZN(n4344) );
  AND2_X1 U3012 ( .A1(n2481), .A2(n2480), .ZN(n2411) );
  AND2_X1 U3013 ( .A1(n3157), .A2(n3156), .ZN(n2412) );
  AND2_X1 U3014 ( .A1(n3555), .A2(n3554), .ZN(n2413) );
  OR2_X1 U3015 ( .A1(n3594), .A2(n3501), .ZN(n2414) );
  OAI21_X1 U3016 ( .B1(n3551), .B2(n3552), .A(n3553), .ZN(n3548) );
  NAND2_X1 U3017 ( .A1(n3617), .A2(n3616), .ZN(n3618) );
  OR2_X1 U3018 ( .A1(n4255), .A2(n2732), .ZN(n3958) );
  AND2_X1 U3019 ( .A1(n3712), .A2(n3514), .ZN(n2968) );
  INV_X1 U3020 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U3021 ( .A1(n2437), .A2(n2822), .ZN(n2448) );
  NOR2_X1 U3022 ( .A1(n2584), .A2(n2583), .ZN(n2592) );
  NAND2_X1 U3023 ( .A1(n3115), .A2(n4582), .ZN(n3919) );
  INV_X1 U3024 ( .A(IR_REG_31__SCAN_IN), .ZN(n2431) );
  NAND2_X1 U3025 ( .A1(n2802), .A2(n2444), .ZN(n2445) );
  NAND2_X1 U3026 ( .A1(n2499), .A2(REG3_REG_6__SCAN_IN), .ZN(n2507) );
  AND2_X1 U3027 ( .A1(n2683), .A2(REG3_REG_25__SCAN_IN), .ZN(n2691) );
  OR2_X1 U3028 ( .A1(n2629), .A2(n2628), .ZN(n2640) );
  INV_X1 U3029 ( .A(IR_REG_13__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U3030 ( .A1(n3993), .A2(n4205), .ZN(n2666) );
  NOR2_X1 U3031 ( .A1(n2640), .A2(n2639), .ZN(n2650) );
  OR2_X1 U3032 ( .A1(n2524), .A2(n4865), .ZN(n2538) );
  INV_X1 U3033 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4623) );
  INV_X1 U3034 ( .A(n4245), .ZN(n2787) );
  AND2_X1 U3035 ( .A1(n4431), .A2(n2937), .ZN(n4362) );
  AND2_X1 U3036 ( .A1(n2533), .A2(n2532), .ZN(n2545) );
  AND2_X1 U3037 ( .A1(n2691), .A2(REG3_REG_26__SCAN_IN), .ZN(n2697) );
  OR2_X1 U3038 ( .A1(n2667), .A2(n3702), .ZN(n2675) );
  OR2_X1 U3039 ( .A1(n2538), .A2(n2537), .ZN(n2549) );
  OR2_X1 U3040 ( .A1(n3672), .A2(n3671), .ZN(n3673) );
  OAI21_X1 U3041 ( .B1(n3531), .B2(n3533), .A(n3532), .ZN(n3385) );
  AND2_X1 U3042 ( .A1(n3659), .A2(n2909), .ZN(n3988) );
  OR2_X1 U3043 ( .A1(n2697), .A2(n2692), .ZN(n4134) );
  INV_X1 U3044 ( .A(n4436), .ZN(n2858) );
  INV_X1 U3045 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4865) );
  INV_X1 U3046 ( .A(n4120), .ZN(n4311) );
  OR2_X1 U3047 ( .A1(n4097), .A2(n2142), .ZN(n2442) );
  INV_X1 U3048 ( .A(n4162), .ZN(n4204) );
  INV_X1 U3049 ( .A(n3873), .ZN(n2610) );
  OR2_X1 U3050 ( .A1(n4289), .A2(n4375), .ZN(n4443) );
  AND2_X1 U3051 ( .A1(n2783), .A2(n2828), .ZN(n2784) );
  INV_X1 U3052 ( .A(n4221), .ZN(n4340) );
  NAND2_X1 U3053 ( .A1(n2979), .A2(n2905), .ZN(n4367) );
  INV_X1 U3054 ( .A(n4363), .ZN(n4573) );
  INV_X1 U3055 ( .A(n4117), .ZN(n4307) );
  INV_X1 U3056 ( .A(n3288), .ZN(n3536) );
  XOR2_X1 U3057 ( .A(n3567), .B(n3566), .Z(n3737) );
  OAI21_X1 U3058 ( .B1(n2156), .B2(n3081), .A(n3080), .ZN(n3082) );
  NAND2_X1 U3059 ( .A1(n2703), .A2(n2702), .ZN(n4129) );
  AND2_X1 U3060 ( .A1(n2617), .A2(n2616), .ZN(n4374) );
  INV_X1 U3061 ( .A(n4574), .ZN(n3164) );
  XNOR2_X1 U3062 ( .A(n2717), .B(IR_REG_28__SCAN_IN), .ZN(n2911) );
  INV_X1 U3063 ( .A(n4150), .ZN(n4223) );
  INV_X1 U3064 ( .A(n4443), .ZN(n4536) );
  AOI21_X1 U3065 ( .B1(n2785), .B2(n2831), .A(n2784), .ZN(n2902) );
  OR2_X1 U3066 ( .A1(n4542), .A2(n4429), .ZN(n4353) );
  NAND2_X1 U3067 ( .A1(n2771), .A2(n4427), .ZN(n2825) );
  INV_X1 U3068 ( .A(n2834), .ZN(n2917) );
  AND2_X1 U3069 ( .A1(n2835), .A2(n2839), .ZN(n4523) );
  OR2_X1 U3070 ( .A1(n2916), .A2(n2908), .ZN(n3806) );
  OAI21_X1 U3071 ( .B1(n3761), .B2(n2142), .A(n2680), .ZN(n4320) );
  INV_X1 U3072 ( .A(n4344), .ZN(n3993) );
  NAND4_X1 U3073 ( .A1(n2597), .A2(n2596), .A3(n2595), .A4(n2594), .ZN(n4379)
         );
  OR2_X1 U3074 ( .A1(n2891), .A2(n4551), .ZN(n4002) );
  INV_X1 U3075 ( .A(n4480), .ZN(n4519) );
  INV_X1 U3076 ( .A(n4220), .ZN(n4293) );
  OR2_X1 U3077 ( .A1(n4088), .A2(n4372), .ZN(n2809) );
  NAND2_X1 U3078 ( .A1(n4604), .A2(n4584), .ZN(n4372) );
  AND2_X2 U3079 ( .A1(n2790), .A2(n2902), .ZN(n4604) );
  NAND2_X1 U3080 ( .A1(n4600), .A2(n4584), .ZN(n4423) );
  INV_X1 U3081 ( .A(n4600), .ZN(n4598) );
  INV_X1 U3082 ( .A(n4549), .ZN(n4550) );
  AND2_X1 U3083 ( .A1(n2521), .A2(n2515), .ZN(n4432) );
  INV_X1 U3084 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2786) );
  NAND2_X1 U3085 ( .A1(n2517), .A2(REG3_REG_8__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U3086 ( .A1(n2570), .A2(REG3_REG_12__SCAN_IN), .ZN(n2571) );
  AND2_X1 U3087 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2415) );
  INV_X1 U3088 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2628) );
  INV_X1 U3089 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2639) );
  INV_X1 U3090 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4868) );
  INV_X1 U3091 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3702) );
  INV_X1 U3092 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4702) );
  AND2_X1 U3093 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2416) );
  NAND2_X1 U3094 ( .A1(n2697), .A2(n2416), .ZN(n4087) );
  INV_X1 U3095 ( .A(n2697), .ZN(n2418) );
  INV_X1 U3096 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4704) );
  INV_X1 U3097 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2417) );
  OAI21_X1 U3098 ( .B1(n2418), .B2(n4704), .A(n2417), .ZN(n2419) );
  NAND2_X1 U3099 ( .A1(n4087), .A2(n2419), .ZN(n4097) );
  NOR2_X2 U3100 ( .A1(n2492), .A2(n2422), .ZN(n2565) );
  NAND2_X1 U3101 ( .A1(n2430), .A2(n2429), .ZN(n2444) );
  INV_X1 U3102 ( .A(n2434), .ZN(n3689) );
  INV_X1 U3103 ( .A(n2822), .ZN(n2436) );
  INV_X1 U3104 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4780) );
  NAND2_X1 U3105 ( .A1(n2944), .A2(REG1_REG_28__SCAN_IN), .ZN(n2439) );
  NAND2_X1 U3106 ( .A1(n2798), .A2(REG2_REG_28__SCAN_IN), .ZN(n2438) );
  OAI211_X1 U3107 ( .C1(n2948), .C2(n4780), .A(n2439), .B(n2438), .ZN(n2440)
         );
  INV_X1 U3108 ( .A(n2440), .ZN(n2441) );
  NAND2_X1 U3109 ( .A1(n2636), .A2(DATAI_28_), .ZN(n3674) );
  INV_X1 U3110 ( .A(n3674), .ZN(n4096) );
  NAND2_X1 U3111 ( .A1(n4311), .A2(n4096), .ZN(n3851) );
  NAND2_X1 U3112 ( .A1(n4120), .A2(n3674), .ZN(n3848) );
  NAND2_X1 U3113 ( .A1(n3851), .A2(n3848), .ZN(n3860) );
  INV_X1 U3114 ( .A(n2447), .ZN(n2469) );
  NAND2_X1 U3115 ( .A1(n2945), .A2(REG2_REG_1__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U3116 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2449)
         );
  INV_X1 U3117 ( .A(n2450), .ZN(n2451) );
  INV_X1 U3118 ( .A(n4006), .ZN(n4438) );
  MUX2_X1 U3119 ( .A(n4438), .B(DATAI_1_), .S(n2458), .Z(n3712) );
  INV_X1 U3120 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U3121 ( .A1(n2798), .A2(REG2_REG_0__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U3122 ( .A1(n2469), .A2(REG0_REG_0__SCAN_IN), .ZN(n2455) );
  MUX2_X1 U3123 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2458), .Z(n2985) );
  NAND2_X1 U3124 ( .A1(n2718), .A2(n2991), .ZN(n2993) );
  NAND2_X1 U3125 ( .A1(n2969), .A2(n3712), .ZN(n2459) );
  INV_X1 U3126 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2460) );
  INV_X1 U3127 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U3128 ( .A1(n2462), .A2(REG1_REG_2__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U3129 ( .A1(n2945), .A2(REG2_REG_2__SCAN_IN), .ZN(n2463) );
  MUX2_X1 U3130 ( .A(n4437), .B(DATAI_2_), .S(n2636), .Z(n2981) );
  NAND2_X1 U3131 ( .A1(n3711), .A2(n3056), .ZN(n3916) );
  NAND2_X1 U3132 ( .A1(n3916), .A2(n3913), .ZN(n2719) );
  NAND2_X1 U3133 ( .A1(n2964), .A2(n3056), .ZN(n3062) );
  INV_X1 U3134 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U3135 ( .A1(n2945), .A2(REG2_REG_3__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U3136 ( .A1(n2469), .A2(REG0_REG_3__SCAN_IN), .ZN(n2470) );
  NOR2_X1 U3137 ( .A1(n2157), .A2(n2472), .ZN(n2474) );
  NAND2_X1 U3138 ( .A1(n2944), .A2(REG1_REG_3__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3139 ( .A1(n2475), .A2(IR_REG_31__SCAN_IN), .ZN(n2476) );
  NAND2_X1 U3140 ( .A1(n2476), .A2(n4721), .ZN(n2485) );
  OR2_X1 U3141 ( .A1(n2476), .A2(n4721), .ZN(n2477) );
  MUX2_X1 U3142 ( .A(n4436), .B(DATAI_3_), .S(n2636), .Z(n3092) );
  INV_X1 U3143 ( .A(n3092), .ZN(n3065) );
  NAND2_X1 U3144 ( .A1(n3055), .A2(n3065), .ZN(n2478) );
  NAND2_X1 U3145 ( .A1(n4580), .A2(n3092), .ZN(n4588) );
  NAND2_X1 U3146 ( .A1(n2944), .A2(REG1_REG_4__SCAN_IN), .ZN(n2484) );
  INV_X1 U3147 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2479) );
  XNOR2_X1 U31480 ( .A(n2479), .B(REG3_REG_3__SCAN_IN), .ZN(n4662) );
  NAND2_X1 U31490 ( .A1(n2698), .A2(n4662), .ZN(n2481) );
  NAND2_X1 U3150 ( .A1(n2945), .A2(REG2_REG_4__SCAN_IN), .ZN(n2480) );
  INV_X1 U3151 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2482) );
  NAND2_X1 U3152 ( .A1(n2485), .A2(IR_REG_31__SCAN_IN), .ZN(n2486) );
  XNOR2_X1 U3153 ( .A(n2486), .B(IR_REG_4__SCAN_IN), .ZN(n4435) );
  MUX2_X1 U3154 ( .A(n4435), .B(DATAI_4_), .S(n2636), .Z(n4582) );
  NAND2_X1 U3155 ( .A1(n4001), .A2(n4582), .ZN(n2488) );
  AND2_X1 U3156 ( .A1(n4588), .A2(n2488), .ZN(n2487) );
  INV_X1 U3157 ( .A(n4582), .ZN(n4572) );
  AOI22_X1 U3158 ( .A1(n2746), .A2(REG0_REG_5__SCAN_IN), .B1(n2944), .B2(
        REG1_REG_5__SCAN_IN), .ZN(n2491) );
  AOI21_X1 U3159 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2489) );
  NOR2_X1 U3160 ( .A1(n2489), .A2(n2499), .ZN(n3104) );
  AOI22_X1 U3161 ( .A1(n2698), .A2(n3104), .B1(n2798), .B2(REG2_REG_5__SCAN_IN), .ZN(n2490) );
  INV_X1 U3162 ( .A(n2533), .ZN(n2495) );
  NAND2_X1 U3163 ( .A1(n2492), .A2(IR_REG_31__SCAN_IN), .ZN(n2493) );
  MUX2_X1 U3164 ( .A(IR_REG_31__SCAN_IN), .B(n2493), .S(IR_REG_5__SCAN_IN), 
        .Z(n2494) );
  NAND2_X1 U3165 ( .A1(n2495), .A2(n2494), .ZN(n2872) );
  INV_X1 U3166 ( .A(DATAI_5_), .ZN(n4696) );
  MUX2_X1 U3167 ( .A(n2872), .B(n4696), .S(n2636), .Z(n3127) );
  NAND2_X1 U3168 ( .A1(n4574), .A2(n3127), .ZN(n2496) );
  NAND2_X1 U3169 ( .A1(n3101), .A2(n2496), .ZN(n2498) );
  INV_X1 U3170 ( .A(n3127), .ZN(n3130) );
  NAND2_X1 U3171 ( .A1(n3164), .A2(n3130), .ZN(n2497) );
  NAND2_X1 U3172 ( .A1(n2746), .A2(REG0_REG_6__SCAN_IN), .ZN(n2504) );
  OAI21_X1 U3173 ( .B1(n2499), .B2(REG3_REG_6__SCAN_IN), .A(n2507), .ZN(n3167)
         );
  INV_X1 U3174 ( .A(n3167), .ZN(n2500) );
  NAND2_X1 U3175 ( .A1(n2698), .A2(n2500), .ZN(n2503) );
  NAND2_X1 U3176 ( .A1(n2944), .A2(REG1_REG_6__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U3177 ( .A1(n2945), .A2(REG2_REG_6__SCAN_IN), .ZN(n2501) );
  NAND4_X1 U3178 ( .A1(n2504), .A2(n2503), .A3(n2502), .A4(n2501), .ZN(n4000)
         );
  OR2_X1 U3179 ( .A1(n2533), .A2(n2431), .ZN(n2505) );
  XNOR2_X1 U3180 ( .A(n2505), .B(IR_REG_6__SCAN_IN), .ZN(n4433) );
  MUX2_X1 U3181 ( .A(n4433), .B(DATAI_6_), .S(n2636), .Z(n3163) );
  AND2_X1 U3182 ( .A1(n4000), .A2(n3163), .ZN(n2506) );
  NAND2_X1 U3183 ( .A1(n2746), .A2(REG0_REG_7__SCAN_IN), .ZN(n2512) );
  AND2_X1 U3184 ( .A1(n2507), .A2(n2880), .ZN(n2508) );
  NOR2_X1 U3185 ( .A1(n2517), .A2(n2508), .ZN(n3178) );
  NAND2_X1 U3186 ( .A1(n2698), .A2(n3178), .ZN(n2511) );
  NAND2_X1 U3187 ( .A1(n2944), .A2(REG1_REG_7__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U3188 ( .A1(n2945), .A2(REG2_REG_7__SCAN_IN), .ZN(n2509) );
  NAND4_X1 U3189 ( .A1(n2512), .A2(n2511), .A3(n2510), .A4(n2509), .ZN(n3537)
         );
  INV_X1 U3190 ( .A(n3537), .ZN(n3230) );
  NAND2_X1 U3191 ( .A1(n2533), .A2(n4720), .ZN(n2513) );
  NAND2_X1 U3192 ( .A1(n2513), .A2(IR_REG_31__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U3193 ( .A1(n2514), .A2(n2531), .ZN(n2521) );
  OR2_X1 U3194 ( .A1(n2514), .A2(n2531), .ZN(n2515) );
  MUX2_X1 U3195 ( .A(n4432), .B(DATAI_7_), .S(n2636), .Z(n3232) );
  NAND2_X1 U3196 ( .A1(n3230), .A2(n3232), .ZN(n2722) );
  INV_X1 U3197 ( .A(n3232), .ZN(n3229) );
  NAND2_X1 U3198 ( .A1(n3537), .A2(n3229), .ZN(n3928) );
  NAND2_X1 U3199 ( .A1(n3537), .A2(n3232), .ZN(n2516) );
  AOI22_X1 U3200 ( .A1(n2746), .A2(REG0_REG_8__SCAN_IN), .B1(n2944), .B2(
        REG1_REG_8__SCAN_IN), .ZN(n2520) );
  OR2_X1 U3201 ( .A1(n2517), .A2(REG3_REG_8__SCAN_IN), .ZN(n2518) );
  AND2_X1 U3202 ( .A1(n2524), .A2(n2518), .ZN(n3538) );
  AOI22_X1 U3203 ( .A1(n2698), .A2(n3538), .B1(n2798), .B2(REG2_REG_8__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U3204 ( .A1(n2521), .A2(IR_REG_31__SCAN_IN), .ZN(n2522) );
  XNOR2_X1 U3205 ( .A(n2522), .B(n4713), .ZN(n3258) );
  INV_X1 U3206 ( .A(DATAI_8_), .ZN(n2523) );
  MUX2_X1 U3207 ( .A(n3258), .B(n2523), .S(n2636), .Z(n3288) );
  NAND2_X1 U3208 ( .A1(n2746), .A2(REG0_REG_9__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U3209 ( .A1(n2524), .A2(n4865), .ZN(n2525) );
  NAND2_X1 U32100 ( .A1(n2538), .A2(n2525), .ZN(n3299) );
  INV_X1 U32110 ( .A(n3299), .ZN(n2526) );
  NAND2_X1 U32120 ( .A1(n2698), .A2(n2526), .ZN(n2529) );
  NAND2_X1 U32130 ( .A1(n2944), .A2(REG1_REG_9__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U32140 ( .A1(n2945), .A2(REG2_REG_9__SCAN_IN), .ZN(n2527) );
  NAND4_X1 U32150 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .ZN(n3998)
         );
  OR2_X1 U32160 ( .A1(n2545), .A2(n2431), .ZN(n2534) );
  XNOR2_X1 U32170 ( .A(n2534), .B(IR_REG_9__SCAN_IN), .ZN(n3257) );
  MUX2_X1 U32180 ( .A(n3257), .B(DATAI_9_), .S(n2636), .Z(n3296) );
  AND2_X1 U32190 ( .A1(n3998), .A2(n3296), .ZN(n2536) );
  NAND2_X1 U32200 ( .A1(n3607), .A2(n3292), .ZN(n2535) );
  NAND2_X1 U32210 ( .A1(n2746), .A2(REG0_REG_10__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U32220 ( .A1(n2538), .A2(n2537), .ZN(n2539) );
  AND2_X1 U32230 ( .A1(n2549), .A2(n2539), .ZN(n3610) );
  NAND2_X1 U32240 ( .A1(n2698), .A2(n3610), .ZN(n2542) );
  NAND2_X1 U32250 ( .A1(n2944), .A2(REG1_REG_10__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32260 ( .A1(n2798), .A2(REG2_REG_10__SCAN_IN), .ZN(n2540) );
  INV_X1 U32270 ( .A(IR_REG_9__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U32280 ( .A1(n2545), .A2(n2544), .ZN(n2555) );
  NAND2_X1 U32290 ( .A1(n2555), .A2(IR_REG_31__SCAN_IN), .ZN(n2546) );
  XNOR2_X1 U32300 ( .A(n2546), .B(IR_REG_10__SCAN_IN), .ZN(n4561) );
  MUX2_X1 U32310 ( .A(n4561), .B(DATAI_10_), .S(n2636), .Z(n3389) );
  NOR2_X1 U32320 ( .A1(n3997), .A2(n3389), .ZN(n2547) );
  INV_X1 U32330 ( .A(n3389), .ZN(n3605) );
  NAND2_X1 U32340 ( .A1(n2746), .A2(REG0_REG_11__SCAN_IN), .ZN(n2554) );
  AND2_X1 U32350 ( .A1(n2549), .A2(n2548), .ZN(n2550) );
  NOR2_X1 U32360 ( .A1(n2570), .A2(n2550), .ZN(n3320) );
  NAND2_X1 U32370 ( .A1(n2698), .A2(n3320), .ZN(n2553) );
  NAND2_X1 U32380 ( .A1(n2944), .A2(REG1_REG_11__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32390 ( .A1(n2798), .A2(REG2_REG_11__SCAN_IN), .ZN(n2551) );
  NAND4_X1 U32400 ( .A1(n2554), .A2(n2553), .A3(n2552), .A4(n2551), .ZN(n3996)
         );
  NAND2_X1 U32410 ( .A1(n2556), .A2(IR_REG_31__SCAN_IN), .ZN(n2558) );
  INV_X1 U32420 ( .A(IR_REG_11__SCAN_IN), .ZN(n2557) );
  OR2_X1 U32430 ( .A1(n2558), .A2(n2557), .ZN(n2559) );
  NAND2_X1 U32440 ( .A1(n2558), .A2(n2557), .ZN(n2577) );
  MUX2_X1 U32450 ( .A(n3256), .B(DATAI_11_), .S(n2636), .Z(n3398) );
  NAND2_X1 U32460 ( .A1(n3437), .A2(n3398), .ZN(n3364) );
  INV_X1 U32470 ( .A(n3398), .ZN(n3396) );
  NAND2_X1 U32480 ( .A1(n3996), .A2(n3396), .ZN(n3366) );
  NAND2_X1 U32490 ( .A1(n3437), .A2(n3396), .ZN(n3355) );
  NAND2_X1 U32500 ( .A1(n2746), .A2(REG0_REG_13__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U32510 ( .A1(n2571), .A2(n4623), .ZN(n2560) );
  AND2_X1 U32520 ( .A1(n2584), .A2(n2560), .ZN(n3500) );
  NAND2_X1 U32530 ( .A1(n2698), .A2(n3500), .ZN(n2563) );
  NAND2_X1 U32540 ( .A1(n2944), .A2(REG1_REG_13__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32550 ( .A1(n2798), .A2(REG2_REG_13__SCAN_IN), .ZN(n2561) );
  BUF_X1 U32560 ( .A(n2565), .Z(n2568) );
  NOR2_X1 U32570 ( .A1(n2568), .A2(n2431), .ZN(n2566) );
  MUX2_X1 U32580 ( .A(n2431), .B(n2566), .S(IR_REG_13__SCAN_IN), .Z(n2569) );
  OR2_X1 U32590 ( .A1(n2569), .A2(n2621), .ZN(n3255) );
  INV_X1 U32600 ( .A(n3255), .ZN(n4052) );
  MUX2_X1 U32610 ( .A(n4052), .B(DATAI_13_), .S(n2636), .Z(n3501) );
  NAND2_X1 U32620 ( .A1(n2746), .A2(REG0_REG_12__SCAN_IN), .ZN(n2576) );
  OR2_X1 U32630 ( .A1(n2570), .A2(REG3_REG_12__SCAN_IN), .ZN(n2572) );
  AND2_X1 U32640 ( .A1(n2572), .A2(n2571), .ZN(n3360) );
  NAND2_X1 U32650 ( .A1(n2698), .A2(n3360), .ZN(n2575) );
  NAND2_X1 U32660 ( .A1(n2944), .A2(REG1_REG_12__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U32670 ( .A1(n2945), .A2(REG2_REG_12__SCAN_IN), .ZN(n2573) );
  NAND4_X1 U32680 ( .A1(n2576), .A2(n2575), .A3(n2574), .A4(n2573), .ZN(n3502)
         );
  INV_X1 U32690 ( .A(n3502), .ZN(n2728) );
  NAND2_X1 U32700 ( .A1(n2577), .A2(IR_REG_31__SCAN_IN), .ZN(n2578) );
  XNOR2_X1 U32710 ( .A(n2578), .B(IR_REG_12__SCAN_IN), .ZN(n3264) );
  MUX2_X1 U32720 ( .A(n3264), .B(DATAI_12_), .S(n2636), .Z(n3593) );
  NAND2_X1 U32730 ( .A1(n2728), .A2(n3357), .ZN(n3407) );
  AND2_X1 U32740 ( .A1(n2414), .A2(n3407), .ZN(n2579) );
  INV_X1 U32750 ( .A(n2579), .ZN(n2580) );
  NAND2_X1 U32760 ( .A1(n3502), .A2(n3593), .ZN(n3405) );
  NOR2_X1 U32770 ( .A1(n2580), .A2(n3405), .ZN(n2582) );
  AND2_X1 U32780 ( .A1(n3594), .A2(n3501), .ZN(n2581) );
  AND2_X1 U32790 ( .A1(n2584), .A2(n2583), .ZN(n2585) );
  NOR2_X1 U32800 ( .A1(n2592), .A2(n2585), .ZN(n3524) );
  NAND2_X1 U32810 ( .A1(n2698), .A2(n3524), .ZN(n2589) );
  NAND2_X1 U32820 ( .A1(n2944), .A2(REG1_REG_14__SCAN_IN), .ZN(n2588) );
  INV_X1 U32830 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4774) );
  OR2_X1 U32840 ( .A1(n2948), .A2(n4774), .ZN(n2587) );
  NAND2_X1 U32850 ( .A1(n2798), .A2(REG2_REG_14__SCAN_IN), .ZN(n2586) );
  OR2_X1 U32860 ( .A1(n2621), .A2(n2431), .ZN(n2590) );
  XNOR2_X1 U32870 ( .A(n2590), .B(IR_REG_14__SCAN_IN), .ZN(n4557) );
  MUX2_X1 U32880 ( .A(n4557), .B(DATAI_14_), .S(n2636), .Z(n3523) );
  NAND2_X1 U32890 ( .A1(n3518), .A2(n3523), .ZN(n3824) );
  INV_X1 U32900 ( .A(n3518), .ZN(n3811) );
  NAND2_X1 U32910 ( .A1(n3811), .A2(n3517), .ZN(n3825) );
  NAND2_X1 U32920 ( .A1(n3824), .A2(n3825), .ZN(n3331) );
  NAND2_X1 U32930 ( .A1(n3518), .A2(n3517), .ZN(n2591) );
  NAND2_X1 U32940 ( .A1(n2746), .A2(REG0_REG_15__SCAN_IN), .ZN(n2597) );
  NOR2_X1 U32950 ( .A1(n2592), .A2(REG3_REG_15__SCAN_IN), .ZN(n2593) );
  OR2_X1 U32960 ( .A1(n2612), .A2(n2593), .ZN(n3816) );
  INV_X1 U32970 ( .A(n3816), .ZN(n3348) );
  NAND2_X1 U32980 ( .A1(n2698), .A2(n3348), .ZN(n2596) );
  NAND2_X1 U32990 ( .A1(n2944), .A2(REG1_REG_15__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U33000 ( .A1(n2798), .A2(REG2_REG_15__SCAN_IN), .ZN(n2594) );
  INV_X1 U33010 ( .A(IR_REG_14__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U33020 ( .A1(n2621), .A2(n2598), .ZN(n2599) );
  NAND2_X1 U33030 ( .A1(n2599), .A2(IR_REG_31__SCAN_IN), .ZN(n2600) );
  INV_X1 U33040 ( .A(IR_REG_15__SCAN_IN), .ZN(n4611) );
  NAND2_X1 U33050 ( .A1(n2600), .A2(n4611), .ZN(n2608) );
  OR2_X1 U33060 ( .A1(n2600), .A2(n4611), .ZN(n2601) );
  MUX2_X1 U33070 ( .A(n4056), .B(DATAI_15_), .S(n2636), .Z(n3810) );
  NAND2_X1 U33080 ( .A1(n4379), .A2(n3810), .ZN(n2602) );
  INV_X1 U33090 ( .A(n3810), .ZN(n3557) );
  INV_X1 U33100 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2603) );
  XNOR2_X1 U33110 ( .A(n2612), .B(n2603), .ZN(n3739) );
  NAND2_X1 U33120 ( .A1(n2698), .A2(n3739), .ZN(n2607) );
  NAND2_X1 U33130 ( .A1(n2944), .A2(REG1_REG_16__SCAN_IN), .ZN(n2606) );
  INV_X1 U33140 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4773) );
  OR2_X1 U33150 ( .A1(n2948), .A2(n4773), .ZN(n2605) );
  NAND2_X1 U33160 ( .A1(n2945), .A2(REG2_REG_16__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U33170 ( .A1(n2608), .A2(IR_REG_31__SCAN_IN), .ZN(n2609) );
  XNOR2_X1 U33180 ( .A(n2609), .B(IR_REG_16__SCAN_IN), .ZN(n4057) );
  MUX2_X1 U33190 ( .A(n4057), .B(DATAI_16_), .S(n2636), .Z(n3738) );
  NAND2_X1 U33200 ( .A1(n4368), .A2(n3738), .ZN(n3959) );
  NAND2_X1 U33210 ( .A1(n3995), .A2(n4373), .ZN(n3955) );
  NAND2_X1 U33220 ( .A1(n3463), .A2(n2610), .ZN(n3464) );
  NAND2_X1 U33230 ( .A1(n3995), .A2(n3738), .ZN(n2611) );
  AOI22_X1 U33240 ( .A1(n2746), .A2(REG0_REG_17__SCAN_IN), .B1(n2944), .B2(
        REG1_REG_17__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U33250 ( .A1(n2612), .A2(REG3_REG_16__SCAN_IN), .ZN(n2614) );
  INV_X1 U33260 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U33270 ( .A1(n2614), .A2(n2613), .ZN(n2615) );
  AND2_X1 U33280 ( .A1(n2615), .A2(n2629), .ZN(n3750) );
  AOI22_X1 U33290 ( .A1(n2698), .A2(n3750), .B1(n2798), .B2(
        REG2_REG_17__SCAN_IN), .ZN(n2616) );
  INV_X1 U33300 ( .A(n2618), .ZN(n2619) );
  NOR2_X1 U33310 ( .A1(n2619), .A2(IR_REG_14__SCAN_IN), .ZN(n2620) );
  NAND2_X1 U33320 ( .A1(n2623), .A2(IR_REG_31__SCAN_IN), .ZN(n2622) );
  MUX2_X1 U33330 ( .A(IR_REG_31__SCAN_IN), .B(n2622), .S(IR_REG_17__SCAN_IN), 
        .Z(n2624) );
  NAND2_X1 U33340 ( .A1(n2624), .A2(n2646), .ZN(n4063) );
  INV_X1 U33350 ( .A(DATAI_17_), .ZN(n2625) );
  MUX2_X1 U33360 ( .A(n4063), .B(n2625), .S(n2636), .Z(n3572) );
  NAND2_X1 U33370 ( .A1(n4374), .A2(n3572), .ZN(n2627) );
  INV_X1 U33380 ( .A(n3572), .ZN(n4361) );
  AND2_X1 U33390 ( .A1(n3994), .A2(n4361), .ZN(n2626) );
  NAND2_X1 U33400 ( .A1(n2746), .A2(REG0_REG_18__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U33410 ( .A1(n2629), .A2(n2628), .ZN(n2630) );
  AND2_X1 U33420 ( .A1(n2640), .A2(n2630), .ZN(n4287) );
  NAND2_X1 U33430 ( .A1(n2698), .A2(n4287), .ZN(n2633) );
  NAND2_X1 U33440 ( .A1(n2944), .A2(REG1_REG_18__SCAN_IN), .ZN(n2632) );
  NAND2_X1 U33450 ( .A1(n2798), .A2(REG2_REG_18__SCAN_IN), .ZN(n2631) );
  NAND4_X1 U33460 ( .A1(n2634), .A2(n2633), .A3(n2632), .A4(n2631), .ZN(n4364)
         );
  NAND2_X1 U33470 ( .A1(n2646), .A2(IR_REG_31__SCAN_IN), .ZN(n2635) );
  XNOR2_X1 U33480 ( .A(n2635), .B(IR_REG_18__SCAN_IN), .ZN(n4074) );
  MUX2_X1 U33490 ( .A(n4074), .B(DATAI_18_), .S(n2636), .Z(n4284) );
  NAND2_X1 U33500 ( .A1(n4265), .A2(n4284), .ZN(n4257) );
  INV_X1 U33510 ( .A(n4284), .ZN(n2637) );
  NAND2_X1 U33520 ( .A1(n4364), .A2(n2637), .ZN(n4258) );
  NAND2_X1 U3353 ( .A1(n4257), .A2(n4258), .ZN(n4278) );
  NAND2_X1 U33540 ( .A1(n4265), .A2(n2637), .ZN(n2638) );
  AND2_X1 U3355 ( .A1(n2640), .A2(n2639), .ZN(n2641) );
  OR2_X1 U3356 ( .A1(n2641), .A2(n2650), .ZN(n4269) );
  NAND2_X1 U3357 ( .A1(n2798), .A2(REG2_REG_19__SCAN_IN), .ZN(n2642) );
  OAI21_X1 U3358 ( .B1(n4269), .B2(n2142), .A(n2642), .ZN(n2643) );
  INV_X1 U3359 ( .A(n2643), .ZN(n2645) );
  AOI22_X1 U3360 ( .A1(n2746), .A2(REG0_REG_19__SCAN_IN), .B1(n2944), .B2(
        REG1_REG_19__SCAN_IN), .ZN(n2644) );
  OAI21_X2 U3361 ( .B1(n2646), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2647) );
  NAND2_X1 U3362 ( .A1(n2647), .A2(n4730), .ZN(n2705) );
  OR2_X1 U3363 ( .A1(n2647), .A2(n4730), .ZN(n2648) );
  MUX2_X1 U3364 ( .A(n4667), .B(DATAI_19_), .S(n2636), .Z(n4266) );
  NAND2_X1 U3365 ( .A1(n4279), .A2(n4266), .ZN(n2649) );
  NOR2_X1 U3366 ( .A1(n2650), .A2(REG3_REG_20__SCAN_IN), .ZN(n2651) );
  OR2_X1 U3367 ( .A1(n2654), .A2(n2651), .ZN(n4247) );
  AOI22_X1 U3368 ( .A1(n2746), .A2(REG0_REG_20__SCAN_IN), .B1(n2944), .B2(
        REG1_REG_20__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U3369 ( .A1(n2798), .A2(REG2_REG_20__SCAN_IN), .ZN(n2652) );
  AND2_X1 U3370 ( .A1(n4341), .A2(n4245), .ZN(n3897) );
  OR2_X1 U3371 ( .A1(n4341), .A2(n4245), .ZN(n3898) );
  OR2_X1 U3372 ( .A1(n2654), .A2(REG3_REG_21__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3373 ( .A1(n2659), .A2(n2655), .ZN(n4224) );
  AOI22_X1 U3374 ( .A1(n2746), .A2(REG0_REG_21__SCAN_IN), .B1(n2944), .B2(
        REG1_REG_21__SCAN_IN), .ZN(n2657) );
  NAND2_X1 U3375 ( .A1(n2798), .A2(REG2_REG_21__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U3376 ( .A1(n2636), .A2(DATAI_21_), .ZN(n4221) );
  NAND2_X1 U3377 ( .A1(n4201), .A2(n4340), .ZN(n2658) );
  INV_X1 U3378 ( .A(n4201), .ZN(n4238) );
  NAND2_X1 U3379 ( .A1(n2659), .A2(n4868), .ZN(n2660) );
  NAND2_X1 U3380 ( .A1(n2667), .A2(n2660), .ZN(n3778) );
  OR2_X1 U3381 ( .A1(n3778), .A2(n2142), .ZN(n2665) );
  INV_X1 U3382 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4407) );
  NAND2_X1 U3383 ( .A1(n2944), .A2(REG1_REG_22__SCAN_IN), .ZN(n2662) );
  NAND2_X1 U3384 ( .A1(n2798), .A2(REG2_REG_22__SCAN_IN), .ZN(n2661) );
  OAI211_X1 U3385 ( .C1(n2948), .C2(n4407), .A(n2662), .B(n2661), .ZN(n2663)
         );
  INV_X1 U3386 ( .A(n2663), .ZN(n2664) );
  NAND2_X1 U3387 ( .A1(n4344), .A2(n4205), .ZN(n4180) );
  NAND2_X1 U3388 ( .A1(n3993), .A2(n3638), .ZN(n2739) );
  NAND2_X1 U3389 ( .A1(n4180), .A2(n2739), .ZN(n4210) );
  NAND2_X1 U3390 ( .A1(n2667), .A2(n3702), .ZN(n2668) );
  AND2_X1 U3391 ( .A1(n2675), .A2(n2668), .ZN(n4191) );
  NAND2_X1 U3392 ( .A1(n4191), .A2(n2698), .ZN(n2673) );
  INV_X1 U3393 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4403) );
  NAND2_X1 U3394 ( .A1(n2944), .A2(REG1_REG_23__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U3395 ( .A1(n2945), .A2(REG2_REG_23__SCAN_IN), .ZN(n2669) );
  OAI211_X1 U3396 ( .C1(n2948), .C2(n4403), .A(n2670), .B(n2669), .ZN(n2671)
         );
  INV_X1 U3397 ( .A(n2671), .ZN(n2672) );
  NAND2_X1 U3398 ( .A1(n2636), .A2(DATAI_23_), .ZN(n4189) );
  NAND2_X1 U3399 ( .A1(n4204), .A2(n4189), .ZN(n2674) );
  AND2_X1 U3400 ( .A1(n2675), .A2(n4702), .ZN(n2676) );
  OR2_X1 U3401 ( .A1(n2676), .A2(n2683), .ZN(n3761) );
  INV_X1 U3402 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4778) );
  NAND2_X1 U3403 ( .A1(n2944), .A2(REG1_REG_24__SCAN_IN), .ZN(n2678) );
  NAND2_X1 U3404 ( .A1(n2798), .A2(REG2_REG_24__SCAN_IN), .ZN(n2677) );
  OAI211_X1 U3405 ( .C1(n2948), .C2(n4778), .A(n2678), .B(n2677), .ZN(n2679)
         );
  INV_X1 U3406 ( .A(n2679), .ZN(n2680) );
  INV_X1 U3407 ( .A(n4320), .ZN(n4151) );
  NAND2_X1 U3408 ( .A1(n2636), .A2(DATAI_24_), .ZN(n4170) );
  NAND2_X1 U3409 ( .A1(n2682), .A2(n2681), .ZN(n4142) );
  NOR2_X1 U3410 ( .A1(n2683), .A2(REG3_REG_25__SCAN_IN), .ZN(n2684) );
  INV_X1 U3411 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U3412 ( .A1(n2944), .A2(REG1_REG_25__SCAN_IN), .ZN(n2686) );
  NAND2_X1 U3413 ( .A1(n2945), .A2(REG2_REG_25__SCAN_IN), .ZN(n2685) );
  OAI211_X1 U3414 ( .C1(n2948), .C2(n4396), .A(n2686), .B(n2685), .ZN(n2687)
         );
  INV_X1 U3415 ( .A(n2687), .ZN(n2688) );
  INV_X1 U3416 ( .A(n4165), .ZN(n3799) );
  NAND2_X1 U3417 ( .A1(n2636), .A2(DATAI_25_), .ZN(n4145) );
  INV_X1 U3418 ( .A(n4145), .ZN(n4319) );
  NOR2_X1 U3419 ( .A1(n2691), .A2(REG3_REG_26__SCAN_IN), .ZN(n2692) );
  INV_X1 U3420 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4777) );
  NAND2_X1 U3421 ( .A1(n2944), .A2(REG1_REG_26__SCAN_IN), .ZN(n2694) );
  NAND2_X1 U3422 ( .A1(n2798), .A2(REG2_REG_26__SCAN_IN), .ZN(n2693) );
  OAI211_X1 U3423 ( .C1(n2948), .C2(n4777), .A(n2694), .B(n2693), .ZN(n2695)
         );
  INV_X1 U3424 ( .A(n2695), .ZN(n2696) );
  NAND2_X1 U3425 ( .A1(n2636), .A2(DATAI_26_), .ZN(n4133) );
  NOR2_X1 U3426 ( .A1(n4308), .A2(n3802), .ZN(n3890) );
  XNOR2_X1 U3427 ( .A(n2697), .B(n4704), .ZN(n4112) );
  NAND2_X1 U3428 ( .A1(n4112), .A2(n2698), .ZN(n2703) );
  INV_X1 U3429 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4389) );
  NAND2_X1 U3430 ( .A1(n2944), .A2(REG1_REG_27__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U3431 ( .A1(n2798), .A2(REG2_REG_27__SCAN_IN), .ZN(n2699) );
  OAI211_X1 U3432 ( .C1(n2948), .C2(n4389), .A(n2700), .B(n2699), .ZN(n2701)
         );
  INV_X1 U3433 ( .A(n2701), .ZN(n2702) );
  NAND2_X1 U3434 ( .A1(n2636), .A2(DATAI_27_), .ZN(n4117) );
  INV_X1 U3435 ( .A(n4129), .ZN(n4102) );
  INV_X1 U3436 ( .A(n2708), .ZN(n2709) );
  NAND2_X1 U3437 ( .A1(n2709), .A2(IR_REG_31__SCAN_IN), .ZN(n2710) );
  MUX2_X1 U3438 ( .A(IR_REG_31__SCAN_IN), .B(n2710), .S(IR_REG_21__SCAN_IN), 
        .Z(n2712) );
  NAND2_X1 U3439 ( .A1(n2712), .A2(n2711), .ZN(n2752) );
  NAND2_X1 U3440 ( .A1(n2711), .A2(IR_REG_31__SCAN_IN), .ZN(n2713) );
  XNOR2_X1 U3441 ( .A(n3045), .B(n4429), .ZN(n2714) );
  NAND2_X1 U3442 ( .A1(n2714), .A2(n4081), .ZN(n4241) );
  NAND2_X1 U3443 ( .A1(n3980), .A2(n4667), .ZN(n4542) );
  NAND2_X1 U3444 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U3445 ( .A1(n2802), .A2(n2716), .ZN(n2717) );
  INV_X1 U3446 ( .A(n2896), .ZN(n2895) );
  NAND2_X1 U3447 ( .A1(n2895), .A2(n2985), .ZN(n3908) );
  NAND2_X1 U3448 ( .A1(n2999), .A2(n3912), .ZN(n2720) );
  NAND2_X1 U3449 ( .A1(n2720), .A2(n3880), .ZN(n3001) );
  NAND2_X1 U3450 ( .A1(n3001), .A2(n3913), .ZN(n3067) );
  NAND2_X1 U3451 ( .A1(n3055), .A2(n3092), .ZN(n3918) );
  NAND2_X1 U3452 ( .A1(n4580), .A2(n3065), .ZN(n3915) );
  INV_X1 U3453 ( .A(n3919), .ZN(n2721) );
  AND2_X1 U3454 ( .A1(n3164), .A2(n3127), .ZN(n3100) );
  NAND2_X1 U3455 ( .A1(n4574), .A2(n3130), .ZN(n3934) );
  INV_X1 U3456 ( .A(n3163), .ZN(n3159) );
  NAND2_X1 U3457 ( .A1(n4000), .A2(n3159), .ZN(n3936) );
  INV_X1 U34580 ( .A(n4000), .ZN(n3160) );
  NAND2_X1 U34590 ( .A1(n3160), .A2(n3163), .ZN(n3924) );
  INV_X1 U3460 ( .A(n2722), .ZN(n2723) );
  NAND2_X1 U3461 ( .A1(n3289), .A2(n3536), .ZN(n3929) );
  NAND2_X1 U3462 ( .A1(n3208), .A2(n3929), .ZN(n2724) );
  NAND2_X1 U3463 ( .A1(n3999), .A2(n3288), .ZN(n3927) );
  AND2_X1 U3464 ( .A1(n3998), .A2(n3292), .ZN(n3932) );
  NAND2_X1 U3465 ( .A1(n3607), .A2(n3296), .ZN(n3930) );
  NAND2_X1 U3466 ( .A1(n3997), .A2(n3605), .ZN(n3945) );
  NAND2_X1 U34670 ( .A1(n3372), .A2(n3389), .ZN(n3940) );
  NAND2_X1 U3468 ( .A1(n2725), .A2(n3940), .ZN(n3367) );
  NAND2_X1 U34690 ( .A1(n3502), .A2(n3357), .ZN(n3410) );
  NAND2_X1 U3470 ( .A1(n3594), .A2(n3418), .ZN(n2726) );
  NAND2_X1 U34710 ( .A1(n3410), .A2(n2726), .ZN(n3946) );
  INV_X1 U3472 ( .A(n3366), .ZN(n3948) );
  NOR2_X1 U34730 ( .A1(n3946), .A2(n3948), .ZN(n2727) );
  NAND2_X1 U3474 ( .A1(n2728), .A2(n3593), .ZN(n3412) );
  NAND2_X1 U34750 ( .A1(n3364), .A2(n3412), .ZN(n2731) );
  INV_X1 U3476 ( .A(n3946), .ZN(n2730) );
  NOR2_X1 U34770 ( .A1(n3594), .A2(n3418), .ZN(n2729) );
  AOI21_X1 U3478 ( .B1(n2731), .B2(n2730), .A(n2729), .ZN(n3954) );
  INV_X1 U34790 ( .A(n3331), .ZN(n3881) );
  NAND2_X1 U3480 ( .A1(n3558), .A2(n3810), .ZN(n3827) );
  NAND2_X1 U34810 ( .A1(n4379), .A2(n3557), .ZN(n3826) );
  NAND2_X1 U3482 ( .A1(n3827), .A2(n3826), .ZN(n3872) );
  NAND2_X1 U34830 ( .A1(n3343), .A2(n3826), .ZN(n3466) );
  NAND2_X1 U3484 ( .A1(n3466), .A2(n3873), .ZN(n3465) );
  NAND2_X1 U34850 ( .A1(n3465), .A2(n3955), .ZN(n4256) );
  AND2_X1 U3486 ( .A1(n3994), .A2(n3572), .ZN(n4255) );
  INV_X1 U34870 ( .A(n4266), .ZN(n2735) );
  NAND2_X1 U3488 ( .A1(n4279), .A2(n2735), .ZN(n3899) );
  NAND2_X1 U34890 ( .A1(n3899), .A2(n4258), .ZN(n2732) );
  OR2_X2 U3490 ( .A1(n4256), .A2(n3958), .ZN(n4233) );
  INV_X1 U34910 ( .A(n2732), .ZN(n2734) );
  NAND2_X1 U3492 ( .A1(n4374), .A2(n4361), .ZN(n4254) );
  NAND2_X1 U34930 ( .A1(n4257), .A2(n4254), .ZN(n2733) );
  NAND2_X1 U3494 ( .A1(n2734), .A2(n2733), .ZN(n2736) );
  OR2_X1 U34950 ( .A1(n4279), .A2(n2735), .ZN(n3900) );
  NAND2_X1 U3496 ( .A1(n2736), .A2(n3900), .ZN(n4234) );
  NOR2_X1 U34970 ( .A1(n4341), .A2(n2787), .ZN(n2737) );
  NOR2_X1 U3498 ( .A1(n4234), .A2(n2737), .ZN(n3831) );
  NAND2_X1 U34990 ( .A1(n4233), .A2(n3831), .ZN(n2738) );
  NAND2_X1 U3500 ( .A1(n4925), .A2(n2787), .ZN(n3962) );
  NAND2_X1 U35010 ( .A1(n2738), .A2(n3962), .ZN(n4216) );
  OR2_X1 U3502 ( .A1(n4201), .A2(n4221), .ZN(n4197) );
  NAND2_X1 U35030 ( .A1(n4180), .A2(n4197), .ZN(n3969) );
  INV_X1 U3504 ( .A(n3969), .ZN(n3834) );
  NAND2_X1 U35050 ( .A1(n4216), .A2(n3834), .ZN(n2741) );
  NAND2_X1 U35060 ( .A1(n4162), .A2(n4189), .ZN(n3896) );
  NAND2_X1 U35070 ( .A1(n3896), .A2(n2739), .ZN(n3838) );
  AND2_X1 U35080 ( .A1(n4201), .A2(n4221), .ZN(n4177) );
  AND2_X1 U35090 ( .A1(n4180), .A2(n4177), .ZN(n3836) );
  NOR2_X1 U35100 ( .A1(n3838), .A2(n3836), .ZN(n2740) );
  NAND2_X1 U35110 ( .A1(n2741), .A2(n2740), .ZN(n4158) );
  OR2_X1 U35120 ( .A1(n4320), .A2(n4170), .ZN(n3894) );
  NAND2_X1 U35130 ( .A1(n4204), .A2(n3701), .ZN(n4157) );
  NAND2_X1 U35140 ( .A1(n4158), .A2(n3965), .ZN(n2742) );
  AND2_X1 U35150 ( .A1(n4320), .A2(n4170), .ZN(n3837) );
  INV_X1 U35160 ( .A(n3837), .ZN(n3895) );
  NAND2_X1 U35170 ( .A1(n2742), .A2(n3895), .ZN(n4140) );
  AND2_X1 U35180 ( .A1(n4165), .A2(n4145), .ZN(n3861) );
  OR2_X2 U35190 ( .A1(n4140), .A2(n3861), .ZN(n2743) );
  OR2_X1 U35200 ( .A1(n4165), .A2(n4145), .ZN(n3862) );
  OR2_X1 U35210 ( .A1(n4308), .A2(n4133), .ZN(n3839) );
  AND2_X1 U35220 ( .A1(n4308), .A2(n4133), .ZN(n3850) );
  XNOR2_X1 U35230 ( .A(n4129), .B(n4307), .ZN(n4110) );
  OR2_X1 U35240 ( .A1(n4129), .A2(n4117), .ZN(n3842) );
  INV_X1 U35250 ( .A(n3842), .ZN(n3852) );
  XNOR2_X1 U35260 ( .A(n2795), .B(n3860), .ZN(n2745) );
  INV_X1 U35270 ( .A(n3980), .ZN(n4431) );
  NAND2_X1 U35280 ( .A1(n4431), .A2(n4430), .ZN(n3984) );
  INV_X1 U35290 ( .A(n4429), .ZN(n2753) );
  OR2_X1 U35300 ( .A1(n4081), .A2(n2753), .ZN(n2744) );
  NAND2_X1 U35310 ( .A1(n2745), .A2(n4282), .ZN(n4107) );
  OR2_X1 U35320 ( .A1(n4087), .A2(n2142), .ZN(n2751) );
  INV_X1 U35330 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4093) );
  NAND2_X1 U35340 ( .A1(n2944), .A2(REG1_REG_29__SCAN_IN), .ZN(n2748) );
  NAND2_X1 U35350 ( .A1(n2746), .A2(REG0_REG_29__SCAN_IN), .ZN(n2747) );
  OAI211_X1 U35360 ( .C1(n4093), .C2(n2448), .A(n2748), .B(n2747), .ZN(n2749)
         );
  INV_X1 U35370 ( .A(n2749), .ZN(n2750) );
  NAND2_X1 U35380 ( .A1(n2751), .A2(n2750), .ZN(n4098) );
  AOI22_X1 U35390 ( .A1(n4098), .A2(n4363), .B1(n4362), .B2(n4096), .ZN(n2754)
         );
  OAI211_X1 U35400 ( .C1(n4102), .C2(n4367), .A(n4107), .B(n2754), .ZN(n2755)
         );
  AOI21_X1 U35410 ( .B1(n4094), .B2(n4593), .A(n2755), .ZN(n2791) );
  OR2_X1 U35420 ( .A1(n2757), .A2(n2756), .ZN(n2759) );
  NAND2_X1 U35430 ( .A1(n2162), .A2(IR_REG_31__SCAN_IN), .ZN(n2766) );
  NAND2_X1 U35440 ( .A1(n2766), .A2(n4607), .ZN(n2768) );
  NOR2_X1 U35450 ( .A1(n2772), .A2(n2828), .ZN(n2765) );
  XNOR2_X2 U35460 ( .A(n2764), .B(IR_REG_26__SCAN_IN), .ZN(n4427) );
  OR2_X1 U35470 ( .A1(n2766), .A2(n4607), .ZN(n2767) );
  NAND2_X1 U35480 ( .A1(n2768), .A2(n2767), .ZN(n3032) );
  INV_X1 U35490 ( .A(n4551), .ZN(n2769) );
  NAND2_X1 U35500 ( .A1(n2891), .A2(n2769), .ZN(n2834) );
  NAND2_X1 U35510 ( .A1(n3980), .A2(n4081), .ZN(n2904) );
  AND2_X1 U35520 ( .A1(n2904), .A2(n2905), .ZN(n3031) );
  OR2_X1 U35530 ( .A1(n2834), .A2(n3031), .ZN(n3040) );
  NOR2_X1 U35540 ( .A1(n4353), .A2(n4430), .ZN(n2918) );
  NOR2_X1 U35550 ( .A1(n3040), .A2(n2918), .ZN(n2782) );
  NAND2_X1 U35560 ( .A1(n2772), .A2(n2828), .ZN(n2770) );
  MUX2_X1 U35570 ( .A(n2828), .B(n2770), .S(B_REG_SCAN_IN), .Z(n2771) );
  INV_X1 U35580 ( .A(n2772), .ZN(n4428) );
  OAI22_X1 U35590 ( .A1(n2825), .A2(D_REG_1__SCAN_IN), .B1(n4428), .B2(n4427), 
        .ZN(n2901) );
  INV_X1 U35600 ( .A(D_REG_22__SCAN_IN), .ZN(n4750) );
  INV_X1 U35610 ( .A(D_REG_27__SCAN_IN), .ZN(n4753) );
  INV_X1 U35620 ( .A(D_REG_8__SCAN_IN), .ZN(n4867) );
  INV_X1 U35630 ( .A(D_REG_9__SCAN_IN), .ZN(n4864) );
  NAND4_X1 U35640 ( .A1(n4750), .A2(n4753), .A3(n4867), .A4(n4864), .ZN(n4616)
         );
  NOR4_X1 U35650 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2776) );
  NOR4_X1 U35660 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2775) );
  NOR4_X1 U35670 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2774) );
  NOR4_X1 U35680 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2773) );
  NAND4_X1 U35690 ( .A1(n2776), .A2(n2775), .A3(n2774), .A4(n2773), .ZN(n2777)
         );
  NOR4_X1 U35700 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(n4616), 
        .A4(n2777), .ZN(n2780) );
  INV_X1 U35710 ( .A(D_REG_2__SCAN_IN), .ZN(n4740) );
  INV_X1 U35720 ( .A(D_REG_17__SCAN_IN), .ZN(n4747) );
  NAND2_X1 U35730 ( .A1(n4740), .A2(n4747), .ZN(n4617) );
  INV_X1 U35740 ( .A(D_REG_31__SCAN_IN), .ZN(n4761) );
  INV_X1 U35750 ( .A(D_REG_3__SCAN_IN), .ZN(n4744) );
  INV_X1 U35760 ( .A(D_REG_14__SCAN_IN), .ZN(n4748) );
  INV_X1 U35770 ( .A(D_REG_26__SCAN_IN), .ZN(n4754) );
  NAND4_X1 U35780 ( .A1(n4761), .A2(n4744), .A3(n4748), .A4(n4754), .ZN(n2778)
         );
  NOR4_X1 U35790 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(n4617), 
        .A4(n2778), .ZN(n2779) );
  NAND2_X1 U35800 ( .A1(n2780), .A2(n2779), .ZN(n2781) );
  NAND2_X1 U35810 ( .A1(n2785), .A2(n2781), .ZN(n3041) );
  INV_X1 U3582 ( .A(D_REG_0__SCAN_IN), .ZN(n2831) );
  INV_X1 U3583 ( .A(n4427), .ZN(n2783) );
  MUX2_X1 U3584 ( .A(n2786), .B(n2791), .S(n4604), .Z(n2789) );
  INV_X1 U3585 ( .A(n2985), .ZN(n2939) );
  NAND2_X1 U3586 ( .A1(n4586), .A2(n3127), .ZN(n3142) );
  OAI21_X1 U3587 ( .B1(n4115), .B2(n3674), .A(n2807), .ZN(n4095) );
  NAND2_X1 U3588 ( .A1(n2789), .A2(n2788), .ZN(U3546) );
  INV_X1 U3589 ( .A(n2902), .ZN(n3043) );
  MUX2_X1 U3590 ( .A(n4780), .B(n2791), .S(n4600), .Z(n2793) );
  NAND2_X1 U3591 ( .A1(n2793), .A2(n2792), .ZN(U3514) );
  INV_X1 U3592 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2806) );
  NAND2_X1 U3593 ( .A1(n2636), .A2(DATAI_29_), .ZN(n3847) );
  XNOR2_X1 U3594 ( .A(n4098), .B(n3847), .ZN(n3904) );
  XOR2_X1 U3595 ( .A(n3904), .B(n2796), .Z(n2797) );
  NAND2_X1 U3596 ( .A1(n2797), .A2(n4282), .ZN(n2805) );
  INV_X1 U3597 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2801) );
  NAND2_X1 U3598 ( .A1(n2944), .A2(REG1_REG_30__SCAN_IN), .ZN(n2800) );
  NAND2_X1 U3599 ( .A1(n2798), .A2(REG2_REG_30__SCAN_IN), .ZN(n2799) );
  OAI211_X1 U3600 ( .C1(n2948), .C2(n2801), .A(n2800), .B(n2799), .ZN(n3846)
         );
  XNOR2_X1 U3601 ( .A(n2802), .B(IR_REG_27__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U3602 ( .A1(n4426), .A2(B_REG_SCAN_IN), .ZN(n2803) );
  AND2_X1 U3603 ( .A1(n4363), .A2(n2803), .ZN(n4294) );
  INV_X1 U3604 ( .A(n3847), .ZN(n3840) );
  AOI22_X1 U3605 ( .A1(n3846), .A2(n4294), .B1(n3840), .B2(n4362), .ZN(n2804)
         );
  OAI211_X1 U3606 ( .C1(n4311), .C2(n4367), .A(n2805), .B(n2804), .ZN(n4090)
         );
  MUX2_X1 U3607 ( .A(n2806), .B(n2811), .S(n4604), .Z(n2810) );
  INV_X1 U3608 ( .A(n2807), .ZN(n2808) );
  OAI21_X1 U3609 ( .B1(n2808), .B2(n3847), .A(n4300), .ZN(n4088) );
  NAND2_X1 U3610 ( .A1(n2810), .A2(n2809), .ZN(U3547) );
  INV_X1 U3611 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2812) );
  NAND2_X1 U3612 ( .A1(n2814), .A2(n2813), .ZN(U3515) );
  INV_X2 U3613 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  MUX2_X1 U3614 ( .A(n2523), .B(n3258), .S(STATE_REG_SCAN_IN), .Z(n2815) );
  INV_X1 U3615 ( .A(n2815), .ZN(U3344) );
  INV_X1 U3616 ( .A(DATAI_13_), .ZN(n4687) );
  NAND2_X1 U3617 ( .A1(n4052), .A2(STATE_REG_SCAN_IN), .ZN(n2816) );
  OAI21_X1 U3618 ( .B1(STATE_REG_SCAN_IN), .B2(n4687), .A(n2816), .ZN(U3339)
         );
  INV_X1 U3619 ( .A(n4063), .ZN(n4072) );
  NAND2_X1 U3620 ( .A1(n4072), .A2(STATE_REG_SCAN_IN), .ZN(n2817) );
  OAI21_X1 U3621 ( .B1(STATE_REG_SCAN_IN), .B2(n2625), .A(n2817), .ZN(U3335)
         );
  INV_X1 U3622 ( .A(DATAI_24_), .ZN(n4678) );
  MUX2_X1 U3623 ( .A(n4678), .B(n2828), .S(STATE_REG_SCAN_IN), .Z(n2818) );
  INV_X1 U3624 ( .A(n2818), .ZN(U3328) );
  INV_X1 U3625 ( .A(DATAI_29_), .ZN(n4671) );
  NAND2_X1 U3626 ( .A1(n2819), .A2(STATE_REG_SCAN_IN), .ZN(n2820) );
  OAI21_X1 U3627 ( .B1(STATE_REG_SCAN_IN), .B2(n4671), .A(n2820), .ZN(U3323)
         );
  INV_X1 U3628 ( .A(DATAI_28_), .ZN(n4675) );
  NAND2_X1 U3629 ( .A1(n2979), .A2(STATE_REG_SCAN_IN), .ZN(n2821) );
  OAI21_X1 U3630 ( .B1(STATE_REG_SCAN_IN), .B2(n4675), .A(n2821), .ZN(U3324)
         );
  INV_X1 U3631 ( .A(DATAI_30_), .ZN(n2824) );
  NAND2_X1 U3632 ( .A1(n2822), .A2(STATE_REG_SCAN_IN), .ZN(n2823) );
  OAI21_X1 U3633 ( .B1(STATE_REG_SCAN_IN), .B2(n2824), .A(n2823), .ZN(U3322)
         );
  INV_X1 U3634 ( .A(D_REG_1__SCAN_IN), .ZN(n2827) );
  NOR3_X1 U3635 ( .A1(n4428), .A2(n4427), .A3(n4551), .ZN(n2826) );
  AOI21_X1 U3636 ( .B1(n4549), .B2(n2827), .A(n2826), .ZN(U3459) );
  INV_X1 U3637 ( .A(n2828), .ZN(n2829) );
  NOR3_X1 U3638 ( .A1(n4427), .A2(n2829), .A3(n4551), .ZN(n2830) );
  AOI21_X1 U3639 ( .B1(n4549), .B2(n2831), .A(n2830), .ZN(U3458) );
  NAND2_X1 U3640 ( .A1(n2905), .A2(n3032), .ZN(n2832) );
  AND2_X1 U3641 ( .A1(n2458), .A2(n2832), .ZN(n2838) );
  INV_X1 U3642 ( .A(n2838), .ZN(n2835) );
  INV_X1 U3643 ( .A(n3032), .ZN(n2833) );
  NAND2_X1 U3644 ( .A1(n2833), .A2(STATE_REG_SCAN_IN), .ZN(n3991) );
  NAND2_X1 U3645 ( .A1(n2834), .A2(n3991), .ZN(n2839) );
  INV_X1 U3646 ( .A(n4523), .ZN(n2883) );
  INV_X1 U3647 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n2843) );
  INV_X1 U3648 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4547) );
  AOI21_X1 U3649 ( .B1(n4426), .B2(n4547), .A(n2911), .ZN(n2925) );
  OAI21_X1 U3650 ( .B1(n4426), .B2(REG1_REG_0__SCAN_IN), .A(n2364), .ZN(n2837)
         );
  NOR2_X1 U3651 ( .A1(n2925), .A2(IR_REG_0__SCAN_IN), .ZN(n2836) );
  AOI21_X1 U3652 ( .B1(n2925), .B2(n2837), .A(n2836), .ZN(n2840) );
  AOI22_X1 U3653 ( .A1(n2840), .A2(n2853), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2842) );
  INV_X1 U3654 ( .A(n4426), .ZN(n2922) );
  INV_X1 U3655 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2897) );
  NAND3_X1 U3656 ( .A1(n4525), .A2(IR_REG_0__SCAN_IN), .A3(n2897), .ZN(n2841)
         );
  OAI211_X1 U3657 ( .C1(n2883), .C2(n2843), .A(n2842), .B(n2841), .ZN(U3240)
         );
  NOR2_X1 U3658 ( .A1(n4523), .A2(U4043), .ZN(U3148) );
  INV_X1 U3659 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U3660 ( .A1(n3537), .A2(U4043), .ZN(n2844) );
  OAI21_X1 U3661 ( .B1(U4043), .B2(n4881), .A(n2844), .ZN(U3557) );
  INV_X1 U3662 ( .A(n2872), .ZN(n4434) );
  INV_X1 U3663 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4017) );
  INV_X1 U3664 ( .A(n4437), .ZN(n4015) );
  INV_X1 U3665 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2845) );
  AND2_X1 U3666 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2846)
         );
  NAND2_X1 U3667 ( .A1(n4438), .A2(REG2_REG_1__SCAN_IN), .ZN(n4019) );
  NAND2_X1 U3668 ( .A1(n4020), .A2(n4019), .ZN(n2849) );
  MUX2_X1 U3669 ( .A(REG2_REG_2__SCAN_IN), .B(n4017), .S(n4437), .Z(n2848) );
  NAND2_X1 U3670 ( .A1(n2849), .A2(n2848), .ZN(n4022) );
  OAI21_X1 U3671 ( .B1(n4017), .B2(n4015), .A(n4022), .ZN(n2850) );
  XNOR2_X1 U3672 ( .A(n2850), .B(n2858), .ZN(n4034) );
  INV_X1 U3673 ( .A(n4435), .ZN(n2932) );
  INV_X1 U3674 ( .A(n2851), .ZN(n2852) );
  INV_X1 U3675 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4823) );
  MUX2_X1 U3676 ( .A(REG2_REG_5__SCAN_IN), .B(n4823), .S(n2872), .Z(n2869) );
  XNOR2_X1 U3677 ( .A(n2884), .B(REG2_REG_6__SCAN_IN), .ZN(n2865) );
  NOR2_X1 U3678 ( .A1(n2922), .A2(n2911), .ZN(n3987) );
  NAND2_X1 U3679 ( .A1(n2853), .A2(n2911), .ZN(n4530) );
  INV_X1 U3680 ( .A(n4530), .ZN(n4030) );
  NAND2_X1 U3681 ( .A1(n4523), .A2(ADDR_REG_6__SCAN_IN), .ZN(n2854) );
  NAND2_X1 U3682 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U3683 ( .A1(n2854), .A2(n3166), .ZN(n2863) );
  XNOR2_X1 U3684 ( .A(n4006), .B(REG1_REG_1__SCAN_IN), .ZN(n4005) );
  AND2_X1 U3685 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4004)
         );
  NAND2_X1 U3686 ( .A1(n4005), .A2(n4004), .ZN(n4003) );
  NAND2_X1 U3687 ( .A1(n4438), .A2(REG1_REG_1__SCAN_IN), .ZN(n2855) );
  NAND2_X1 U3688 ( .A1(n4003), .A2(n2855), .ZN(n4024) );
  INV_X1 U3689 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2856) );
  NAND2_X1 U3690 ( .A1(n4024), .A2(n4025), .ZN(n4023) );
  NAND2_X1 U3691 ( .A1(n4437), .A2(REG1_REG_2__SCAN_IN), .ZN(n2857) );
  NAND2_X1 U3692 ( .A1(n4023), .A2(n2857), .ZN(n2859) );
  XNOR2_X1 U3693 ( .A(n2859), .B(n2858), .ZN(n4032) );
  NAND2_X1 U3694 ( .A1(n4032), .A2(REG1_REG_3__SCAN_IN), .ZN(n4031) );
  NAND2_X1 U3695 ( .A1(n2859), .A2(n4436), .ZN(n2860) );
  XOR2_X1 U3696 ( .A(REG1_REG_5__SCAN_IN), .B(n2872), .Z(n2867) );
  AOI21_X1 U3697 ( .B1(REG1_REG_5__SCAN_IN), .B2(n4434), .A(n2866), .ZN(n2876)
         );
  INV_X1 U3698 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4797) );
  INV_X1 U3699 ( .A(n4525), .ZN(n4068) );
  AOI211_X1 U3700 ( .C1(n2861), .C2(n4797), .A(n4068), .B(n2877), .ZN(n2862)
         );
  AOI211_X1 U3701 ( .C1(n4030), .C2(n4433), .A(n2863), .B(n2862), .ZN(n2864)
         );
  OAI21_X1 U3702 ( .B1(n2865), .B2(n4519), .A(n2864), .ZN(U3246) );
  AOI211_X1 U3703 ( .C1(n2159), .C2(n2867), .A(n2866), .B(n4068), .ZN(n2875)
         );
  AOI211_X1 U3704 ( .C1(n2870), .C2(n2869), .A(n2868), .B(n4519), .ZN(n2874)
         );
  AND2_X1 U3705 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3131) );
  AOI21_X1 U3706 ( .B1(n4523), .B2(ADDR_REG_5__SCAN_IN), .A(n3131), .ZN(n2871)
         );
  OAI21_X1 U3707 ( .B1(n2872), .B2(n4530), .A(n2871), .ZN(n2873) );
  OR3_X1 U3708 ( .A1(n2875), .A2(n2874), .A3(n2873), .ZN(U3245) );
  INV_X1 U3709 ( .A(n2876), .ZN(n2878) );
  INV_X1 U3710 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4793) );
  MUX2_X1 U3711 ( .A(REG1_REG_7__SCAN_IN), .B(n4793), .S(n4432), .Z(n2879) );
  XNOR2_X1 U3712 ( .A(n3011), .B(n2879), .ZN(n2890) );
  INV_X1 U3713 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n2882) );
  NOR2_X1 U3714 ( .A1(STATE_REG_SCAN_IN), .A2(n2880), .ZN(n3233) );
  INV_X1 U3715 ( .A(n3233), .ZN(n2881) );
  OAI21_X1 U3716 ( .B1(n2883), .B2(n2882), .A(n2881), .ZN(n2888) );
  INV_X1 U3717 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3179) );
  MUX2_X1 U3718 ( .A(n3179), .B(REG2_REG_7__SCAN_IN), .S(n4432), .Z(n2885) );
  NOR2_X1 U3719 ( .A1(n2886), .A2(n2885), .ZN(n3014) );
  AOI211_X1 U3720 ( .C1(n2886), .C2(n2885), .A(n4519), .B(n3014), .ZN(n2887)
         );
  AOI211_X1 U3721 ( .C1(n4030), .C2(n4432), .A(n2888), .B(n2887), .ZN(n2889)
         );
  OAI21_X1 U3722 ( .B1(n2890), .B2(n4068), .A(n2889), .ZN(U3247) );
  INV_X1 U3723 ( .A(n3045), .ZN(n2892) );
  OAI22_X1 U3724 ( .A1(n2939), .A2(n3676), .B1(n2364), .B2(n2891), .ZN(n2893)
         );
  OR2_X1 U3725 ( .A1(n2897), .A2(n2891), .ZN(n2898) );
  NAND2_X1 U3726 ( .A1(n2970), .A2(n2898), .ZN(n2900) );
  NAND2_X1 U3727 ( .A1(n2900), .A2(n2899), .ZN(n2971) );
  OAI21_X1 U3728 ( .B1(n2899), .B2(n2900), .A(n2971), .ZN(n2923) );
  INV_X1 U3729 ( .A(n2901), .ZN(n3042) );
  NAND3_X1 U3730 ( .A1(n3042), .A2(n2902), .A3(n3041), .ZN(n2914) );
  INV_X1 U3731 ( .A(n2914), .ZN(n2903) );
  NAND2_X1 U3732 ( .A1(n2903), .A2(n2917), .ZN(n2916) );
  NAND2_X1 U3733 ( .A1(n2904), .A2(n2937), .ZN(n2907) );
  INV_X1 U3734 ( .A(n2905), .ZN(n2906) );
  NAND2_X1 U3735 ( .A1(n2907), .A2(n2906), .ZN(n2908) );
  NAND2_X1 U3736 ( .A1(n4081), .A2(n4429), .ZN(n2962) );
  NOR2_X1 U3737 ( .A1(n2962), .A2(n4551), .ZN(n2909) );
  INV_X1 U3738 ( .A(n3988), .ZN(n2910) );
  NOR2_X1 U3739 ( .A1(n2914), .A2(n2910), .ZN(n2980) );
  AND2_X2 U3740 ( .A1(n2980), .A2(n2911), .ZN(n3813) );
  INV_X1 U3741 ( .A(n2965), .ZN(n3005) );
  NAND2_X1 U3742 ( .A1(n2937), .A2(n4667), .ZN(n2912) );
  OR2_X1 U3743 ( .A1(n4362), .A2(n2912), .ZN(n2913) );
  NAND2_X1 U3744 ( .A1(n2914), .A2(n2913), .ZN(n3034) );
  INV_X1 U3745 ( .A(n3040), .ZN(n2915) );
  NAND2_X1 U3746 ( .A1(n3034), .A2(n2915), .ZN(n3710) );
  AOI22_X1 U3747 ( .A1(n3813), .A2(n3005), .B1(REG3_REG_0__SCAN_IN), .B2(n3710), .ZN(n2921) );
  OR2_X1 U3748 ( .A1(n2916), .A2(n4571), .ZN(n2919) );
  NAND2_X1 U3749 ( .A1(n3801), .A2(n2985), .ZN(n2920) );
  OAI211_X1 U3750 ( .C1(n2923), .C2(n3806), .A(n2921), .B(n2920), .ZN(U3229)
         );
  NAND3_X1 U3751 ( .A1(n2923), .A2(n2979), .A3(n2922), .ZN(n2927) );
  NAND2_X1 U3752 ( .A1(n3987), .A2(REG2_REG_0__SCAN_IN), .ZN(n2924) );
  MUX2_X1 U3753 ( .A(n2925), .B(n2924), .S(IR_REG_0__SCAN_IN), .Z(n2926) );
  NAND3_X1 U3754 ( .A1(n2927), .A2(U4043), .A3(n2926), .ZN(n4029) );
  XNOR2_X1 U3755 ( .A(n2928), .B(REG2_REG_4__SCAN_IN), .ZN(n2934) );
  OAI211_X1 U3756 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2929), .A(n4525), .B(n2345), 
        .ZN(n2931) );
  AND2_X1 U3757 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4609) );
  AOI21_X1 U3758 ( .B1(n4523), .B2(ADDR_REG_4__SCAN_IN), .A(n4609), .ZN(n2930)
         );
  OAI211_X1 U3759 ( .C1(n4530), .C2(n2932), .A(n2931), .B(n2930), .ZN(n2933)
         );
  AOI21_X1 U3760 ( .B1(n4480), .B2(n2934), .A(n2933), .ZN(n2935) );
  NAND2_X1 U3761 ( .A1(n4029), .A2(n2935), .ZN(U3244) );
  INV_X1 U3762 ( .A(n4353), .ZN(n2941) );
  NAND2_X1 U3763 ( .A1(n2936), .A2(n2939), .ZN(n3910) );
  AND2_X1 U3764 ( .A1(n3908), .A2(n3910), .ZN(n3874) );
  INV_X1 U3765 ( .A(n3874), .ZN(n4545) );
  INV_X1 U3766 ( .A(n2937), .ZN(n2938) );
  NOR2_X1 U3767 ( .A1(n2939), .A2(n2938), .ZN(n4543) );
  INV_X1 U3768 ( .A(n4241), .ZN(n3213) );
  NOR2_X1 U3769 ( .A1(n3213), .A2(n4282), .ZN(n2940) );
  OAI22_X1 U3770 ( .A1(n3874), .A2(n2940), .B1(n2965), .B2(n4573), .ZN(n4541)
         );
  AOI211_X1 U3771 ( .C1(n2941), .C2(n4545), .A(n4543), .B(n4541), .ZN(n4564)
         );
  NAND2_X1 U3772 ( .A1(n4602), .A2(REG1_REG_0__SCAN_IN), .ZN(n2942) );
  OAI21_X1 U3773 ( .B1(n4564), .B2(n4602), .A(n2942), .ZN(U3518) );
  INV_X1 U3774 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4892) );
  NAND2_X1 U3775 ( .A1(n4162), .A2(U4043), .ZN(n2943) );
  OAI21_X1 U3776 ( .B1(U4043), .B2(n4892), .A(n2943), .ZN(U3573) );
  INV_X1 U3777 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n2950) );
  INV_X1 U3778 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4386) );
  NAND2_X1 U3779 ( .A1(n2944), .A2(REG1_REG_31__SCAN_IN), .ZN(n2947) );
  NAND2_X1 U3780 ( .A1(n2945), .A2(REG2_REG_31__SCAN_IN), .ZN(n2946) );
  OAI211_X1 U3781 ( .C1(n2948), .C2(n4386), .A(n2947), .B(n2946), .ZN(n4295)
         );
  NAND2_X1 U3782 ( .A1(n4295), .A2(U4043), .ZN(n2949) );
  OAI21_X1 U3783 ( .B1(U4043), .B2(n2950), .A(n2949), .ZN(U3581) );
  INV_X1 U3784 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4902) );
  NAND2_X1 U3785 ( .A1(n3846), .A2(U4043), .ZN(n2951) );
  OAI21_X1 U3786 ( .B1(U4043), .B2(n4902), .A(n2951), .ZN(U3580) );
  INV_X1 U3787 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U3788 ( .A1(n3594), .A2(U4043), .ZN(n2952) );
  OAI21_X1 U3789 ( .B1(U4043), .B2(n4885), .A(n2952), .ZN(U3563) );
  INV_X1 U3790 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4886) );
  NAND2_X1 U3791 ( .A1(n3811), .A2(U4043), .ZN(n2953) );
  OAI21_X1 U3792 ( .B1(U4043), .B2(n4886), .A(n2953), .ZN(U3564) );
  INV_X1 U3793 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4883) );
  NAND2_X1 U3794 ( .A1(n3164), .A2(U4043), .ZN(n2954) );
  OAI21_X1 U3795 ( .B1(U4043), .B2(n4883), .A(n2954), .ZN(U3555) );
  INV_X1 U3796 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U3797 ( .A1(n3502), .A2(U4043), .ZN(n2955) );
  OAI21_X1 U3798 ( .B1(U4043), .B2(n4880), .A(n2955), .ZN(U3562) );
  INV_X1 U3799 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U3800 ( .A1(n3711), .A2(U4043), .ZN(n2956) );
  OAI21_X1 U3801 ( .B1(U4043), .B2(n4884), .A(n2956), .ZN(U3552) );
  INV_X1 U3802 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4878) );
  NAND2_X1 U3803 ( .A1(n3005), .A2(U4043), .ZN(n2957) );
  OAI21_X1 U3804 ( .B1(U4043), .B2(n4878), .A(n2957), .ZN(U3551) );
  INV_X1 U3805 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4893) );
  NAND2_X1 U3806 ( .A1(n4925), .A2(U4043), .ZN(n2958) );
  OAI21_X1 U3807 ( .B1(U4043), .B2(n4893), .A(n2958), .ZN(U3570) );
  INV_X1 U3808 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4640) );
  NAND2_X1 U3809 ( .A1(n4165), .A2(U4043), .ZN(n2959) );
  OAI21_X1 U3810 ( .B1(U4043), .B2(n4640), .A(n2959), .ZN(U3575) );
  INV_X1 U3811 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4901) );
  NAND2_X1 U3812 ( .A1(n4098), .A2(U4043), .ZN(n2960) );
  OAI21_X1 U3813 ( .B1(U4043), .B2(n4901), .A(n2960), .ZN(U3579) );
  INV_X1 U3814 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4899) );
  NAND2_X1 U3815 ( .A1(n4129), .A2(U4043), .ZN(n2961) );
  OAI21_X1 U3816 ( .B1(U4043), .B2(n4899), .A(n2961), .ZN(U3577) );
  INV_X1 U3817 ( .A(n3514), .ZN(n3676) );
  OAI22_X1 U3818 ( .A1(n2964), .A2(n3676), .B1(n3056), .B2(n3675), .ZN(n2963)
         );
  XNOR2_X1 U3819 ( .A(n2963), .B(n3656), .ZN(n3024) );
  INV_X2 U3820 ( .A(n3514), .ZN(n3516) );
  OAI22_X1 U3821 ( .A1(n2964), .A2(n2967), .B1(n3056), .B2(n3516), .ZN(n3023)
         );
  XNOR2_X1 U3822 ( .A(n3024), .B(n3023), .ZN(n2977) );
  OAI22_X1 U3823 ( .A1(n2965), .A2(n3676), .B1(n2236), .B2(n3675), .ZN(n2966)
         );
  XNOR2_X1 U3824 ( .A(n2966), .B(n3656), .ZN(n2973) );
  XNOR2_X1 U3825 ( .A(n2973), .B(n2975), .ZN(n3707) );
  INV_X1 U3826 ( .A(n2970), .ZN(n2972) );
  OAI21_X1 U3827 ( .B1(n2972), .B2(n3656), .A(n2971), .ZN(n3709) );
  NAND2_X1 U3828 ( .A1(n3707), .A2(n3709), .ZN(n3708) );
  INV_X1 U3829 ( .A(n2973), .ZN(n2974) );
  OR2_X1 U3830 ( .A1(n2975), .A2(n2974), .ZN(n2976) );
  NAND2_X1 U3831 ( .A1(n3708), .A2(n2976), .ZN(n2978) );
  AOI22_X1 U3832 ( .A1(n3813), .A2(n4580), .B1(REG3_REG_2__SCAN_IN), .B2(n3710), .ZN(n2983) );
  AOI22_X1 U3833 ( .A1(n3812), .A2(n3005), .B1(n3801), .B2(n2981), .ZN(n2982)
         );
  OAI211_X1 U3834 ( .C1(n2984), .C2(n3806), .A(n2983), .B(n2982), .ZN(U3234)
         );
  AOI21_X1 U3835 ( .B1(n2985), .B2(n3712), .A(n3007), .ZN(n3052) );
  NAND2_X1 U3836 ( .A1(n2999), .A2(n2986), .ZN(n2990) );
  NAND2_X1 U3837 ( .A1(n2936), .A2(n4581), .ZN(n2988) );
  NAND2_X1 U3838 ( .A1(n3711), .A2(n4363), .ZN(n2987) );
  OAI211_X1 U3839 ( .C1(n4571), .C2(n2236), .A(n2988), .B(n2987), .ZN(n2989)
         );
  AOI21_X1 U3840 ( .B1(n2990), .B2(n4282), .A(n2989), .ZN(n2995) );
  AND2_X1 U3841 ( .A1(n2993), .A2(n2992), .ZN(n2996) );
  NAND2_X1 U3842 ( .A1(n2996), .A2(n3213), .ZN(n2994) );
  NAND2_X1 U3843 ( .A1(n2995), .A2(n2994), .ZN(n3049) );
  INV_X1 U3844 ( .A(n2996), .ZN(n3048) );
  NOR2_X1 U3845 ( .A1(n3048), .A2(n4353), .ZN(n2997) );
  AOI211_X1 U3846 ( .C1(n4584), .C2(n3052), .A(n3049), .B(n2997), .ZN(n4566)
         );
  NAND2_X1 U3847 ( .A1(n4602), .A2(REG1_REG_1__SCAN_IN), .ZN(n2998) );
  OAI21_X1 U3848 ( .B1(n4566), .B2(n4602), .A(n2998), .ZN(U3519) );
  OAI21_X1 U3849 ( .B1(n2146), .B2(n2719), .A(n3063), .ZN(n3003) );
  INV_X1 U3850 ( .A(n3003), .ZN(n3061) );
  NAND3_X1 U3851 ( .A1(n2719), .A2(n3912), .A3(n2999), .ZN(n3000) );
  AOI21_X1 U3852 ( .B1(n3001), .B2(n3000), .A(n4576), .ZN(n3002) );
  AOI21_X1 U3853 ( .B1(n3003), .B2(n3213), .A(n3002), .ZN(n3054) );
  OAI22_X1 U3854 ( .A1(n3055), .A2(n4573), .B1(n3056), .B2(n4571), .ZN(n3004)
         );
  AOI21_X1 U3855 ( .B1(n4581), .B2(n3005), .A(n3004), .ZN(n3006) );
  OAI211_X1 U3856 ( .C1(n3061), .C2(n4353), .A(n3054), .B(n3006), .ZN(n4569)
         );
  INV_X1 U3857 ( .A(n4569), .ZN(n3010) );
  OR2_X1 U3858 ( .A1(n3007), .A2(n3056), .ZN(n3008) );
  AOI22_X1 U3859 ( .A1(n3310), .A2(n4567), .B1(REG1_REG_2__SCAN_IN), .B2(n4602), .ZN(n3009) );
  OAI21_X1 U3860 ( .B1(n3010), .B2(n4602), .A(n3009), .ZN(U3520) );
  OAI21_X1 U3861 ( .B1(n3011), .B2(REG1_REG_7__SCAN_IN), .A(n4432), .ZN(n3012)
         );
  OAI21_X1 U3862 ( .B1(n3013), .B2(n4793), .A(n3012), .ZN(n3240) );
  XNOR2_X1 U3863 ( .A(n3240), .B(n3258), .ZN(n3242) );
  XNOR2_X1 U3864 ( .A(n3242), .B(REG1_REG_8__SCAN_IN), .ZN(n3020) );
  AOI21_X1 U3865 ( .B1(n4432), .B2(REG2_REG_7__SCAN_IN), .A(n3014), .ZN(n3259)
         );
  XNOR2_X1 U3866 ( .A(REG2_REG_8__SCAN_IN), .B(n3260), .ZN(n3015) );
  NAND2_X1 U3867 ( .A1(n4480), .A2(n3015), .ZN(n3016) );
  NAND2_X1 U3868 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3540) );
  NAND2_X1 U3869 ( .A1(n3016), .A2(n3540), .ZN(n3018) );
  NOR2_X1 U3870 ( .A1(n4530), .A2(n3258), .ZN(n3017) );
  AOI211_X1 U3871 ( .C1(n4523), .C2(ADDR_REG_8__SCAN_IN), .A(n3018), .B(n3017), 
        .ZN(n3019) );
  OAI21_X1 U3872 ( .B1(n3020), .B2(n4068), .A(n3019), .ZN(U3248) );
  INV_X1 U3873 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n4898) );
  NAND2_X1 U3874 ( .A1(n4120), .A2(U4043), .ZN(n3021) );
  OAI21_X1 U3875 ( .B1(U4043), .B2(n4898), .A(n3021), .ZN(U3578) );
  INV_X1 U3876 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4896) );
  NAND2_X1 U3877 ( .A1(n4308), .A2(U4043), .ZN(n3022) );
  OAI21_X1 U3878 ( .B1(U4043), .B2(n4896), .A(n3022), .ZN(U3576) );
  INV_X1 U3879 ( .A(n3023), .ZN(n3026) );
  INV_X1 U3880 ( .A(n3024), .ZN(n3025) );
  NAND2_X1 U3881 ( .A1(n4580), .A2(n3514), .ZN(n3029) );
  NAND2_X1 U3882 ( .A1(n3092), .A2(n3620), .ZN(n3028) );
  NAND2_X1 U3883 ( .A1(n3029), .A2(n3028), .ZN(n3030) );
  XNOR2_X1 U3884 ( .A(n3030), .B(n3656), .ZN(n3079) );
  OAI22_X1 U3885 ( .A1(n3055), .A2(n2967), .B1(n3065), .B2(n3516), .ZN(n3078)
         );
  XNOR2_X1 U3886 ( .A(n3079), .B(n3078), .ZN(n3081) );
  XOR2_X1 U3887 ( .A(n2156), .B(n3081), .Z(n3039) );
  INV_X1 U3888 ( .A(n3812), .ZN(n3798) );
  INV_X1 U3889 ( .A(n3813), .ZN(n3779) );
  OAI22_X1 U3890 ( .A1(n2964), .A2(n3798), .B1(n3779), .B2(n3115), .ZN(n3037)
         );
  INV_X1 U3891 ( .A(n3031), .ZN(n3033) );
  NAND4_X1 U3892 ( .A1(n3034), .A2(n3033), .A3(n3032), .A4(n2891), .ZN(n3035)
         );
  NAND2_X1 U3893 ( .A1(n3035), .A2(STATE_REG_SCAN_IN), .ZN(n3817) );
  INV_X1 U3894 ( .A(n3817), .ZN(n3781) );
  MUX2_X1 U3895 ( .A(n3781), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n3036) );
  AOI211_X1 U3896 ( .C1(n3092), .C2(n3801), .A(n3037), .B(n3036), .ZN(n3038)
         );
  OAI21_X1 U3897 ( .B1(n3039), .B2(n3806), .A(n3038), .ZN(U3215) );
  NAND4_X1 U3898 ( .A1(n3043), .A2(n3042), .A3(n2915), .A4(n3041), .ZN(n3044)
         );
  NAND2_X1 U3899 ( .A1(n2143), .A2(n4081), .ZN(n4289) );
  OR2_X1 U3900 ( .A1(n3045), .A2(n4081), .ZN(n3089) );
  INV_X1 U3901 ( .A(n3089), .ZN(n3046) );
  AND2_X1 U3902 ( .A1(n2143), .A2(n3046), .ZN(n4544) );
  INV_X1 U3903 ( .A(n4544), .ZN(n3329) );
  INV_X1 U3904 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3047) );
  OAI22_X1 U3905 ( .A1(n3048), .A2(n3329), .B1(n3047), .B2(n4531), .ZN(n3051)
         );
  MUX2_X1 U3906 ( .A(n3049), .B(REG2_REG_1__SCAN_IN), .S(n4661), .Z(n3050) );
  AOI211_X1 U3907 ( .C1(n4536), .C2(n3052), .A(n3051), .B(n3050), .ZN(n3053)
         );
  INV_X1 U3908 ( .A(n3053), .ZN(U3289) );
  MUX2_X1 U3909 ( .A(n4017), .B(n3054), .S(n2143), .Z(n3060) );
  INV_X1 U3910 ( .A(n4146), .ZN(n4228) );
  OAI22_X1 U3911 ( .A1(n4228), .A2(n3055), .B1(n2460), .B2(n4531), .ZN(n3058)
         );
  INV_X1 U3912 ( .A(n4222), .ZN(n3336) );
  NAND2_X1 U3913 ( .A1(n2143), .A2(n4581), .ZN(n4150) );
  OAI22_X1 U3914 ( .A1(n3336), .A2(n3056), .B1(n2965), .B2(n4150), .ZN(n3057)
         );
  AOI211_X1 U3915 ( .C1(n4536), .C2(n4567), .A(n3058), .B(n3057), .ZN(n3059)
         );
  OAI211_X1 U3916 ( .C1(n3061), .C2(n3329), .A(n3060), .B(n3059), .ZN(U3288)
         );
  NAND2_X1 U3917 ( .A1(n3063), .A2(n3062), .ZN(n3064) );
  XOR2_X1 U3918 ( .A(n3879), .B(n3064), .Z(n3090) );
  OAI22_X1 U3919 ( .A1(n3115), .A2(n4573), .B1(n4571), .B2(n3065), .ZN(n3070)
         );
  OAI21_X1 U3920 ( .B1(n3879), .B2(n3067), .A(n3066), .ZN(n3068) );
  AOI22_X1 U3921 ( .A1(n3068), .A2(n4282), .B1(n4581), .B2(n3711), .ZN(n3069)
         );
  INV_X1 U3922 ( .A(n3069), .ZN(n3097) );
  AOI211_X1 U3923 ( .C1(n4593), .C2(n3090), .A(n3070), .B(n3097), .ZN(n3074)
         );
  INV_X1 U3924 ( .A(n4423), .ZN(n4568) );
  AND2_X1 U3925 ( .A1(n4583), .A2(n3071), .ZN(n3093) );
  AOI22_X1 U3926 ( .A1(n4568), .A2(n3093), .B1(REG0_REG_3__SCAN_IN), .B2(n4598), .ZN(n3072) );
  OAI21_X1 U3927 ( .B1(n3074), .B2(n4598), .A(n3072), .ZN(U3473) );
  AOI22_X1 U3928 ( .A1(n3310), .A2(n3093), .B1(REG1_REG_3__SCAN_IN), .B2(n4602), .ZN(n3073) );
  OAI21_X1 U3929 ( .B1(n3074), .B2(n4602), .A(n3073), .ZN(U3521) );
  AND2_X1 U3930 ( .A1(n4582), .A2(n3514), .ZN(n3075) );
  AOI21_X1 U3931 ( .B1(n4001), .B2(n3670), .A(n3075), .ZN(n3122) );
  NAND2_X1 U3932 ( .A1(n4582), .A2(n3620), .ZN(n3076) );
  XNOR2_X1 U3933 ( .A(n3077), .B(n3656), .ZN(n3124) );
  XOR2_X1 U3934 ( .A(n3122), .B(n3124), .Z(n3083) );
  NOR2_X1 U3935 ( .A1(n3082), .A2(n3083), .ZN(n3125) );
  AOI211_X1 U3936 ( .C1(n3083), .C2(n3082), .A(n3806), .B(n3125), .ZN(n3088)
         );
  INV_X1 U3937 ( .A(n4662), .ZN(n3086) );
  AOI22_X1 U3938 ( .A1(n3812), .A2(n4580), .B1(n3801), .B2(n4582), .ZN(n3085)
         );
  AOI21_X1 U3939 ( .B1(n3813), .B2(n3164), .A(n4609), .ZN(n3084) );
  OAI211_X1 U3940 ( .C1(n3817), .C2(n3086), .A(n3085), .B(n3084), .ZN(n3087)
         );
  OR2_X1 U3941 ( .A1(n3088), .A2(n3087), .ZN(U3227) );
  NAND2_X1 U3942 ( .A1(n4241), .A2(n3089), .ZN(n4658) );
  INV_X1 U3943 ( .A(n3090), .ZN(n3099) );
  INV_X1 U3944 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4033) );
  OAI22_X1 U3945 ( .A1(n2143), .A2(n4033), .B1(REG3_REG_3__SCAN_IN), .B2(n4531), .ZN(n3091) );
  AOI21_X1 U3946 ( .B1(n3092), .B2(n4222), .A(n3091), .ZN(n3095) );
  NAND2_X1 U3947 ( .A1(n4536), .A2(n3093), .ZN(n3094) );
  OAI211_X1 U3948 ( .C1(n3115), .C2(n4228), .A(n3095), .B(n3094), .ZN(n3096)
         );
  AOI21_X1 U3949 ( .B1(n3097), .B2(n2143), .A(n3096), .ZN(n3098) );
  OAI21_X1 U3950 ( .B1(n4293), .B2(n3099), .A(n3098), .ZN(U3287) );
  INV_X1 U3951 ( .A(n3100), .ZN(n3921) );
  AND2_X1 U3952 ( .A1(n3921), .A2(n3934), .ZN(n3882) );
  XNOR2_X1 U3953 ( .A(n3101), .B(n3882), .ZN(n3117) );
  XOR2_X1 U3954 ( .A(n3882), .B(n3102), .Z(n3103) );
  NAND2_X1 U3955 ( .A1(n3103), .A2(n4282), .ZN(n3114) );
  INV_X1 U3956 ( .A(n3104), .ZN(n3134) );
  OAI22_X1 U3957 ( .A1(n2143), .A2(n4823), .B1(n3134), .B2(n4531), .ZN(n3106)
         );
  OAI22_X1 U3958 ( .A1(n3336), .A2(n3127), .B1(n3115), .B2(n4150), .ZN(n3105)
         );
  AOI211_X1 U3959 ( .C1(n4146), .C2(n4000), .A(n3106), .B(n3105), .ZN(n3110)
         );
  INV_X1 U3960 ( .A(n4586), .ZN(n3108) );
  INV_X1 U3961 ( .A(n3142), .ZN(n3107) );
  AOI21_X1 U3962 ( .B1(n3130), .B2(n3108), .A(n3107), .ZN(n3119) );
  NAND2_X1 U3963 ( .A1(n3119), .A2(n4536), .ZN(n3109) );
  OAI211_X1 U3964 ( .C1(n3114), .C2(n4661), .A(n3110), .B(n3109), .ZN(n3111)
         );
  AOI21_X1 U3965 ( .B1(n4220), .B2(n3117), .A(n3111), .ZN(n3112) );
  INV_X1 U3966 ( .A(n3112), .ZN(U3285) );
  AOI22_X1 U3967 ( .A1(n4000), .A2(n4363), .B1(n4362), .B2(n3130), .ZN(n3113)
         );
  OAI211_X1 U3968 ( .C1(n3115), .C2(n4367), .A(n3114), .B(n3113), .ZN(n3116)
         );
  AOI21_X1 U3969 ( .B1(n3117), .B2(n4593), .A(n3116), .ZN(n3121) );
  AOI22_X1 U3970 ( .A1(n3119), .A2(n3310), .B1(REG1_REG_5__SCAN_IN), .B2(n4602), .ZN(n3118) );
  OAI21_X1 U3971 ( .B1(n3121), .B2(n4602), .A(n3118), .ZN(U3523) );
  AOI22_X1 U3972 ( .A1(n3119), .A2(n4568), .B1(REG0_REG_5__SCAN_IN), .B2(n4598), .ZN(n3120) );
  OAI21_X1 U3973 ( .B1(n3121), .B2(n4598), .A(n3120), .ZN(U3477) );
  INV_X1 U3974 ( .A(n3122), .ZN(n3123) );
  OAI22_X1 U3975 ( .A1(n4574), .A2(n3676), .B1(n3127), .B2(n3675), .ZN(n3126)
         );
  XNOR2_X1 U3976 ( .A(n3126), .B(n3656), .ZN(n3157) );
  OAI22_X1 U3977 ( .A1(n4574), .A2(n2967), .B1(n3127), .B2(n3516), .ZN(n3156)
         );
  XNOR2_X1 U3978 ( .A(n3157), .B(n3156), .ZN(n3128) );
  AOI211_X1 U3979 ( .C1(n3129), .C2(n3128), .A(n3806), .B(n3158), .ZN(n3136)
         );
  AOI22_X1 U3980 ( .A1(n3812), .A2(n4001), .B1(n3801), .B2(n3130), .ZN(n3133)
         );
  AOI21_X1 U3981 ( .B1(n3813), .B2(n4000), .A(n3131), .ZN(n3132) );
  OAI211_X1 U3982 ( .C1(n3817), .C2(n3134), .A(n3133), .B(n3132), .ZN(n3135)
         );
  OR2_X1 U3983 ( .A1(n3136), .A2(n3135), .ZN(U3224) );
  AND2_X1 U3984 ( .A1(n3924), .A2(n3936), .ZN(n3883) );
  XNOR2_X1 U3985 ( .A(n3137), .B(n3883), .ZN(n3151) );
  XOR2_X1 U3986 ( .A(n3883), .B(n3138), .Z(n3149) );
  NAND2_X1 U3987 ( .A1(n2143), .A2(n4282), .ZN(n3341) );
  INV_X1 U3988 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3139) );
  OAI22_X1 U3989 ( .A1(n2143), .A2(n3139), .B1(n3167), .B2(n4531), .ZN(n3141)
         );
  OAI22_X1 U3990 ( .A1(n4228), .A2(n3230), .B1(n4574), .B2(n4150), .ZN(n3140)
         );
  AOI211_X1 U3991 ( .C1(n3163), .C2(n4222), .A(n3141), .B(n3140), .ZN(n3144)
         );
  AOI21_X1 U3992 ( .B1(n3163), .B2(n3142), .A(n2331), .ZN(n3153) );
  NAND2_X1 U3993 ( .A1(n3153), .A2(n4536), .ZN(n3143) );
  OAI211_X1 U3994 ( .C1(n3149), .C2(n3341), .A(n3144), .B(n3143), .ZN(n3145)
         );
  AOI21_X1 U3995 ( .B1(n3151), .B2(n4220), .A(n3145), .ZN(n3146) );
  INV_X1 U3996 ( .A(n3146), .ZN(U3284) );
  OAI22_X1 U3997 ( .A1(n3230), .A2(n4573), .B1(n4571), .B2(n3159), .ZN(n3147)
         );
  AOI21_X1 U3998 ( .B1(n4581), .B2(n3164), .A(n3147), .ZN(n3148) );
  OAI21_X1 U3999 ( .B1(n3149), .B2(n4576), .A(n3148), .ZN(n3150) );
  AOI21_X1 U4000 ( .B1(n3151), .B2(n4593), .A(n3150), .ZN(n3155) );
  AOI22_X1 U4001 ( .A1(n3153), .A2(n3310), .B1(n4602), .B2(REG1_REG_6__SCAN_IN), .ZN(n3152) );
  OAI21_X1 U4002 ( .B1(n3155), .B2(n4602), .A(n3152), .ZN(U3524) );
  AOI22_X1 U4003 ( .A1(n3153), .A2(n4568), .B1(n4598), .B2(REG0_REG_6__SCAN_IN), .ZN(n3154) );
  OAI21_X1 U4004 ( .B1(n3155), .B2(n4598), .A(n3154), .ZN(U3479) );
  OAI22_X1 U4005 ( .A1(n3160), .A2(n3676), .B1(n3159), .B2(n3675), .ZN(n3161)
         );
  XOR2_X1 U4006 ( .A(n3656), .B(n3161), .Z(n3225) );
  AOI22_X1 U4007 ( .A1(n4000), .A2(n3670), .B1(n3163), .B2(n3659), .ZN(n3226)
         );
  XNOR2_X1 U4008 ( .A(n3225), .B(n3226), .ZN(n3162) );
  XNOR2_X1 U4009 ( .A(n2182), .B(n3162), .ZN(n3171) );
  AOI22_X1 U4010 ( .A1(n3812), .A2(n3164), .B1(n3801), .B2(n3163), .ZN(n3170)
         );
  NAND2_X1 U4011 ( .A1(n3813), .A2(n3537), .ZN(n3165) );
  OAI211_X1 U4012 ( .C1(n3817), .C2(n3167), .A(n3166), .B(n3165), .ZN(n3168)
         );
  INV_X1 U4013 ( .A(n3168), .ZN(n3169) );
  OAI211_X1 U4014 ( .C1(n3171), .C2(n3806), .A(n3170), .B(n3169), .ZN(U3236)
         );
  OAI22_X1 U4015 ( .A1(n3289), .A2(n4573), .B1(n3229), .B2(n4571), .ZN(n3175)
         );
  XOR2_X1 U4016 ( .A(n3925), .B(n3172), .Z(n3173) );
  NOR2_X1 U4017 ( .A1(n3173), .A2(n4576), .ZN(n3174) );
  AOI211_X1 U4018 ( .C1(n4581), .C2(n4000), .A(n3175), .B(n3174), .ZN(n4597)
         );
  AOI21_X1 U4019 ( .B1(n3176), .B2(n3232), .A(n4375), .ZN(n3177) );
  NAND2_X1 U4020 ( .A1(n3177), .A2(n3215), .ZN(n4596) );
  INV_X1 U4021 ( .A(n4596), .ZN(n3182) );
  INV_X1 U4022 ( .A(n4289), .ZN(n3181) );
  INV_X1 U4023 ( .A(n3178), .ZN(n3236) );
  OAI22_X1 U4024 ( .A1(n2143), .A2(n3179), .B1(n3236), .B2(n4531), .ZN(n3180)
         );
  AOI21_X1 U4025 ( .B1(n3182), .B2(n3181), .A(n3180), .ZN(n3186) );
  NAND2_X1 U4026 ( .A1(n3184), .A2(n3925), .ZN(n4594) );
  NAND3_X1 U4027 ( .A1(n3183), .A2(n4594), .A3(n4220), .ZN(n3185) );
  OAI211_X1 U4028 ( .C1(n4597), .C2(n4661), .A(n3186), .B(n3185), .ZN(U3283)
         );
  INV_X1 U4029 ( .A(n3932), .ZN(n3937) );
  AND2_X1 U4030 ( .A1(n3937), .A2(n3930), .ZN(n3885) );
  INV_X1 U4031 ( .A(n3885), .ZN(n3187) );
  XNOR2_X1 U4032 ( .A(n3188), .B(n3187), .ZN(n3189) );
  NAND2_X1 U4033 ( .A1(n3189), .A2(n4282), .ZN(n3273) );
  XNOR2_X1 U4034 ( .A(n3190), .B(n3885), .ZN(n3271) );
  NAND2_X1 U4035 ( .A1(n3271), .A2(n4220), .ZN(n3196) );
  OAI21_X1 U4036 ( .B1(n3217), .B2(n3292), .A(n3199), .ZN(n3281) );
  INV_X1 U4037 ( .A(n3281), .ZN(n3194) );
  INV_X1 U4038 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4825) );
  OAI22_X1 U4039 ( .A1(n3299), .A2(n4531), .B1(n4825), .B2(n2143), .ZN(n3193)
         );
  AOI22_X1 U4040 ( .A1(n4223), .A2(n3999), .B1(n4146), .B2(n3997), .ZN(n3191)
         );
  OAI21_X1 U4041 ( .B1(n3292), .B2(n3336), .A(n3191), .ZN(n3192) );
  AOI211_X1 U4042 ( .C1(n3194), .C2(n4536), .A(n3193), .B(n3192), .ZN(n3195)
         );
  OAI211_X1 U40430 ( .C1(n3273), .C2(n4661), .A(n3196), .B(n3195), .ZN(U3281)
         );
  NAND2_X1 U4044 ( .A1(n3940), .A2(n3945), .ZN(n3865) );
  XNOR2_X1 U4045 ( .A(n3197), .B(n3865), .ZN(n3305) );
  XNOR2_X1 U4046 ( .A(n3198), .B(n3865), .ZN(n3307) );
  NAND2_X1 U4047 ( .A1(n3307), .A2(n4220), .ZN(n3206) );
  INV_X1 U4048 ( .A(n3199), .ZN(n3200) );
  OAI21_X1 U4049 ( .B1(n3200), .B2(n3605), .A(n3322), .ZN(n3314) );
  INV_X1 U4050 ( .A(n3314), .ZN(n3204) );
  AOI22_X1 U4051 ( .A1(n4223), .A2(n3998), .B1(n4146), .B2(n3996), .ZN(n3202)
         );
  INV_X1 U4052 ( .A(n4531), .ZN(n4663) );
  AOI22_X1 U4053 ( .A1(n4661), .A2(REG2_REG_10__SCAN_IN), .B1(n3610), .B2(
        n4663), .ZN(n3201) );
  OAI211_X1 U4054 ( .C1(n3605), .C2(n3336), .A(n3202), .B(n3201), .ZN(n3203)
         );
  AOI21_X1 U4055 ( .B1(n3204), .B2(n4536), .A(n3203), .ZN(n3205) );
  OAI211_X1 U4056 ( .C1(n3305), .C2(n3341), .A(n3206), .B(n3205), .ZN(U3280)
         );
  INV_X1 U4057 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3220) );
  AND2_X1 U4058 ( .A1(n3929), .A2(n3927), .ZN(n3884) );
  XNOR2_X1 U4059 ( .A(n3207), .B(n3884), .ZN(n4537) );
  INV_X1 U4060 ( .A(n4537), .ZN(n3214) );
  XNOR2_X1 U4061 ( .A(n3208), .B(n3884), .ZN(n3211) );
  OAI22_X1 U4062 ( .A1(n3230), .A2(n4367), .B1(n4571), .B2(n3288), .ZN(n3209)
         );
  AOI21_X1 U4063 ( .B1(n4363), .B2(n3998), .A(n3209), .ZN(n3210) );
  OAI21_X1 U4064 ( .B1(n3211), .B2(n4576), .A(n3210), .ZN(n3212) );
  AOI21_X1 U4065 ( .B1(n3213), .B2(n4537), .A(n3212), .ZN(n4540) );
  OAI21_X1 U4066 ( .B1(n4353), .B2(n3214), .A(n4540), .ZN(n3221) );
  NAND2_X1 U4067 ( .A1(n3221), .A2(n4600), .ZN(n3219) );
  AND2_X1 U4068 ( .A1(n3215), .A2(n3536), .ZN(n3216) );
  NOR2_X1 U4069 ( .A1(n3217), .A2(n3216), .ZN(n4535) );
  NAND2_X1 U4070 ( .A1(n4535), .A2(n4568), .ZN(n3218) );
  OAI211_X1 U4071 ( .C1(n4600), .C2(n3220), .A(n3219), .B(n3218), .ZN(U3483)
         );
  INV_X1 U4072 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3224) );
  NAND2_X1 U4073 ( .A1(n3221), .A2(n4604), .ZN(n3223) );
  NAND2_X1 U4074 ( .A1(n4535), .A2(n3310), .ZN(n3222) );
  OAI211_X1 U4075 ( .C1(n4604), .C2(n3224), .A(n3223), .B(n3222), .ZN(U3526)
         );
  INV_X1 U4076 ( .A(n3226), .ZN(n3227) );
  AND2_X1 U4077 ( .A1(n3232), .A2(n3659), .ZN(n3228) );
  AOI21_X1 U4078 ( .B1(n3537), .B2(n3670), .A(n3228), .ZN(n3284) );
  OAI22_X1 U4079 ( .A1(n3230), .A2(n3516), .B1(n3675), .B2(n3229), .ZN(n3231)
         );
  XNOR2_X1 U4080 ( .A(n3231), .B(n3656), .ZN(n3282) );
  XOR2_X1 U4081 ( .A(n3284), .B(n3282), .Z(n3285) );
  XOR2_X1 U4082 ( .A(n3286), .B(n3285), .Z(n3238) );
  AOI22_X1 U4083 ( .A1(n3812), .A2(n4000), .B1(n3801), .B2(n3232), .ZN(n3235)
         );
  AOI21_X1 U4084 ( .B1(n3813), .B2(n3999), .A(n3233), .ZN(n3234) );
  OAI211_X1 U4085 ( .C1(n3817), .C2(n3236), .A(n3235), .B(n3234), .ZN(n3237)
         );
  AOI21_X1 U4086 ( .B1(n3238), .B2(n3819), .A(n3237), .ZN(n3239) );
  INV_X1 U4087 ( .A(n3239), .ZN(U3210) );
  NAND2_X1 U4088 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3256), .ZN(n3247) );
  INV_X1 U4089 ( .A(n3256), .ZN(n4560) );
  INV_X1 U4090 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4790) );
  AOI22_X1 U4091 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3256), .B1(n4560), .B2(
        n4790), .ZN(n4470) );
  NAND2_X1 U4092 ( .A1(n3257), .A2(REG1_REG_9__SCAN_IN), .ZN(n3244) );
  INV_X1 U4093 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4794) );
  INV_X1 U4094 ( .A(n3257), .ZN(n4563) );
  AOI22_X1 U4095 ( .A1(n3257), .A2(REG1_REG_9__SCAN_IN), .B1(n4794), .B2(n4563), .ZN(n4449) );
  INV_X1 U4096 ( .A(n3258), .ZN(n3241) );
  AOI22_X1 U4097 ( .A1(n3242), .A2(REG1_REG_8__SCAN_IN), .B1(n3241), .B2(n3240), .ZN(n3243) );
  INV_X1 U4098 ( .A(n3243), .ZN(n4448) );
  NAND2_X1 U4099 ( .A1(n4449), .A2(n4448), .ZN(n4447) );
  NAND2_X1 U4100 ( .A1(n3244), .A2(n4447), .ZN(n3245) );
  NAND2_X1 U4101 ( .A1(n4561), .A2(n3245), .ZN(n3246) );
  INV_X1 U4102 ( .A(n4561), .ZN(n4467) );
  XNOR2_X1 U4103 ( .A(n3245), .B(n4467), .ZN(n4464) );
  NAND2_X1 U4104 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4464), .ZN(n4463) );
  NAND2_X1 U4105 ( .A1(n3246), .A2(n4463), .ZN(n4469) );
  NAND2_X1 U4106 ( .A1(n4470), .A2(n4469), .ZN(n4468) );
  NAND2_X1 U4107 ( .A1(n3247), .A2(n4468), .ZN(n3248) );
  NAND2_X1 U4108 ( .A1(n3264), .A2(n3248), .ZN(n3249) );
  INV_X1 U4109 ( .A(n3264), .ZN(n4559) );
  XNOR2_X1 U4110 ( .A(n3248), .B(n4559), .ZN(n4486) );
  NAND2_X1 U4111 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4486), .ZN(n4485) );
  NAND2_X1 U4112 ( .A1(n3249), .A2(n4485), .ZN(n3251) );
  INV_X1 U4113 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4791) );
  NOR2_X1 U4114 ( .A1(n3255), .A2(n4791), .ZN(n4040) );
  AOI21_X1 U4115 ( .B1(n4791), .B2(n3255), .A(n4040), .ZN(n3250) );
  NAND2_X1 U4116 ( .A1(n3250), .A2(n3251), .ZN(n4041) );
  OAI211_X1 U4117 ( .C1(n3251), .C2(n3250), .A(n4525), .B(n4041), .ZN(n3253)
         );
  NOR2_X1 U4118 ( .A1(STATE_REG_SCAN_IN), .A2(n4623), .ZN(n3503) );
  AOI21_X1 U4119 ( .B1(n4523), .B2(ADDR_REG_13__SCAN_IN), .A(n3503), .ZN(n3252) );
  OAI211_X1 U4120 ( .C1(n4530), .C2(n3255), .A(n3253), .B(n3252), .ZN(n3270)
         );
  NOR2_X1 U4121 ( .A1(n3255), .A2(n2213), .ZN(n3254) );
  AOI21_X1 U4122 ( .B1(n2213), .B2(n3255), .A(n3254), .ZN(n3268) );
  NAND2_X1 U4123 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3256), .ZN(n3263) );
  INV_X1 U4124 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4125 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3256), .B1(n4560), .B2(
        n3321), .ZN(n4473) );
  AOI22_X1 U4126 ( .A1(n3257), .A2(REG2_REG_9__SCAN_IN), .B1(n4825), .B2(n4563), .ZN(n4452) );
  INV_X1 U4127 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4533) );
  NAND2_X1 U4128 ( .A1(n4561), .A2(n3261), .ZN(n3262) );
  XNOR2_X1 U4129 ( .A(n3261), .B(n4467), .ZN(n4459) );
  NAND2_X1 U4130 ( .A1(n3264), .A2(n3265), .ZN(n3266) );
  XNOR2_X1 U4131 ( .A(n3265), .B(n4559), .ZN(n4481) );
  OAI21_X1 U4132 ( .B1(n3268), .B2(n4051), .A(n4480), .ZN(n3267) );
  AOI21_X1 U4133 ( .B1(n3268), .B2(n4051), .A(n3267), .ZN(n3269) );
  OR2_X1 U4134 ( .A1(n3270), .A2(n3269), .ZN(U3253) );
  NAND2_X1 U4135 ( .A1(n3271), .A2(n4593), .ZN(n3275) );
  AOI22_X1 U4136 ( .A1(n3997), .A2(n4363), .B1(n4362), .B2(n3296), .ZN(n3274)
         );
  OR2_X1 U4137 ( .A1(n3289), .A2(n4367), .ZN(n3272) );
  NAND4_X1 U4138 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .ZN(n3278)
         );
  MUX2_X1 U4139 ( .A(REG0_REG_9__SCAN_IN), .B(n3278), .S(n4600), .Z(n3276) );
  INV_X1 U4140 ( .A(n3276), .ZN(n3277) );
  OAI21_X1 U4141 ( .B1(n3281), .B2(n4423), .A(n3277), .ZN(U3485) );
  MUX2_X1 U4142 ( .A(REG1_REG_9__SCAN_IN), .B(n3278), .S(n4604), .Z(n3279) );
  INV_X1 U4143 ( .A(n3279), .ZN(n3280) );
  OAI21_X1 U4144 ( .B1(n4372), .B2(n3281), .A(n3280), .ZN(U3527) );
  INV_X1 U4145 ( .A(n3282), .ZN(n3283) );
  OAI22_X1 U4146 ( .A1(n3289), .A2(n3516), .B1(n3675), .B2(n3288), .ZN(n3287)
         );
  XNOR2_X1 U4147 ( .A(n3287), .B(n3656), .ZN(n3291) );
  OAI22_X1 U4148 ( .A1(n3289), .A2(n2967), .B1(n3516), .B2(n3288), .ZN(n3290)
         );
  AND2_X1 U4149 ( .A1(n3291), .A2(n3290), .ZN(n3533) );
  OR2_X1 U4150 ( .A1(n3291), .A2(n3290), .ZN(n3532) );
  OAI22_X1 U4151 ( .A1(n3607), .A2(n2967), .B1(n3292), .B2(n3516), .ZN(n3381)
         );
  NAND2_X1 U4152 ( .A1(n3998), .A2(n3659), .ZN(n3294) );
  NAND2_X1 U4153 ( .A1(n3296), .A2(n3620), .ZN(n3293) );
  NAND2_X1 U4154 ( .A1(n3294), .A2(n3293), .ZN(n3295) );
  XNOR2_X1 U4155 ( .A(n3295), .B(n3656), .ZN(n3382) );
  XOR2_X1 U4156 ( .A(n3381), .B(n3382), .Z(n3384) );
  XNOR2_X1 U4157 ( .A(n3385), .B(n3384), .ZN(n3301) );
  AOI22_X1 U4158 ( .A1(n3812), .A2(n3999), .B1(n3801), .B2(n3296), .ZN(n3298)
         );
  NOR2_X1 U4159 ( .A1(STATE_REG_SCAN_IN), .A2(n4865), .ZN(n4456) );
  AOI21_X1 U4160 ( .B1(n3813), .B2(n3997), .A(n4456), .ZN(n3297) );
  OAI211_X1 U4161 ( .C1(n3817), .C2(n3299), .A(n3298), .B(n3297), .ZN(n3300)
         );
  AOI21_X1 U4162 ( .B1(n3301), .B2(n3819), .A(n3300), .ZN(n3302) );
  INV_X1 U4163 ( .A(n3302), .ZN(U3228) );
  INV_X1 U4164 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3308) );
  OAI22_X1 U4165 ( .A1(n3437), .A2(n4573), .B1(n4571), .B2(n3605), .ZN(n3303)
         );
  AOI21_X1 U4166 ( .B1(n4581), .B2(n3998), .A(n3303), .ZN(n3304) );
  OAI21_X1 U4167 ( .B1(n3305), .B2(n4576), .A(n3304), .ZN(n3306) );
  AOI21_X1 U4168 ( .B1(n4593), .B2(n3307), .A(n3306), .ZN(n3311) );
  MUX2_X1 U4169 ( .A(n3308), .B(n3311), .S(n4600), .Z(n3309) );
  OAI21_X1 U4170 ( .B1(n3314), .B2(n4423), .A(n3309), .ZN(U3487) );
  INV_X1 U4171 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3312) );
  MUX2_X1 U4172 ( .A(n3312), .B(n3311), .S(n4604), .Z(n3313) );
  OAI21_X1 U4173 ( .B1(n3314), .B2(n4372), .A(n3313), .ZN(U3528) );
  INV_X1 U4174 ( .A(n3356), .ZN(n3315) );
  AOI21_X1 U4175 ( .B1(n3875), .B2(n3316), .A(n3315), .ZN(n3373) );
  AOI22_X1 U4176 ( .A1(n3502), .A2(n4363), .B1(n3398), .B2(n4362), .ZN(n3319)
         );
  XNOR2_X1 U4177 ( .A(n3367), .B(n3875), .ZN(n3317) );
  NAND2_X1 U4178 ( .A1(n3317), .A2(n4282), .ZN(n3318) );
  OAI211_X1 U4179 ( .C1(n3373), .C2(n4241), .A(n3319), .B(n3318), .ZN(n3375)
         );
  NAND2_X1 U4180 ( .A1(n3375), .A2(n2143), .ZN(n3328) );
  INV_X1 U4181 ( .A(n3320), .ZN(n3401) );
  OAI22_X1 U4182 ( .A1(n2143), .A2(n3321), .B1(n3401), .B2(n4531), .ZN(n3326)
         );
  INV_X1 U4183 ( .A(n3322), .ZN(n3324) );
  INV_X1 U4184 ( .A(n3358), .ZN(n3323) );
  OAI21_X1 U4185 ( .B1(n3324), .B2(n3396), .A(n3323), .ZN(n3380) );
  NOR2_X1 U4186 ( .A1(n3380), .A2(n4443), .ZN(n3325) );
  AOI211_X1 U4187 ( .C1(n4223), .C2(n3997), .A(n3326), .B(n3325), .ZN(n3327)
         );
  OAI211_X1 U4188 ( .C1(n3373), .C2(n3329), .A(n3328), .B(n3327), .ZN(U3279)
         );
  XNOR2_X1 U4189 ( .A(n3828), .B(n3331), .ZN(n3428) );
  OAI21_X1 U4190 ( .B1(n3332), .B2(n3331), .A(n3330), .ZN(n3430) );
  NAND2_X1 U4191 ( .A1(n3430), .A2(n4220), .ZN(n3340) );
  INV_X1 U4192 ( .A(n3421), .ZN(n3333) );
  OAI21_X1 U4193 ( .B1(n3333), .B2(n3517), .A(n3346), .ZN(n3434) );
  INV_X1 U4194 ( .A(n3434), .ZN(n3338) );
  AOI22_X1 U4195 ( .A1(n4223), .A2(n3594), .B1(n4146), .B2(n4379), .ZN(n3335)
         );
  AOI22_X1 U4196 ( .A1(n4661), .A2(REG2_REG_14__SCAN_IN), .B1(n3524), .B2(
        n4663), .ZN(n3334) );
  OAI211_X1 U4197 ( .C1(n3517), .C2(n3336), .A(n3335), .B(n3334), .ZN(n3337)
         );
  AOI21_X1 U4198 ( .B1(n3338), .B2(n4536), .A(n3337), .ZN(n3339) );
  OAI211_X1 U4199 ( .C1(n3428), .C2(n3341), .A(n3340), .B(n3339), .ZN(U3276)
         );
  AOI21_X1 U4200 ( .B1(n3342), .B2(n3872), .A(n4576), .ZN(n3344) );
  NAND2_X1 U4201 ( .A1(n3344), .A2(n3343), .ZN(n3454) );
  XNOR2_X1 U4202 ( .A(n3345), .B(n3872), .ZN(n3456) );
  NAND2_X1 U4203 ( .A1(n3456), .A2(n4220), .ZN(n3354) );
  INV_X1 U4204 ( .A(n3346), .ZN(n3347) );
  OAI21_X1 U4205 ( .B1(n3347), .B2(n3557), .A(n2335), .ZN(n3462) );
  INV_X1 U4206 ( .A(n3462), .ZN(n3352) );
  AOI22_X1 U4207 ( .A1(n4223), .A2(n3811), .B1(n4222), .B2(n3810), .ZN(n3350)
         );
  AOI22_X1 U4208 ( .A1(n4661), .A2(REG2_REG_15__SCAN_IN), .B1(n3348), .B2(
        n4663), .ZN(n3349) );
  OAI211_X1 U4209 ( .C1(n4368), .C2(n4228), .A(n3350), .B(n3349), .ZN(n3351)
         );
  AOI21_X1 U4210 ( .B1(n3352), .B2(n4536), .A(n3351), .ZN(n3353) );
  OAI211_X1 U4211 ( .C1(n4661), .C2(n3454), .A(n3354), .B(n3353), .ZN(U3275)
         );
  NAND2_X1 U4212 ( .A1(n3356), .A2(n3355), .ZN(n3406) );
  NAND2_X1 U4213 ( .A1(n3412), .A2(n3410), .ZN(n3866) );
  XNOR2_X1 U4214 ( .A(n3406), .B(n3866), .ZN(n3439) );
  NOR2_X1 U4215 ( .A1(n3358), .A2(n3357), .ZN(n3359) );
  OR2_X1 U4216 ( .A1(n3419), .A2(n3359), .ZN(n3445) );
  INV_X1 U4217 ( .A(n3360), .ZN(n3596) );
  OAI22_X1 U4218 ( .A1(n2143), .A2(n2214), .B1(n3596), .B2(n4531), .ZN(n3361)
         );
  AOI21_X1 U4219 ( .B1(n4146), .B2(n3594), .A(n3361), .ZN(n3363) );
  AOI22_X1 U4220 ( .A1(n4223), .A2(n3996), .B1(n4222), .B2(n3593), .ZN(n3362)
         );
  OAI211_X1 U4221 ( .C1(n3445), .C2(n4443), .A(n3363), .B(n3362), .ZN(n3370)
         );
  INV_X1 U4222 ( .A(n3364), .ZN(n3365) );
  AOI21_X1 U4223 ( .B1(n3367), .B2(n3366), .A(n3365), .ZN(n3413) );
  XNOR2_X1 U4224 ( .A(n3413), .B(n3866), .ZN(n3368) );
  NAND2_X1 U4225 ( .A1(n3368), .A2(n4282), .ZN(n3436) );
  NOR2_X1 U4226 ( .A1(n3436), .A2(n4661), .ZN(n3369) );
  AOI211_X1 U4227 ( .C1(n4220), .C2(n3439), .A(n3370), .B(n3369), .ZN(n3371)
         );
  INV_X1 U4228 ( .A(n3371), .ZN(U3278) );
  OAI22_X1 U4229 ( .A1(n3373), .A2(n4353), .B1(n3372), .B2(n4367), .ZN(n3374)
         );
  NOR2_X1 U4230 ( .A1(n3375), .A2(n3374), .ZN(n3377) );
  MUX2_X1 U4231 ( .A(n4790), .B(n3377), .S(n4604), .Z(n3376) );
  OAI21_X1 U4232 ( .B1(n4372), .B2(n3380), .A(n3376), .ZN(U3529) );
  INV_X1 U4233 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3378) );
  MUX2_X1 U4234 ( .A(n3378), .B(n3377), .S(n4600), .Z(n3379) );
  OAI21_X1 U4235 ( .B1(n3380), .B2(n4423), .A(n3379), .ZN(U3489) );
  NOR2_X1 U4236 ( .A1(n3382), .A2(n3381), .ZN(n3383) );
  AOI21_X1 U4237 ( .B1(n3385), .B2(n3384), .A(n3383), .ZN(n3603) );
  NAND2_X1 U4238 ( .A1(n3997), .A2(n3659), .ZN(n3387) );
  NAND2_X1 U4239 ( .A1(n3389), .A2(n3620), .ZN(n3386) );
  NAND2_X1 U4240 ( .A1(n3387), .A2(n3386), .ZN(n3388) );
  XNOR2_X1 U4241 ( .A(n3388), .B(n3656), .ZN(n3393) );
  AND2_X1 U4242 ( .A1(n3389), .A2(n3659), .ZN(n3390) );
  AOI21_X1 U4243 ( .B1(n3997), .B2(n3670), .A(n3390), .ZN(n3391) );
  XNOR2_X1 U4244 ( .A(n3393), .B(n3391), .ZN(n3602) );
  NAND2_X1 U4245 ( .A1(n3603), .A2(n3602), .ZN(n3601) );
  INV_X1 U4246 ( .A(n3391), .ZN(n3392) );
  NAND2_X1 U4247 ( .A1(n3393), .A2(n3392), .ZN(n3394) );
  OAI22_X1 U4248 ( .A1(n3437), .A2(n3516), .B1(n3675), .B2(n3396), .ZN(n3395)
         );
  XNOR2_X1 U4249 ( .A(n3395), .B(n3656), .ZN(n3485) );
  OAI22_X1 U4250 ( .A1(n3437), .A2(n2967), .B1(n3516), .B2(n3396), .ZN(n3486)
         );
  XNOR2_X1 U4251 ( .A(n3485), .B(n3486), .ZN(n3397) );
  XNOR2_X1 U4252 ( .A(n3487), .B(n3397), .ZN(n3403) );
  AOI22_X1 U4253 ( .A1(n3812), .A2(n3997), .B1(n3801), .B2(n3398), .ZN(n3400)
         );
  AND2_X1 U4254 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4477) );
  AOI21_X1 U4255 ( .B1(n3813), .B2(n3502), .A(n4477), .ZN(n3399) );
  OAI211_X1 U4256 ( .C1(n3817), .C2(n3401), .A(n3400), .B(n3399), .ZN(n3402)
         );
  AOI21_X1 U4257 ( .B1(n3403), .B2(n3819), .A(n3402), .ZN(n3404) );
  INV_X1 U4258 ( .A(n3404), .ZN(U3233) );
  XNOR2_X1 U4259 ( .A(n3594), .B(n3501), .ZN(n3868) );
  NAND2_X1 U4260 ( .A1(n3406), .A2(n3405), .ZN(n3408) );
  NAND2_X1 U4261 ( .A1(n3408), .A2(n3407), .ZN(n3409) );
  XOR2_X1 U4262 ( .A(n3868), .B(n3409), .Z(n3447) );
  INV_X1 U4263 ( .A(n3447), .ZN(n3425) );
  INV_X1 U4264 ( .A(n3410), .ZN(n3411) );
  AOI21_X1 U4265 ( .B1(n3413), .B2(n3412), .A(n3411), .ZN(n3414) );
  XOR2_X1 U4266 ( .A(n3868), .B(n3414), .Z(n3417) );
  OAI22_X1 U4267 ( .A1(n3518), .A2(n4573), .B1(n4571), .B2(n3418), .ZN(n3415)
         );
  AOI21_X1 U4268 ( .B1(n4581), .B2(n3502), .A(n3415), .ZN(n3416) );
  OAI21_X1 U4269 ( .B1(n3417), .B2(n4576), .A(n3416), .ZN(n3446) );
  OR2_X1 U4270 ( .A1(n3419), .A2(n3418), .ZN(n3420) );
  NAND2_X1 U4271 ( .A1(n3421), .A2(n3420), .ZN(n3452) );
  AOI22_X1 U4272 ( .A1(n4661), .A2(REG2_REG_13__SCAN_IN), .B1(n3500), .B2(
        n4663), .ZN(n3422) );
  OAI21_X1 U4273 ( .B1(n3452), .B2(n4443), .A(n3422), .ZN(n3423) );
  AOI21_X1 U4274 ( .B1(n3446), .B2(n2143), .A(n3423), .ZN(n3424) );
  OAI21_X1 U4275 ( .B1(n3425), .B2(n4293), .A(n3424), .ZN(U3277) );
  OAI22_X1 U4276 ( .A1(n3558), .A2(n4573), .B1(n3517), .B2(n4571), .ZN(n3426)
         );
  AOI21_X1 U4277 ( .B1(n4581), .B2(n3594), .A(n3426), .ZN(n3427) );
  OAI21_X1 U4278 ( .B1(n3428), .B2(n4576), .A(n3427), .ZN(n3429) );
  AOI21_X1 U4279 ( .B1(n3430), .B2(n4593), .A(n3429), .ZN(n3432) );
  MUX2_X1 U4280 ( .A(n3432), .B(n4774), .S(n4598), .Z(n3431) );
  OAI21_X1 U4281 ( .B1(n3434), .B2(n4423), .A(n3431), .ZN(U3495) );
  INV_X1 U4282 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4806) );
  MUX2_X1 U4283 ( .A(n3432), .B(n4806), .S(n4602), .Z(n3433) );
  OAI21_X1 U4284 ( .B1(n4372), .B2(n3434), .A(n3433), .ZN(U3532) );
  INV_X1 U4285 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4286 ( .A1(n3594), .A2(n4363), .B1(n4362), .B2(n3593), .ZN(n3435)
         );
  OAI211_X1 U4287 ( .C1(n3437), .C2(n4367), .A(n3436), .B(n3435), .ZN(n3438)
         );
  AOI21_X1 U4288 ( .B1(n4593), .B2(n3439), .A(n3438), .ZN(n3442) );
  MUX2_X1 U4289 ( .A(n3440), .B(n3442), .S(n4600), .Z(n3441) );
  OAI21_X1 U4290 ( .B1(n3445), .B2(n4423), .A(n3441), .ZN(U3491) );
  INV_X1 U4291 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3443) );
  MUX2_X1 U4292 ( .A(n3443), .B(n3442), .S(n4604), .Z(n3444) );
  OAI21_X1 U4293 ( .B1(n4372), .B2(n3445), .A(n3444), .ZN(U3530) );
  INV_X1 U4294 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3448) );
  AOI21_X1 U4295 ( .B1(n4593), .B2(n3447), .A(n3446), .ZN(n3450) );
  MUX2_X1 U4296 ( .A(n3448), .B(n3450), .S(n4600), .Z(n3449) );
  OAI21_X1 U4297 ( .B1(n3452), .B2(n4423), .A(n3449), .ZN(U3493) );
  MUX2_X1 U4298 ( .A(n4791), .B(n3450), .S(n4604), .Z(n3451) );
  OAI21_X1 U4299 ( .B1(n4372), .B2(n3452), .A(n3451), .ZN(U3531) );
  AOI22_X1 U4300 ( .A1(n3995), .A2(n4363), .B1(n4362), .B2(n3810), .ZN(n3453)
         );
  OAI211_X1 U4301 ( .C1(n3518), .C2(n4367), .A(n3454), .B(n3453), .ZN(n3455)
         );
  AOI21_X1 U4302 ( .B1(n3456), .B2(n4593), .A(n3455), .ZN(n3460) );
  INV_X1 U4303 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3457) );
  MUX2_X1 U4304 ( .A(n3460), .B(n3457), .S(n4598), .Z(n3458) );
  OAI21_X1 U4305 ( .B1(n3462), .B2(n4423), .A(n3458), .ZN(U3497) );
  INV_X1 U4306 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3459) );
  MUX2_X1 U4307 ( .A(n3460), .B(n3459), .S(n4602), .Z(n3461) );
  OAI21_X1 U4308 ( .B1(n4372), .B2(n3462), .A(n3461), .ZN(U3533) );
  OAI21_X1 U4309 ( .B1(n3463), .B2(n2610), .A(n3464), .ZN(n4383) );
  OAI211_X1 U4310 ( .C1(n3466), .C2(n3873), .A(n3465), .B(n4282), .ZN(n4380)
         );
  INV_X1 U4311 ( .A(n4380), .ZN(n3473) );
  NOR2_X1 U4312 ( .A1(n3467), .A2(n4373), .ZN(n3468) );
  OR2_X1 U4313 ( .A1(n3478), .A2(n3468), .ZN(n4376) );
  NOR2_X1 U4314 ( .A1(n4376), .A2(n4443), .ZN(n3472) );
  AOI22_X1 U4315 ( .A1(n4223), .A2(n4379), .B1(n4222), .B2(n3738), .ZN(n3470)
         );
  AOI22_X1 U4316 ( .A1(n4661), .A2(REG2_REG_16__SCAN_IN), .B1(n3739), .B2(
        n4663), .ZN(n3469) );
  OAI211_X1 U4317 ( .C1(n4374), .C2(n4228), .A(n3470), .B(n3469), .ZN(n3471)
         );
  AOI211_X1 U4318 ( .C1(n3473), .C2(n2143), .A(n3472), .B(n3471), .ZN(n3474)
         );
  OAI21_X1 U4319 ( .B1(n4383), .B2(n4293), .A(n3474), .ZN(U3274) );
  INV_X1 U4320 ( .A(n4255), .ZN(n3475) );
  NAND2_X1 U4321 ( .A1(n3475), .A2(n4254), .ZN(n3901) );
  XNOR2_X1 U4322 ( .A(n4256), .B(n3901), .ZN(n3476) );
  NAND2_X1 U4323 ( .A1(n3476), .A2(n4282), .ZN(n4366) );
  XOR2_X1 U4324 ( .A(n3901), .B(n3477), .Z(n4370) );
  NAND2_X1 U4325 ( .A1(n4370), .A2(n4220), .ZN(n3484) );
  OAI21_X1 U4326 ( .B1(n3478), .B2(n3572), .A(n4285), .ZN(n4424) );
  INV_X1 U4327 ( .A(n4424), .ZN(n3482) );
  AOI22_X1 U4328 ( .A1(n4223), .A2(n3995), .B1(n4222), .B2(n4361), .ZN(n3480)
         );
  AOI22_X1 U4329 ( .A1(n4661), .A2(REG2_REG_17__SCAN_IN), .B1(n3750), .B2(
        n4663), .ZN(n3479) );
  OAI211_X1 U4330 ( .C1(n4265), .C2(n4228), .A(n3480), .B(n3479), .ZN(n3481)
         );
  AOI21_X1 U4331 ( .B1(n3482), .B2(n4536), .A(n3481), .ZN(n3483) );
  OAI211_X1 U4332 ( .C1(n4661), .C2(n4366), .A(n3484), .B(n3483), .ZN(U3273)
         );
  NAND2_X1 U4333 ( .A1(n3502), .A2(n3659), .ZN(n3489) );
  NAND2_X1 U4334 ( .A1(n3593), .A2(n3620), .ZN(n3488) );
  NAND2_X1 U4335 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  XNOR2_X1 U4336 ( .A(n3490), .B(n2150), .ZN(n3493) );
  AND2_X1 U4337 ( .A1(n3593), .A2(n3659), .ZN(n3491) );
  AOI21_X1 U4338 ( .B1(n3502), .B2(n3670), .A(n3491), .ZN(n3492) );
  NOR2_X1 U4339 ( .A1(n3493), .A2(n3492), .ZN(n3590) );
  NAND2_X1 U4340 ( .A1(n3493), .A2(n3492), .ZN(n3588) );
  NAND2_X1 U4341 ( .A1(n3594), .A2(n3659), .ZN(n3495) );
  NAND2_X1 U4342 ( .A1(n3501), .A2(n3620), .ZN(n3494) );
  NAND2_X1 U4343 ( .A1(n3495), .A2(n3494), .ZN(n3496) );
  XNOR2_X1 U4344 ( .A(n3496), .B(n2150), .ZN(n3551) );
  INV_X1 U4345 ( .A(n3551), .ZN(n3512) );
  NAND2_X1 U4346 ( .A1(n3594), .A2(n3670), .ZN(n3498) );
  NAND2_X1 U4347 ( .A1(n3501), .A2(n3659), .ZN(n3497) );
  XNOR2_X1 U4348 ( .A(n3512), .B(n3552), .ZN(n3499) );
  XNOR2_X1 U4349 ( .A(n3510), .B(n3499), .ZN(n3508) );
  INV_X1 U4350 ( .A(n3500), .ZN(n3506) );
  AOI22_X1 U4351 ( .A1(n3812), .A2(n3502), .B1(n3801), .B2(n3501), .ZN(n3505)
         );
  AOI21_X1 U4352 ( .B1(n3813), .B2(n3811), .A(n3503), .ZN(n3504) );
  OAI211_X1 U4353 ( .C1(n3817), .C2(n3506), .A(n3505), .B(n3504), .ZN(n3507)
         );
  AOI21_X1 U4354 ( .B1(n3508), .B2(n3819), .A(n3507), .ZN(n3509) );
  INV_X1 U4355 ( .A(n3509), .ZN(U3231) );
  INV_X1 U4356 ( .A(n3510), .ZN(n3513) );
  AOI21_X1 U4357 ( .B1(n3510), .B2(n3551), .A(n3552), .ZN(n3511) );
  AOI21_X1 U4358 ( .B1(n3513), .B2(n3512), .A(n3511), .ZN(n3522) );
  OAI22_X1 U4359 ( .A1(n3518), .A2(n3516), .B1(n3517), .B2(n3675), .ZN(n3515)
         );
  XNOR2_X1 U4360 ( .A(n3515), .B(n3656), .ZN(n3520) );
  OAI22_X1 U4361 ( .A1(n3518), .A2(n2967), .B1(n3517), .B2(n3516), .ZN(n3519)
         );
  NAND2_X1 U4362 ( .A1(n3520), .A2(n3519), .ZN(n3553) );
  OR2_X1 U4363 ( .A1(n3520), .A2(n3519), .ZN(n3554) );
  NAND2_X1 U4364 ( .A1(n3553), .A2(n3554), .ZN(n3521) );
  XNOR2_X1 U4365 ( .A(n3522), .B(n3521), .ZN(n3530) );
  AOI22_X1 U4366 ( .A1(n3812), .A2(n3594), .B1(n3801), .B2(n3523), .ZN(n3529)
         );
  INV_X1 U4367 ( .A(n3524), .ZN(n3526) );
  NAND2_X1 U4368 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4489) );
  NAND2_X1 U4369 ( .A1(n3813), .A2(n4379), .ZN(n3525) );
  OAI211_X1 U4370 ( .C1(n3817), .C2(n3526), .A(n4489), .B(n3525), .ZN(n3527)
         );
  INV_X1 U4371 ( .A(n3527), .ZN(n3528) );
  OAI211_X1 U4372 ( .C1(n3530), .C2(n3806), .A(n3529), .B(n3528), .ZN(U3212)
         );
  INV_X1 U4373 ( .A(n3532), .ZN(n3534) );
  NOR2_X1 U4374 ( .A1(n3534), .A2(n3533), .ZN(n3535) );
  XNOR2_X1 U4375 ( .A(n3531), .B(n3535), .ZN(n3544) );
  AOI22_X1 U4376 ( .A1(n3812), .A2(n3537), .B1(n3801), .B2(n3536), .ZN(n3543)
         );
  INV_X1 U4377 ( .A(n3538), .ZN(n4532) );
  NAND2_X1 U4378 ( .A1(n3813), .A2(n3998), .ZN(n3539) );
  OAI211_X1 U4379 ( .C1(n3817), .C2(n4532), .A(n3540), .B(n3539), .ZN(n3541)
         );
  INV_X1 U4380 ( .A(n3541), .ZN(n3542) );
  OAI211_X1 U4381 ( .C1(n3544), .C2(n3806), .A(n3543), .B(n3542), .ZN(U3218)
         );
  NAND2_X1 U4382 ( .A1(n4279), .A2(n3659), .ZN(n3546) );
  NAND2_X1 U4383 ( .A1(n4266), .A2(n3620), .ZN(n3545) );
  NAND2_X1 U4384 ( .A1(n3546), .A2(n3545), .ZN(n3547) );
  XNOR2_X1 U4385 ( .A(n3547), .B(n3656), .ZN(n3615) );
  AOI22_X1 U4386 ( .A1(n4279), .A2(n3670), .B1(n3659), .B2(n4266), .ZN(n3616)
         );
  XNOR2_X1 U4387 ( .A(n3615), .B(n3616), .ZN(n3613) );
  NAND2_X1 U4388 ( .A1(n3550), .A2(n3549), .ZN(n3556) );
  NAND3_X1 U4389 ( .A1(n3553), .A2(n3552), .A3(n3551), .ZN(n3555) );
  NAND2_X1 U4390 ( .A1(n3556), .A2(n2413), .ZN(n3561) );
  OAI22_X1 U4391 ( .A1(n3558), .A2(n3516), .B1(n3675), .B2(n3557), .ZN(n3559)
         );
  XOR2_X1 U4392 ( .A(n3656), .B(n3559), .Z(n3560) );
  NAND2_X1 U4393 ( .A1(n3561), .A2(n3560), .ZN(n3734) );
  NAND2_X1 U4394 ( .A1(n4379), .A2(n3670), .ZN(n3563) );
  NAND2_X1 U4395 ( .A1(n3810), .A2(n3659), .ZN(n3562) );
  NAND2_X1 U4396 ( .A1(n3563), .A2(n3562), .ZN(n3808) );
  NAND2_X1 U4397 ( .A1(n3734), .A2(n3808), .ZN(n3565) );
  OAI22_X1 U4398 ( .A1(n4368), .A2(n2967), .B1(n3516), .B2(n4373), .ZN(n3567)
         );
  OAI22_X1 U4399 ( .A1(n4368), .A2(n3676), .B1(n3675), .B2(n4373), .ZN(n3564)
         );
  XNOR2_X1 U4400 ( .A(n3564), .B(n3656), .ZN(n3566) );
  OAI22_X1 U4401 ( .A1(n4374), .A2(n3516), .B1(n3675), .B2(n3572), .ZN(n3571)
         );
  XNOR2_X1 U4402 ( .A(n3571), .B(n3656), .ZN(n3747) );
  OR2_X1 U4403 ( .A1(n4374), .A2(n2967), .ZN(n3574) );
  OR2_X1 U4404 ( .A1(n3572), .A2(n3516), .ZN(n3573) );
  NAND2_X1 U4405 ( .A1(n3574), .A2(n3573), .ZN(n3748) );
  NOR2_X1 U4406 ( .A1(n3747), .A2(n3748), .ZN(n3576) );
  NAND2_X1 U4407 ( .A1(n3747), .A2(n3748), .ZN(n3575) );
  NAND2_X1 U4408 ( .A1(n4364), .A2(n3659), .ZN(n3578) );
  NAND2_X1 U4409 ( .A1(n4284), .A2(n3620), .ZN(n3577) );
  NAND2_X1 U4410 ( .A1(n3578), .A2(n3577), .ZN(n3579) );
  XNOR2_X1 U4411 ( .A(n3579), .B(n2150), .ZN(n3582) );
  AND2_X1 U4412 ( .A1(n4284), .A2(n3659), .ZN(n3580) );
  AOI21_X1 U4413 ( .B1(n4364), .B2(n3670), .A(n3580), .ZN(n3581) );
  NAND2_X1 U4414 ( .A1(n3582), .A2(n3581), .ZN(n3785) );
  XOR2_X1 U4415 ( .A(n3613), .B(n3614), .Z(n3587) );
  AOI22_X1 U4416 ( .A1(n3812), .A2(n4364), .B1(n3801), .B2(n4266), .ZN(n3586)
         );
  NAND2_X1 U4417 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4080) );
  NAND2_X1 U4418 ( .A1(n3813), .A2(n4925), .ZN(n3583) );
  OAI211_X1 U4419 ( .C1(n3817), .C2(n4269), .A(n4080), .B(n3583), .ZN(n3584)
         );
  INV_X1 U4420 ( .A(n3584), .ZN(n3585) );
  OAI211_X1 U4421 ( .C1(n3587), .C2(n3806), .A(n3586), .B(n3585), .ZN(U3216)
         );
  INV_X1 U4422 ( .A(n3588), .ZN(n3589) );
  NOR2_X1 U4423 ( .A1(n3590), .A2(n3589), .ZN(n3591) );
  XNOR2_X1 U4424 ( .A(n3592), .B(n3591), .ZN(n3600) );
  AOI22_X1 U4425 ( .A1(n3812), .A2(n3996), .B1(n3801), .B2(n3593), .ZN(n3599)
         );
  NAND2_X1 U4426 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4482) );
  NAND2_X1 U4427 ( .A1(n3813), .A2(n3594), .ZN(n3595) );
  OAI211_X1 U4428 ( .C1(n3817), .C2(n3596), .A(n4482), .B(n3595), .ZN(n3597)
         );
  INV_X1 U4429 ( .A(n3597), .ZN(n3598) );
  OAI211_X1 U4430 ( .C1(n3600), .C2(n3806), .A(n3599), .B(n3598), .ZN(U3221)
         );
  OAI211_X1 U4431 ( .C1(n3603), .C2(n3602), .A(n3601), .B(n3819), .ZN(n3612)
         );
  NAND2_X1 U4432 ( .A1(n3813), .A2(n3996), .ZN(n3604) );
  NAND2_X1 U4433 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4461) );
  NAND2_X1 U4434 ( .A1(n3604), .A2(n4461), .ZN(n3609) );
  INV_X1 U4435 ( .A(n3801), .ZN(n3606) );
  OAI22_X1 U4436 ( .A1(n3607), .A2(n3798), .B1(n3606), .B2(n3605), .ZN(n3608)
         );
  AOI211_X1 U4437 ( .C1(n3610), .C2(n3781), .A(n3609), .B(n3608), .ZN(n3611)
         );
  NAND2_X1 U4438 ( .A1(n3612), .A2(n3611), .ZN(U3214) );
  NAND2_X1 U4439 ( .A1(n3614), .A2(n3613), .ZN(n3619) );
  INV_X1 U4440 ( .A(n3615), .ZN(n3617) );
  NAND2_X1 U4441 ( .A1(n4925), .A2(n3659), .ZN(n3622) );
  NAND2_X1 U4442 ( .A1(n4245), .A2(n3620), .ZN(n3621) );
  NAND2_X1 U4443 ( .A1(n3622), .A2(n3621), .ZN(n3623) );
  XNOR2_X1 U4444 ( .A(n3623), .B(n3656), .ZN(n3626) );
  NAND2_X1 U4445 ( .A1(n4925), .A2(n3670), .ZN(n3625) );
  NAND2_X1 U4446 ( .A1(n4245), .A2(n3659), .ZN(n3624) );
  NAND2_X1 U4447 ( .A1(n3625), .A2(n3624), .ZN(n3627) );
  NAND2_X1 U4448 ( .A1(n3626), .A2(n3627), .ZN(n3767) );
  INV_X1 U4449 ( .A(n3626), .ZN(n3629) );
  INV_X1 U4450 ( .A(n3627), .ZN(n3628) );
  NAND2_X1 U4451 ( .A1(n3629), .A2(n3628), .ZN(n3769) );
  NAND2_X1 U4452 ( .A1(n4201), .A2(n3659), .ZN(n3631) );
  OR2_X1 U4453 ( .A1(n4221), .A2(n3675), .ZN(n3630) );
  NAND2_X1 U4454 ( .A1(n3631), .A2(n3630), .ZN(n3632) );
  XNOR2_X1 U4455 ( .A(n3632), .B(n3656), .ZN(n3718) );
  NAND2_X1 U4456 ( .A1(n4201), .A2(n3670), .ZN(n3634) );
  OR2_X1 U4457 ( .A1(n4221), .A2(n3516), .ZN(n3633) );
  NAND2_X1 U4458 ( .A1(n3634), .A2(n3633), .ZN(n3635) );
  INV_X1 U4459 ( .A(n3718), .ZN(n3636) );
  INV_X1 U4460 ( .A(n3635), .ZN(n3717) );
  OAI22_X1 U4461 ( .A1(n4344), .A2(n3516), .B1(n3675), .B2(n3638), .ZN(n3637)
         );
  XNOR2_X1 U4462 ( .A(n3637), .B(n3656), .ZN(n3644) );
  OAI22_X1 U4463 ( .A1(n4344), .A2(n2967), .B1(n3516), .B2(n3638), .ZN(n3643)
         );
  XNOR2_X1 U4464 ( .A(n3644), .B(n3643), .ZN(n3777) );
  NAND2_X1 U4465 ( .A1(n4162), .A2(n3659), .ZN(n3640) );
  OR2_X1 U4466 ( .A1(n4189), .A2(n3675), .ZN(n3639) );
  NAND2_X1 U4467 ( .A1(n3640), .A2(n3639), .ZN(n3641) );
  XNOR2_X1 U4468 ( .A(n3641), .B(n2150), .ZN(n3647) );
  NOR2_X1 U4469 ( .A1(n4189), .A2(n3516), .ZN(n3642) );
  AOI21_X1 U4470 ( .B1(n4162), .B2(n3670), .A(n3642), .ZN(n3646) );
  XNOR2_X1 U4471 ( .A(n3647), .B(n3646), .ZN(n3697) );
  NOR2_X1 U4472 ( .A1(n3644), .A2(n3643), .ZN(n3698) );
  NOR2_X1 U4473 ( .A1(n3697), .A2(n3698), .ZN(n3645) );
  OR2_X1 U4474 ( .A1(n3647), .A2(n3646), .ZN(n3650) );
  NOR2_X1 U4475 ( .A1(n4170), .A2(n3516), .ZN(n3648) );
  AOI21_X1 U4476 ( .B1(n4320), .B2(n3670), .A(n3648), .ZN(n3651) );
  OAI22_X1 U4477 ( .A1(n4151), .A2(n3516), .B1(n3675), .B2(n4170), .ZN(n3649)
         );
  XNOR2_X1 U4478 ( .A(n3649), .B(n3656), .ZN(n3760) );
  NAND2_X1 U4479 ( .A1(n3758), .A2(n3760), .ZN(n3654) );
  NAND2_X1 U4480 ( .A1(n3699), .A2(n3650), .ZN(n3653) );
  INV_X1 U4481 ( .A(n3651), .ZN(n3652) );
  OAI22_X1 U4482 ( .A1(n3799), .A2(n3516), .B1(n4145), .B2(n3675), .ZN(n3655)
         );
  XOR2_X1 U4483 ( .A(n3656), .B(n3655), .Z(n3658) );
  AOI22_X1 U4484 ( .A1(n4165), .A2(n3670), .B1(n4319), .B2(n3659), .ZN(n3657)
         );
  NOR2_X1 U4485 ( .A1(n3658), .A2(n3657), .ZN(n3725) );
  NAND2_X1 U4486 ( .A1(n4308), .A2(n3659), .ZN(n3661) );
  OR2_X1 U4487 ( .A1(n4133), .A2(n3675), .ZN(n3660) );
  NAND2_X1 U4488 ( .A1(n3661), .A2(n3660), .ZN(n3662) );
  XNOR2_X1 U4489 ( .A(n3662), .B(n2150), .ZN(n3665) );
  NOR2_X1 U4490 ( .A1(n4133), .A2(n3516), .ZN(n3663) );
  AOI21_X1 U4491 ( .B1(n4308), .B2(n3670), .A(n3663), .ZN(n3664) );
  NAND2_X1 U4492 ( .A1(n3665), .A2(n3664), .ZN(n3795) );
  NAND2_X1 U4493 ( .A1(n4129), .A2(n3659), .ZN(n3667) );
  OR2_X1 U4494 ( .A1(n4117), .A2(n3675), .ZN(n3666) );
  NAND2_X1 U4495 ( .A1(n3667), .A2(n3666), .ZN(n3668) );
  XNOR2_X1 U4496 ( .A(n3668), .B(n2150), .ZN(n3672) );
  NOR2_X1 U4497 ( .A1(n4117), .A2(n3516), .ZN(n3669) );
  AOI21_X1 U4498 ( .B1(n4129), .B2(n3670), .A(n3669), .ZN(n3671) );
  XNOR2_X1 U4499 ( .A(n3672), .B(n3671), .ZN(n3691) );
  OAI22_X1 U4500 ( .A1(n4311), .A2(n2967), .B1(n3516), .B2(n3674), .ZN(n3679)
         );
  OAI22_X1 U4501 ( .A1(n4311), .A2(n3676), .B1(n3675), .B2(n3674), .ZN(n3677)
         );
  XNOR2_X1 U4502 ( .A(n3677), .B(n3656), .ZN(n3678) );
  XOR2_X1 U4503 ( .A(n3679), .B(n3678), .Z(n3680) );
  XNOR2_X1 U4504 ( .A(n3681), .B(n3680), .ZN(n3687) );
  NAND2_X1 U4505 ( .A1(n4129), .A2(n3812), .ZN(n3685) );
  AOI22_X1 U4506 ( .A1(n4098), .A2(n3813), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3684) );
  OR2_X1 U4507 ( .A1(n4097), .A2(n3817), .ZN(n3683) );
  NAND2_X1 U4508 ( .A1(n3801), .A2(n4096), .ZN(n3682) );
  AND4_X1 U4509 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3686)
         );
  OAI21_X1 U4510 ( .B1(n3687), .B2(n3806), .A(n3686), .ZN(U3217) );
  INV_X1 U4511 ( .A(IR_REG_30__SCAN_IN), .ZN(n4605) );
  NAND3_X1 U4512 ( .A1(n4605), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3688) );
  INV_X1 U4513 ( .A(DATAI_31_), .ZN(n4672) );
  OAI22_X1 U4514 ( .A1(n3689), .A2(n3688), .B1(STATE_REG_SCAN_IN), .B2(n4672), 
        .ZN(U3321) );
  XNOR2_X1 U4515 ( .A(n3690), .B(n3691), .ZN(n3695) );
  INV_X1 U4516 ( .A(n4308), .ZN(n4323) );
  OAI22_X1 U4517 ( .A1(n4323), .A2(n3798), .B1(STATE_REG_SCAN_IN), .B2(n4704), 
        .ZN(n3692) );
  AOI21_X1 U4518 ( .B1(n4307), .B2(n3801), .A(n3692), .ZN(n3694) );
  AOI22_X1 U4519 ( .A1(n4120), .A2(n3813), .B1(n4112), .B2(n3781), .ZN(n3693)
         );
  OAI211_X1 U4520 ( .C1(n3695), .C2(n3806), .A(n3694), .B(n3693), .ZN(U3211)
         );
  INV_X1 U4521 ( .A(n3696), .ZN(n3775) );
  OAI21_X1 U4522 ( .B1(n3775), .B2(n3698), .A(n3697), .ZN(n3700) );
  NAND3_X1 U4523 ( .A1(n3700), .A2(n3819), .A3(n3699), .ZN(n3706) );
  AOI22_X1 U4524 ( .A1(n3993), .A2(n3812), .B1(n3701), .B2(n3801), .ZN(n3705)
         );
  OAI22_X1 U4525 ( .A1(n4151), .A2(n3779), .B1(STATE_REG_SCAN_IN), .B2(n3702), 
        .ZN(n3703) );
  AOI21_X1 U4526 ( .B1(n4191), .B2(n3781), .A(n3703), .ZN(n3704) );
  NAND3_X1 U4527 ( .A1(n3706), .A2(n3705), .A3(n3704), .ZN(U3213) );
  OAI211_X1 U4528 ( .C1(n3707), .C2(n3709), .A(n3708), .B(n3819), .ZN(n3715)
         );
  AOI22_X1 U4529 ( .A1(n3813), .A2(n3711), .B1(REG3_REG_1__SCAN_IN), .B2(n3710), .ZN(n3714) );
  AOI22_X1 U4530 ( .A1(n3812), .A2(n2936), .B1(n3801), .B2(n3712), .ZN(n3713)
         );
  NAND3_X1 U4531 ( .A1(n3715), .A2(n3714), .A3(n3713), .ZN(U3219) );
  XNOR2_X1 U4532 ( .A(n3718), .B(n3717), .ZN(n3719) );
  XNOR2_X1 U4533 ( .A(n3716), .B(n3719), .ZN(n3723) );
  AOI22_X1 U4534 ( .A1(n3993), .A2(n3813), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3721) );
  AOI22_X1 U4535 ( .A1(n3812), .A2(n4925), .B1(n3801), .B2(n4340), .ZN(n3720)
         );
  OAI211_X1 U4536 ( .C1(n3817), .C2(n4224), .A(n3721), .B(n3720), .ZN(n3722)
         );
  AOI21_X1 U4537 ( .B1(n3723), .B2(n3819), .A(n3722), .ZN(n3724) );
  INV_X1 U4538 ( .A(n3724), .ZN(U3220) );
  NOR2_X1 U4539 ( .A1(n3725), .A2(n2171), .ZN(n3726) );
  XNOR2_X1 U4540 ( .A(n3727), .B(n3726), .ZN(n3733) );
  AOI22_X1 U4541 ( .A1(n4308), .A2(n3813), .B1(n4319), .B2(n3801), .ZN(n3732)
         );
  INV_X1 U4542 ( .A(n3728), .ZN(n4147) );
  INV_X1 U4543 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3729) );
  OAI22_X1 U4544 ( .A1(n4151), .A2(n3798), .B1(STATE_REG_SCAN_IN), .B2(n3729), 
        .ZN(n3730) );
  AOI21_X1 U4545 ( .B1(n4147), .B2(n3781), .A(n3730), .ZN(n3731) );
  OAI211_X1 U4546 ( .C1(n3733), .C2(n3806), .A(n3732), .B(n3731), .ZN(U3222)
         );
  INV_X1 U4547 ( .A(n2152), .ZN(n3735) );
  OAI21_X1 U4548 ( .B1(n3735), .B2(n3808), .A(n3734), .ZN(n3736) );
  XOR2_X1 U4549 ( .A(n3737), .B(n3736), .Z(n3745) );
  AOI22_X1 U4550 ( .A1(n3812), .A2(n4379), .B1(n3801), .B2(n3738), .ZN(n3744)
         );
  INV_X1 U4551 ( .A(n3739), .ZN(n3741) );
  NAND2_X1 U4552 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4509) );
  NAND2_X1 U4553 ( .A1(n3813), .A2(n3994), .ZN(n3740) );
  OAI211_X1 U4554 ( .C1(n3817), .C2(n3741), .A(n4509), .B(n3740), .ZN(n3742)
         );
  INV_X1 U4555 ( .A(n3742), .ZN(n3743) );
  OAI211_X1 U4556 ( .C1(n3745), .C2(n3806), .A(n3744), .B(n3743), .ZN(U3223)
         );
  XOR2_X1 U4557 ( .A(n3748), .B(n3747), .Z(n3749) );
  XNOR2_X1 U4558 ( .A(n3746), .B(n3749), .ZN(n3755) );
  INV_X1 U4559 ( .A(n3750), .ZN(n3753) );
  AOI22_X1 U4560 ( .A1(n3812), .A2(n3995), .B1(n3801), .B2(n4361), .ZN(n3752)
         );
  AND2_X1 U4561 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4065) );
  AOI21_X1 U4562 ( .B1(n3813), .B2(n4364), .A(n4065), .ZN(n3751) );
  OAI211_X1 U4563 ( .C1(n3817), .C2(n3753), .A(n3752), .B(n3751), .ZN(n3754)
         );
  AOI21_X1 U4564 ( .B1(n3755), .B2(n3819), .A(n3754), .ZN(n3756) );
  INV_X1 U4565 ( .A(n3756), .ZN(U3225) );
  NAND2_X1 U4566 ( .A1(n3757), .A2(n3758), .ZN(n3759) );
  XOR2_X1 U4567 ( .A(n3760), .B(n3759), .Z(n3765) );
  AOI22_X1 U4568 ( .A1(n4162), .A2(n3812), .B1(n2340), .B2(n3801), .ZN(n3764)
         );
  INV_X1 U4569 ( .A(n3761), .ZN(n4171) );
  OAI22_X1 U4570 ( .A1(n3799), .A2(n3779), .B1(STATE_REG_SCAN_IN), .B2(n4702), 
        .ZN(n3762) );
  AOI21_X1 U4571 ( .B1(n4171), .B2(n3781), .A(n3762), .ZN(n3763) );
  OAI211_X1 U4572 ( .C1(n3765), .C2(n3806), .A(n3764), .B(n3763), .ZN(U3226)
         );
  AOI21_X1 U4573 ( .B1(n3769), .B2(n3767), .A(n3766), .ZN(n3768) );
  AOI21_X1 U4574 ( .B1(n2158), .B2(n3769), .A(n3768), .ZN(n3774) );
  AOI22_X1 U4575 ( .A1(n3812), .A2(n4279), .B1(n3801), .B2(n4245), .ZN(n3771)
         );
  AOI22_X1 U4576 ( .A1(n3813), .A2(n4201), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3770) );
  OAI211_X1 U4577 ( .C1(n3817), .C2(n4247), .A(n3771), .B(n3770), .ZN(n3772)
         );
  INV_X1 U4578 ( .A(n3772), .ZN(n3773) );
  OAI21_X1 U4579 ( .B1(n3774), .B2(n3806), .A(n3773), .ZN(U3230) );
  AOI21_X1 U4580 ( .B1(n3777), .B2(n3776), .A(n3775), .ZN(n3784) );
  AOI22_X1 U4581 ( .A1(n3812), .A2(n4201), .B1(n3801), .B2(n4205), .ZN(n3783)
         );
  INV_X1 U4582 ( .A(n3778), .ZN(n4208) );
  OAI22_X1 U4583 ( .A1(n4204), .A2(n3779), .B1(STATE_REG_SCAN_IN), .B2(n4868), 
        .ZN(n3780) );
  AOI21_X1 U4584 ( .B1(n4208), .B2(n3781), .A(n3780), .ZN(n3782) );
  OAI211_X1 U4585 ( .C1(n3784), .C2(n3806), .A(n3783), .B(n3782), .ZN(U3232)
         );
  NAND2_X1 U4586 ( .A1(n2183), .A2(n3785), .ZN(n3786) );
  XNOR2_X1 U4587 ( .A(n3787), .B(n3786), .ZN(n3792) );
  INV_X1 U4588 ( .A(n4287), .ZN(n3790) );
  AOI22_X1 U4589 ( .A1(n3812), .A2(n3994), .B1(n3801), .B2(n4284), .ZN(n3789)
         );
  AND2_X1 U4590 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4522) );
  AOI21_X1 U4591 ( .B1(n3813), .B2(n4279), .A(n4522), .ZN(n3788) );
  OAI211_X1 U4592 ( .C1(n3817), .C2(n3790), .A(n3789), .B(n3788), .ZN(n3791)
         );
  AOI21_X1 U4593 ( .B1(n3792), .B2(n3819), .A(n3791), .ZN(n3793) );
  INV_X1 U4594 ( .A(n3793), .ZN(U3235) );
  NAND2_X1 U4595 ( .A1(n3796), .A2(n3795), .ZN(n3797) );
  XNOR2_X1 U4596 ( .A(n3794), .B(n3797), .ZN(n3807) );
  INV_X1 U4597 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4871) );
  OAI22_X1 U4598 ( .A1(n3799), .A2(n3798), .B1(STATE_REG_SCAN_IN), .B2(n4871), 
        .ZN(n3800) );
  AOI21_X1 U4599 ( .B1(n3802), .B2(n3801), .A(n3800), .ZN(n3803) );
  OAI21_X1 U4600 ( .B1(n3817), .B2(n4134), .A(n3803), .ZN(n3804) );
  AOI21_X1 U4601 ( .B1(n3813), .B2(n4129), .A(n3804), .ZN(n3805) );
  OAI21_X1 U4602 ( .B1(n3807), .B2(n3806), .A(n3805), .ZN(U3237) );
  NAND2_X1 U4603 ( .A1(n2152), .A2(n3734), .ZN(n3809) );
  XNOR2_X1 U4604 ( .A(n3809), .B(n3808), .ZN(n3820) );
  AOI22_X1 U4605 ( .A1(n3812), .A2(n3811), .B1(n3801), .B2(n3810), .ZN(n3815)
         );
  AND2_X1 U4606 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4503) );
  AOI21_X1 U4607 ( .B1(n3813), .B2(n3995), .A(n4503), .ZN(n3814) );
  OAI211_X1 U4608 ( .C1(n3817), .C2(n3816), .A(n3815), .B(n3814), .ZN(n3818)
         );
  AOI21_X1 U4609 ( .B1(n3820), .B2(n3819), .A(n3818), .ZN(n3821) );
  INV_X1 U4610 ( .A(n3821), .ZN(U3238) );
  AND2_X1 U4611 ( .A1(n2636), .A2(DATAI_30_), .ZN(n4303) );
  NAND2_X1 U4612 ( .A1(n2636), .A2(DATAI_31_), .ZN(n4296) );
  INV_X1 U4613 ( .A(n3846), .ZN(n3822) );
  NAND2_X1 U4614 ( .A1(n3822), .A2(n4303), .ZN(n3823) );
  NAND2_X1 U4615 ( .A1(n4295), .A2(n4296), .ZN(n3975) );
  AND2_X1 U4616 ( .A1(n3823), .A2(n3975), .ZN(n3869) );
  NAND2_X1 U4617 ( .A1(n3827), .A2(n3824), .ZN(n3950) );
  NAND2_X1 U4618 ( .A1(n3826), .A2(n3825), .ZN(n3933) );
  NAND2_X1 U4619 ( .A1(n3933), .A2(n3827), .ZN(n3951) );
  OAI21_X1 U4620 ( .B1(n3828), .B2(n3950), .A(n3951), .ZN(n3830) );
  INV_X1 U4621 ( .A(n3955), .ZN(n3829) );
  AOI211_X1 U4622 ( .C1(n3959), .C2(n3830), .A(n3829), .B(n3958), .ZN(n3832)
         );
  INV_X1 U4623 ( .A(n3831), .ZN(n3963) );
  OAI21_X1 U4624 ( .B1(n3832), .B2(n3963), .A(n3962), .ZN(n3833) );
  AND2_X1 U4625 ( .A1(n3834), .A2(n3833), .ZN(n3835) );
  OAI21_X1 U4626 ( .B1(n3836), .B2(n3835), .A(n3965), .ZN(n3844) );
  AOI211_X1 U4627 ( .C1(n3965), .C2(n3838), .A(n3861), .B(n3837), .ZN(n3967)
         );
  AND2_X1 U4628 ( .A1(n3839), .A2(n3862), .ZN(n3974) );
  INV_X1 U4629 ( .A(n4098), .ZN(n3841) );
  NAND2_X1 U4630 ( .A1(n3841), .A2(n3840), .ZN(n3853) );
  NAND4_X1 U4631 ( .A1(n3974), .A2(n3853), .A3(n3851), .A4(n3842), .ZN(n3843)
         );
  AOI21_X1 U4632 ( .B1(n3844), .B2(n3967), .A(n3843), .ZN(n3858) );
  INV_X1 U4633 ( .A(n4303), .ZN(n3845) );
  NAND2_X1 U4634 ( .A1(n3846), .A2(n3845), .ZN(n3864) );
  AOI21_X1 U4635 ( .B1(n3864), .B2(n4295), .A(n4296), .ZN(n3857) );
  NAND2_X1 U4636 ( .A1(n4098), .A2(n3847), .ZN(n3849) );
  NAND2_X1 U4637 ( .A1(n3849), .A2(n3848), .ZN(n3854) );
  NOR2_X1 U4638 ( .A1(n3850), .A2(n3854), .ZN(n3970) );
  NOR2_X1 U4639 ( .A1(n2317), .A2(n3852), .ZN(n3855) );
  OAI211_X1 U4640 ( .C1(n3855), .C2(n3854), .A(n3869), .B(n3853), .ZN(n3978)
         );
  AOI21_X1 U4641 ( .B1(n4110), .B2(n3970), .A(n3978), .ZN(n3856) );
  AOI211_X1 U4642 ( .C1(n3869), .C2(n3858), .A(n3857), .B(n3856), .ZN(n3859)
         );
  AOI21_X1 U4643 ( .B1(n4303), .B2(n4296), .A(n3859), .ZN(n3985) );
  INV_X1 U4644 ( .A(n3860), .ZN(n3893) );
  INV_X1 U4645 ( .A(n3861), .ZN(n3863) );
  NAND2_X1 U4646 ( .A1(n3863), .A2(n3862), .ZN(n4143) );
  INV_X1 U4647 ( .A(n4143), .ZN(n3892) );
  OAI21_X1 U4648 ( .B1(n4295), .B2(n4296), .A(n3864), .ZN(n3976) );
  NOR4_X1 U4649 ( .A1(n3866), .A2(n3865), .A3(n4430), .A4(n3976), .ZN(n3871)
         );
  INV_X1 U4650 ( .A(n4197), .ZN(n3867) );
  OR2_X1 U4651 ( .A1(n3867), .A2(n4177), .ZN(n4218) );
  INV_X1 U4652 ( .A(n4218), .ZN(n3870) );
  NAND4_X1 U4653 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3889)
         );
  INV_X1 U4654 ( .A(n4210), .ZN(n4178) );
  INV_X1 U4655 ( .A(n3872), .ZN(n3877) );
  AND4_X1 U4656 ( .A1(n3875), .A2(n3874), .A3(n3925), .A4(n3873), .ZN(n3876)
         );
  NAND4_X1 U4657 ( .A1(n4178), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3888)
         );
  NAND4_X1 U4658 ( .A1(n3882), .A2(n3881), .A3(n3880), .A4(n3879), .ZN(n3887)
         );
  NAND4_X1 U4659 ( .A1(n3885), .A2(n4590), .A3(n3884), .A4(n3883), .ZN(n3886)
         );
  NOR4_X1 U4660 ( .A1(n3889), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n3891)
         );
  OR2_X1 U4661 ( .A1(n3890), .A2(n2155), .ZN(n4123) );
  NAND4_X1 U4662 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n4123), .ZN(n3907)
         );
  AND2_X1 U4663 ( .A1(n3895), .A2(n3894), .ZN(n4159) );
  AND2_X1 U4664 ( .A1(n4157), .A2(n3896), .ZN(n4181) );
  AND2_X1 U4665 ( .A1(n3900), .A2(n3899), .ZN(n4261) );
  INV_X1 U4666 ( .A(n4261), .ZN(n3902) );
  NOR4_X1 U4667 ( .A1(n4239), .A2(n4278), .A3(n3902), .A4(n3901), .ZN(n3903)
         );
  NAND3_X1 U4668 ( .A1(n4159), .A2(n4181), .A3(n3903), .ZN(n3906) );
  INV_X1 U4669 ( .A(n4110), .ZN(n3905) );
  OR4_X1 U4670 ( .A1(n3907), .A2(n3906), .A3(n3905), .A4(n3904), .ZN(n3982) );
  INV_X1 U4671 ( .A(n3908), .ZN(n3911) );
  OAI211_X1 U4672 ( .C1(n3911), .C2(n4430), .A(n3910), .B(n3909), .ZN(n3914)
         );
  NAND3_X1 U4673 ( .A1(n3914), .A2(n3913), .A3(n3912), .ZN(n3917) );
  NAND3_X1 U4674 ( .A1(n3917), .A2(n3916), .A3(n3915), .ZN(n3920) );
  NAND3_X1 U4675 ( .A1(n3920), .A2(n3919), .A3(n3918), .ZN(n3923) );
  NAND4_X1 U4676 ( .A1(n3923), .A2(n3922), .A3(n3921), .A4(n3936), .ZN(n3926)
         );
  AND3_X1 U4677 ( .A1(n3926), .A2(n3925), .A3(n3924), .ZN(n3931) );
  NAND2_X1 U4678 ( .A1(n3928), .A2(n3927), .ZN(n3935) );
  OAI211_X1 U4679 ( .C1(n3931), .C2(n3935), .A(n3930), .B(n3929), .ZN(n3944)
         );
  NOR2_X1 U4680 ( .A1(n3933), .A2(n3932), .ZN(n3943) );
  INV_X1 U4681 ( .A(n3934), .ZN(n3939) );
  INV_X1 U4682 ( .A(n3935), .ZN(n3938) );
  NAND4_X1 U4683 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3941)
         );
  NAND2_X1 U4684 ( .A1(n3941), .A2(n3940), .ZN(n3942) );
  AOI22_X1 U4685 ( .A1(n3944), .A2(n3943), .B1(n3951), .B2(n3942), .ZN(n3949)
         );
  INV_X1 U4686 ( .A(n3945), .ZN(n3947) );
  NOR4_X1 U4687 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3957)
         );
  INV_X1 U4688 ( .A(n3950), .ZN(n3953) );
  INV_X1 U4689 ( .A(n3951), .ZN(n3952) );
  AOI21_X1 U4690 ( .B1(n3954), .B2(n3953), .A(n3952), .ZN(n3956) );
  OAI21_X1 U4691 ( .B1(n3957), .B2(n3956), .A(n3955), .ZN(n3960) );
  AOI21_X1 U4692 ( .B1(n3960), .B2(n3959), .A(n3958), .ZN(n3964) );
  INV_X1 U4693 ( .A(n4177), .ZN(n3961) );
  OAI211_X1 U4694 ( .C1(n3964), .C2(n3963), .A(n3962), .B(n3961), .ZN(n3966)
         );
  NAND2_X1 U4695 ( .A1(n3966), .A2(n3965), .ZN(n3968) );
  OAI21_X1 U4696 ( .B1(n3969), .B2(n3968), .A(n3967), .ZN(n3973) );
  NOR2_X1 U4697 ( .A1(n4102), .A2(n4307), .ZN(n3972) );
  INV_X1 U4698 ( .A(n3970), .ZN(n3971) );
  AOI211_X1 U4699 ( .C1(n3974), .C2(n3973), .A(n3972), .B(n3971), .ZN(n3979)
         );
  NAND2_X1 U4700 ( .A1(n3976), .A2(n3975), .ZN(n3977) );
  OAI21_X1 U4701 ( .B1(n3979), .B2(n3978), .A(n3977), .ZN(n3981) );
  MUX2_X1 U4702 ( .A(n3982), .B(n3981), .S(n3980), .Z(n3983) );
  OAI21_X1 U4703 ( .B1(n3985), .B2(n3984), .A(n3983), .ZN(n3986) );
  XNOR2_X1 U4704 ( .A(n3986), .B(n4667), .ZN(n3992) );
  NAND2_X1 U4705 ( .A1(n3988), .A2(n3987), .ZN(n3989) );
  OAI211_X1 U4706 ( .C1(n4429), .C2(n3991), .A(n3989), .B(B_REG_SCAN_IN), .ZN(
        n3990) );
  OAI21_X1 U4707 ( .B1(n3992), .B2(n3991), .A(n3990), .ZN(U3239) );
  MUX2_X1 U4708 ( .A(n4320), .B(DATAO_REG_24__SCAN_IN), .S(n4002), .Z(U3574)
         );
  MUX2_X1 U4709 ( .A(n3993), .B(DATAO_REG_22__SCAN_IN), .S(n4002), .Z(U3572)
         );
  MUX2_X1 U4710 ( .A(n4201), .B(DATAO_REG_21__SCAN_IN), .S(n4002), .Z(U3571)
         );
  MUX2_X1 U4711 ( .A(n4279), .B(DATAO_REG_19__SCAN_IN), .S(n4002), .Z(U3569)
         );
  MUX2_X1 U4712 ( .A(n4364), .B(DATAO_REG_18__SCAN_IN), .S(n4002), .Z(U3568)
         );
  MUX2_X1 U4713 ( .A(DATAO_REG_17__SCAN_IN), .B(n3994), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4714 ( .A(DATAO_REG_16__SCAN_IN), .B(n3995), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4715 ( .A(n4379), .B(DATAO_REG_15__SCAN_IN), .S(n4002), .Z(U3565)
         );
  MUX2_X1 U4716 ( .A(n3996), .B(DATAO_REG_11__SCAN_IN), .S(n4002), .Z(U3561)
         );
  MUX2_X1 U4717 ( .A(n3997), .B(DATAO_REG_10__SCAN_IN), .S(n4002), .Z(U3560)
         );
  MUX2_X1 U4718 ( .A(n3998), .B(DATAO_REG_9__SCAN_IN), .S(n4002), .Z(U3559) );
  MUX2_X1 U4719 ( .A(DATAO_REG_8__SCAN_IN), .B(n3999), .S(U4043), .Z(U3558) );
  MUX2_X1 U4720 ( .A(n4000), .B(DATAO_REG_6__SCAN_IN), .S(n4002), .Z(U3556) );
  MUX2_X1 U4721 ( .A(n4001), .B(DATAO_REG_4__SCAN_IN), .S(n4002), .Z(U3554) );
  MUX2_X1 U4722 ( .A(n4580), .B(DATAO_REG_3__SCAN_IN), .S(n4002), .Z(U3553) );
  MUX2_X1 U4723 ( .A(n2936), .B(DATAO_REG_0__SCAN_IN), .S(n4002), .Z(U3550) );
  NAND2_X1 U4724 ( .A1(n4030), .A2(n4438), .ZN(n4012) );
  OAI211_X1 U4725 ( .C1(n4005), .C2(n4004), .A(n4525), .B(n4003), .ZN(n4011)
         );
  AOI22_X1 U4726 ( .A1(n4523), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4010) );
  MUX2_X1 U4727 ( .A(REG2_REG_1__SCAN_IN), .B(n2845), .S(n4006), .Z(n4007) );
  OAI21_X1 U4728 ( .B1(n4547), .B2(n2364), .A(n4007), .ZN(n4008) );
  NAND3_X1 U4729 ( .A1(n4480), .A2(n4020), .A3(n4008), .ZN(n4009) );
  NAND4_X1 U4730 ( .A1(n4012), .A2(n4011), .A3(n4010), .A4(n4009), .ZN(U3241)
         );
  NAND2_X1 U4731 ( .A1(U3149), .A2(REG3_REG_2__SCAN_IN), .ZN(n4014) );
  NAND2_X1 U4732 ( .A1(n4523), .A2(ADDR_REG_2__SCAN_IN), .ZN(n4013) );
  OAI211_X1 U4733 ( .C1(n4530), .C2(n4015), .A(n4014), .B(n4013), .ZN(n4016)
         );
  INV_X1 U4734 ( .A(n4016), .ZN(n4028) );
  MUX2_X1 U4735 ( .A(n4017), .B(REG2_REG_2__SCAN_IN), .S(n4437), .Z(n4018) );
  NAND3_X1 U4736 ( .A1(n4020), .A2(n4019), .A3(n4018), .ZN(n4021) );
  NAND3_X1 U4737 ( .A1(n4480), .A2(n4022), .A3(n4021), .ZN(n4027) );
  OAI211_X1 U4738 ( .C1(n4025), .C2(n4024), .A(n4525), .B(n4023), .ZN(n4026)
         );
  NAND4_X1 U4739 ( .A1(n4029), .A2(n4028), .A3(n4027), .A4(n4026), .ZN(U3242)
         );
  NAND2_X1 U4740 ( .A1(n4030), .A2(n4436), .ZN(n4039) );
  OAI211_X1 U4741 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4032), .A(n4525), .B(n4031), 
        .ZN(n4038) );
  AOI22_X1 U4742 ( .A1(n4523), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n4037) );
  XNOR2_X1 U4743 ( .A(n4034), .B(n4033), .ZN(n4035) );
  NAND2_X1 U4744 ( .A1(n4480), .A2(n4035), .ZN(n4036) );
  NAND4_X1 U4745 ( .A1(n4039), .A2(n4038), .A3(n4037), .A4(n4036), .ZN(U3243)
         );
  NAND2_X1 U4746 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4056), .ZN(n4045) );
  INV_X1 U4747 ( .A(n4056), .ZN(n4556) );
  AOI22_X1 U4748 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4056), .B1(n4556), .B2(
        n3459), .ZN(n4506) );
  INV_X1 U4749 ( .A(n4040), .ZN(n4042) );
  NAND2_X1 U4750 ( .A1(n4042), .A2(n4041), .ZN(n4043) );
  NAND2_X1 U4751 ( .A1(n4557), .A2(n4043), .ZN(n4044) );
  INV_X1 U4752 ( .A(n4557), .ZN(n4498) );
  XNOR2_X1 U4753 ( .A(n4043), .B(n4498), .ZN(n4495) );
  NAND2_X1 U4754 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4495), .ZN(n4494) );
  NAND2_X1 U4755 ( .A1(n4044), .A2(n4494), .ZN(n4505) );
  NAND2_X1 U4756 ( .A1(n4506), .A2(n4505), .ZN(n4504) );
  NOR2_X1 U4757 ( .A1(n4057), .A2(n4046), .ZN(n4047) );
  INV_X1 U4758 ( .A(n4057), .ZN(n4555) );
  INV_X1 U4759 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4809) );
  NOR2_X1 U4760 ( .A1(n4072), .A2(REG1_REG_17__SCAN_IN), .ZN(n4076) );
  INV_X1 U4761 ( .A(n4076), .ZN(n4048) );
  OAI21_X1 U4762 ( .B1(n4809), .B2(n4063), .A(n4048), .ZN(n4049) );
  NOR2_X1 U4763 ( .A1(n4050), .A2(n4049), .ZN(n4075) );
  AOI21_X1 U4764 ( .B1(n4050), .B2(n4049), .A(n4075), .ZN(n4069) );
  XNOR2_X1 U4765 ( .A(n4063), .B(REG2_REG_17__SCAN_IN), .ZN(n4061) );
  NOR2_X1 U4766 ( .A1(n4498), .A2(n4053), .ZN(n4054) );
  INV_X1 U4767 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4833) );
  NOR2_X1 U4768 ( .A1(n4833), .A2(n4491), .ZN(n4490) );
  NAND2_X1 U4769 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4056), .ZN(n4055) );
  OAI21_X1 U4770 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4056), .A(n4055), .ZN(n4500) );
  NAND2_X1 U4771 ( .A1(n4058), .A2(n4555), .ZN(n4059) );
  INV_X1 U4772 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U4773 ( .A1(n4059), .A2(n4511), .ZN(n4060) );
  NAND2_X1 U4774 ( .A1(n4060), .A2(n4061), .ZN(n4071) );
  AOI221_X1 U4775 ( .B1(n4061), .B2(n4071), .C1(n4060), .C2(n4071), .A(n4519), 
        .ZN(n4062) );
  INV_X1 U4776 ( .A(n4062), .ZN(n4067) );
  NOR2_X1 U4777 ( .A1(n4530), .A2(n4063), .ZN(n4064) );
  AOI211_X1 U4778 ( .C1(n4523), .C2(ADDR_REG_17__SCAN_IN), .A(n4065), .B(n4064), .ZN(n4066) );
  OAI211_X1 U4779 ( .C1(n4069), .C2(n4068), .A(n4067), .B(n4066), .ZN(U3257)
         );
  INV_X1 U4780 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4836) );
  MUX2_X1 U4781 ( .A(n4836), .B(REG2_REG_19__SCAN_IN), .S(n4081), .Z(n4073) );
  INV_X1 U4782 ( .A(n4074), .ZN(n4554) );
  INV_X1 U4783 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U4784 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4554), .B1(n4074), .B2(
        n4070), .ZN(n4521) );
  INV_X1 U4785 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U4786 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4074), .B1(n4554), .B2(
        n4077), .ZN(n4527) );
  INV_X1 U4787 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4811) );
  MUX2_X1 U4788 ( .A(REG1_REG_19__SCAN_IN), .B(n4811), .S(n4081), .Z(n4078) );
  NAND2_X1 U4789 ( .A1(n4523), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4079) );
  OAI211_X1 U4790 ( .C1(n4530), .C2(n4081), .A(n4080), .B(n4079), .ZN(n4082)
         );
  AOI21_X1 U4791 ( .B1(n4083), .B2(n4525), .A(n4082), .ZN(n4084) );
  OAI21_X1 U4792 ( .B1(n4085), .B2(n4519), .A(n4084), .ZN(U3259) );
  NAND2_X1 U4793 ( .A1(n4086), .A2(n4220), .ZN(n4092) );
  OAI22_X1 U4794 ( .A1(n4088), .A2(n4443), .B1(n4087), .B2(n4531), .ZN(n4089)
         );
  OAI21_X1 U4795 ( .B1(n4090), .B2(n4089), .A(n2143), .ZN(n4091) );
  OAI211_X1 U4796 ( .C1(n2143), .C2(n4093), .A(n4092), .B(n4091), .ZN(U3354)
         );
  NAND2_X1 U4797 ( .A1(n4094), .A2(n4220), .ZN(n4106) );
  INV_X1 U4798 ( .A(n4095), .ZN(n4104) );
  AOI22_X1 U4799 ( .A1(n4222), .A2(n4096), .B1(n4661), .B2(
        REG2_REG_28__SCAN_IN), .ZN(n4101) );
  INV_X1 U4800 ( .A(n4097), .ZN(n4099) );
  AOI22_X1 U4801 ( .A1(n4663), .A2(n4099), .B1(n4098), .B2(n4146), .ZN(n4100)
         );
  OAI211_X1 U4802 ( .C1(n4102), .C2(n4150), .A(n4101), .B(n4100), .ZN(n4103)
         );
  AOI21_X1 U4803 ( .B1(n4104), .B2(n4536), .A(n4103), .ZN(n4105) );
  OAI211_X1 U4804 ( .C1(n4661), .C2(n4107), .A(n4106), .B(n4105), .ZN(U3262)
         );
  XNOR2_X1 U4805 ( .A(n4108), .B(n4110), .ZN(n4109) );
  NAND2_X1 U4806 ( .A1(n4109), .A2(n4282), .ZN(n4310) );
  XNOR2_X1 U4807 ( .A(n4111), .B(n4110), .ZN(n4313) );
  NAND2_X1 U4808 ( .A1(n4313), .A2(n4220), .ZN(n4122) );
  AOI22_X1 U4809 ( .A1(n4222), .A2(n4307), .B1(n4661), .B2(
        REG2_REG_27__SCAN_IN), .ZN(n4114) );
  NAND2_X1 U4810 ( .A1(n4112), .A2(n4663), .ZN(n4113) );
  OAI211_X1 U4811 ( .C1(n4323), .C2(n4150), .A(n4114), .B(n4113), .ZN(n4119)
         );
  INV_X1 U4812 ( .A(n4115), .ZN(n4116) );
  OAI21_X1 U4813 ( .B1(n2341), .B2(n4117), .A(n4116), .ZN(n4391) );
  NOR2_X1 U4814 ( .A1(n4391), .A2(n4443), .ZN(n4118) );
  AOI211_X1 U4815 ( .C1(n4146), .C2(n4120), .A(n4119), .B(n4118), .ZN(n4121)
         );
  OAI211_X1 U4816 ( .C1(n4661), .C2(n4310), .A(n4122), .B(n4121), .ZN(U3263)
         );
  XOR2_X1 U4817 ( .A(n4123), .B(n2165), .Z(n4317) );
  INV_X1 U4818 ( .A(n4317), .ZN(n4139) );
  INV_X1 U4819 ( .A(n4123), .ZN(n4124) );
  XNOR2_X1 U4820 ( .A(n4125), .B(n4124), .ZN(n4126) );
  NAND2_X1 U4821 ( .A1(n4126), .A2(n4282), .ZN(n4131) );
  NAND2_X1 U4822 ( .A1(n4165), .A2(n4581), .ZN(n4127) );
  OAI21_X1 U4823 ( .B1(n4571), .B2(n4133), .A(n4127), .ZN(n4128) );
  AOI21_X1 U4824 ( .B1(n4129), .B2(n4363), .A(n4128), .ZN(n4130) );
  NAND2_X1 U4825 ( .A1(n4131), .A2(n4130), .ZN(n4316) );
  OAI21_X1 U4826 ( .B1(n2338), .B2(n4133), .A(n4132), .ZN(n4394) );
  INV_X1 U4827 ( .A(n4134), .ZN(n4135) );
  AOI22_X1 U4828 ( .A1(n4135), .A2(n4663), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4661), .ZN(n4136) );
  OAI21_X1 U4829 ( .B1(n4394), .B2(n4443), .A(n4136), .ZN(n4137) );
  AOI21_X1 U4830 ( .B1(n4316), .B2(n2143), .A(n4137), .ZN(n4138) );
  OAI21_X1 U4831 ( .B1(n4139), .B2(n4293), .A(n4138), .ZN(U3264) );
  XNOR2_X1 U4832 ( .A(n4140), .B(n4143), .ZN(n4141) );
  NAND2_X1 U4833 ( .A1(n4141), .A2(n4282), .ZN(n4322) );
  XNOR2_X1 U4834 ( .A(n4142), .B(n4143), .ZN(n4325) );
  NAND2_X1 U4835 ( .A1(n4325), .A2(n4220), .ZN(n4155) );
  OAI21_X1 U4836 ( .B1(n4168), .B2(n4145), .A(n4144), .ZN(n4398) );
  INV_X1 U4837 ( .A(n4398), .ZN(n4153) );
  AOI22_X1 U4838 ( .A1(n4308), .A2(n4146), .B1(n4222), .B2(n4319), .ZN(n4149)
         );
  AOI22_X1 U4839 ( .A1(n4147), .A2(n4663), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4661), .ZN(n4148) );
  OAI211_X1 U4840 ( .C1(n4151), .C2(n4150), .A(n4149), .B(n4148), .ZN(n4152)
         );
  AOI21_X1 U4841 ( .B1(n4153), .B2(n4536), .A(n4152), .ZN(n4154) );
  OAI211_X1 U4842 ( .C1(n4661), .C2(n4322), .A(n4155), .B(n4154), .ZN(U3265)
         );
  XOR2_X1 U4843 ( .A(n4159), .B(n4156), .Z(n4329) );
  INV_X1 U4844 ( .A(n4329), .ZN(n4175) );
  NAND2_X1 U4845 ( .A1(n4158), .A2(n4157), .ZN(n4160) );
  XNOR2_X1 U4846 ( .A(n4160), .B(n4159), .ZN(n4161) );
  NAND2_X1 U4847 ( .A1(n4161), .A2(n4282), .ZN(n4167) );
  NAND2_X1 U4848 ( .A1(n4162), .A2(n4581), .ZN(n4163) );
  OAI21_X1 U4849 ( .B1(n4571), .B2(n4170), .A(n4163), .ZN(n4164) );
  AOI21_X1 U4850 ( .B1(n4165), .B2(n4363), .A(n4164), .ZN(n4166) );
  NAND2_X1 U4851 ( .A1(n4167), .A2(n4166), .ZN(n4328) );
  INV_X1 U4852 ( .A(n4168), .ZN(n4169) );
  OAI21_X1 U4853 ( .B1(n4187), .B2(n4170), .A(n4169), .ZN(n4401) );
  AOI22_X1 U4854 ( .A1(n4171), .A2(n4663), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4661), .ZN(n4172) );
  OAI21_X1 U4855 ( .B1(n4401), .B2(n4443), .A(n4172), .ZN(n4173) );
  AOI21_X1 U4856 ( .B1(n4328), .B2(n2143), .A(n4173), .ZN(n4174) );
  OAI21_X1 U4857 ( .B1(n4175), .B2(n4293), .A(n4174), .ZN(U3266) );
  XNOR2_X1 U4858 ( .A(n4176), .B(n4181), .ZN(n4332) );
  INV_X1 U4859 ( .A(n4332), .ZN(n4195) );
  OR2_X1 U4860 ( .A1(n4216), .A2(n4177), .ZN(n4198) );
  NAND2_X1 U4861 ( .A1(n4198), .A2(n4197), .ZN(n4179) );
  NAND2_X1 U4862 ( .A1(n4179), .A2(n4178), .ZN(n4196) );
  NAND2_X1 U4863 ( .A1(n4196), .A2(n4180), .ZN(n4182) );
  XNOR2_X1 U4864 ( .A(n4182), .B(n4181), .ZN(n4183) );
  NAND2_X1 U4865 ( .A1(n4183), .A2(n4282), .ZN(n4186) );
  OAI22_X1 U4866 ( .A1(n4344), .A2(n4367), .B1(n4571), .B2(n4189), .ZN(n4184)
         );
  AOI21_X1 U4867 ( .B1(n4320), .B2(n4363), .A(n4184), .ZN(n4185) );
  NAND2_X1 U4868 ( .A1(n4186), .A2(n4185), .ZN(n4331) );
  INV_X1 U4869 ( .A(n4207), .ZN(n4190) );
  INV_X1 U4870 ( .A(n4187), .ZN(n4188) );
  OAI21_X1 U4871 ( .B1(n4190), .B2(n4189), .A(n4188), .ZN(n4405) );
  AOI22_X1 U4872 ( .A1(n4191), .A2(n4663), .B1(n4661), .B2(
        REG2_REG_23__SCAN_IN), .ZN(n4192) );
  OAI21_X1 U4873 ( .B1(n4405), .B2(n4443), .A(n4192), .ZN(n4193) );
  AOI21_X1 U4874 ( .B1(n4331), .B2(n2143), .A(n4193), .ZN(n4194) );
  OAI21_X1 U4875 ( .B1(n4195), .B2(n4293), .A(n4194), .ZN(U3267) );
  INV_X1 U4876 ( .A(n4196), .ZN(n4200) );
  AND3_X1 U4877 ( .A1(n4198), .A2(n4210), .A3(n4197), .ZN(n4199) );
  OAI21_X1 U4878 ( .B1(n4200), .B2(n4199), .A(n4282), .ZN(n4203) );
  AOI22_X1 U4879 ( .A1(n4201), .A2(n4581), .B1(n4205), .B2(n4362), .ZN(n4202)
         );
  OAI211_X1 U4880 ( .C1(n4204), .C2(n4573), .A(n4203), .B(n4202), .ZN(n4336)
         );
  NAND2_X1 U4881 ( .A1(n2145), .A2(n4205), .ZN(n4206) );
  NAND2_X1 U4882 ( .A1(n4207), .A2(n4206), .ZN(n4409) );
  AOI22_X1 U4883 ( .A1(n4661), .A2(REG2_REG_22__SCAN_IN), .B1(n4208), .B2(
        n4663), .ZN(n4209) );
  OAI21_X1 U4884 ( .B1(n4409), .B2(n4443), .A(n4209), .ZN(n4214) );
  NOR2_X1 U4885 ( .A1(n4211), .A2(n4210), .ZN(n4335) );
  INV_X1 U4886 ( .A(n4337), .ZN(n4212) );
  NOR3_X1 U4887 ( .A1(n4335), .A2(n4212), .A3(n4293), .ZN(n4213) );
  AOI211_X1 U4888 ( .C1(n2143), .C2(n4336), .A(n4214), .B(n4213), .ZN(n4215)
         );
  INV_X1 U4889 ( .A(n4215), .ZN(U3268) );
  XNOR2_X1 U4890 ( .A(n4216), .B(n4218), .ZN(n4217) );
  NAND2_X1 U4891 ( .A1(n4217), .A2(n4282), .ZN(n4343) );
  XNOR2_X1 U4892 ( .A(n4219), .B(n4218), .ZN(n4346) );
  NAND2_X1 U4893 ( .A1(n4346), .A2(n4220), .ZN(n4232) );
  OAI21_X1 U4894 ( .B1(n2336), .B2(n4221), .A(n2145), .ZN(n4413) );
  INV_X1 U4895 ( .A(n4413), .ZN(n4230) );
  AOI22_X1 U4896 ( .A1(n4223), .A2(n4925), .B1(n4222), .B2(n4340), .ZN(n4227)
         );
  INV_X1 U4897 ( .A(n4224), .ZN(n4225) );
  AOI22_X1 U4898 ( .A1(n4661), .A2(REG2_REG_21__SCAN_IN), .B1(n4225), .B2(
        n4663), .ZN(n4226) );
  OAI211_X1 U4899 ( .C1(n4344), .C2(n4228), .A(n4227), .B(n4226), .ZN(n4229)
         );
  AOI21_X1 U4900 ( .B1(n4230), .B2(n4536), .A(n4229), .ZN(n4231) );
  OAI211_X1 U4901 ( .C1(n4661), .C2(n4343), .A(n4232), .B(n4231), .ZN(U3269)
         );
  INV_X1 U4902 ( .A(n4233), .ZN(n4235) );
  NOR2_X1 U4903 ( .A1(n4235), .A2(n4234), .ZN(n4236) );
  XNOR2_X1 U4904 ( .A(n4236), .B(n4239), .ZN(n4244) );
  AOI22_X1 U4905 ( .A1(n4279), .A2(n4581), .B1(n4245), .B2(n4362), .ZN(n4237)
         );
  OAI21_X1 U4906 ( .B1(n4238), .B2(n4573), .A(n4237), .ZN(n4243) );
  XNOR2_X1 U4907 ( .A(n4240), .B(n4239), .ZN(n4354) );
  NOR2_X1 U4908 ( .A1(n4354), .A2(n4241), .ZN(n4242) );
  AOI211_X1 U4909 ( .C1(n4282), .C2(n4244), .A(n4243), .B(n4242), .ZN(n4352)
         );
  INV_X1 U4910 ( .A(n4354), .ZN(n4251) );
  INV_X1 U4911 ( .A(n4267), .ZN(n4246) );
  NAND2_X1 U4912 ( .A1(n4246), .A2(n4245), .ZN(n4350) );
  AND3_X1 U4913 ( .A1(n4350), .A2(n4536), .A3(n4349), .ZN(n4250) );
  INV_X1 U4914 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4248) );
  OAI22_X1 U4915 ( .A1(n2143), .A2(n4248), .B1(n4247), .B2(n4531), .ZN(n4249)
         );
  AOI211_X1 U4916 ( .C1(n4251), .C2(n4544), .A(n4250), .B(n4249), .ZN(n4252)
         );
  OAI21_X1 U4917 ( .B1(n4352), .B2(n4661), .A(n4252), .ZN(U3270) );
  XOR2_X1 U4918 ( .A(n4261), .B(n4253), .Z(n4356) );
  INV_X1 U4919 ( .A(n4356), .ZN(n4273) );
  OAI21_X1 U4920 ( .B1(n4256), .B2(n4255), .A(n4254), .ZN(n4277) );
  INV_X1 U4921 ( .A(n4257), .ZN(n4259) );
  OAI21_X1 U4922 ( .B1(n4277), .B2(n4259), .A(n4258), .ZN(n4260) );
  XOR2_X1 U4923 ( .A(n4261), .B(n4260), .Z(n4262) );
  NAND2_X1 U4924 ( .A1(n4262), .A2(n4282), .ZN(n4264) );
  AOI22_X1 U4925 ( .A1(n4925), .A2(n4363), .B1(n4362), .B2(n4266), .ZN(n4263)
         );
  OAI211_X1 U4926 ( .C1(n4265), .C2(n4367), .A(n4264), .B(n4263), .ZN(n4355)
         );
  AND2_X1 U4927 ( .A1(n2173), .A2(n4266), .ZN(n4268) );
  OR2_X1 U4928 ( .A1(n4268), .A2(n4267), .ZN(n4418) );
  NOR2_X1 U4929 ( .A1(n4418), .A2(n4443), .ZN(n4271) );
  OAI22_X1 U4930 ( .A1(n2143), .A2(n4836), .B1(n4269), .B2(n4531), .ZN(n4270)
         );
  AOI211_X1 U4931 ( .C1(n4355), .C2(n2143), .A(n4271), .B(n4270), .ZN(n4272)
         );
  OAI21_X1 U4932 ( .B1(n4273), .B2(n4293), .A(n4272), .ZN(U3271) );
  OAI21_X1 U4933 ( .B1(n4275), .B2(n4278), .A(n4274), .ZN(n4276) );
  INV_X1 U4934 ( .A(n4276), .ZN(n4360) );
  XOR2_X1 U4935 ( .A(n4278), .B(n4277), .Z(n4283) );
  AOI22_X1 U4936 ( .A1(n4279), .A2(n4363), .B1(n4284), .B2(n4362), .ZN(n4280)
         );
  OAI21_X1 U4937 ( .B1(n4374), .B2(n4367), .A(n4280), .ZN(n4281) );
  AOI21_X1 U4938 ( .B1(n4283), .B2(n4282), .A(n4281), .ZN(n4359) );
  INV_X1 U4939 ( .A(n4359), .ZN(n4291) );
  AOI21_X1 U4940 ( .B1(n4285), .B2(n4284), .A(n4375), .ZN(n4286) );
  NAND2_X1 U4941 ( .A1(n4286), .A2(n2173), .ZN(n4358) );
  AOI22_X1 U4942 ( .A1(n4661), .A2(REG2_REG_18__SCAN_IN), .B1(n4287), .B2(
        n4663), .ZN(n4288) );
  OAI21_X1 U4943 ( .B1(n4358), .B2(n4289), .A(n4288), .ZN(n4290) );
  AOI21_X1 U4944 ( .B1(n4291), .B2(n2143), .A(n4290), .ZN(n4292) );
  OAI21_X1 U4945 ( .B1(n4360), .B2(n4293), .A(n4292), .ZN(U3272) );
  INV_X1 U4946 ( .A(n4440), .ZN(n4299) );
  NAND2_X1 U4947 ( .A1(n4295), .A2(n4294), .ZN(n4305) );
  OAI21_X1 U4948 ( .B1(n4296), .B2(n4571), .A(n4305), .ZN(n4439) );
  NAND2_X1 U4949 ( .A1(n4604), .A2(n4439), .ZN(n4298) );
  NAND2_X1 U4950 ( .A1(n4602), .A2(REG1_REG_31__SCAN_IN), .ZN(n4297) );
  OAI211_X1 U4951 ( .C1(n4299), .C2(n4372), .A(n4298), .B(n4297), .ZN(U3549)
         );
  AND2_X1 U4952 ( .A1(n4300), .A2(n4303), .ZN(n4302) );
  INV_X1 U4953 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U4954 ( .A1(n4303), .A2(n4362), .ZN(n4304) );
  AND2_X1 U4955 ( .A1(n4305), .A2(n4304), .ZN(n4442) );
  MUX2_X1 U4956 ( .A(n4820), .B(n4442), .S(n4604), .Z(n4306) );
  OAI21_X1 U4957 ( .B1(n4444), .B2(n4372), .A(n4306), .ZN(U3548) );
  INV_X1 U4958 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4314) );
  AOI22_X1 U4959 ( .A1(n4308), .A2(n4581), .B1(n4307), .B2(n4362), .ZN(n4309)
         );
  OAI211_X1 U4960 ( .C1(n4311), .C2(n4573), .A(n4310), .B(n4309), .ZN(n4312)
         );
  AOI21_X1 U4961 ( .B1(n4313), .B2(n4593), .A(n4312), .ZN(n4388) );
  MUX2_X1 U4962 ( .A(n4314), .B(n4388), .S(n4604), .Z(n4315) );
  OAI21_X1 U4963 ( .B1(n4372), .B2(n4391), .A(n4315), .ZN(U3545) );
  INV_X1 U4964 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4821) );
  AOI21_X1 U4965 ( .B1(n4317), .B2(n4593), .A(n4316), .ZN(n4392) );
  MUX2_X1 U4966 ( .A(n4821), .B(n4392), .S(n4604), .Z(n4318) );
  OAI21_X1 U4967 ( .B1(n4372), .B2(n4394), .A(n4318), .ZN(U3544) );
  INV_X1 U4968 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4326) );
  AOI22_X1 U4969 ( .A1(n4320), .A2(n4581), .B1(n4319), .B2(n4362), .ZN(n4321)
         );
  OAI211_X1 U4970 ( .C1(n4323), .C2(n4573), .A(n4322), .B(n4321), .ZN(n4324)
         );
  AOI21_X1 U4971 ( .B1(n4325), .B2(n4593), .A(n4324), .ZN(n4395) );
  MUX2_X1 U4972 ( .A(n4326), .B(n4395), .S(n4604), .Z(n4327) );
  OAI21_X1 U4973 ( .B1(n4372), .B2(n4398), .A(n4327), .ZN(U3543) );
  INV_X1 U4974 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4813) );
  AOI21_X1 U4975 ( .B1(n4329), .B2(n4593), .A(n4328), .ZN(n4399) );
  MUX2_X1 U4976 ( .A(n4813), .B(n4399), .S(n4604), .Z(n4330) );
  OAI21_X1 U4977 ( .B1(n4372), .B2(n4401), .A(n4330), .ZN(U3542) );
  INV_X1 U4978 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4333) );
  AOI21_X1 U4979 ( .B1(n4332), .B2(n4593), .A(n4331), .ZN(n4402) );
  MUX2_X1 U4980 ( .A(n4333), .B(n4402), .S(n4604), .Z(n4334) );
  OAI21_X1 U4981 ( .B1(n4372), .B2(n4405), .A(n4334), .ZN(U3541) );
  INV_X1 U4982 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4814) );
  INV_X1 U4983 ( .A(n4593), .ZN(n4382) );
  NOR2_X1 U4984 ( .A1(n4335), .A2(n4382), .ZN(n4338) );
  AOI21_X1 U4985 ( .B1(n4338), .B2(n4337), .A(n4336), .ZN(n4406) );
  MUX2_X1 U4986 ( .A(n4814), .B(n4406), .S(n4604), .Z(n4339) );
  OAI21_X1 U4987 ( .B1(n4372), .B2(n4409), .A(n4339), .ZN(U3540) );
  INV_X1 U4988 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4347) );
  AOI22_X1 U4989 ( .A1(n4925), .A2(n4581), .B1(n4362), .B2(n4340), .ZN(n4342)
         );
  OAI211_X1 U4990 ( .C1(n4344), .C2(n4573), .A(n4343), .B(n4342), .ZN(n4345)
         );
  AOI21_X1 U4991 ( .B1(n4346), .B2(n4593), .A(n4345), .ZN(n4410) );
  MUX2_X1 U4992 ( .A(n4347), .B(n4410), .S(n4604), .Z(n4348) );
  OAI21_X1 U4993 ( .B1(n4372), .B2(n4413), .A(n4348), .ZN(U3539) );
  NAND3_X1 U4994 ( .A1(n4350), .A2(n4584), .A3(n4349), .ZN(n4351) );
  OAI211_X1 U4995 ( .C1(n4354), .C2(n4353), .A(n4352), .B(n4351), .ZN(n4414)
         );
  MUX2_X1 U4996 ( .A(REG1_REG_20__SCAN_IN), .B(n4414), .S(n4604), .Z(U3538) );
  AOI21_X1 U4997 ( .B1(n4356), .B2(n4593), .A(n4355), .ZN(n4415) );
  MUX2_X1 U4998 ( .A(n4811), .B(n4415), .S(n4604), .Z(n4357) );
  OAI21_X1 U4999 ( .B1(n4372), .B2(n4418), .A(n4357), .ZN(U3537) );
  OAI211_X1 U5000 ( .C1(n4360), .C2(n4382), .A(n4359), .B(n4358), .ZN(n4419)
         );
  MUX2_X1 U5001 ( .A(REG1_REG_18__SCAN_IN), .B(n4419), .S(n4604), .Z(U3536) );
  AOI22_X1 U5002 ( .A1(n4364), .A2(n4363), .B1(n4362), .B2(n4361), .ZN(n4365)
         );
  OAI211_X1 U5003 ( .C1(n4368), .C2(n4367), .A(n4366), .B(n4365), .ZN(n4369)
         );
  AOI21_X1 U5004 ( .B1(n4370), .B2(n4593), .A(n4369), .ZN(n4421) );
  MUX2_X1 U5005 ( .A(n4421), .B(n4809), .S(n4602), .Z(n4371) );
  OAI21_X1 U5006 ( .B1(n4372), .B2(n4424), .A(n4371), .ZN(U3535) );
  OAI22_X1 U5007 ( .A1(n4374), .A2(n4573), .B1(n4373), .B2(n4571), .ZN(n4378)
         );
  NOR2_X1 U5008 ( .A1(n4376), .A2(n4375), .ZN(n4377) );
  AOI211_X1 U5009 ( .C1(n4581), .C2(n4379), .A(n4378), .B(n4377), .ZN(n4381)
         );
  OAI211_X1 U5010 ( .C1(n4383), .C2(n4382), .A(n4381), .B(n4380), .ZN(n4425)
         );
  MUX2_X1 U5011 ( .A(REG1_REG_16__SCAN_IN), .B(n4425), .S(n4604), .Z(U3534) );
  NAND2_X1 U5012 ( .A1(n4440), .A2(n4568), .ZN(n4385) );
  NAND2_X1 U5013 ( .A1(n4600), .A2(n4439), .ZN(n4384) );
  OAI211_X1 U5014 ( .C1(n4600), .C2(n4386), .A(n4385), .B(n4384), .ZN(U3517)
         );
  MUX2_X1 U5015 ( .A(n2801), .B(n4442), .S(n4600), .Z(n4387) );
  OAI21_X1 U5016 ( .B1(n4444), .B2(n4423), .A(n4387), .ZN(U3516) );
  MUX2_X1 U5017 ( .A(n4389), .B(n4388), .S(n4600), .Z(n4390) );
  OAI21_X1 U5018 ( .B1(n4391), .B2(n4423), .A(n4390), .ZN(U3513) );
  MUX2_X1 U5019 ( .A(n4777), .B(n4392), .S(n4600), .Z(n4393) );
  OAI21_X1 U5020 ( .B1(n4394), .B2(n4423), .A(n4393), .ZN(U3512) );
  MUX2_X1 U5021 ( .A(n4396), .B(n4395), .S(n4600), .Z(n4397) );
  OAI21_X1 U5022 ( .B1(n4398), .B2(n4423), .A(n4397), .ZN(U3511) );
  MUX2_X1 U5023 ( .A(n4778), .B(n4399), .S(n4600), .Z(n4400) );
  OAI21_X1 U5024 ( .B1(n4401), .B2(n4423), .A(n4400), .ZN(U3510) );
  MUX2_X1 U5025 ( .A(n4403), .B(n4402), .S(n4600), .Z(n4404) );
  OAI21_X1 U5026 ( .B1(n4405), .B2(n4423), .A(n4404), .ZN(U3509) );
  MUX2_X1 U5027 ( .A(n4407), .B(n4406), .S(n4600), .Z(n4408) );
  OAI21_X1 U5028 ( .B1(n4409), .B2(n4423), .A(n4408), .ZN(U3508) );
  INV_X1 U5029 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4411) );
  MUX2_X1 U5030 ( .A(n4411), .B(n4410), .S(n4600), .Z(n4412) );
  OAI21_X1 U5031 ( .B1(n4413), .B2(n4423), .A(n4412), .ZN(U3507) );
  MUX2_X1 U5032 ( .A(REG0_REG_20__SCAN_IN), .B(n4414), .S(n4600), .Z(U3506) );
  INV_X1 U5033 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4416) );
  MUX2_X1 U5034 ( .A(n4416), .B(n4415), .S(n4600), .Z(n4417) );
  OAI21_X1 U5035 ( .B1(n4418), .B2(n4423), .A(n4417), .ZN(U3505) );
  MUX2_X1 U5036 ( .A(REG0_REG_18__SCAN_IN), .B(n4419), .S(n4600), .Z(U3503) );
  INV_X1 U5037 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4420) );
  MUX2_X1 U5038 ( .A(n4421), .B(n4420), .S(n4598), .Z(n4422) );
  OAI21_X1 U5039 ( .B1(n4424), .B2(n4423), .A(n4422), .ZN(U3501) );
  MUX2_X1 U5040 ( .A(REG0_REG_16__SCAN_IN), .B(n4425), .S(n4600), .Z(U3499) );
  MUX2_X1 U5041 ( .A(DATAI_27_), .B(n4426), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5042 ( .A(n4427), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5043 ( .A(n4428), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5044 ( .A(DATAI_22_), .B(n4429), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5045 ( .A(n4430), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5046 ( .A(DATAI_20_), .B(n4431), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5047 ( .A(DATAI_19_), .B(n4667), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5048 ( .A(n4432), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5049 ( .A(n4433), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5050 ( .A(n4434), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5051 ( .A(DATAI_4_), .B(n4435), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5052 ( .A(n4436), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5053 ( .A(n4437), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5054 ( .A(n4438), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5055 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X1 U5056 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4858) );
  AOI22_X1 U5057 ( .A1(n4440), .A2(n4536), .B1(n2143), .B2(n4439), .ZN(n4441)
         );
  OAI21_X1 U5058 ( .B1(n2143), .B2(n4858), .A(n4441), .ZN(U3260) );
  INV_X1 U5059 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4841) );
  OAI22_X1 U5060 ( .A1(n4444), .A2(n4443), .B1(n4661), .B2(n4442), .ZN(n4445)
         );
  INV_X1 U5061 ( .A(n4445), .ZN(n4446) );
  OAI21_X1 U5062 ( .B1(n4841), .B2(n2143), .A(n4446), .ZN(U3261) );
  OAI211_X1 U5063 ( .C1(n4449), .C2(n4448), .A(n4525), .B(n4447), .ZN(n4454)
         );
  OAI211_X1 U5064 ( .C1(n4452), .C2(n4451), .A(n4480), .B(n4450), .ZN(n4453)
         );
  OAI211_X1 U5065 ( .C1(n4530), .C2(n4563), .A(n4454), .B(n4453), .ZN(n4455)
         );
  AOI211_X1 U5066 ( .C1(n4523), .C2(ADDR_REG_9__SCAN_IN), .A(n4456), .B(n4455), 
        .ZN(n4457) );
  INV_X1 U5067 ( .A(n4457), .ZN(U3249) );
  OAI211_X1 U5068 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4459), .A(n4480), .B(n4458), .ZN(n4460) );
  NAND2_X1 U5069 ( .A1(n4461), .A2(n4460), .ZN(n4462) );
  AOI21_X1 U5070 ( .B1(n4523), .B2(ADDR_REG_10__SCAN_IN), .A(n4462), .ZN(n4466) );
  OAI211_X1 U5071 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4464), .A(n4525), .B(n4463), .ZN(n4465) );
  OAI211_X1 U5072 ( .C1(n4530), .C2(n4467), .A(n4466), .B(n4465), .ZN(U3250)
         );
  OAI211_X1 U5073 ( .C1(n4470), .C2(n4469), .A(n4525), .B(n4468), .ZN(n4475)
         );
  OAI211_X1 U5074 ( .C1(n4473), .C2(n4472), .A(n4480), .B(n4471), .ZN(n4474)
         );
  OAI211_X1 U5075 ( .C1(n4530), .C2(n4560), .A(n4475), .B(n4474), .ZN(n4476)
         );
  AOI211_X1 U5076 ( .C1(n4523), .C2(ADDR_REG_11__SCAN_IN), .A(n4477), .B(n4476), .ZN(n4478) );
  INV_X1 U5077 ( .A(n4478), .ZN(U3251) );
  OAI211_X1 U5078 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4481), .A(n4480), .B(n4479), .ZN(n4483) );
  NAND2_X1 U5079 ( .A1(n4483), .A2(n4482), .ZN(n4484) );
  AOI21_X1 U5080 ( .B1(n4523), .B2(ADDR_REG_12__SCAN_IN), .A(n4484), .ZN(n4488) );
  OAI211_X1 U5081 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4486), .A(n4525), .B(n4485), .ZN(n4487) );
  OAI211_X1 U5082 ( .C1(n4530), .C2(n4559), .A(n4488), .B(n4487), .ZN(U3252)
         );
  INV_X1 U5083 ( .A(n4489), .ZN(n4493) );
  AOI211_X1 U5084 ( .C1(n4833), .C2(n4491), .A(n4490), .B(n4519), .ZN(n4492)
         );
  AOI211_X1 U5085 ( .C1(n4523), .C2(ADDR_REG_14__SCAN_IN), .A(n4493), .B(n4492), .ZN(n4497) );
  OAI211_X1 U5086 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4495), .A(n4525), .B(n4494), .ZN(n4496) );
  OAI211_X1 U5087 ( .C1(n4530), .C2(n4498), .A(n4497), .B(n4496), .ZN(U3254)
         );
  AOI211_X1 U5088 ( .C1(n4501), .C2(n4500), .A(n4499), .B(n4519), .ZN(n4502)
         );
  AOI211_X1 U5089 ( .C1(n4523), .C2(ADDR_REG_15__SCAN_IN), .A(n4503), .B(n4502), .ZN(n4508) );
  OAI211_X1 U5090 ( .C1(n4506), .C2(n4505), .A(n4525), .B(n4504), .ZN(n4507)
         );
  OAI211_X1 U5091 ( .C1(n4530), .C2(n4556), .A(n4508), .B(n4507), .ZN(U3255)
         );
  INV_X1 U5092 ( .A(n4509), .ZN(n4514) );
  AOI221_X1 U5093 ( .B1(n4512), .B2(n4511), .C1(n4510), .C2(n4511), .A(n4519), 
        .ZN(n4513) );
  AOI211_X1 U5094 ( .C1(n4523), .C2(ADDR_REG_16__SCAN_IN), .A(n4514), .B(n4513), .ZN(n4518) );
  OAI221_X1 U5095 ( .B1(n4516), .B2(REG1_REG_16__SCAN_IN), .C1(n4516), .C2(
        n4515), .A(n4525), .ZN(n4517) );
  OAI211_X1 U5096 ( .C1(n4530), .C2(n4555), .A(n4518), .B(n4517), .ZN(U3256)
         );
  OAI211_X1 U5097 ( .C1(n4527), .C2(n4526), .A(n4525), .B(n4524), .ZN(n4528)
         );
  OAI211_X1 U5098 ( .C1(n4530), .C2(n4554), .A(n4529), .B(n4528), .ZN(U3258)
         );
  OAI22_X1 U5099 ( .A1(n2143), .A2(n4533), .B1(n4532), .B2(n4531), .ZN(n4534)
         );
  INV_X1 U5100 ( .A(n4534), .ZN(n4539) );
  AOI22_X1 U5101 ( .A1(n4537), .A2(n4544), .B1(n4536), .B2(n4535), .ZN(n4538)
         );
  OAI211_X1 U5102 ( .C1(n4661), .C2(n4540), .A(n4539), .B(n4538), .ZN(U3282)
         );
  AOI21_X1 U5103 ( .B1(n4543), .B2(n4542), .A(n4541), .ZN(n4548) );
  AOI22_X1 U5104 ( .A1(n4545), .A2(n4544), .B1(REG3_REG_0__SCAN_IN), .B2(n4663), .ZN(n4546) );
  OAI221_X1 U5105 ( .B1(n4661), .B2(n4548), .C1(n2143), .C2(n4547), .A(n4546), 
        .ZN(U3290) );
  NOR2_X1 U5106 ( .A1(n4550), .A2(n4761), .ZN(U3291) );
  AND2_X1 U5107 ( .A1(D_REG_30__SCAN_IN), .A2(n4549), .ZN(U3292) );
  INV_X1 U5108 ( .A(D_REG_29__SCAN_IN), .ZN(n4760) );
  NOR2_X1 U5109 ( .A1(n4550), .A2(n4760), .ZN(U3293) );
  AND2_X1 U5110 ( .A1(D_REG_28__SCAN_IN), .A2(n4549), .ZN(U3294) );
  NOR2_X1 U5111 ( .A1(n4550), .A2(n4753), .ZN(U3295) );
  NOR2_X1 U5112 ( .A1(n4550), .A2(n4754), .ZN(U3296) );
  AND2_X1 U5113 ( .A1(D_REG_25__SCAN_IN), .A2(n4549), .ZN(U3297) );
  AND2_X1 U5114 ( .A1(D_REG_24__SCAN_IN), .A2(n4549), .ZN(U3298) );
  AND2_X1 U5115 ( .A1(D_REG_23__SCAN_IN), .A2(n4549), .ZN(U3299) );
  NOR2_X1 U5116 ( .A1(n4550), .A2(n4750), .ZN(U3300) );
  INV_X1 U5117 ( .A(D_REG_21__SCAN_IN), .ZN(n4751) );
  NOR2_X1 U5118 ( .A1(n4550), .A2(n4751), .ZN(U3301) );
  AND2_X1 U5119 ( .A1(D_REG_20__SCAN_IN), .A2(n4549), .ZN(U3302) );
  AND2_X1 U5120 ( .A1(D_REG_19__SCAN_IN), .A2(n4549), .ZN(U3303) );
  AND2_X1 U5121 ( .A1(D_REG_18__SCAN_IN), .A2(n4549), .ZN(U3304) );
  NOR2_X1 U5122 ( .A1(n4550), .A2(n4747), .ZN(U3305) );
  AND2_X1 U5123 ( .A1(D_REG_16__SCAN_IN), .A2(n4549), .ZN(U3306) );
  AND2_X1 U5124 ( .A1(D_REG_15__SCAN_IN), .A2(n4549), .ZN(U3307) );
  NOR2_X1 U5125 ( .A1(n4550), .A2(n4748), .ZN(U3308) );
  AND2_X1 U5126 ( .A1(D_REG_13__SCAN_IN), .A2(n4549), .ZN(U3309) );
  AND2_X1 U5127 ( .A1(D_REG_12__SCAN_IN), .A2(n4549), .ZN(U3310) );
  AND2_X1 U5128 ( .A1(D_REG_11__SCAN_IN), .A2(n4549), .ZN(U3311) );
  AND2_X1 U5129 ( .A1(D_REG_10__SCAN_IN), .A2(n4549), .ZN(U3312) );
  NOR2_X1 U5130 ( .A1(n4550), .A2(n4864), .ZN(U3313) );
  NOR2_X1 U5131 ( .A1(n4550), .A2(n4867), .ZN(U3314) );
  AND2_X1 U5132 ( .A1(D_REG_7__SCAN_IN), .A2(n4549), .ZN(U3315) );
  INV_X1 U5133 ( .A(D_REG_6__SCAN_IN), .ZN(n4745) );
  NOR2_X1 U5134 ( .A1(n4550), .A2(n4745), .ZN(U3316) );
  AND2_X1 U5135 ( .A1(D_REG_5__SCAN_IN), .A2(n4549), .ZN(U3317) );
  AND2_X1 U5136 ( .A1(D_REG_4__SCAN_IN), .A2(n4549), .ZN(U3318) );
  NOR2_X1 U5137 ( .A1(n4550), .A2(n4744), .ZN(U3319) );
  NOR2_X1 U5138 ( .A1(n4550), .A2(n4740), .ZN(U3320) );
  OAI21_X1 U5139 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4551), .ZN(
        n4552) );
  INV_X1 U5140 ( .A(n4552), .ZN(U3329) );
  INV_X1 U5141 ( .A(DATAI_18_), .ZN(n4553) );
  AOI22_X1 U5142 ( .A1(STATE_REG_SCAN_IN), .A2(n4554), .B1(n4553), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5143 ( .A(DATAI_16_), .ZN(n4680) );
  AOI22_X1 U5144 ( .A1(STATE_REG_SCAN_IN), .A2(n4555), .B1(n4680), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5145 ( .A(DATAI_15_), .ZN(n4681) );
  AOI22_X1 U5146 ( .A1(STATE_REG_SCAN_IN), .A2(n4556), .B1(n4681), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5147 ( .A1(U3149), .A2(n4557), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4558) );
  INV_X1 U5148 ( .A(n4558), .ZN(U3338) );
  INV_X1 U5149 ( .A(DATAI_12_), .ZN(n4688) );
  AOI22_X1 U5150 ( .A1(STATE_REG_SCAN_IN), .A2(n4559), .B1(n4688), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5151 ( .A(DATAI_11_), .ZN(n4691) );
  AOI22_X1 U5152 ( .A1(STATE_REG_SCAN_IN), .A2(n4560), .B1(n4691), .B2(U3149), 
        .ZN(U3341) );
  OAI22_X1 U5153 ( .A1(U3149), .A2(n4561), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4562) );
  INV_X1 U5154 ( .A(n4562), .ZN(U3342) );
  INV_X1 U5155 ( .A(DATAI_9_), .ZN(n4690) );
  AOI22_X1 U5156 ( .A1(STATE_REG_SCAN_IN), .A2(n4563), .B1(n4690), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5157 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4763) );
  AOI22_X1 U5158 ( .A1(n4600), .A2(n4564), .B1(n4763), .B2(n4598), .ZN(U3467)
         );
  INV_X1 U5159 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4565) );
  AOI22_X1 U5160 ( .A1(n4600), .A2(n4566), .B1(n4565), .B2(n4598), .ZN(U3469)
         );
  AOI22_X1 U5161 ( .A1(n4569), .A2(n4600), .B1(n4568), .B2(n4567), .ZN(n4570)
         );
  OAI21_X1 U5162 ( .B1(n4600), .B2(n2461), .A(n4570), .ZN(U3471) );
  OAI22_X1 U5163 ( .A1(n4574), .A2(n4573), .B1(n4572), .B2(n4571), .ZN(n4579)
         );
  XOR2_X1 U5164 ( .A(n4590), .B(n4575), .Z(n4577) );
  NOR2_X1 U5165 ( .A1(n4577), .A2(n4576), .ZN(n4578) );
  AOI211_X1 U5166 ( .C1(n4581), .C2(n4580), .A(n4579), .B(n4578), .ZN(n4657)
         );
  NAND2_X1 U5167 ( .A1(n4583), .A2(n4582), .ZN(n4585) );
  NAND2_X1 U5168 ( .A1(n4585), .A2(n4584), .ZN(n4587) );
  OR2_X1 U5169 ( .A1(n4587), .A2(n4586), .ZN(n4666) );
  AND2_X1 U5170 ( .A1(n4589), .A2(n4588), .ZN(n4591) );
  OR2_X1 U5171 ( .A1(n4591), .A2(n4590), .ZN(n4660) );
  NAND2_X1 U5172 ( .A1(n4591), .A2(n4590), .ZN(n4659) );
  NAND3_X1 U5173 ( .A1(n4660), .A2(n4659), .A3(n4593), .ZN(n4592) );
  AND3_X1 U5174 ( .A1(n4657), .A2(n4666), .A3(n4592), .ZN(n4601) );
  AOI22_X1 U5175 ( .A1(n4600), .A2(n4601), .B1(n2482), .B2(n4598), .ZN(U3475)
         );
  NAND3_X1 U5176 ( .A1(n3183), .A2(n4594), .A3(n4593), .ZN(n4595) );
  AND3_X1 U5177 ( .A1(n4597), .A2(n4596), .A3(n4595), .ZN(n4603) );
  INV_X1 U5178 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4599) );
  AOI22_X1 U5179 ( .A1(n4600), .A2(n4603), .B1(n4599), .B2(n4598), .ZN(U3481)
         );
  INV_X1 U5180 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4798) );
  AOI22_X1 U5181 ( .A1(n4604), .A2(n4601), .B1(n4798), .B2(n4602), .ZN(U3522)
         );
  AOI22_X1 U5182 ( .A1(n4604), .A2(n4603), .B1(n4793), .B2(n4602), .ZN(U3525)
         );
  NAND4_X1 U5183 ( .A1(n4606), .A2(n4605), .A3(IR_REG_22__SCAN_IN), .A4(
        REG1_REG_4__SCAN_IN), .ZN(n4608) );
  NOR3_X1 U5184 ( .A1(n4608), .A2(n2482), .A3(n4607), .ZN(n4621) );
  OR4_X1 U5185 ( .A1(REG0_REG_5__SCAN_IN), .A2(REG0_REG_0__SCAN_IN), .A3(
        REG1_REG_0__SCAN_IN), .A4(n4033), .ZN(n4619) );
  INV_X1 U5186 ( .A(n4609), .ZN(n4613) );
  NOR4_X1 U5187 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .A3(
        IR_REG_6__SCAN_IN), .A4(IR_REG_0__SCAN_IN), .ZN(n4610) );
  NAND3_X1 U5188 ( .A1(n4713), .A2(n4610), .A3(REG0_REG_2__SCAN_IN), .ZN(n4612) );
  NOR4_X1 U5189 ( .A1(n4613), .A2(n4612), .A3(DATAI_4_), .A4(n4611), .ZN(n4615) );
  NOR2_X1 U5190 ( .A1(n4721), .A2(DATAI_3_), .ZN(n4614) );
  NAND4_X1 U5191 ( .A1(n4615), .A2(DATAI_0_), .A3(n4614), .A4(
        IR_REG_12__SCAN_IN), .ZN(n4618) );
  NOR4_X1 U5192 ( .A1(n4619), .A2(n4618), .A3(n4617), .A4(n4616), .ZN(n4620)
         );
  NAND4_X1 U5193 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .A3(n4621), .A4(n4620), .ZN(n4656) );
  INV_X1 U5194 ( .A(DATAI_6_), .ZN(n4693) );
  NOR4_X1 U5195 ( .A1(DATAI_9_), .A2(n2523), .A3(n4693), .A4(n4696), .ZN(n4627) );
  NOR4_X1 U5196 ( .A1(DATAI_16_), .A2(DATAI_13_), .A3(n4688), .A4(n4691), .ZN(
        n4626) );
  INV_X1 U5197 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4622) );
  NOR4_X1 U5198 ( .A1(REG0_REG_13__SCAN_IN), .A2(REG0_REG_6__SCAN_IN), .A3(
        n4623), .A4(n4622), .ZN(n4625) );
  NOR4_X1 U5199 ( .A1(REG3_REG_28__SCAN_IN), .A2(REG3_REG_24__SCAN_IN), .A3(
        REG3_REG_23__SCAN_IN), .A4(n4704), .ZN(n4624) );
  NAND4_X1 U5200 ( .A1(n4627), .A2(n4626), .A3(n4625), .A4(n4624), .ZN(n4655)
         );
  NOR4_X1 U5201 ( .A1(n4761), .A2(n4744), .A3(n4748), .A4(n4754), .ZN(n4631)
         );
  NOR4_X1 U5202 ( .A1(D_REG_21__SCAN_IN), .A2(REG2_REG_5__SCAN_IN), .A3(
        REG1_REG_5__SCAN_IN), .A4(n4760), .ZN(n4630) );
  NOR4_X1 U5203 ( .A1(DATAI_29_), .A2(DATAI_27_), .A3(n4675), .A4(n4678), .ZN(
        n4629) );
  INV_X1 U5204 ( .A(DATAI_21_), .ZN(n4677) );
  NOR4_X1 U5205 ( .A1(n4677), .A2(n4745), .A3(n4672), .A4(DATAI_15_), .ZN(
        n4628) );
  NAND4_X1 U5206 ( .A1(n4631), .A2(n4630), .A3(n4629), .A4(n4628), .ZN(n4654)
         );
  NAND4_X1 U5207 ( .A1(REG1_REG_24__SCAN_IN), .A2(n4821), .A3(n3139), .A4(
        n4820), .ZN(n4635) );
  INV_X1 U5208 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4808) );
  NAND4_X1 U5209 ( .A1(REG1_REG_21__SCAN_IN), .A2(n4814), .A3(n4811), .A4(
        n4808), .ZN(n4634) );
  INV_X1 U5210 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4839) );
  NAND4_X1 U5211 ( .A1(REG2_REG_19__SCAN_IN), .A2(REG2_REG_15__SCAN_IN), .A3(
        n4839), .A4(n4833), .ZN(n4633) );
  INV_X1 U5212 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4827) );
  NAND4_X1 U5213 ( .A1(REG2_REG_12__SCAN_IN), .A2(n2213), .A3(n4827), .A4(
        n4825), .ZN(n4632) );
  NOR4_X1 U5214 ( .A1(n4635), .A2(n4634), .A3(n4633), .A4(n4632), .ZN(n4652)
         );
  NAND4_X1 U5215 ( .A1(REG0_REG_24__SCAN_IN), .A2(REG0_REG_30__SCAN_IN), .A3(
        n4780), .A4(n4777), .ZN(n4639) );
  NAND4_X1 U5216 ( .A1(REG0_REG_19__SCAN_IN), .A2(REG0_REG_23__SCAN_IN), .A3(
        REG0_REG_16__SCAN_IN), .A4(n4774), .ZN(n4638) );
  NAND4_X1 U5217 ( .A1(n4809), .A2(n3459), .A3(n4806), .A4(n4790), .ZN(n4637)
         );
  NAND4_X1 U5218 ( .A1(REG1_REG_13__SCAN_IN), .A2(REG1_REG_7__SCAN_IN), .A3(
        n4797), .A4(n4794), .ZN(n4636) );
  NOR4_X1 U5219 ( .A1(n4639), .A2(n4638), .A3(n4637), .A4(n4636), .ZN(n4651)
         );
  NAND4_X1 U5220 ( .A1(DATAO_REG_23__SCAN_IN), .A2(DATAO_REG_27__SCAN_IN), 
        .A3(n4640), .A4(n4896), .ZN(n4644) );
  NAND4_X1 U5221 ( .A1(DATAO_REG_13__SCAN_IN), .A2(DATAO_REG_14__SCAN_IN), 
        .A3(DATAO_REG_20__SCAN_IN), .A4(n4880), .ZN(n4643) );
  NAND4_X1 U5222 ( .A1(REG3_REG_22__SCAN_IN), .A2(DATAO_REG_31__SCAN_IN), .A3(
        n3729), .A4(n4865), .ZN(n4642) );
  NAND4_X1 U5223 ( .A1(REG3_REG_26__SCAN_IN), .A2(DATAO_REG_30__SCAN_IN), .A3(
        n4898), .A4(n4901), .ZN(n4641) );
  NOR4_X1 U5224 ( .A1(n4644), .A2(n4643), .A3(n4642), .A4(n4641), .ZN(n4650)
         );
  INV_X1 U5225 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4857) );
  NAND4_X1 U5226 ( .A1(ADDR_REG_15__SCAN_IN), .A2(ADDR_REG_13__SCAN_IN), .A3(
        ADDR_REG_7__SCAN_IN), .A4(n4857), .ZN(n4648) );
  INV_X1 U5227 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4838) );
  NAND4_X1 U5228 ( .A1(REG2_REG_29__SCAN_IN), .A2(REG2_REG_31__SCAN_IN), .A3(
        n4841), .A4(n4838), .ZN(n4647) );
  NAND4_X1 U5229 ( .A1(DATAO_REG_1__SCAN_IN), .A2(DATAO_REG_5__SCAN_IN), .A3(
        n4884), .A4(n4881), .ZN(n4646) );
  INV_X1 U5230 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4852) );
  INV_X1 U5231 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4851) );
  OR4_X1 U5232 ( .A1(n4852), .A2(n4851), .A3(ADDR_REG_10__SCAN_IN), .A4(
        ADDR_REG_0__SCAN_IN), .ZN(n4645) );
  NOR4_X1 U5233 ( .A1(n4648), .A2(n4647), .A3(n4646), .A4(n4645), .ZN(n4649)
         );
  NAND4_X1 U5234 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), .ZN(n4653)
         );
  NOR4_X1 U5235 ( .A1(n4656), .A2(n4655), .A3(n4654), .A4(n4653), .ZN(n4922)
         );
  INV_X1 U5236 ( .A(n4657), .ZN(n4669) );
  NAND3_X1 U5237 ( .A1(n4660), .A2(n4659), .A3(n4658), .ZN(n4665) );
  AOI21_X1 U5238 ( .B1(n4663), .B2(n4662), .A(n4661), .ZN(n4664) );
  OAI211_X1 U5239 ( .C1(n4667), .C2(n4666), .A(n4665), .B(n4664), .ZN(n4668)
         );
  OAI22_X1 U5240 ( .A1(n4669), .A2(n4668), .B1(REG2_REG_4__SCAN_IN), .B2(n2143), .ZN(n4920) );
  AOI22_X1 U5241 ( .A1(n4672), .A2(keyinput117), .B1(n4671), .B2(keyinput21), 
        .ZN(n4670) );
  OAI221_X1 U5242 ( .B1(n4672), .B2(keyinput117), .C1(n4671), .C2(keyinput21), 
        .A(n4670), .ZN(n4685) );
  INV_X1 U5243 ( .A(DATAI_27_), .ZN(n4674) );
  AOI22_X1 U5244 ( .A1(n4675), .A2(keyinput29), .B1(keyinput48), .B2(n4674), 
        .ZN(n4673) );
  OAI221_X1 U5245 ( .B1(n4675), .B2(keyinput29), .C1(n4674), .C2(keyinput48), 
        .A(n4673), .ZN(n4684) );
  AOI22_X1 U5246 ( .A1(n4678), .A2(keyinput81), .B1(n4677), .B2(keyinput84), 
        .ZN(n4676) );
  OAI221_X1 U5247 ( .B1(n4678), .B2(keyinput81), .C1(n4677), .C2(keyinput84), 
        .A(n4676), .ZN(n4683) );
  AOI22_X1 U5248 ( .A1(n4681), .A2(keyinput98), .B1(n4680), .B2(keyinput92), 
        .ZN(n4679) );
  OAI221_X1 U5249 ( .B1(n4681), .B2(keyinput98), .C1(n4680), .C2(keyinput92), 
        .A(n4679), .ZN(n4682) );
  NOR4_X1 U5250 ( .A1(n4685), .A2(n4684), .A3(n4683), .A4(n4682), .ZN(n4729)
         );
  AOI22_X1 U5251 ( .A1(n4688), .A2(keyinput45), .B1(n4687), .B2(keyinput61), 
        .ZN(n4686) );
  OAI221_X1 U5252 ( .B1(n4688), .B2(keyinput45), .C1(n4687), .C2(keyinput61), 
        .A(n4686), .ZN(n4700) );
  AOI22_X1 U5253 ( .A1(n4691), .A2(keyinput18), .B1(keyinput116), .B2(n4690), 
        .ZN(n4689) );
  OAI221_X1 U5254 ( .B1(n4691), .B2(keyinput18), .C1(n4690), .C2(keyinput116), 
        .A(n4689), .ZN(n4699) );
  AOI22_X1 U5255 ( .A1(n4693), .A2(keyinput22), .B1(n2523), .B2(keyinput35), 
        .ZN(n4692) );
  OAI221_X1 U5256 ( .B1(n4693), .B2(keyinput22), .C1(n2523), .C2(keyinput35), 
        .A(n4692), .ZN(n4698) );
  INV_X1 U5257 ( .A(DATAI_4_), .ZN(n4695) );
  AOI22_X1 U5258 ( .A1(n4696), .A2(keyinput53), .B1(keyinput34), .B2(n4695), 
        .ZN(n4694) );
  OAI221_X1 U5259 ( .B1(n4696), .B2(keyinput53), .C1(n4695), .C2(keyinput34), 
        .A(n4694), .ZN(n4697) );
  NOR4_X1 U5260 ( .A1(n4700), .A2(n4699), .A3(n4698), .A4(n4697), .ZN(n4728)
         );
  AOI22_X1 U5261 ( .A1(n2417), .A2(keyinput15), .B1(keyinput23), .B2(n4702), 
        .ZN(n4701) );
  OAI221_X1 U5262 ( .B1(n2417), .B2(keyinput15), .C1(n4702), .C2(keyinput23), 
        .A(n4701), .ZN(n4711) );
  AOI22_X1 U5263 ( .A1(U3149), .A2(keyinput31), .B1(keyinput60), .B2(n4704), 
        .ZN(n4703) );
  OAI221_X1 U5264 ( .B1(U3149), .B2(keyinput31), .C1(n4704), .C2(keyinput60), 
        .A(n4703), .ZN(n4710) );
  XNOR2_X1 U5265 ( .A(DATAI_3_), .B(keyinput73), .ZN(n4708) );
  XNOR2_X1 U5266 ( .A(DATAI_0_), .B(keyinput68), .ZN(n4707) );
  XNOR2_X1 U5267 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput6), .ZN(n4706) );
  XNOR2_X1 U5268 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput78), .ZN(n4705) );
  NAND4_X1 U5269 ( .A1(n4708), .A2(n4707), .A3(n4706), .A4(n4705), .ZN(n4709)
         );
  NOR3_X1 U5270 ( .A1(n4711), .A2(n4710), .A3(n4709), .ZN(n4727) );
  INV_X1 U5271 ( .A(IR_REG_12__SCAN_IN), .ZN(n4714) );
  AOI22_X1 U5272 ( .A1(n4714), .A2(keyinput82), .B1(n4713), .B2(keyinput121), 
        .ZN(n4712) );
  OAI221_X1 U5273 ( .B1(n4714), .B2(keyinput82), .C1(n4713), .C2(keyinput121), 
        .A(n4712), .ZN(n4725) );
  XNOR2_X1 U5274 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput75), .ZN(n4719) );
  XNOR2_X1 U5275 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput47), .ZN(n4718) );
  XNOR2_X1 U5276 ( .A(IR_REG_0__SCAN_IN), .B(keyinput126), .ZN(n4717) );
  XNOR2_X1 U5277 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput40), .ZN(n4716) );
  NAND4_X1 U5278 ( .A1(n4719), .A2(n4718), .A3(n4717), .A4(n4716), .ZN(n4724)
         );
  XNOR2_X1 U5279 ( .A(n4720), .B(keyinput115), .ZN(n4723) );
  XNOR2_X1 U5280 ( .A(n4721), .B(keyinput57), .ZN(n4722) );
  NOR4_X1 U5281 ( .A1(n4725), .A2(n4724), .A3(n4723), .A4(n4722), .ZN(n4726)
         );
  NAND4_X1 U5282 ( .A1(n4729), .A2(n4728), .A3(n4727), .A4(n4726), .ZN(n4918)
         );
  XOR2_X1 U5283 ( .A(IR_REG_17__SCAN_IN), .B(keyinput96), .Z(n4735) );
  XOR2_X1 U5284 ( .A(IR_REG_22__SCAN_IN), .B(keyinput74), .Z(n4734) );
  XNOR2_X1 U5285 ( .A(n4730), .B(keyinput100), .ZN(n4733) );
  XNOR2_X1 U5286 ( .A(n4731), .B(keyinput12), .ZN(n4732) );
  NOR4_X1 U5287 ( .A1(n4735), .A2(n4734), .A3(n4733), .A4(n4732), .ZN(n4739)
         );
  XNOR2_X1 U5288 ( .A(IR_REG_23__SCAN_IN), .B(keyinput67), .ZN(n4738) );
  XNOR2_X1 U5289 ( .A(IR_REG_15__SCAN_IN), .B(keyinput58), .ZN(n4737) );
  XNOR2_X1 U5290 ( .A(IR_REG_13__SCAN_IN), .B(keyinput88), .ZN(n4736) );
  NAND4_X1 U5291 ( .A1(n4739), .A2(n4738), .A3(n4737), .A4(n4736), .ZN(n4742)
         );
  XNOR2_X1 U5292 ( .A(n4740), .B(keyinput46), .ZN(n4741) );
  NOR2_X1 U5293 ( .A1(n4742), .A2(n4741), .ZN(n4788) );
  AOI22_X1 U5294 ( .A1(n4745), .A2(keyinput108), .B1(n4744), .B2(keyinput91), 
        .ZN(n4743) );
  OAI221_X1 U5295 ( .B1(n4745), .B2(keyinput108), .C1(n4744), .C2(keyinput91), 
        .A(n4743), .ZN(n4758) );
  AOI22_X1 U5296 ( .A1(n4748), .A2(keyinput41), .B1(n4747), .B2(keyinput43), 
        .ZN(n4746) );
  OAI221_X1 U5297 ( .B1(n4748), .B2(keyinput41), .C1(n4747), .C2(keyinput43), 
        .A(n4746), .ZN(n4757) );
  AOI22_X1 U5298 ( .A1(n4751), .A2(keyinput66), .B1(n4750), .B2(keyinput8), 
        .ZN(n4749) );
  OAI221_X1 U5299 ( .B1(n4751), .B2(keyinput66), .C1(n4750), .C2(keyinput8), 
        .A(n4749), .ZN(n4756) );
  AOI22_X1 U5300 ( .A1(n4754), .A2(keyinput76), .B1(n4753), .B2(keyinput65), 
        .ZN(n4752) );
  OAI221_X1 U5301 ( .B1(n4754), .B2(keyinput76), .C1(n4753), .C2(keyinput65), 
        .A(n4752), .ZN(n4755) );
  NOR4_X1 U5302 ( .A1(n4758), .A2(n4757), .A3(n4756), .A4(n4755), .ZN(n4787)
         );
  AOI22_X1 U5303 ( .A1(n4761), .A2(keyinput112), .B1(n4760), .B2(keyinput89), 
        .ZN(n4759) );
  OAI221_X1 U5304 ( .B1(n4761), .B2(keyinput112), .C1(n4760), .C2(keyinput89), 
        .A(n4759), .ZN(n4771) );
  AOI22_X1 U5305 ( .A1(n2461), .A2(keyinput1), .B1(keyinput44), .B2(n4763), 
        .ZN(n4762) );
  OAI221_X1 U5306 ( .B1(n2461), .B2(keyinput1), .C1(n4763), .C2(keyinput44), 
        .A(n4762), .ZN(n4770) );
  INV_X1 U5307 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4765) );
  AOI22_X1 U5308 ( .A1(n2482), .A2(keyinput13), .B1(n4765), .B2(keyinput49), 
        .ZN(n4764) );
  OAI221_X1 U5309 ( .B1(n2482), .B2(keyinput13), .C1(n4765), .C2(keyinput49), 
        .A(n4764), .ZN(n4769) );
  INV_X1 U5310 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4767) );
  AOI22_X1 U5311 ( .A1(n3448), .A2(keyinput36), .B1(keyinput28), .B2(n4767), 
        .ZN(n4766) );
  OAI221_X1 U5312 ( .B1(n3448), .B2(keyinput36), .C1(n4767), .C2(keyinput28), 
        .A(n4766), .ZN(n4768) );
  NOR4_X1 U5313 ( .A1(n4771), .A2(n4770), .A3(n4769), .A4(n4768), .ZN(n4786)
         );
  AOI22_X1 U5314 ( .A1(n4774), .A2(keyinput30), .B1(n4773), .B2(keyinput7), 
        .ZN(n4772) );
  OAI221_X1 U5315 ( .B1(n4774), .B2(keyinput30), .C1(n4773), .C2(keyinput7), 
        .A(n4772), .ZN(n4784) );
  AOI22_X1 U5316 ( .A1(n4416), .A2(keyinput119), .B1(n4403), .B2(keyinput3), 
        .ZN(n4775) );
  OAI221_X1 U5317 ( .B1(n4416), .B2(keyinput119), .C1(n4403), .C2(keyinput3), 
        .A(n4775), .ZN(n4783) );
  AOI22_X1 U5318 ( .A1(n4778), .A2(keyinput17), .B1(n4777), .B2(keyinput85), 
        .ZN(n4776) );
  OAI221_X1 U5319 ( .B1(n4778), .B2(keyinput17), .C1(n4777), .C2(keyinput85), 
        .A(n4776), .ZN(n4782) );
  AOI22_X1 U5320 ( .A1(n4780), .A2(keyinput80), .B1(keyinput111), .B2(n2801), 
        .ZN(n4779) );
  OAI221_X1 U5321 ( .B1(n4780), .B2(keyinput80), .C1(n2801), .C2(keyinput111), 
        .A(n4779), .ZN(n4781) );
  NOR4_X1 U5322 ( .A1(n4784), .A2(n4783), .A3(n4782), .A4(n4781), .ZN(n4785)
         );
  NAND4_X1 U5323 ( .A1(n4788), .A2(n4787), .A3(n4786), .A4(n4785), .ZN(n4917)
         );
  AOI22_X1 U5324 ( .A1(n4791), .A2(keyinput79), .B1(keyinput54), .B2(n4790), 
        .ZN(n4789) );
  OAI221_X1 U5325 ( .B1(n4791), .B2(keyinput79), .C1(n4790), .C2(keyinput54), 
        .A(n4789), .ZN(n4804) );
  AOI22_X1 U5326 ( .A1(n4794), .A2(keyinput114), .B1(keyinput11), .B2(n4793), 
        .ZN(n4792) );
  OAI221_X1 U5327 ( .B1(n4794), .B2(keyinput114), .C1(n4793), .C2(keyinput11), 
        .A(n4792), .ZN(n4803) );
  INV_X1 U5328 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4796) );
  AOI22_X1 U5329 ( .A1(n4797), .A2(keyinput37), .B1(keyinput127), .B2(n4796), 
        .ZN(n4795) );
  OAI221_X1 U5330 ( .B1(n4797), .B2(keyinput37), .C1(n4796), .C2(keyinput127), 
        .A(n4795), .ZN(n4802) );
  XOR2_X1 U5331 ( .A(n4798), .B(keyinput104), .Z(n4800) );
  XNOR2_X1 U5332 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput122), .ZN(n4799) );
  NAND2_X1 U5333 ( .A1(n4800), .A2(n4799), .ZN(n4801) );
  NOR4_X1 U5334 ( .A1(n4804), .A2(n4803), .A3(n4802), .A4(n4801), .ZN(n4849)
         );
  AOI22_X1 U5335 ( .A1(n3459), .A2(keyinput123), .B1(keyinput32), .B2(n4806), 
        .ZN(n4805) );
  OAI221_X1 U5336 ( .B1(n3459), .B2(keyinput123), .C1(n4806), .C2(keyinput32), 
        .A(n4805), .ZN(n4818) );
  AOI22_X1 U5337 ( .A1(n4809), .A2(keyinput86), .B1(keyinput39), .B2(n4808), 
        .ZN(n4807) );
  OAI221_X1 U5338 ( .B1(n4809), .B2(keyinput86), .C1(n4808), .C2(keyinput39), 
        .A(n4807), .ZN(n4817) );
  AOI22_X1 U5339 ( .A1(n4811), .A2(keyinput125), .B1(n4347), .B2(keyinput95), 
        .ZN(n4810) );
  OAI221_X1 U5340 ( .B1(n4811), .B2(keyinput125), .C1(n4347), .C2(keyinput95), 
        .A(n4810), .ZN(n4816) );
  AOI22_X1 U5341 ( .A1(n4814), .A2(keyinput72), .B1(keyinput102), .B2(n4813), 
        .ZN(n4812) );
  OAI221_X1 U5342 ( .B1(n4814), .B2(keyinput72), .C1(n4813), .C2(keyinput102), 
        .A(n4812), .ZN(n4815) );
  NOR4_X1 U5343 ( .A1(n4818), .A2(n4817), .A3(n4816), .A4(n4815), .ZN(n4848)
         );
  AOI22_X1 U5344 ( .A1(n4821), .A2(keyinput19), .B1(keyinput109), .B2(n4820), 
        .ZN(n4819) );
  OAI221_X1 U5345 ( .B1(n4821), .B2(keyinput19), .C1(n4820), .C2(keyinput109), 
        .A(n4819), .ZN(n4831) );
  AOI22_X1 U5346 ( .A1(n4033), .A2(keyinput27), .B1(n4823), .B2(keyinput50), 
        .ZN(n4822) );
  OAI221_X1 U5347 ( .B1(n4033), .B2(keyinput27), .C1(n4823), .C2(keyinput50), 
        .A(n4822), .ZN(n4830) );
  AOI22_X1 U5348 ( .A1(n3139), .A2(keyinput120), .B1(n4825), .B2(keyinput124), 
        .ZN(n4824) );
  OAI221_X1 U5349 ( .B1(n3139), .B2(keyinput120), .C1(n4825), .C2(keyinput124), 
        .A(n4824), .ZN(n4829) );
  AOI22_X1 U5350 ( .A1(n4827), .A2(keyinput5), .B1(n2214), .B2(keyinput24), 
        .ZN(n4826) );
  OAI221_X1 U5351 ( .B1(n4827), .B2(keyinput5), .C1(n2214), .C2(keyinput24), 
        .A(n4826), .ZN(n4828) );
  NOR4_X1 U5352 ( .A1(n4831), .A2(n4830), .A3(n4829), .A4(n4828), .ZN(n4847)
         );
  AOI22_X1 U5353 ( .A1(n2213), .A2(keyinput62), .B1(n4833), .B2(keyinput20), 
        .ZN(n4832) );
  OAI221_X1 U5354 ( .B1(n2213), .B2(keyinput62), .C1(n4833), .C2(keyinput20), 
        .A(n4832), .ZN(n4845) );
  INV_X1 U5355 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4835) );
  AOI22_X1 U5356 ( .A1(n4836), .A2(keyinput38), .B1(keyinput101), .B2(n4835), 
        .ZN(n4834) );
  OAI221_X1 U5357 ( .B1(n4836), .B2(keyinput38), .C1(n4835), .C2(keyinput101), 
        .A(n4834), .ZN(n4844) );
  AOI22_X1 U5358 ( .A1(n4839), .A2(keyinput51), .B1(keyinput42), .B2(n4838), 
        .ZN(n4837) );
  OAI221_X1 U5359 ( .B1(n4839), .B2(keyinput51), .C1(n4838), .C2(keyinput42), 
        .A(n4837), .ZN(n4843) );
  AOI22_X1 U5360 ( .A1(n4093), .A2(keyinput55), .B1(keyinput0), .B2(n4841), 
        .ZN(n4840) );
  OAI221_X1 U5361 ( .B1(n4093), .B2(keyinput55), .C1(n4841), .C2(keyinput0), 
        .A(n4840), .ZN(n4842) );
  NOR4_X1 U5362 ( .A1(n4845), .A2(n4844), .A3(n4843), .A4(n4842), .ZN(n4846)
         );
  NAND4_X1 U5363 ( .A1(n4849), .A2(n4848), .A3(n4847), .A4(n4846), .ZN(n4916)
         );
  OAI22_X1 U5364 ( .A1(keyinput83), .A2(n4852), .B1(n4851), .B2(keyinput16), 
        .ZN(n4850) );
  AOI221_X1 U5365 ( .B1(n4852), .B2(keyinput83), .C1(n4851), .C2(keyinput16), 
        .A(n4850), .ZN(n4914) );
  XOR2_X1 U5366 ( .A(keyinput4), .B(ADDR_REG_7__SCAN_IN), .Z(n4862) );
  XOR2_X1 U5367 ( .A(keyinput64), .B(ADDR_REG_10__SCAN_IN), .Z(n4861) );
  INV_X1 U5368 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4855) );
  INV_X1 U5369 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4854) );
  AOI22_X1 U5370 ( .A1(n4855), .A2(keyinput10), .B1(keyinput99), .B2(n4854), 
        .ZN(n4853) );
  OAI221_X1 U5371 ( .B1(n4855), .B2(keyinput10), .C1(n4854), .C2(keyinput99), 
        .A(n4853), .ZN(n4860) );
  AOI22_X1 U5372 ( .A1(n4858), .A2(keyinput33), .B1(keyinput105), .B2(n4857), 
        .ZN(n4856) );
  OAI221_X1 U5373 ( .B1(n4858), .B2(keyinput33), .C1(n4857), .C2(keyinput105), 
        .A(n4856), .ZN(n4859) );
  NOR4_X1 U5374 ( .A1(n4862), .A2(n4861), .A3(n4860), .A4(n4859), .ZN(n4913)
         );
  AOI22_X1 U5375 ( .A1(n4865), .A2(keyinput71), .B1(n4864), .B2(keyinput26), 
        .ZN(n4863) );
  OAI221_X1 U5376 ( .B1(n4865), .B2(keyinput71), .C1(n4864), .C2(keyinput26), 
        .A(n4863), .ZN(n4877) );
  AOI22_X1 U5377 ( .A1(n4868), .A2(keyinput59), .B1(n4867), .B2(keyinput25), 
        .ZN(n4866) );
  OAI221_X1 U5378 ( .B1(n4868), .B2(keyinput59), .C1(n4867), .C2(keyinput25), 
        .A(n4866), .ZN(n4876) );
  INV_X1 U5379 ( .A(keyinput14), .ZN(n4870) );
  AOI22_X1 U5380 ( .A1(n4871), .A2(keyinput106), .B1(DATAO_REG_31__SCAN_IN), 
        .B2(n4870), .ZN(n4869) );
  OAI221_X1 U5381 ( .B1(n4871), .B2(keyinput106), .C1(n4870), .C2(
        DATAO_REG_31__SCAN_IN), .A(n4869), .ZN(n4875) );
  XOR2_X1 U5382 ( .A(n3729), .B(keyinput118), .Z(n4873) );
  XNOR2_X1 U5383 ( .A(IR_REG_30__SCAN_IN), .B(keyinput113), .ZN(n4872) );
  NAND2_X1 U5384 ( .A1(n4873), .A2(n4872), .ZN(n4874) );
  NOR4_X1 U5385 ( .A1(n4877), .A2(n4876), .A3(n4875), .A4(n4874), .ZN(n4912)
         );
  XOR2_X1 U5386 ( .A(keyinput52), .B(ADDR_REG_0__SCAN_IN), .Z(n4910) );
  XNOR2_X1 U5387 ( .A(keyinput69), .B(n4878), .ZN(n4909) );
  OAI22_X1 U5388 ( .A1(keyinput70), .A2(n4881), .B1(n4880), .B2(keyinput2), 
        .ZN(n4879) );
  AOI221_X1 U5389 ( .B1(n4881), .B2(keyinput70), .C1(n4880), .C2(keyinput2), 
        .A(n4879), .ZN(n4890) );
  OAI22_X1 U5390 ( .A1(keyinput87), .A2(n4884), .B1(n4883), .B2(keyinput97), 
        .ZN(n4882) );
  AOI221_X1 U5391 ( .B1(n4884), .B2(keyinput87), .C1(n4883), .C2(keyinput97), 
        .A(n4882), .ZN(n4889) );
  XOR2_X1 U5392 ( .A(keyinput56), .B(n4885), .Z(n4888) );
  XOR2_X1 U5393 ( .A(keyinput107), .B(n4886), .Z(n4887) );
  NAND4_X1 U5394 ( .A1(n4890), .A2(n4889), .A3(n4888), .A4(n4887), .ZN(n4908)
         );
  OAI22_X1 U5395 ( .A1(n4893), .A2(keyinput93), .B1(n4892), .B2(keyinput90), 
        .ZN(n4891) );
  AOI221_X1 U5396 ( .B1(n4893), .B2(keyinput93), .C1(keyinput90), .C2(n4892), 
        .A(n4891), .ZN(n4906) );
  INV_X1 U5397 ( .A(keyinput94), .ZN(n4895) );
  OAI22_X1 U5398 ( .A1(keyinput103), .A2(n4896), .B1(n4895), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4894) );
  AOI221_X1 U5399 ( .B1(n4896), .B2(keyinput103), .C1(n4895), .C2(
        DATAO_REG_25__SCAN_IN), .A(n4894), .ZN(n4905) );
  OAI22_X1 U5400 ( .A1(keyinput110), .A2(n4899), .B1(n4898), .B2(keyinput77), 
        .ZN(n4897) );
  AOI221_X1 U5401 ( .B1(n4899), .B2(keyinput110), .C1(n4898), .C2(keyinput77), 
        .A(n4897), .ZN(n4904) );
  OAI22_X1 U5402 ( .A1(keyinput9), .A2(n4902), .B1(n4901), .B2(keyinput63), 
        .ZN(n4900) );
  AOI221_X1 U5403 ( .B1(n4902), .B2(keyinput9), .C1(n4901), .C2(keyinput63), 
        .A(n4900), .ZN(n4903) );
  NAND4_X1 U5404 ( .A1(n4906), .A2(n4905), .A3(n4904), .A4(n4903), .ZN(n4907)
         );
  NOR4_X1 U5405 ( .A1(n4910), .A2(n4909), .A3(n4908), .A4(n4907), .ZN(n4911)
         );
  NAND4_X1 U5406 ( .A1(n4914), .A2(n4913), .A3(n4912), .A4(n4911), .ZN(n4915)
         );
  NOR4_X1 U5407 ( .A1(n4918), .A2(n4917), .A3(n4916), .A4(n4915), .ZN(n4919)
         );
  XOR2_X1 U5408 ( .A(n4920), .B(n4919), .Z(n4921) );
  XNOR2_X1 U5409 ( .A(n4922), .B(n4921), .ZN(U3286) );
  CLKBUF_X1 U2394 ( .A(n3027), .Z(n3620) );
  CLKBUF_X1 U2421 ( .A(n2447), .Z(n2948) );
  OAI211_X1 U2456 ( .C1(n2449), .C2(n2363), .A(n2451), .B(n2362), .ZN(n4006)
         );
  OAI211_X1 U2611 ( .C1(n4247), .C2(n2142), .A(n2653), .B(n2652), .ZN(n4925)
         );
  BUF_X2 U2993 ( .A(n2468), .Z(n2142) );
endmodule

