

module b17_C_gen_AntiSAT_k_256_2 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, 
        keyinput_f65, keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, 
        keyinput_f70, keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, 
        keyinput_f75, keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, 
        keyinput_f80, keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, 
        keyinput_f85, keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, 
        keyinput_f90, keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, 
        keyinput_f95, keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, 
        keyinput_f100, keyinput_f101, keyinput_f102, keyinput_f103, 
        keyinput_f104, keyinput_f105, keyinput_f106, keyinput_f107, 
        keyinput_f108, keyinput_f109, keyinput_f110, keyinput_f111, 
        keyinput_f112, keyinput_f113, keyinput_f114, keyinput_f115, 
        keyinput_f116, keyinput_f117, keyinput_f118, keyinput_f119, 
        keyinput_f120, keyinput_f121, keyinput_f122, keyinput_f123, 
        keyinput_f124, keyinput_f125, keyinput_f126, keyinput_f127, 
        keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, 
        keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, 
        keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, 
        keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, 
        keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, 
        keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, 
        keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, 
        keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, 
        keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, 
        keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, 
        keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, 
        keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, 
        keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, keyinput_g64, 
        keyinput_g65, keyinput_g66, keyinput_g67, keyinput_g68, keyinput_g69, 
        keyinput_g70, keyinput_g71, keyinput_g72, keyinput_g73, keyinput_g74, 
        keyinput_g75, keyinput_g76, keyinput_g77, keyinput_g78, keyinput_g79, 
        keyinput_g80, keyinput_g81, keyinput_g82, keyinput_g83, keyinput_g84, 
        keyinput_g85, keyinput_g86, keyinput_g87, keyinput_g88, keyinput_g89, 
        keyinput_g90, keyinput_g91, keyinput_g92, keyinput_g93, keyinput_g94, 
        keyinput_g95, keyinput_g96, keyinput_g97, keyinput_g98, keyinput_g99, 
        keyinput_g100, keyinput_g101, keyinput_g102, keyinput_g103, 
        keyinput_g104, keyinput_g105, keyinput_g106, keyinput_g107, 
        keyinput_g108, keyinput_g109, keyinput_g110, keyinput_g111, 
        keyinput_g112, keyinput_g113, keyinput_g114, keyinput_g115, 
        keyinput_g116, keyinput_g117, keyinput_g118, keyinput_g119, 
        keyinput_g120, keyinput_g121, keyinput_g122, keyinput_g123, 
        keyinput_g124, keyinput_g125, keyinput_g126, keyinput_g127, U355, U356, 
        U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, 
        U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, 
        U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, 
        U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, 
        U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, 
        U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, 
        U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, 
        U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, 
        P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, 
        P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, 
        P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, 
        P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, 
        P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, 
        P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, 
        P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, 
        P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, 
        P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, 
        P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, 
        P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, 
        P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, 
        P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, 
        P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, 
        P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, 
        P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, 
        P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, 
        P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, 
        P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, 
        P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, 
        P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, 
        P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, 
        P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, 
        P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, 
        P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, 
        P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, 
        P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, 
        P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, 
        P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, 
        P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, 
        P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, 
        P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, 
        P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, 
        P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, 
        P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, 
        P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, 
        P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, 
        P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, 
        P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, 
        P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, 
        P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, 
        P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, 
        P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, 
        P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, 
        P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, 
        P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, 
        P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, 
        P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, 
        P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, 
        P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, 
        P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, 
        P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, 
        P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, 
        P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, 
        P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, 
        P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, 
        P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, 
        P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, 
        P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, 
        P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, 
        P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, 
        P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, 
        P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, 
        P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, 
        P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, 
        P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, 
        P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, 
        P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, 
        P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, 
        P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, 
        P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, 
        P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, 
        P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, 
        P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, 
        P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, 
        P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, 
        P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, 
        P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, 
        P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, 
        P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, 
        P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, 
        P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, 
        P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, 
        P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, 
        P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, 
        P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, 
        P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, 
        P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, 
        P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, 
        P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, 
        P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, 
        P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, 
        P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, 
        P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, 
        P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, 
        P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, 
        P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, 
        P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, 
        P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, 
        P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, 
        P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, 
        P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, 
        P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, 
        P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, 
        P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, 
        P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, 
        P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, 
        P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, 
        P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, 
        P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, 
        P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, 
        P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, 
        P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, 
        P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, 
        P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, 
        P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, 
        P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, 
        P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, 
        P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, 
        P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, 
        P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, 
        P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, 
        P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, 
        P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, 
        P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, 
        P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, 
        P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, 
        P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, 
        P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, 
        P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, 
        P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, 
        P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, 
        P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, 
        P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, 
        P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, 
        P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, 
        P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, 
        P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, 
        P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, 
        P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, 
        P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, 
        P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, 
        P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, 
        P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, 
        P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, 
        P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, 
        P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, 
        P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, 
        P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, 
        P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, 
        P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, 
        P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, 
        P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, 
        P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, 
        P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, 
        P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, 
        P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, 
        P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, 
        P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, 
        P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, 
        P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, 
        P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, 
        P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, 
        P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, 
        P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, 
        P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, 
        P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, 
        P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, 
        P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, 
        P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, 
        P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, 
        P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, 
        P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, 
        P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, 
        P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, 
        P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, 
        P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, 
        P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, 
        P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, 
        P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
         n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
         n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168,
         n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,
         n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
         n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192,
         n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,
         n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
         n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216,
         n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,
         n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,
         n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240,
         n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
         n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,
         n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264,
         n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
         n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
         n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288,
         n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,
         n21297, n21298, n21299, n21300, n21301, n21302, n21303;

  NOR2_X1 U11241 ( .A1(n14626), .A2(n14625), .ZN(n14897) );
  BUF_X1 U11242 ( .A(n14610), .Z(n14626) );
  OR2_X2 U11243 ( .A1(n12704), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12853) );
  CLKBUF_X1 U11244 ( .A(n17096), .Z(n9807) );
  INV_X1 U11245 ( .A(n18002), .ZN(n17969) );
  INV_X2 U11246 ( .A(n9844), .ZN(n16068) );
  CLKBUF_X2 U11247 ( .A(n9846), .Z(n9804) );
  OR2_X1 U11248 ( .A1(n10658), .A2(n10651), .ZN(n19472) );
  OR2_X1 U11249 ( .A1(n10660), .A2(n10659), .ZN(n19668) );
  NAND2_X1 U11250 ( .A1(n9950), .A2(n9953), .ZN(n19736) );
  NAND2_X1 U11251 ( .A1(n9954), .A2(n9953), .ZN(n19622) );
  OR2_X2 U11252 ( .A1(n10658), .A2(n10659), .ZN(n13669) );
  BUF_X1 U11253 ( .A(n10641), .Z(n12888) );
  NAND2_X1 U11254 ( .A1(n12966), .A2(n12967), .ZN(n13576) );
  INV_X1 U11255 ( .A(n11496), .ZN(n14036) );
  AND2_X1 U11258 ( .A1(n12066), .A2(n12883), .ZN(n10776) );
  BUF_X1 U11259 ( .A(n11399), .Z(n11882) );
  AND2_X1 U11260 ( .A1(n12063), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10774) );
  AND2_X1 U11261 ( .A1(n12065), .A2(n12883), .ZN(n10798) );
  NAND4_X1 U11262 ( .A1(n13005), .A2(n12440), .A3(n13007), .A4(n13019), .ZN(
        n12449) );
  INV_X4 U11263 ( .A(n17321), .ZN(n11667) );
  CLKBUF_X2 U11264 ( .A(n11477), .Z(n17433) );
  BUF_X1 U11265 ( .A(n12387), .Z(n15164) );
  OR2_X1 U11266 ( .A1(n20254), .A2(n13364), .ZN(n20905) );
  CLKBUF_X2 U11267 ( .A(n12261), .Z(n12492) );
  NAND3_X1 U11268 ( .A1(n17094), .A2(n10145), .A3(n19050), .ZN(n17441) );
  AND2_X1 U11270 ( .A1(n19451), .A2(n10461), .ZN(n10550) );
  INV_X2 U11272 ( .A(n17426), .ZN(n11629) );
  INV_X2 U11273 ( .A(n10412), .ZN(n17442) );
  CLKBUF_X2 U11275 ( .A(n12250), .Z(n20280) );
  AND2_X1 U11276 ( .A1(n15173), .A2(n12193), .ZN(n12648) );
  AND2_X1 U11277 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13192) );
  NAND2_X1 U11278 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10226) );
  CLKBUF_X1 U11279 ( .A(n14491), .Z(n9797) );
  AOI21_X1 U11280 ( .B1(n15439), .B2(n11751), .A(n10167), .ZN(n14491) );
  NAND2_X1 U11281 ( .A1(n12443), .A2(n15164), .ZN(n12461) );
  INV_X1 U11282 ( .A(n20260), .ZN(n12993) );
  AND2_X1 U11283 ( .A1(n12490), .A2(n12488), .ZN(n12740) );
  CLKBUF_X1 U11284 ( .A(n10668), .Z(n9802) );
  AND2_X1 U11285 ( .A1(n12199), .A2(n12205), .ZN(n12647) );
  CLKBUF_X2 U11286 ( .A(n10616), .Z(n14468) );
  OR2_X1 U11287 ( .A1(n10652), .A2(n10659), .ZN(n19795) );
  BUF_X1 U11288 ( .A(n10842), .Z(n9799) );
  INV_X2 U11289 ( .A(n17441), .ZN(n11665) );
  AOI21_X1 U11290 ( .B1(n14607), .B2(n9798), .A(n14702), .ZN(n14649) );
  INV_X1 U11291 ( .A(n20133), .ZN(n15998) );
  NAND2_X1 U11292 ( .A1(n13113), .A2(n20285), .ZN(n14446) );
  NAND2_X1 U11293 ( .A1(n12907), .A2(n13118), .ZN(n10569) );
  INV_X2 U11294 ( .A(n10990), .ZN(n11251) );
  OR2_X1 U11295 ( .A1(n10652), .A2(n10651), .ZN(n13124) );
  INV_X2 U11296 ( .A(n12181), .ZN(n13118) );
  INV_X1 U11297 ( .A(n17848), .ZN(n17814) );
  INV_X1 U11298 ( .A(n20140), .ZN(n20158) );
  INV_X1 U11300 ( .A(n11253), .ZN(n12907) );
  INV_X2 U11301 ( .A(n17372), .ZN(n17437) );
  NAND2_X1 U11302 ( .A1(n11729), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18295) );
  NOR2_X2 U11303 ( .A1(n18448), .A2(n18334), .ZN(n18867) );
  INV_X1 U11304 ( .A(n10430), .ZN(n18478) );
  INV_X1 U11305 ( .A(n13098), .ZN(n13097) );
  OAI21_X1 U11306 ( .B1(n14626), .B2(n14612), .A(n14611), .ZN(n14888) );
  INV_X1 U11307 ( .A(n17092), .ZN(n17127) );
  NAND2_X2 U11308 ( .A1(n13169), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12733) );
  NOR2_X4 U11309 ( .A1(n10952), .A2(n10925), .ZN(n10940) );
  INV_X2 U11310 ( .A(n15492), .ZN(n15476) );
  INV_X2 U11311 ( .A(n17096), .ZN(n17116) );
  NAND2_X2 U11312 ( .A1(n10098), .A2(n11649), .ZN(n17637) );
  AND2_X2 U11313 ( .A1(n13617), .A2(n13783), .ZN(n9844) );
  AND2_X4 U11314 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11055) );
  AOI211_X4 U11315 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n11659), .B(n11658), .ZN(n17625) );
  OAI21_X2 U11316 ( .B1(n15829), .B2(n10310), .A(n10307), .ZN(n15598) );
  NOR2_X2 U11317 ( .A1(n18107), .A2(n17613), .ZN(n18012) );
  AOI211_X2 U11318 ( .C1(n15703), .C2(n15725), .A(n15731), .B(n15702), .ZN(
        n15720) );
  BUF_X4 U11319 ( .A(n12262), .Z(n9800) );
  INV_X1 U11320 ( .A(n14408), .ZN(n12262) );
  NOR2_X2 U11321 ( .A1(n18104), .A2(n18089), .ZN(n17819) );
  INV_X1 U11322 ( .A(n18103), .ZN(n18089) );
  BUF_X1 U11323 ( .A(n10668), .Z(n9801) );
  OAI21_X1 U11324 ( .B1(n10139), .B2(n9836), .A(n10417), .ZN(n14892) );
  OR2_X1 U11325 ( .A1(n12004), .A2(n12003), .ZN(n9993) );
  NAND2_X1 U11326 ( .A1(n15309), .A2(n15311), .ZN(n15310) );
  NOR2_X1 U11327 ( .A1(n19557), .A2(n19596), .ZN(n19612) );
  OR2_X1 U11328 ( .A1(n16090), .A2(n16141), .ZN(n16066) );
  INV_X2 U11329 ( .A(n18249), .ZN(n17897) );
  NAND2_X1 U11330 ( .A1(n18016), .A2(n11701), .ZN(n11729) );
  NAND2_X1 U11331 ( .A1(n19079), .A2(n18920), .ZN(n16753) );
  NOR2_X2 U11333 ( .A1(n18878), .A2(n18890), .ZN(n18317) );
  INV_X4 U11334 ( .A(n18304), .ZN(n18898) );
  OAI21_X1 U11335 ( .B1(n9873), .B2(n10156), .A(n11577), .ZN(n18304) );
  NAND2_X1 U11336 ( .A1(n20356), .A2(n12740), .ZN(n12743) );
  CLKBUF_X1 U11337 ( .A(n12415), .Z(n12424) );
  NOR2_X1 U11338 ( .A1(n16794), .A2(n16608), .ZN(n16607) );
  BUF_X1 U11339 ( .A(n17685), .Z(n9810) );
  INV_X1 U11340 ( .A(n10595), .ZN(n11168) );
  CLKBUF_X1 U11341 ( .A(n12426), .Z(n12455) );
  INV_X1 U11342 ( .A(n18441), .ZN(n17081) );
  AOI211_X1 U11343 ( .C1(n11667), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n11696), .B(n11695), .ZN(n17618) );
  NAND2_X1 U11344 ( .A1(n10569), .A2(n13477), .ZN(n11116) );
  BUF_X1 U11345 ( .A(n10567), .Z(n12079) );
  INV_X1 U11346 ( .A(n11048), .ZN(n10558) );
  CLKBUF_X1 U11347 ( .A(n11752), .Z(n10495) );
  NAND2_X1 U11348 ( .A1(n10447), .A2(n10448), .ZN(n10496) );
  NAND2_X1 U11349 ( .A1(n10511), .A2(n10510), .ZN(n12181) );
  INV_X4 U11350 ( .A(n17438), .ZN(n17415) );
  AND2_X2 U11351 ( .A1(n12058), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11818) );
  NAND2_X1 U11352 ( .A1(n11464), .A2(n10078), .ZN(n17416) );
  CLKBUF_X2 U11353 ( .A(n10529), .Z(n12058) );
  CLKBUF_X2 U11354 ( .A(n14420), .Z(n14352) );
  CLKBUF_X2 U11355 ( .A(n12648), .Z(n14419) );
  INV_X1 U11356 ( .A(n12733), .ZN(n9809) );
  AND2_X1 U11357 ( .A1(n12192), .A2(n13193), .ZN(n12267) );
  CLKBUF_X2 U11358 ( .A(n10530), .Z(n12063) );
  INV_X4 U11359 ( .A(n11517), .ZN(n9803) );
  CLKBUF_X2 U11360 ( .A(n10669), .Z(n12059) );
  CLKBUF_X2 U11361 ( .A(n12236), .Z(n14240) );
  AND2_X1 U11362 ( .A1(n10105), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10145) );
  NOR2_X1 U11363 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12205) );
  OAI211_X1 U11364 ( .C1(n12025), .C2(n10390), .A(n10387), .B(n10385), .ZN(
        n12124) );
  NOR2_X1 U11365 ( .A1(n14882), .A2(n10137), .ZN(n14883) );
  NAND2_X1 U11366 ( .A1(n12025), .A2(n10388), .ZN(n10387) );
  NOR2_X1 U11367 ( .A1(n10139), .A2(n9905), .ZN(n10137) );
  AND2_X1 U11368 ( .A1(n10139), .A2(n10138), .ZN(n14882) );
  NAND2_X1 U11369 ( .A1(n9993), .A2(n15295), .ZN(n9992) );
  AND2_X1 U11370 ( .A1(n14623), .A2(n14624), .ZN(n14625) );
  NAND2_X1 U11371 ( .A1(n12004), .A2(n12003), .ZN(n15288) );
  AOI21_X1 U11372 ( .B1(n15450), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15452) );
  NAND2_X1 U11373 ( .A1(n15302), .A2(n10423), .ZN(n12004) );
  NOR2_X1 U11374 ( .A1(n14948), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14933) );
  OR2_X1 U11375 ( .A1(n11980), .A2(n11979), .ZN(n10423) );
  INV_X1 U11376 ( .A(n14070), .ZN(n10017) );
  NOR2_X1 U11377 ( .A1(n15584), .A2(n15689), .ZN(n15570) );
  NAND2_X1 U11378 ( .A1(n15310), .A2(n11954), .ZN(n11978) );
  NAND2_X1 U11379 ( .A1(n10018), .A2(n9865), .ZN(n14070) );
  NAND2_X1 U11380 ( .A1(n14065), .A2(n14066), .ZN(n10144) );
  NAND2_X1 U11381 ( .A1(n16443), .A2(n9935), .ZN(n15723) );
  INV_X1 U11382 ( .A(n9986), .ZN(n11952) );
  CLKBUF_X1 U11383 ( .A(n14999), .Z(n16089) );
  OAI21_X1 U11384 ( .B1(n10023), .B2(n10021), .A(n10019), .ZN(n14999) );
  AND2_X1 U11385 ( .A1(n14072), .A2(n13917), .ZN(n13919) );
  AND2_X1 U11386 ( .A1(n16790), .A2(n9807), .ZN(n16781) );
  AND2_X1 U11387 ( .A1(n16043), .A2(n14057), .ZN(n14061) );
  OR2_X1 U11388 ( .A1(n16792), .A2(n16793), .ZN(n16790) );
  AND2_X1 U11389 ( .A1(n16066), .A2(n14056), .ZN(n16043) );
  NOR2_X1 U11390 ( .A1(n19733), .A2(n20034), .ZN(n19783) );
  INV_X1 U11391 ( .A(n15430), .ZN(n10262) );
  OAI21_X1 U11392 ( .B1(n13154), .B2(n13153), .A(n11086), .ZN(n13509) );
  NAND2_X1 U11393 ( .A1(n10786), .A2(n11102), .ZN(n11076) );
  OR2_X1 U11394 ( .A1(n14736), .A2(n14541), .ZN(n14702) );
  INV_X2 U11395 ( .A(n9844), .ZN(n16090) );
  NOR2_X1 U11396 ( .A1(n10960), .A2(n15522), .ZN(n10053) );
  OR2_X1 U11397 ( .A1(n10785), .A2(n10784), .ZN(n10786) );
  NAND2_X1 U11398 ( .A1(n17927), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18246) );
  OAI21_X1 U11399 ( .B1(n20883), .B2(n10037), .A(n13335), .ZN(n13336) );
  NAND2_X1 U11400 ( .A1(n13254), .A2(n13433), .ZN(n20883) );
  NAND2_X1 U11401 ( .A1(n14652), .A2(n14637), .ZN(n14639) );
  NOR2_X2 U11402 ( .A1(n19042), .A2(n18098), .ZN(n17952) );
  AOI21_X1 U11403 ( .B1(n13409), .B2(n14128), .A(n13408), .ZN(n13452) );
  NAND4_X1 U11404 ( .A1(n10703), .A2(n10702), .A3(n10701), .A4(n10700), .ZN(
        n10739) );
  INV_X1 U11405 ( .A(n18012), .ZN(n17943) );
  NOR2_X2 U11406 ( .A1(n18295), .A2(n18239), .ZN(n17924) );
  INV_X1 U11407 ( .A(n18040), .ZN(n18108) );
  OAI21_X2 U11408 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19078), .A(n16753), 
        .ZN(n18103) );
  NAND2_X1 U11409 ( .A1(n13253), .A2(n9864), .ZN(n13572) );
  NAND2_X1 U11410 ( .A1(n10973), .A2(n10974), .ZN(n10985) );
  AND2_X1 U11411 ( .A1(n12687), .A2(n11778), .ZN(n9983) );
  AOI21_X1 U11412 ( .B1(n18004), .B2(n9845), .A(n10106), .ZN(n18278) );
  OAI22_X1 U11413 ( .A1(n11908), .A2(n13124), .B1(n19881), .B2(n10696), .ZN(
        n10699) );
  OR2_X2 U11414 ( .A1(n10649), .A2(n10651), .ZN(n19592) );
  NAND2_X1 U11415 ( .A1(n18017), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18016) );
  NAND2_X1 U11416 ( .A1(n11758), .A2(n11757), .ZN(n11768) );
  XNOR2_X1 U11417 ( .A(n17967), .B(n11700), .ZN(n18017) );
  AOI21_X1 U11418 ( .B1(n12682), .B2(n12681), .A(n11767), .ZN(n12598) );
  AND2_X1 U11419 ( .A1(n12746), .A2(n12745), .ZN(n12972) );
  NOR2_X1 U11420 ( .A1(n20396), .A2(n20281), .ZN(n20779) );
  NOR2_X1 U11421 ( .A1(n20396), .A2(n20274), .ZN(n20774) );
  NOR2_X1 U11422 ( .A1(n20396), .A2(n20262), .ZN(n20762) );
  NOR2_X1 U11423 ( .A1(n20396), .A2(n20255), .ZN(n20756) );
  XNOR2_X1 U11424 ( .A(n15846), .B(n11765), .ZN(n12682) );
  NAND2_X1 U11425 ( .A1(n13251), .A2(n13250), .ZN(n20233) );
  NOR2_X1 U11426 ( .A1(n20396), .A2(n20297), .ZN(n20795) );
  NAND2_X1 U11427 ( .A1(n11761), .A2(n11760), .ZN(n15846) );
  NAND2_X1 U11428 ( .A1(n13348), .A2(n13347), .ZN(n13595) );
  AND2_X1 U11429 ( .A1(n12583), .A2(n12381), .ZN(n13348) );
  NAND2_X1 U11430 ( .A1(n18044), .A2(n11719), .ZN(n18035) );
  CLKBUF_X1 U11431 ( .A(n13216), .Z(n20702) );
  NOR2_X2 U11432 ( .A1(n19452), .A2(n19888), .ZN(n19453) );
  NOR2_X2 U11433 ( .A1(n19463), .A2(n19888), .ZN(n19464) );
  NAND2_X1 U11434 ( .A1(n18045), .A2(n18046), .ZN(n18044) );
  NOR2_X2 U11435 ( .A1(n19331), .A2(n19888), .ZN(n13305) );
  OR2_X1 U11436 ( .A1(n12975), .A2(n12974), .ZN(n12976) );
  NOR2_X2 U11437 ( .A1(n14459), .A2(n19459), .ZN(n13312) );
  NOR2_X2 U11438 ( .A1(n19322), .A2(n19888), .ZN(n13101) );
  NOR2_X2 U11439 ( .A1(n13682), .A2(n19459), .ZN(n13683) );
  NOR2_X2 U11440 ( .A1(n19440), .A2(n19888), .ZN(n19441) );
  XNOR2_X1 U11441 ( .A(n12720), .B(n12719), .ZN(n20329) );
  NOR2_X2 U11442 ( .A1(n19358), .A2(n19888), .ZN(n13681) );
  NOR2_X2 U11443 ( .A1(n19446), .A2(n19888), .ZN(n19447) );
  NOR2_X2 U11444 ( .A1(n19368), .A2(n19888), .ZN(n13117) );
  NAND2_X1 U11445 ( .A1(n12722), .A2(n12721), .ZN(n12975) );
  NAND2_X1 U11446 ( .A1(n10584), .A2(n10583), .ZN(n10622) );
  NAND2_X1 U11447 ( .A1(n12743), .A2(n12470), .ZN(n12954) );
  NAND2_X1 U11448 ( .A1(n18062), .A2(n11718), .ZN(n18045) );
  OAI211_X1 U11449 ( .C1(n20246), .C2(n12704), .A(n12477), .B(n12476), .ZN(
        n12953) );
  AND2_X1 U11450 ( .A1(n10586), .A2(n10585), .ZN(n10624) );
  NOR2_X2 U11451 ( .A1(n11739), .A2(n16645), .ZN(n18002) );
  AOI21_X1 U11452 ( .B1(n10630), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10633), .ZN(n11151) );
  NOR2_X2 U11453 ( .A1(n19084), .A2(n17747), .ZN(n17739) );
  OAI211_X1 U11454 ( .C1(n11566), .C2(n11574), .A(n13955), .B(n13954), .ZN(
        n11570) );
  OR2_X2 U11455 ( .A1(n18923), .A2(n17683), .ZN(n17749) );
  OR2_X1 U11456 ( .A1(n15270), .A2(n15269), .ZN(n15272) );
  AND2_X1 U11457 ( .A1(n10088), .A2(n10085), .ZN(n13955) );
  NAND2_X1 U11458 ( .A1(n10554), .A2(n10553), .ZN(n10598) );
  INV_X1 U11459 ( .A(n10589), .ZN(n10590) );
  NOR2_X1 U11460 ( .A1(n10829), .A2(n9975), .ZN(n10895) );
  NAND2_X1 U11461 ( .A1(n10134), .A2(n9829), .ZN(n12439) );
  OR2_X1 U11462 ( .A1(n11562), .A2(n11563), .ZN(n10088) );
  NAND2_X1 U11463 ( .A1(n12916), .A2(n11129), .ZN(n11249) );
  NAND2_X1 U11464 ( .A1(n18478), .A2(n18457), .ZN(n11573) );
  NAND3_X1 U11465 ( .A1(n13962), .A2(n11560), .A3(n11601), .ZN(n11567) );
  NAND2_X1 U11466 ( .A1(n10547), .A2(n10549), .ZN(n12910) );
  NAND2_X1 U11467 ( .A1(n10228), .A2(n12635), .ZN(n12764) );
  NAND2_X1 U11468 ( .A1(n10556), .A2(n13118), .ZN(n12909) );
  AND2_X1 U11469 ( .A1(n11049), .A2(n10601), .ZN(n10616) );
  AOI211_X2 U11470 ( .C1(n17413), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n11535), .B(n11534), .ZN(n13962) );
  INV_X1 U11471 ( .A(n10576), .ZN(n12076) );
  INV_X1 U11472 ( .A(n11559), .ZN(n18467) );
  INV_X1 U11473 ( .A(n18448), .ZN(n19084) );
  AND2_X1 U11474 ( .A1(n14597), .A2(n14614), .ZN(n14586) );
  AND2_X1 U11475 ( .A1(n10133), .A2(n20238), .ZN(n9829) );
  AND2_X1 U11476 ( .A1(n13106), .A2(n14614), .ZN(n12457) );
  AND2_X1 U11477 ( .A1(n17820), .A2(n10272), .ZN(n16584) );
  BUF_X2 U11478 ( .A(n13735), .Z(n14593) );
  OAI211_X1 U11479 ( .C1(n17415), .C2(n17361), .A(n11516), .B(n11515), .ZN(
        n18462) );
  NAND3_X1 U11480 ( .A1(n10343), .A2(n12096), .A3(n19451), .ZN(n10546) );
  AND2_X2 U11481 ( .A1(n10550), .A2(n9955), .ZN(n11049) );
  AOI211_X1 U11482 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n11546), .B(n11545), .ZN(n11559) );
  OR3_X2 U11483 ( .A1(n12659), .A2(n13364), .A3(n20237), .ZN(n13579) );
  INV_X1 U11484 ( .A(n20905), .ZN(n13786) );
  CLKBUF_X3 U11485 ( .A(n10558), .Z(n19439) );
  AND2_X1 U11486 ( .A1(n10558), .A2(n10557), .ZN(n11129) );
  NAND2_X1 U11487 ( .A1(n10496), .A2(n10461), .ZN(n10567) );
  INV_X1 U11489 ( .A(n11121), .ZN(n10557) );
  NAND2_X1 U11490 ( .A1(n10496), .A2(n11752), .ZN(n10539) );
  NAND2_X1 U11491 ( .A1(n12181), .A2(n11253), .ZN(n13477) );
  INV_X2 U11492 ( .A(U212), .ZN(n16692) );
  INV_X1 U11493 ( .A(n13002), .ZN(n12659) );
  INV_X1 U11494 ( .A(n10496), .ZN(n10990) );
  NAND3_X1 U11495 ( .A1(n10012), .A2(n9859), .A3(n9825), .ZN(n20260) );
  OR2_X2 U11496 ( .A1(n12249), .A2(n12248), .ZN(n13113) );
  NAND3_X1 U11497 ( .A1(n12232), .A2(n12231), .A3(n12230), .ZN(n13002) );
  NAND2_X2 U11498 ( .A1(n10523), .A2(n10522), .ZN(n11253) );
  OR2_X2 U11499 ( .A1(n16702), .A2(n16659), .ZN(n16704) );
  NAND2_X2 U11500 ( .A1(n9956), .A2(n9958), .ZN(n12096) );
  AND2_X2 U11501 ( .A1(n10494), .A2(n10493), .ZN(n11121) );
  AND4_X1 U11502 ( .A1(n12266), .A2(n12265), .A3(n12264), .A4(n12263), .ZN(
        n12274) );
  NAND2_X1 U11503 ( .A1(n9957), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9956) );
  NAND2_X1 U11504 ( .A1(n9959), .A2(n12883), .ZN(n9958) );
  AND4_X1 U11505 ( .A1(n12271), .A2(n12270), .A3(n12269), .A4(n12268), .ZN(
        n12272) );
  AND4_X1 U11506 ( .A1(n12225), .A2(n12224), .A3(n12223), .A4(n12222), .ZN(
        n12232) );
  NAND2_X1 U11507 ( .A1(n10504), .A2(n12883), .ZN(n10511) );
  NAND2_X1 U11508 ( .A1(n10509), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10510) );
  BUF_X2 U11509 ( .A(n11626), .Z(n17443) );
  AND4_X1 U11510 ( .A1(n12215), .A2(n12214), .A3(n12213), .A4(n12212), .ZN(
        n12221) );
  AND3_X1 U11511 ( .A1(n12257), .A2(n12254), .A3(n10007), .ZN(n9998) );
  AND4_X1 U11512 ( .A1(n12219), .A2(n12218), .A3(n12217), .A4(n12216), .ZN(
        n12220) );
  AND4_X1 U11513 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n10471) );
  NAND2_X2 U11514 ( .A1(n19026), .A2(n18959), .ZN(n19022) );
  INV_X2 U11515 ( .A(n18963), .ZN(n9805) );
  INV_X2 U11516 ( .A(n17416), .ZN(n14033) );
  INV_X2 U11517 ( .A(n14411), .ZN(n14235) );
  AND4_X1 U11518 ( .A1(n10465), .A2(n10464), .A3(n10463), .A4(n10462), .ZN(
        n10466) );
  INV_X4 U11519 ( .A(n17230), .ZN(n17413) );
  INV_X2 U11520 ( .A(n20843), .ZN(n9806) );
  OR2_X1 U11521 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11467), .ZN(
        n17230) );
  INV_X1 U11522 ( .A(n11684), .ZN(n11496) );
  NAND2_X2 U11523 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20015), .ZN(n20017) );
  AND2_X1 U11524 ( .A1(n12184), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10563) );
  NAND2_X1 U11525 ( .A1(n11459), .A2(n11458), .ZN(n17258) );
  INV_X2 U11526 ( .A(n9926), .ZN(n17397) );
  NAND2_X2 U11527 ( .A1(n20015), .A2(n19957), .ZN(n20021) );
  INV_X2 U11528 ( .A(n12733), .ZN(n9808) );
  INV_X2 U11529 ( .A(n14408), .ZN(n12252) );
  INV_X1 U11530 ( .A(n12733), .ZN(n14389) );
  CLKBUF_X1 U11531 ( .A(n10671), .Z(n12065) );
  NOR2_X1 U11532 ( .A1(n11466), .A2(n11465), .ZN(n11684) );
  AND3_X2 U11533 ( .A1(n13332), .A2(n10224), .A3(n15166), .ZN(n14418) );
  AND3_X2 U11534 ( .A1(n20885), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(n20237), 
        .ZN(n16105) );
  NAND2_X1 U11535 ( .A1(n10145), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11467) );
  OR2_X1 U11536 ( .A1(n17126), .A2(n11460), .ZN(n10416) );
  OR2_X2 U11537 ( .A1(n11465), .A2(n18886), .ZN(n9926) );
  NOR2_X1 U11538 ( .A1(n19042), .A2(n18104), .ZN(n19081) );
  AND2_X2 U11539 ( .A1(n12204), .A2(n13192), .ZN(n14420) );
  CLKBUF_X1 U11540 ( .A(n10670), .Z(n12064) );
  INV_X2 U11541 ( .A(n16743), .ZN(n16745) );
  NOR2_X2 U11542 ( .A1(n19050), .A2(n19057), .ZN(n18887) );
  NAND2_X1 U11543 ( .A1(n19064), .A2(n19057), .ZN(n17126) );
  AND2_X2 U11544 ( .A1(n12201), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13176) );
  NAND4_X2 U11545 ( .A1(n19050), .A2(n19057), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17426) );
  NAND2_X1 U11546 ( .A1(n19050), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11465) );
  AND2_X1 U11547 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12454), .ZN(
        n12204) );
  NAND2_X1 U11548 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n17094), .ZN(
        n11460) );
  AND2_X1 U11549 ( .A1(n12644), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12199) );
  NAND2_X1 U11550 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18886) );
  INV_X1 U11551 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19064) );
  INV_X1 U11552 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12873) );
  AND2_X1 U11553 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12872) );
  NOR2_X1 U11554 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10436) );
  INV_X2 U11555 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n12749) );
  INV_X2 U11556 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15166) );
  INV_X2 U11557 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13332) );
  INV_X1 U11558 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13175) );
  NAND2_X2 U11559 ( .A1(n18317), .A2(n18898), .ZN(n18334) );
  NAND2_X2 U11560 ( .A1(n17829), .A2(n17814), .ZN(n17868) );
  INV_X2 U11561 ( .A(n10135), .ZN(n14591) );
  AOI221_X2 U11562 ( .B1(n21040), .B2(n9798), .C1(n21200), .C2(n9798), .A(
        n16035), .ZN(n16031) );
  NOR2_X2 U11563 ( .A1(n15332), .A2(n15334), .ZN(n11897) );
  NOR2_X4 U11564 ( .A1(n14671), .A2(n14673), .ZN(n14659) );
  XNOR2_X1 U11565 ( .A(n10269), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17096) );
  NOR4_X1 U11566 ( .A1(n17081), .A2(n11573), .A3(n11567), .A4(n18467), .ZN(
        n17685) );
  AND2_X1 U11567 ( .A1(n20254), .A2(n10136), .ZN(n9846) );
  XNOR2_X1 U11568 ( .A(n12748), .B(n12747), .ZN(n13211) );
  NOR2_X2 U11569 ( .A1(n12148), .A2(n18891), .ZN(n18900) );
  NOR2_X1 U11570 ( .A1(n19084), .A2(n17747), .ZN(n9812) );
  OR2_X1 U11571 ( .A1(n13904), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13902) );
  NAND2_X1 U11572 ( .A1(n11249), .A2(n10574), .ZN(n10614) );
  AND3_X1 U11573 ( .A1(n12909), .A2(n12943), .A3(n10573), .ZN(n10574) );
  INV_X1 U11574 ( .A(n10983), .ZN(n10351) );
  AND2_X2 U11575 ( .A1(n12631), .A2(n11251), .ZN(n11410) );
  NAND2_X1 U11576 ( .A1(n15392), .A2(n9928), .ZN(n11443) );
  OAI21_X1 U11577 ( .B1(n10055), .B2(n10052), .A(n10049), .ZN(n16398) );
  NAND2_X1 U11578 ( .A1(n10053), .A2(n15510), .ZN(n10052) );
  AND2_X1 U11579 ( .A1(n10050), .A2(n10056), .ZN(n10049) );
  INV_X1 U11580 ( .A(n10057), .ZN(n10056) );
  AND2_X1 U11581 ( .A1(n15489), .A2(n12105), .ZN(n12102) );
  NOR3_X1 U11582 ( .A1(n9815), .A2(n10298), .A3(n10297), .ZN(n12112) );
  NAND2_X1 U11583 ( .A1(n11734), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10199) );
  INV_X1 U11584 ( .A(n17613), .ZN(n11739) );
  NAND2_X1 U11585 ( .A1(n11698), .A2(n11705), .ZN(n16645) );
  NOR2_X1 U11586 ( .A1(n9901), .A2(n13432), .ZN(n10366) );
  OR2_X1 U11587 ( .A1(n17632), .A2(n11702), .ZN(n11712) );
  NAND2_X1 U11588 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  INV_X1 U11589 ( .A(n10381), .ZN(n10034) );
  INV_X1 U11590 ( .A(n14765), .ZN(n10035) );
  NAND2_X1 U11591 ( .A1(n13588), .A2(n10038), .ZN(n14072) );
  AND2_X1 U11592 ( .A1(n13589), .A2(n10039), .ZN(n10038) );
  AND2_X1 U11593 ( .A1(n10378), .A2(n10040), .ZN(n10039) );
  AND2_X1 U11594 ( .A1(n9900), .A2(n13917), .ZN(n10378) );
  AOI21_X1 U11595 ( .B1(n13906), .B2(n9862), .A(n10362), .ZN(n14055) );
  OR2_X1 U11596 ( .A1(n12439), .A2(n12508), .ZN(n13005) );
  OAI21_X1 U11597 ( .B1(n12646), .B2(n12672), .A(n10028), .ZN(n12722) );
  AND2_X1 U11598 ( .A1(n10029), .A2(n12719), .ZN(n10028) );
  NOR2_X1 U11599 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n12454), .ZN(
        n12200) );
  INV_X1 U11600 ( .A(n10226), .ZN(n10224) );
  NAND2_X1 U11601 ( .A1(n15166), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10225) );
  NOR2_X1 U11602 ( .A1(n10890), .A2(n10185), .ZN(n10184) );
  INV_X1 U11603 ( .A(n10826), .ZN(n10185) );
  NAND2_X1 U11604 ( .A1(n10183), .A2(n9899), .ZN(n10891) );
  INV_X1 U11605 ( .A(n10829), .ZN(n10183) );
  OR2_X1 U11606 ( .A1(n11952), .A2(n11953), .ZN(n11954) );
  NAND2_X1 U11607 ( .A1(n10403), .A2(n9918), .ZN(n13890) );
  XNOR2_X1 U11608 ( .A(n11153), .B(n11151), .ZN(n11155) );
  NAND2_X1 U11609 ( .A1(n10300), .A2(n10299), .ZN(n10298) );
  INV_X1 U11610 ( .A(n15312), .ZN(n10299) );
  NOR2_X1 U11611 ( .A1(n16358), .A2(n10807), .ZN(n10989) );
  NAND2_X1 U11612 ( .A1(n13830), .A2(n10119), .ZN(n9968) );
  INV_X1 U11613 ( .A(n13137), .ZN(n10281) );
  OR2_X1 U11614 ( .A1(n11103), .A2(n10807), .ZN(n11105) );
  NAND2_X1 U11615 ( .A1(n15827), .A2(n15826), .ZN(n10312) );
  XNOR2_X1 U11616 ( .A(n11105), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15599) );
  OR2_X1 U11617 ( .A1(n15827), .A2(n15826), .ZN(n10311) );
  OAI211_X1 U11618 ( .C1(n11206), .C2(n10619), .A(n10618), .B(n10617), .ZN(
        n10634) );
  OR2_X1 U11619 ( .A1(n10615), .A2(n12410), .ZN(n10618) );
  NOR2_X1 U11620 ( .A1(n13962), .A2(n11559), .ZN(n11563) );
  AOI21_X1 U11621 ( .B1(n11585), .B2(n11584), .A(n11583), .ZN(n11598) );
  INV_X1 U11622 ( .A(n17637), .ZN(n11702) );
  INV_X1 U11623 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17311) );
  AND2_X1 U11624 ( .A1(n13346), .A2(n13345), .ZN(n13347) );
  INV_X2 U11625 ( .A(n9846), .ZN(n14614) );
  NAND2_X1 U11626 ( .A1(n10069), .A2(n10065), .ZN(n12342) );
  INV_X1 U11627 ( .A(n10066), .ZN(n10065) );
  NAND2_X1 U11628 ( .A1(n11049), .A2(n12181), .ZN(n12172) );
  INV_X1 U11629 ( .A(n15469), .ZN(n13465) );
  NAND2_X1 U11630 ( .A1(n12113), .A2(n11246), .ZN(n14467) );
  INV_X1 U11631 ( .A(n10128), .ZN(n15489) );
  NAND2_X1 U11632 ( .A1(n16396), .A2(n10350), .ZN(n10349) );
  OR3_X1 U11633 ( .A1(n15335), .A2(n10302), .A3(n15321), .ZN(n10301) );
  OR2_X1 U11634 ( .A1(n10989), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15500) );
  NAND2_X1 U11635 ( .A1(n9964), .A2(n13150), .ZN(n10841) );
  NAND2_X1 U11636 ( .A1(n9963), .A2(n9962), .ZN(n9964) );
  AOI21_X1 U11637 ( .B1(n14462), .B2(n15249), .A(n11137), .ZN(n9962) );
  NAND2_X1 U11638 ( .A1(n13154), .A2(n15249), .ZN(n9963) );
  NAND2_X1 U11639 ( .A1(n9960), .A2(n9893), .ZN(n10130) );
  AND2_X1 U11640 ( .A1(n11075), .A2(n16570), .ZN(n11450) );
  AND3_X1 U11641 ( .A1(n11289), .A2(n11288), .A3(n11287), .ZN(n13159) );
  AND2_X1 U11642 ( .A1(n11751), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12349) );
  NAND3_X1 U11643 ( .A1(n11464), .A2(n17094), .A3(n19050), .ZN(n17321) );
  NAND2_X1 U11644 ( .A1(n11735), .A2(n18002), .ZN(n11736) );
  OR2_X1 U11645 ( .A1(n11734), .A2(n18114), .ZN(n11735) );
  NOR2_X1 U11646 ( .A1(n15024), .A2(n20162), .ZN(n10076) );
  AND2_X1 U11647 ( .A1(n14476), .A2(n11445), .ZN(n16307) );
  AND2_X2 U11648 ( .A1(n10434), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10435) );
  INV_X1 U11649 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10434) );
  OAI211_X1 U11650 ( .C1(n17447), .C2(n17355), .A(n10152), .B(n10151), .ZN(
        n10150) );
  NAND2_X1 U11651 ( .A1(n17417), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10152) );
  NAND2_X1 U11652 ( .A1(n11665), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10151) );
  INV_X1 U11653 ( .A(n13821), .ZN(n10379) );
  CLKBUF_X1 U11654 ( .A(n14366), .Z(n14198) );
  BUF_X1 U11655 ( .A(n14422), .Z(n14373) );
  NAND2_X1 U11657 ( .A1(n12450), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12466) );
  OR2_X1 U11658 ( .A1(n13249), .A2(n13248), .ZN(n13276) );
  INV_X1 U11659 ( .A(n13579), .ZN(n13530) );
  NOR2_X1 U11660 ( .A1(n12373), .A2(n13682), .ZN(n10601) );
  AND4_X1 U11661 ( .A1(n10793), .A2(n10792), .A3(n10791), .A4(n10790), .ZN(
        n10805) );
  AND2_X1 U11662 ( .A1(n10880), .A2(n10879), .ZN(n11094) );
  NAND2_X1 U11663 ( .A1(n10785), .A2(n10784), .ZN(n11102) );
  OAI22_X1 U11664 ( .A1(n10687), .A2(n19668), .B1(n13696), .B2(n10686), .ZN(
        n10688) );
  NAND2_X1 U11665 ( .A1(n10537), .A2(n10536), .ZN(n11048) );
  NAND2_X1 U11666 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10205) );
  NAND2_X1 U11667 ( .A1(n11629), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10208) );
  NOR2_X1 U11668 ( .A1(n17628), .A2(n11712), .ZN(n11661) );
  OAI21_X1 U11669 ( .B1(n18102), .B2(n11702), .A(n17632), .ZN(n11711) );
  NAND2_X1 U11670 ( .A1(n10246), .A2(n14685), .ZN(n10245) );
  INV_X1 U11671 ( .A(n14708), .ZN(n10246) );
  NAND2_X1 U11672 ( .A1(n10376), .A2(n14660), .ZN(n10375) );
  INV_X1 U11673 ( .A(n14648), .ZN(n10376) );
  NAND2_X1 U11674 ( .A1(n10368), .A2(n14683), .ZN(n10367) );
  INV_X1 U11675 ( .A(n10369), .ZN(n10368) );
  OR2_X1 U11676 ( .A1(n14696), .A2(n10370), .ZN(n10369) );
  AND2_X1 U11677 ( .A1(n13572), .A2(n10030), .ZN(n13610) );
  NAND2_X1 U11678 ( .A1(n10031), .A2(n9901), .ZN(n10030) );
  NAND2_X1 U11679 ( .A1(n13253), .A2(n9828), .ZN(n10031) );
  INV_X1 U11680 ( .A(n14697), .ZN(n10247) );
  NAND2_X1 U11681 ( .A1(n10144), .A2(n9827), .ZN(n10018) );
  OR2_X1 U11682 ( .A1(n14788), .A2(n10238), .ZN(n10237) );
  INV_X1 U11683 ( .A(n14785), .ZN(n10238) );
  AOI21_X1 U11684 ( .B1(n10022), .B2(n10026), .A(n10020), .ZN(n10019) );
  INV_X1 U11685 ( .A(n13780), .ZN(n10021) );
  INV_X1 U11686 ( .A(n14053), .ZN(n10020) );
  INV_X1 U11687 ( .A(n13738), .ZN(n10241) );
  INV_X1 U11688 ( .A(n13616), .ZN(n10360) );
  NAND2_X1 U11689 ( .A1(n10230), .A2(n13292), .ZN(n10233) );
  INV_X1 U11690 ( .A(n13410), .ZN(n10230) );
  INV_X1 U11691 ( .A(n13411), .ZN(n10231) );
  NAND2_X1 U11692 ( .A1(n13253), .A2(n20233), .ZN(n13433) );
  NAND2_X1 U11693 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10015) );
  INV_X1 U11694 ( .A(n12238), .ZN(n10013) );
  NAND2_X1 U11695 ( .A1(n14421), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10011) );
  NAND2_X1 U11696 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10010) );
  AOI22_X1 U11697 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10009) );
  NAND2_X1 U11698 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10007) );
  NAND2_X1 U11699 ( .A1(n14366), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n9999) );
  NAND2_X1 U11700 ( .A1(n14331), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10008) );
  NAND2_X1 U11701 ( .A1(n12660), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10006) );
  NAND2_X1 U11702 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10004) );
  AOI22_X1 U11703 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14418), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10005) );
  NAND2_X1 U11704 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10002) );
  NAND2_X1 U11705 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10003) );
  AND2_X1 U11706 ( .A1(n12283), .A2(n12282), .ZN(n12311) );
  NOR2_X1 U11707 ( .A1(n13579), .A2(n13258), .ZN(n12336) );
  INV_X1 U11708 ( .A(n12298), .ZN(n10133) );
  INV_X1 U11709 ( .A(n10539), .ZN(n10343) );
  NAND2_X1 U11710 ( .A1(n9974), .A2(n9973), .ZN(n10957) );
  INV_X1 U11711 ( .A(n10956), .ZN(n9974) );
  OR2_X1 U11712 ( .A1(n10946), .A2(n10923), .ZN(n10952) );
  NAND2_X1 U11713 ( .A1(n10918), .A2(n9978), .ZN(n10946) );
  NOR2_X1 U11714 ( .A1(n9980), .A2(n9979), .ZN(n9978) );
  INV_X1 U11715 ( .A(n9916), .ZN(n9980) );
  INV_X1 U11716 ( .A(n10917), .ZN(n9979) );
  AND2_X1 U11717 ( .A1(n10895), .A2(n10893), .ZN(n10900) );
  NAND2_X1 U11718 ( .A1(n9874), .A2(n9977), .ZN(n9976) );
  INV_X1 U11719 ( .A(n11947), .ZN(n12001) );
  NAND2_X1 U11720 ( .A1(n12716), .A2(n12349), .ZN(n11776) );
  OAI211_X1 U11721 ( .C1(n15327), .C2(n10394), .A(n9915), .B(n9987), .ZN(n9986) );
  OR2_X1 U11722 ( .A1(n15318), .A2(n15329), .ZN(n10394) );
  NOR2_X1 U11723 ( .A1(n10405), .A2(n13747), .ZN(n10404) );
  INV_X1 U11724 ( .A(n13765), .ZN(n10405) );
  NAND2_X1 U11725 ( .A1(n11168), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10596) );
  AND2_X1 U11726 ( .A1(n10124), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10122) );
  NAND2_X1 U11727 ( .A1(n10350), .A2(n10125), .ZN(n10124) );
  INV_X1 U11728 ( .A(n16397), .ZN(n10125) );
  AND2_X1 U11729 ( .A1(n10347), .A2(n15487), .ZN(n10346) );
  NOR2_X1 U11730 ( .A1(n10264), .A2(n15195), .ZN(n10263) );
  INV_X1 U11731 ( .A(n15409), .ZN(n10264) );
  INV_X1 U11732 ( .A(n13767), .ZN(n10287) );
  INV_X1 U11733 ( .A(n13856), .ZN(n10252) );
  AND2_X1 U11734 ( .A1(n10911), .A2(n15776), .ZN(n9967) );
  INV_X1 U11735 ( .A(n15778), .ZN(n10055) );
  NOR2_X1 U11736 ( .A1(n10044), .A2(n9904), .ZN(n10119) );
  INV_X1 U11737 ( .A(n13388), .ZN(n10280) );
  AOI21_X1 U11738 ( .B1(n10311), .B2(n10309), .A(n10308), .ZN(n10307) );
  INV_X1 U11739 ( .A(n10311), .ZN(n10310) );
  INV_X1 U11740 ( .A(n15599), .ZN(n10308) );
  NAND2_X1 U11741 ( .A1(n10883), .A2(n10345), .ZN(n10044) );
  INV_X1 U11742 ( .A(n15819), .ZN(n10345) );
  INV_X1 U11743 ( .A(n11094), .ZN(n11101) );
  XNOR2_X1 U11744 ( .A(n11102), .B(n11094), .ZN(n11098) );
  NAND2_X1 U11745 ( .A1(n13638), .A2(n10846), .ZN(n13828) );
  OAI21_X1 U11746 ( .B1(n11076), .B2(n11302), .A(n13554), .ZN(n10845) );
  INV_X1 U11747 ( .A(n11168), .ZN(n11206) );
  INV_X1 U11748 ( .A(n11249), .ZN(n12868) );
  OR2_X1 U11749 ( .A1(n12001), .A2(n11762), .ZN(n11765) );
  AND2_X1 U11750 ( .A1(n10384), .A2(n19425), .ZN(n9953) );
  NAND2_X1 U11751 ( .A1(n10516), .A2(n12883), .ZN(n10523) );
  INV_X1 U11752 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13990) );
  INV_X1 U11753 ( .A(n17892), .ZN(n10270) );
  AND2_X1 U11754 ( .A1(n16644), .A2(n10219), .ZN(n10218) );
  NOR2_X1 U11755 ( .A1(n16652), .A2(n17969), .ZN(n10219) );
  AOI21_X1 U11756 ( .B1(n11739), .B2(n16645), .A(n18002), .ZN(n11700) );
  INV_X1 U11757 ( .A(n17618), .ZN(n11705) );
  NOR2_X1 U11758 ( .A1(n11564), .A2(n10086), .ZN(n10085) );
  NAND2_X1 U11759 ( .A1(n11561), .A2(n10087), .ZN(n10086) );
  XNOR2_X1 U11760 ( .A(n17637), .B(n17632), .ZN(n11663) );
  NAND2_X1 U11761 ( .A1(n11629), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10327) );
  INV_X1 U11762 ( .A(n10324), .ZN(n10323) );
  INV_X1 U11763 ( .A(n11672), .ZN(n10328) );
  OR2_X1 U11764 ( .A1(n18891), .A2(n12149), .ZN(n10084) );
  INV_X1 U11765 ( .A(n18871), .ZN(n16750) );
  AND2_X1 U11766 ( .A1(n13364), .A2(n12508), .ZN(n13355) );
  INV_X1 U11767 ( .A(n13593), .ZN(n14540) );
  OR2_X1 U11768 ( .A1(n12997), .A2(n20811), .ZN(n13107) );
  NOR2_X1 U11769 ( .A1(n13585), .A2(n13584), .ZN(n13586) );
  NAND2_X1 U11770 ( .A1(n14753), .A2(n14740), .ZN(n10032) );
  INV_X1 U11771 ( .A(n10144), .ZN(n14995) );
  NAND2_X1 U11772 ( .A1(n13903), .A2(n13902), .ZN(n13906) );
  NOR2_X1 U11773 ( .A1(n13533), .A2(n13535), .ZN(n13581) );
  NAND2_X1 U11774 ( .A1(n13326), .A2(n13325), .ZN(n13337) );
  AOI21_X1 U11775 ( .B1(n13069), .B2(n14128), .A(n10420), .ZN(n13074) );
  NOR2_X1 U11776 ( .A1(n10354), .A2(n15030), .ZN(n10138) );
  OAI21_X1 U11777 ( .B1(n14995), .B2(n10357), .A(n16090), .ZN(n10356) );
  INV_X1 U11778 ( .A(n10358), .ZN(n10357) );
  NAND2_X1 U11779 ( .A1(n13780), .A2(n16100), .ZN(n13903) );
  NAND2_X1 U11780 ( .A1(n9996), .A2(n13609), .ZN(n16108) );
  CLKBUF_X1 U11781 ( .A(n13005), .Z(n13108) );
  INV_X1 U11782 ( .A(n13735), .ZN(n14597) );
  NAND2_X1 U11783 ( .A1(n12763), .A2(n12762), .ZN(n10229) );
  NAND4_X1 U11784 ( .A1(n13355), .A2(n13168), .A3(n12846), .A4(n12641), .ZN(
        n13019) );
  XNOR2_X1 U11785 ( .A(n12975), .B(n12739), .ZN(n12973) );
  NOR2_X1 U11786 ( .A1(n15952), .A2(n20237), .ZN(n13111) );
  AND4_X1 U11787 ( .A1(n12229), .A2(n12228), .A3(n12227), .A4(n12226), .ZN(
        n12231) );
  NOR2_X1 U11788 ( .A1(n20630), .A2(n20396), .ZN(n20559) );
  NOR2_X1 U11789 ( .A1(n20552), .A2(n20396), .ZN(n20708) );
  INV_X1 U11790 ( .A(n20548), .ZN(n20697) );
  AOI21_X1 U11791 ( .B1(n20670), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20396), 
        .ZN(n20752) );
  NAND2_X1 U11792 ( .A1(n20237), .A2(n20236), .ZN(n20396) );
  CLKBUF_X1 U11793 ( .A(n12439), .Z(n12299) );
  NAND2_X1 U11794 ( .A1(n16272), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15952) );
  OR3_X1 U11795 ( .A1(n11114), .A2(n11119), .A3(n11113), .ZN(n12900) );
  OAI22_X1 U11796 ( .A1(n10825), .A2(n10824), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12883), .ZN(n11026) );
  XNOR2_X1 U11797 ( .A(n14458), .B(n14454), .ZN(n16294) );
  NAND2_X1 U11798 ( .A1(n10194), .A2(n10193), .ZN(n10192) );
  NOR2_X1 U11799 ( .A1(n10195), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10193) );
  NAND2_X1 U11800 ( .A1(n10895), .A2(n11251), .ZN(n10995) );
  NOR3_X1 U11801 ( .A1(n10985), .A2(n10984), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n10994) );
  NAND2_X1 U11802 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13317) );
  NAND2_X1 U11803 ( .A1(n10411), .A2(n13136), .ZN(n10410) );
  NOR2_X1 U11804 ( .A1(n15285), .A2(n10393), .ZN(n10392) );
  INV_X1 U11805 ( .A(n15290), .ZN(n10393) );
  NAND2_X1 U11806 ( .A1(n12052), .A2(n10391), .ZN(n10390) );
  AND2_X1 U11807 ( .A1(n15392), .A2(n10267), .ZN(n15376) );
  XNOR2_X1 U11808 ( .A(n11978), .B(n11979), .ZN(n15300) );
  NOR2_X1 U11809 ( .A1(n16473), .A2(n15178), .ZN(n15181) );
  CLKBUF_X1 U11810 ( .A(n11150), .Z(n11156) );
  INV_X1 U11811 ( .A(n15607), .ZN(n10258) );
  NOR2_X1 U11812 ( .A1(n9815), .A2(n10298), .ZN(n15306) );
  NOR2_X1 U11813 ( .A1(n16390), .A2(n10348), .ZN(n10347) );
  INV_X1 U11814 ( .A(n15500), .ZN(n10348) );
  NOR2_X1 U11815 ( .A1(n13659), .A2(n13660), .ZN(n13658) );
  AND3_X1 U11816 ( .A1(n11385), .A2(n11384), .A3(n11383), .ZN(n13227) );
  NAND2_X1 U11817 ( .A1(n10055), .A2(n15775), .ZN(n10054) );
  NOR2_X1 U11818 ( .A1(n13138), .A2(n9818), .ZN(n13395) );
  NAND2_X1 U11819 ( .A1(n13828), .A2(n13827), .ZN(n13830) );
  AND2_X1 U11820 ( .A1(n10295), .A2(n10293), .ZN(n12699) );
  NOR2_X1 U11821 ( .A1(n11154), .A2(n10294), .ZN(n10293) );
  INV_X1 U11822 ( .A(n13511), .ZN(n10129) );
  NAND2_X1 U11823 ( .A1(n9961), .A2(n10807), .ZN(n9960) );
  INV_X1 U11824 ( .A(n13154), .ZN(n9961) );
  NOR2_X1 U11825 ( .A1(n11253), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12631) );
  AND2_X1 U11826 ( .A1(n9923), .A2(n12398), .ZN(n19269) );
  AOI21_X1 U11827 ( .B1(n19425), .B2(n12349), .A(n11764), .ZN(n12681) );
  NAND2_X1 U11828 ( .A1(n20039), .A2(n20069), .ZN(n19557) );
  NAND2_X1 U11829 ( .A1(n20039), .A2(n19364), .ZN(n19597) );
  OAI21_X1 U11830 ( .B1(n20031), .B2(n16562), .A(n12345), .ZN(n19737) );
  OR2_X1 U11831 ( .A1(n20051), .A2(n20038), .ZN(n20034) );
  NAND2_X1 U11832 ( .A1(n20051), .A2(n20038), .ZN(n19596) );
  AND2_X1 U11833 ( .A1(n19326), .A2(n19364), .ZN(n19760) );
  NAND2_X1 U11834 ( .A1(n19326), .A2(n20069), .ZN(n19733) );
  AND2_X1 U11835 ( .A1(n20051), .A2(n20060), .ZN(n19892) );
  AND2_X1 U11836 ( .A1(n19326), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19891) );
  NAND2_X1 U11837 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19737), .ZN(n19459) );
  INV_X1 U11838 ( .A(n19737), .ZN(n19888) );
  AND2_X1 U11839 ( .A1(n11037), .A2(n20076), .ZN(n12896) );
  AOI21_X1 U11840 ( .B1(n17433), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n11488), .ZN(n11489) );
  NOR2_X1 U11841 ( .A1(n17258), .A2(n17459), .ZN(n11488) );
  NOR2_X1 U11842 ( .A1(n11628), .A2(n10207), .ZN(n11630) );
  NAND2_X1 U11843 ( .A1(n10081), .A2(n19079), .ZN(n17494) );
  OR2_X1 U11844 ( .A1(n15989), .A2(n15988), .ZN(n10081) );
  AND2_X1 U11845 ( .A1(n9813), .A2(n9909), .ZN(n10272) );
  AND2_X1 U11846 ( .A1(n17775), .A2(n9906), .ZN(n10198) );
  NAND2_X1 U11847 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17821) );
  NAND2_X1 U11848 ( .A1(n18278), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17928) );
  NOR2_X1 U11849 ( .A1(n16619), .A2(n15970), .ZN(n16575) );
  NAND2_X1 U11850 ( .A1(n9830), .A2(n11738), .ZN(n10222) );
  AND2_X1 U11851 ( .A1(n17868), .A2(n18144), .ZN(n10201) );
  NOR4_X1 U11852 ( .A1(n18181), .A2(n10095), .A3(n11727), .A4(n11730), .ZN(
        n18146) );
  INV_X1 U11853 ( .A(n17927), .ZN(n10095) );
  NAND2_X1 U11854 ( .A1(n10319), .A2(n10320), .ZN(n10318) );
  OR2_X1 U11855 ( .A1(n11732), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10320) );
  NAND2_X1 U11856 ( .A1(n17924), .A2(n9863), .ZN(n10319) );
  NAND2_X1 U11857 ( .A1(n18069), .A2(n11678), .ZN(n18057) );
  AOI211_X1 U11858 ( .C1(n11591), .C2(n11590), .A(n11598), .B(n11595), .ZN(
        n18868) );
  XNOR2_X1 U11859 ( .A(n11663), .B(n10196), .ZN(n18081) );
  INV_X1 U11860 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10196) );
  NAND2_X1 U11861 ( .A1(n18094), .A2(n11673), .ZN(n18080) );
  NAND2_X1 U11862 ( .A1(n18101), .A2(n18095), .ZN(n18094) );
  XNOR2_X1 U11863 ( .A(n17637), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18095) );
  NAND2_X1 U11864 ( .A1(n10073), .A2(n10072), .ZN(n12583) );
  NOR2_X1 U11865 ( .A1(n12299), .A2(n20089), .ZN(n10072) );
  INV_X1 U11866 ( .A(n14608), .ZN(n10235) );
  NOR3_X1 U11867 ( .A1(n14658), .A2(n21102), .A3(n14905), .ZN(n14633) );
  OR2_X1 U11868 ( .A1(n14694), .A2(n14607), .ZN(n14658) );
  OR2_X1 U11869 ( .A1(n14593), .A2(n13361), .ZN(n20162) );
  INV_X1 U11870 ( .A(n14888), .ZN(n10132) );
  NAND2_X1 U11871 ( .A1(n20095), .A2(n12705), .ZN(n16116) );
  OR3_X2 U11872 ( .A1(n15942), .A2(n12997), .A3(n20089), .ZN(n20095) );
  INV_X1 U11873 ( .A(n12853), .ZN(n16255) );
  INV_X1 U11874 ( .A(n16263), .ZN(n16242) );
  INV_X1 U11875 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20631) );
  CLKBUF_X1 U11876 ( .A(n13188), .Z(n13189) );
  INV_X1 U11877 ( .A(n20602), .ZN(n20886) );
  INV_X1 U11878 ( .A(n20499), .ZN(n20520) );
  NAND2_X1 U11879 ( .A1(n13486), .A2(n13485), .ZN(n19293) );
  INV_X1 U11880 ( .A(n19301), .ZN(n19245) );
  NAND2_X1 U11881 ( .A1(n15284), .A2(n15285), .ZN(n15361) );
  NAND2_X1 U11882 ( .A1(n10407), .A2(n13394), .ZN(n10406) );
  INV_X1 U11883 ( .A(n10408), .ZN(n10407) );
  CLKBUF_X1 U11884 ( .A(n15323), .Z(n15352) );
  NOR2_X2 U11885 ( .A1(n15352), .A2(n19460), .ZN(n15346) );
  OAI21_X1 U11886 ( .B1(n12858), .B2(n12867), .A(n16570), .ZN(n15323) );
  XNOR2_X1 U11887 ( .A(n14481), .B(n14480), .ZN(n19303) );
  OAI211_X1 U11888 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n13465), .A(
        n10164), .B(n10162), .ZN(n15439) );
  NAND2_X1 U11889 ( .A1(n10163), .A2(n10168), .ZN(n10162) );
  NAND2_X1 U11890 ( .A1(n13465), .A2(n9930), .ZN(n10164) );
  XNOR2_X1 U11891 ( .A(n14467), .B(n14466), .ZN(n16295) );
  NAND2_X1 U11892 ( .A1(n16392), .A2(n16493), .ZN(n10047) );
  NAND2_X1 U11893 ( .A1(n16520), .A2(n16491), .ZN(n10046) );
  INV_X1 U11894 ( .A(n16488), .ZN(n16475) );
  NAND2_X1 U11895 ( .A1(n12357), .A2(n12348), .ZN(n16498) );
  OR2_X1 U11896 ( .A1(n12357), .A2(n11259), .ZN(n16478) );
  INV_X1 U11897 ( .A(n16486), .ZN(n16491) );
  NAND3_X1 U11898 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20037), .A3(n19737), 
        .ZN(n16486) );
  NOR2_X1 U11899 ( .A1(n14467), .A2(n14466), .ZN(n14474) );
  AOI21_X1 U11900 ( .B1(n16307), .B2(n19420), .A(n11453), .ZN(n11454) );
  XNOR2_X1 U11901 ( .A(n11010), .B(n10421), .ZN(n15466) );
  NAND2_X1 U11902 ( .A1(n10115), .A2(n9981), .ZN(n11010) );
  AOI21_X1 U11903 ( .B1(n12102), .B2(n12107), .A(n10336), .ZN(n10115) );
  OAI21_X1 U11904 ( .B1(n12112), .B2(n12115), .A(n12114), .ZN(n15468) );
  NOR2_X1 U11905 ( .A1(n12119), .A2(n10284), .ZN(n10283) );
  NAND2_X1 U11906 ( .A1(n16319), .A2(n19420), .ZN(n10285) );
  OR2_X1 U11907 ( .A1(n15475), .A2(n19419), .ZN(n12122) );
  XNOR2_X1 U11908 ( .A(n10048), .B(n16391), .ZN(n16521) );
  NAND2_X1 U11909 ( .A1(n10349), .A2(n15500), .ZN(n10048) );
  NAND2_X1 U11910 ( .A1(n11450), .A2(n20080), .ZN(n19436) );
  AND2_X1 U11911 ( .A1(n11450), .A2(n11449), .ZN(n19420) );
  INV_X1 U11912 ( .A(n19436), .ZN(n19414) );
  INV_X1 U11913 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20074) );
  INV_X1 U11914 ( .A(n20038), .ZN(n20060) );
  NAND2_X1 U11915 ( .A1(n19760), .A2(n19771), .ZN(n19832) );
  INV_X1 U11916 ( .A(n16778), .ZN(n10275) );
  NOR2_X1 U11917 ( .A1(n17127), .A2(n16779), .ZN(n10276) );
  NOR2_X1 U11918 ( .A1(n17511), .A2(n17710), .ZN(n17507) );
  NAND2_X1 U11919 ( .A1(n16607), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10269) );
  NAND2_X1 U11920 ( .A1(n16618), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10330) );
  INV_X1 U11921 ( .A(n17821), .ZN(n11741) );
  NOR2_X1 U11922 ( .A1(n18107), .A2(n11739), .ZN(n17997) );
  XNOR2_X1 U11923 ( .A(n15884), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16616) );
  NAND2_X1 U11924 ( .A1(n15971), .A2(n15970), .ZN(n15884) );
  OAI21_X1 U11925 ( .B1(n18128), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n18409), .ZN(n10103) );
  INV_X1 U11926 ( .A(n12647), .ZN(n14411) );
  NAND2_X1 U11927 ( .A1(n13176), .A2(n13174), .ZN(n14408) );
  AND2_X1 U11928 ( .A1(n10539), .A2(n19439), .ZN(n10542) );
  OR2_X1 U11929 ( .A1(n11584), .A2(n11585), .ZN(n11580) );
  OAI21_X1 U11930 ( .B1(n14053), .B2(n10363), .A(n10354), .ZN(n10362) );
  INV_X1 U11931 ( .A(n14054), .ZN(n10363) );
  NAND2_X1 U11932 ( .A1(n13902), .A2(n10025), .ZN(n10024) );
  INV_X1 U11933 ( .A(n16100), .ZN(n10025) );
  OR2_X1 U11934 ( .A1(n13273), .A2(n13272), .ZN(n13280) );
  INV_X1 U11935 ( .A(n12297), .ZN(n12847) );
  OR2_X1 U11936 ( .A1(n12439), .A2(n12438), .ZN(n12440) );
  NAND2_X1 U11937 ( .A1(n12673), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10029) );
  NOR2_X1 U11938 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13193) );
  NOR2_X1 U11939 ( .A1(n12388), .A2(n12298), .ZN(n12429) );
  NAND2_X1 U11940 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12269) );
  NAND2_X1 U11941 ( .A1(n14366), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12268) );
  AOI22_X1 U11942 ( .A1(n12647), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U11943 ( .A1(n14459), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n9977) );
  NOR2_X1 U11944 ( .A1(n15318), .A2(n10396), .ZN(n10395) );
  INV_X1 U11945 ( .A(n11924), .ZN(n10396) );
  INV_X1 U11946 ( .A(n10496), .ZN(n10548) );
  NAND2_X1 U11947 ( .A1(n10499), .A2(n10498), .ZN(n10588) );
  INV_X1 U11948 ( .A(n10312), .ZN(n10309) );
  OR2_X1 U11949 ( .A1(n11102), .A2(n11101), .ZN(n11103) );
  AND3_X1 U11950 ( .A1(n10684), .A2(n10739), .A3(n9910), .ZN(n10785) );
  AOI21_X1 U11951 ( .B1(n10766), .B2(n10043), .A(n9891), .ZN(n10784) );
  AND3_X1 U11952 ( .A1(n10767), .A2(n10768), .A3(n10769), .ZN(n10043) );
  NAND2_X1 U11953 ( .A1(n10629), .A2(n10628), .ZN(n11153) );
  OR2_X1 U11954 ( .A1(n10724), .A2(n10723), .ZN(n11077) );
  AND4_X1 U11955 ( .A1(n10487), .A2(n10486), .A3(n10485), .A4(n10484), .ZN(
        n10488) );
  NAND2_X1 U11956 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20074), .ZN(
        n11011) );
  NAND2_X1 U11957 ( .A1(n18478), .A2(n17081), .ZN(n11565) );
  NAND2_X1 U11958 ( .A1(n11661), .A2(n11660), .ZN(n11683) );
  NAND2_X1 U11959 ( .A1(n11565), .A2(n11566), .ZN(n10087) );
  AOI21_X1 U11960 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18905), .A(
        n11579), .ZN(n11585) );
  NOR2_X1 U11961 ( .A1(n11594), .A2(n11593), .ZN(n11579) );
  AOI22_X1 U11962 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18910), .B2(n19050), .ZN(
        n11584) );
  OAI211_X1 U11963 ( .C1(n17453), .C2(n17435), .A(n10326), .B(n10325), .ZN(
        n10324) );
  NAND2_X1 U11964 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10325) );
  NAND2_X1 U11965 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10326) );
  NAND2_X1 U11966 ( .A1(n11629), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10153) );
  INV_X1 U11967 ( .A(n10150), .ZN(n10149) );
  INV_X1 U11968 ( .A(n11532), .ZN(n10154) );
  NOR2_X1 U11969 ( .A1(n14604), .A2(n10064), .ZN(n10063) );
  INV_X1 U11970 ( .A(n15999), .ZN(n10064) );
  NOR2_X1 U11971 ( .A1(n9911), .A2(n13590), .ZN(n13585) );
  INV_X1 U11972 ( .A(n14624), .ZN(n10372) );
  NOR2_X1 U11973 ( .A1(n10377), .A2(n10375), .ZN(n10374) );
  INV_X1 U11974 ( .A(n14636), .ZN(n10377) );
  NAND2_X1 U11975 ( .A1(n14707), .A2(n10371), .ZN(n10370) );
  OR2_X1 U11976 ( .A1(n15164), .A2(n20237), .ZN(n14434) );
  NAND2_X1 U11977 ( .A1(n10383), .A2(n10382), .ZN(n10381) );
  INV_X1 U11978 ( .A(n14869), .ZN(n10382) );
  INV_X1 U11979 ( .A(n14784), .ZN(n10383) );
  INV_X1 U11980 ( .A(n13726), .ZN(n10380) );
  NOR2_X1 U11981 ( .A1(n12674), .A2(n20237), .ZN(n13782) );
  INV_X1 U11982 ( .A(n13572), .ZN(n13575) );
  NOR2_X1 U11983 ( .A1(n14994), .A2(n9936), .ZN(n10358) );
  INV_X1 U11984 ( .A(n13902), .ZN(n10026) );
  OR2_X1 U11985 ( .A1(n13529), .A2(n13528), .ZN(n13785) );
  OR2_X1 U11986 ( .A1(n12658), .A2(n12657), .ZN(n13784) );
  NAND2_X1 U11987 ( .A1(n12952), .A2(n12951), .ZN(n13234) );
  OR2_X1 U11988 ( .A1(n12671), .A2(n12670), .ZN(n12979) );
  AND3_X1 U11989 ( .A1(n10425), .A2(n12735), .A3(n12734), .ZN(n12978) );
  AND2_X1 U11990 ( .A1(n20595), .A2(n12474), .ZN(n20246) );
  NAND2_X1 U11991 ( .A1(n12742), .A2(n12741), .ZN(n20302) );
  NAND2_X1 U11992 ( .A1(n10141), .A2(n20237), .ZN(n13251) );
  OAI21_X1 U11993 ( .B1(n12340), .B2(n12339), .A(n10067), .ZN(n10066) );
  AND2_X1 U11994 ( .A1(n12341), .A2(n10068), .ZN(n10067) );
  NAND2_X1 U11995 ( .A1(n20237), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10068) );
  NAND2_X1 U11996 ( .A1(n10070), .A2(n9867), .ZN(n10069) );
  OR2_X1 U11997 ( .A1(n12334), .A2(n10071), .ZN(n10070) );
  AND2_X1 U11998 ( .A1(n12336), .A2(n12335), .ZN(n10071) );
  OR2_X1 U11999 ( .A1(n10736), .A2(n10735), .ZN(n11273) );
  NOR2_X1 U12000 ( .A1(n11007), .A2(n10191), .ZN(n10190) );
  NAND2_X1 U12001 ( .A1(n10976), .A2(n10995), .ZN(n10973) );
  AND2_X1 U12002 ( .A1(n10900), .A2(n10898), .ZN(n10902) );
  AND2_X1 U12003 ( .A1(n15382), .A2(n15374), .ZN(n10267) );
  AOI211_X1 U12004 ( .C1(n12005), .C2(n12002), .A(n12001), .B(n12026), .ZN(
        n12003) );
  AND2_X1 U12005 ( .A1(n12629), .A2(n11259), .ZN(n11947) );
  AND2_X1 U12006 ( .A1(n10548), .A2(n12096), .ZN(n11258) );
  AND2_X1 U12007 ( .A1(n10404), .A2(n10402), .ZN(n10401) );
  INV_X1 U12008 ( .A(n13848), .ZN(n10402) );
  INV_X1 U12009 ( .A(n13601), .ZN(n9994) );
  NAND3_X1 U12010 ( .A1(n10497), .A2(n19460), .A3(n10990), .ZN(n10576) );
  AND2_X1 U12011 ( .A1(n19451), .A2(n10495), .ZN(n10497) );
  AOI22_X1 U12012 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10476) );
  NOR2_X1 U12013 ( .A1(n15453), .A2(n10166), .ZN(n10165) );
  NOR2_X1 U12014 ( .A1(n11229), .A2(n10182), .ZN(n10181) );
  INV_X1 U12015 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10182) );
  OAI21_X1 U12016 ( .B1(n10972), .B2(n10058), .A(n15511), .ZN(n10057) );
  NAND2_X1 U12017 ( .A1(n10053), .A2(n10051), .ZN(n10050) );
  NOR2_X1 U12018 ( .A1(n10058), .A2(n15775), .ZN(n10051) );
  NOR2_X1 U12019 ( .A1(n16415), .A2(n10178), .ZN(n10177) );
  INV_X1 U12020 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10178) );
  NOR2_X1 U12021 ( .A1(n16465), .A2(n10174), .ZN(n10173) );
  NAND2_X1 U12022 ( .A1(n10303), .A2(n15325), .ZN(n10302) );
  INV_X1 U12023 ( .A(n15192), .ZN(n10303) );
  INV_X1 U12024 ( .A(n13748), .ZN(n10288) );
  INV_X1 U12025 ( .A(n13061), .ZN(n10251) );
  AND4_X1 U12026 ( .A1(n10802), .A2(n10801), .A3(n10800), .A4(n10799), .ZN(
        n10803) );
  AND4_X1 U12027 ( .A1(n10797), .A2(n10796), .A3(n10795), .A4(n10794), .ZN(
        n10804) );
  INV_X2 U12028 ( .A(n10615), .ZN(n12128) );
  INV_X1 U12029 ( .A(n13477), .ZN(n11014) );
  AND2_X1 U12030 ( .A1(n11266), .A2(n11265), .ZN(n11271) );
  INV_X1 U12031 ( .A(n13159), .ZN(n10260) );
  NAND2_X1 U12032 ( .A1(n9982), .A2(n11756), .ZN(n11758) );
  NAND2_X1 U12033 ( .A1(n10641), .A2(n12349), .ZN(n9982) );
  AND2_X1 U12034 ( .A1(n11947), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11757) );
  NAND2_X1 U12035 ( .A1(n12181), .A2(n16562), .ZN(n12373) );
  OR2_X1 U12036 ( .A1(n19425), .A2(n12928), .ZN(n10659) );
  INV_X1 U12037 ( .A(n10658), .ZN(n9952) );
  INV_X1 U12038 ( .A(n10649), .ZN(n9954) );
  INV_X1 U12039 ( .A(n10652), .ZN(n9951) );
  AOI22_X1 U12040 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10468) );
  NOR2_X1 U12041 ( .A1(n18886), .A2(n11460), .ZN(n11461) );
  INV_X1 U12042 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10105) );
  NOR2_X1 U12043 ( .A1(n17094), .A2(n19050), .ZN(n10078) );
  NOR3_X1 U12044 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n18886), .ZN(n11477) );
  NOR3_X1 U12045 ( .A1(n19050), .A2(n17094), .A3(n17126), .ZN(n11625) );
  NOR2_X1 U12046 ( .A1(n10204), .A2(n10203), .ZN(n10202) );
  NAND2_X1 U12047 ( .A1(n10206), .A2(n10208), .ZN(n10203) );
  NAND2_X1 U12048 ( .A1(n11626), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10206) );
  NOR2_X1 U12049 ( .A1(n18097), .A2(n16612), .ZN(n16587) );
  NAND2_X1 U12050 ( .A1(n17820), .A2(n9813), .ZN(n12155) );
  AND2_X1 U12051 ( .A1(n17950), .A2(n9881), .ZN(n17857) );
  NOR2_X1 U12052 ( .A1(n11727), .A2(n18181), .ZN(n10216) );
  INV_X1 U12053 ( .A(n11733), .ZN(n10214) );
  INV_X1 U12054 ( .A(n10216), .ZN(n10212) );
  OR2_X1 U12055 ( .A1(n17896), .A2(n18002), .ZN(n10209) );
  INV_X1 U12056 ( .A(n18457), .ZN(n11566) );
  NAND2_X1 U12057 ( .A1(n17897), .A2(n18218), .ZN(n17829) );
  NOR2_X1 U12058 ( .A1(n17621), .A2(n11683), .ZN(n11698) );
  NAND2_X1 U12059 ( .A1(n18056), .A2(n11679), .ZN(n11681) );
  AOI22_X1 U12060 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18905), .B2(n19057), .ZN(
        n11594) );
  NOR2_X1 U12061 ( .A1(n11570), .A2(n11568), .ZN(n12148) );
  AOI21_X1 U12062 ( .B1(n14033), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n10090), .ZN(n10089) );
  OAI211_X1 U12063 ( .C1(n17447), .C2(n17414), .A(n10092), .B(n10091), .ZN(
        n10090) );
  NAND2_X1 U12064 ( .A1(n11665), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10092) );
  NAND2_X1 U12065 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10091) );
  AOI22_X1 U12066 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11482) );
  AND2_X1 U12067 ( .A1(n10083), .A2(n10082), .ZN(n15989) );
  INV_X1 U12068 ( .A(n13959), .ZN(n10082) );
  NAND2_X1 U12069 ( .A1(n10084), .A2(n9868), .ZN(n10083) );
  NOR2_X1 U12070 ( .A1(n11576), .A2(n11599), .ZN(n13965) );
  NAND2_X1 U12071 ( .A1(n13953), .A2(n13952), .ZN(n17645) );
  AND2_X1 U12072 ( .A1(n10063), .A2(n10062), .ZN(n10061) );
  INV_X1 U12073 ( .A(n14605), .ZN(n10062) );
  NAND2_X1 U12074 ( .A1(n16027), .A2(n10063), .ZN(n14748) );
  NAND2_X1 U12075 ( .A1(n14089), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14074) );
  NOR2_X1 U12076 ( .A1(n13367), .A2(n13368), .ZN(n13593) );
  NAND2_X1 U12077 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13595), .ZN(n13377) );
  OR3_X1 U12078 ( .A1(n10245), .A2(n10247), .A3(n14674), .ZN(n10244) );
  NAND2_X1 U12079 ( .A1(n16003), .A2(n9931), .ZN(n10236) );
  OR2_X1 U12080 ( .A1(n14799), .A2(n14800), .ZN(n14797) );
  NOR2_X1 U12081 ( .A1(n14344), .A2(n13351), .ZN(n14382) );
  OAI21_X1 U12082 ( .B1(n14363), .B2(n14915), .A(n14362), .ZN(n14648) );
  AND2_X1 U12083 ( .A1(n14659), .A2(n10373), .ZN(n14647) );
  INV_X1 U12084 ( .A(n10375), .ZN(n10373) );
  NAND2_X1 U12085 ( .A1(n14304), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14323) );
  AND2_X1 U12086 ( .A1(n13350), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14304) );
  INV_X1 U12087 ( .A(n14287), .ZN(n13350) );
  NAND2_X1 U12088 ( .A1(n14253), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14287) );
  AND2_X1 U12089 ( .A1(n13349), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14253) );
  INV_X1 U12090 ( .A(n14233), .ZN(n13349) );
  NOR2_X1 U12091 ( .A1(n14196), .A2(n14743), .ZN(n14213) );
  NAND2_X1 U12092 ( .A1(n14213), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14233) );
  CLKBUF_X1 U12093 ( .A(n14717), .Z(n14718) );
  AND2_X1 U12094 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n14164), .ZN(
        n14180) );
  INV_X1 U12095 ( .A(n14150), .ZN(n14164) );
  NOR2_X1 U12096 ( .A1(n14119), .A2(n16008), .ZN(n14151) );
  NAND2_X1 U12097 ( .A1(n14151), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14150) );
  CLKBUF_X1 U12098 ( .A(n14791), .Z(n14792) );
  NAND2_X1 U12099 ( .A1(n14105), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14119) );
  NOR2_X1 U12100 ( .A1(n14074), .A2(n16024), .ZN(n14105) );
  NAND2_X1 U12101 ( .A1(n13922), .A2(n13921), .ZN(n13935) );
  NOR2_X1 U12102 ( .A1(n13805), .A2(n20112), .ZN(n13875) );
  NAND2_X1 U12103 ( .A1(n13720), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13805) );
  AOI21_X1 U12104 ( .B1(n13618), .B2(n14128), .A(n13539), .ZN(n13542) );
  CLKBUF_X1 U12105 ( .A(n13588), .Z(n13541) );
  NAND2_X1 U12106 ( .A1(n13446), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13533) );
  INV_X1 U12107 ( .A(n13452), .ZN(n13453) );
  AND2_X1 U12108 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n13404), .ZN(
        n13446) );
  NAND2_X1 U12109 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13327) );
  NOR2_X1 U12110 ( .A1(n13327), .A2(n13419), .ZN(n13404) );
  NAND2_X1 U12111 ( .A1(n13071), .A2(n13070), .ZN(n13326) );
  INV_X1 U12112 ( .A(n13073), .ZN(n13071) );
  NOR2_X1 U12113 ( .A1(n14639), .A2(n14628), .ZN(n14627) );
  NOR3_X1 U12114 ( .A1(n14722), .A2(n10247), .A3(n14708), .ZN(n14699) );
  NOR2_X1 U12115 ( .A1(n14722), .A2(n14708), .ZN(n14710) );
  NOR2_X1 U12116 ( .A1(n14995), .A2(n14994), .ZN(n14993) );
  OR2_X1 U12117 ( .A1(n9817), .A2(n14754), .ZN(n14756) );
  NOR2_X1 U12118 ( .A1(n14756), .A2(n14742), .ZN(n14741) );
  OR2_X1 U12119 ( .A1(n16206), .A2(n15027), .ZN(n15105) );
  AND2_X1 U12120 ( .A1(n16090), .A2(n14060), .ZN(n16048) );
  NOR2_X1 U12121 ( .A1(n14797), .A2(n14788), .ZN(n16004) );
  NOR3_X1 U12122 ( .A1(n14797), .A2(n10240), .A3(n14788), .ZN(n16006) );
  OR2_X1 U12123 ( .A1(n16090), .A2(n16210), .ZN(n16075) );
  OR2_X1 U12124 ( .A1(n16090), .A2(n14062), .ZN(n16078) );
  INV_X1 U12125 ( .A(n13888), .ZN(n10242) );
  NOR2_X1 U12126 ( .A1(n13939), .A2(n13940), .ZN(n14512) );
  OAI21_X1 U12127 ( .B1(n13780), .B2(n10026), .A(n10022), .ZN(n16088) );
  NAND2_X1 U12128 ( .A1(n13734), .A2(n9822), .ZN(n16240) );
  AND2_X1 U12129 ( .A1(n13734), .A2(n9855), .ZN(n16238) );
  AOI21_X1 U12130 ( .B1(n13770), .B2(n10360), .A(n9871), .ZN(n10359) );
  NAND2_X1 U12131 ( .A1(n13734), .A2(n10424), .ZN(n16254) );
  AND2_X1 U12132 ( .A1(n13733), .A2(n13732), .ZN(n16249) );
  NOR2_X1 U12133 ( .A1(n10233), .A2(n13463), .ZN(n10232) );
  NAND2_X1 U12134 ( .A1(n10231), .A2(n10234), .ZN(n13462) );
  INV_X1 U12135 ( .A(n10233), .ZN(n10234) );
  NAND2_X1 U12136 ( .A1(n13021), .A2(n13172), .ZN(n16130) );
  NAND2_X1 U12137 ( .A1(n13262), .A2(n13261), .ZN(n13607) );
  NOR2_X1 U12138 ( .A1(n13411), .A2(n13410), .ZN(n13413) );
  NAND2_X1 U12139 ( .A1(n12764), .A2(n14597), .ZN(n10227) );
  OR2_X1 U12140 ( .A1(n13028), .A2(n13027), .ZN(n13411) );
  OR2_X1 U12141 ( .A1(n16201), .A2(n13047), .ZN(n16206) );
  XNOR2_X1 U12142 ( .A(n13234), .B(n13023), .ZN(n13233) );
  XNOR2_X1 U12143 ( .A(n12950), .B(n12948), .ZN(n12947) );
  AND2_X1 U12144 ( .A1(n14591), .A2(n14614), .ZN(n14567) );
  NAND2_X1 U12145 ( .A1(n12977), .A2(n12976), .ZN(n13237) );
  CLKBUF_X1 U12146 ( .A(n13174), .Z(n15172) );
  NOR2_X1 U12147 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20625) );
  NOR2_X1 U12148 ( .A1(n10014), .A2(n10013), .ZN(n10012) );
  NAND2_X1 U12149 ( .A1(n12255), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10001) );
  INV_X1 U12150 ( .A(n20295), .ZN(n20286) );
  OR2_X1 U12151 ( .A1(n20883), .A2(n13069), .ZN(n20602) );
  NAND2_X1 U12152 ( .A1(n9811), .A2(n20234), .ZN(n20601) );
  NAND2_X1 U12153 ( .A1(n16105), .A2(n20229), .ZN(n20291) );
  INV_X1 U12154 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16272) );
  AND2_X1 U12155 ( .A1(n11023), .A2(n11022), .ZN(n11066) );
  AND2_X1 U12156 ( .A1(n10558), .A2(n11121), .ZN(n10549) );
  NAND2_X1 U12157 ( .A1(n13465), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15459) );
  NAND2_X1 U12158 ( .A1(n14457), .A2(n10998), .ZN(n11008) );
  NAND2_X1 U12159 ( .A1(n16357), .A2(n10993), .ZN(n10195) );
  NAND2_X1 U12160 ( .A1(n9970), .A2(n9969), .ZN(n16358) );
  INV_X1 U12161 ( .A(n10988), .ZN(n9970) );
  INV_X1 U12162 ( .A(n10994), .ZN(n9969) );
  NAND2_X1 U12163 ( .A1(n9972), .A2(n9971), .ZN(n10976) );
  INV_X1 U12164 ( .A(n10957), .ZN(n9972) );
  NAND2_X1 U12165 ( .A1(n10940), .A2(n10931), .ZN(n10956) );
  NOR2_X1 U12166 ( .A1(n15188), .A2(n15563), .ZN(n15191) );
  NAND2_X1 U12167 ( .A1(n15186), .A2(n9835), .ZN(n15187) );
  AND2_X1 U12168 ( .A1(n10947), .A2(n10951), .ZN(n19187) );
  NAND2_X1 U12169 ( .A1(n10918), .A2(n10917), .ZN(n10954) );
  AND2_X1 U12170 ( .A1(n10902), .A2(n13142), .ZN(n10903) );
  NAND2_X1 U12171 ( .A1(n10919), .A2(n10995), .ZN(n10918) );
  NOR2_X1 U12172 ( .A1(n10829), .A2(n10186), .ZN(n10827) );
  NAND2_X1 U12173 ( .A1(n9799), .A2(n10187), .ZN(n10186) );
  NOR2_X1 U12174 ( .A1(n13317), .A2(n15250), .ZN(n13467) );
  AND2_X1 U12175 ( .A1(n16562), .A2(n14471), .ZN(n10167) );
  NAND2_X1 U12176 ( .A1(n10409), .A2(n9903), .ZN(n10408) );
  INV_X1 U12177 ( .A(n10410), .ZN(n10409) );
  NOR2_X1 U12178 ( .A1(n12693), .A2(n11781), .ZN(n11782) );
  NAND2_X1 U12179 ( .A1(n12712), .A2(n9983), .ZN(n10399) );
  AND2_X1 U12180 ( .A1(n12076), .A2(n10577), .ZN(n12867) );
  INV_X1 U12181 ( .A(n12073), .ZN(n10391) );
  NOR2_X1 U12182 ( .A1(n10389), .A2(n10391), .ZN(n10388) );
  INV_X1 U12183 ( .A(n10392), .ZN(n10389) );
  AND2_X1 U12184 ( .A1(n12024), .A2(n12023), .ZN(n15290) );
  AND2_X1 U12185 ( .A1(n15392), .A2(n15382), .ZN(n15384) );
  NAND2_X1 U12186 ( .A1(n11897), .A2(n11924), .ZN(n10397) );
  CLKBUF_X1 U12187 ( .A(n15332), .Z(n15333) );
  CLKBUF_X1 U12188 ( .A(n13890), .Z(n13891) );
  OR2_X1 U12189 ( .A1(n11805), .A2(n11804), .ZN(n13765) );
  NOR2_X1 U12190 ( .A1(n15222), .A2(n15223), .ZN(n15224) );
  AND2_X1 U12191 ( .A1(n11129), .A2(n10559), .ZN(n12077) );
  AOI22_X1 U12192 ( .A1(n12901), .A2(n12075), .B1(n12074), .B2(n12896), .ZN(
        n12860) );
  AND2_X1 U12193 ( .A1(n12372), .A2(n12371), .ZN(n19369) );
  INV_X1 U12194 ( .A(n12093), .ZN(n13098) );
  INV_X1 U12195 ( .A(n10165), .ZN(n10163) );
  NAND2_X1 U12196 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n15479), .ZN(
        n15469) );
  AND2_X1 U12197 ( .A1(n16282), .A2(n10180), .ZN(n15479) );
  AND2_X1 U12198 ( .A1(n9840), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10180) );
  NAND2_X1 U12199 ( .A1(n16282), .A2(n9840), .ZN(n15493) );
  NAND2_X1 U12200 ( .A1(n16282), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16281) );
  NOR2_X1 U12201 ( .A1(n16405), .A2(n16283), .ZN(n16282) );
  NAND2_X1 U12202 ( .A1(n15514), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16283) );
  NAND2_X1 U12203 ( .A1(n15191), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15190) );
  NOR2_X1 U12204 ( .A1(n15190), .A2(n15538), .ZN(n15514) );
  OR2_X1 U12205 ( .A1(n15355), .A2(n15347), .ZN(n15349) );
  OR2_X1 U12206 ( .A1(n13849), .A2(n15353), .ZN(n15355) );
  AND2_X1 U12207 ( .A1(n15186), .A2(n10176), .ZN(n15189) );
  AND2_X1 U12208 ( .A1(n9835), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10176) );
  NAND2_X1 U12209 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n15189), .ZN(
        n15188) );
  AND2_X1 U12210 ( .A1(n9841), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10313) );
  NAND2_X1 U12211 ( .A1(n15186), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15185) );
  NOR2_X1 U12212 ( .A1(n19197), .A2(n15183), .ZN(n15186) );
  NAND2_X1 U12213 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n15184), .ZN(
        n15183) );
  AND2_X1 U12214 ( .A1(n15181), .A2(n10172), .ZN(n15184) );
  AND2_X1 U12215 ( .A1(n9819), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10172) );
  NAND2_X1 U12216 ( .A1(n15181), .A2(n9819), .ZN(n15182) );
  NAND2_X1 U12217 ( .A1(n15181), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15180) );
  AND2_X1 U12218 ( .A1(n10295), .A2(n9833), .ZN(n14522) );
  INV_X1 U12219 ( .A(n13475), .ZN(n10292) );
  NAND3_X1 U12220 ( .A1(n10171), .A2(n10169), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15178) );
  NOR2_X1 U12221 ( .A1(n16499), .A2(n10170), .ZN(n10169) );
  NAND3_X1 U12222 ( .A1(n10600), .A2(n10599), .A3(n10433), .ZN(n10636) );
  AOI22_X1 U12223 ( .A1(n12868), .A2(n16562), .B1(n12184), .B2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10606) );
  NAND2_X2 U12224 ( .A1(n10636), .A2(n10637), .ZN(n10042) );
  NAND2_X1 U12225 ( .A1(n11001), .A2(n10332), .ZN(n10333) );
  AND2_X1 U12226 ( .A1(n10335), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10332) );
  NAND2_X1 U12227 ( .A1(n10331), .A2(n12102), .ZN(n10189) );
  NOR2_X1 U12228 ( .A1(n10334), .A2(n10127), .ZN(n10331) );
  NAND2_X1 U12229 ( .A1(n10335), .A2(n10336), .ZN(n10188) );
  NOR2_X1 U12230 ( .A1(n9856), .A2(n10339), .ZN(n10338) );
  INV_X1 U12231 ( .A(n15445), .ZN(n10339) );
  NAND2_X1 U12232 ( .A1(n15392), .A2(n10265), .ZN(n14476) );
  AND2_X1 U12233 ( .A1(n9928), .A2(n10266), .ZN(n10265) );
  INV_X1 U12234 ( .A(n11444), .ZN(n10266) );
  NAND2_X1 U12235 ( .A1(n10350), .A2(n10127), .ZN(n10123) );
  NAND2_X1 U12236 ( .A1(n10121), .A2(n10127), .ZN(n10120) );
  AOI21_X1 U12237 ( .B1(n12102), .B2(n10113), .A(n10111), .ZN(n10110) );
  NOR2_X1 U12238 ( .A1(n10114), .A2(n10127), .ZN(n10113) );
  NAND2_X1 U12239 ( .A1(n10112), .A2(n15445), .ZN(n10111) );
  NAND2_X1 U12240 ( .A1(n10336), .A2(n14451), .ZN(n10112) );
  NAND2_X1 U12241 ( .A1(n12104), .A2(n10337), .ZN(n10336) );
  NAND2_X1 U12242 ( .A1(n12107), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10337) );
  NAND2_X1 U12243 ( .A1(n11001), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9981) );
  NOR3_X1 U12244 ( .A1(n9815), .A2(n10296), .A3(n10298), .ZN(n12113) );
  NAND2_X1 U12245 ( .A1(n15296), .A2(n12115), .ZN(n10296) );
  INV_X1 U12246 ( .A(n15471), .ZN(n10284) );
  NOR2_X1 U12247 ( .A1(n12103), .A2(n12102), .ZN(n15477) );
  NOR2_X2 U12248 ( .A1(n15521), .A2(n16530), .ZN(n16400) );
  INV_X1 U12249 ( .A(n9929), .ZN(n10261) );
  NOR3_X1 U12250 ( .A1(n15349), .A2(n15335), .A3(n15192), .ZN(n15336) );
  NOR2_X1 U12251 ( .A1(n15430), .A2(n15195), .ZN(n15410) );
  AND2_X1 U12252 ( .A1(n13658), .A2(n9895), .ZN(n13851) );
  AND2_X1 U12253 ( .A1(n11417), .A2(n11416), .ZN(n13839) );
  NAND2_X1 U12254 ( .A1(n13658), .A2(n13602), .ZN(n13749) );
  NAND2_X1 U12255 ( .A1(n13658), .A2(n9889), .ZN(n13766) );
  AND2_X1 U12256 ( .A1(n16443), .A2(n10313), .ZN(n15721) );
  NAND2_X1 U12257 ( .A1(n9968), .A2(n9967), .ZN(n15527) );
  NAND2_X1 U12258 ( .A1(n16443), .A2(n9841), .ZN(n15760) );
  NOR2_X1 U12259 ( .A1(n9818), .A2(n10279), .ZN(n10278) );
  INV_X1 U12260 ( .A(n13396), .ZN(n10279) );
  NAND2_X1 U12261 ( .A1(n16443), .A2(n15648), .ZN(n16442) );
  OAI211_X1 U12262 ( .C1(n13830), .C2(n10118), .A(n15524), .B(n10116), .ZN(
        n15778) );
  INV_X1 U12263 ( .A(n10911), .ZN(n10118) );
  NAND2_X1 U12264 ( .A1(n10117), .A2(n10911), .ZN(n10116) );
  INV_X1 U12265 ( .A(n10119), .ZN(n10117) );
  NAND2_X1 U12266 ( .A1(n10277), .A2(n9890), .ZN(n13387) );
  NOR2_X1 U12267 ( .A1(n16562), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12184) );
  INV_X1 U12268 ( .A(n12841), .ZN(n11180) );
  NOR2_X1 U12269 ( .A1(n13138), .A2(n13137), .ZN(n13144) );
  NAND2_X1 U12271 ( .A1(n10250), .A2(n13058), .ZN(n10248) );
  OR2_X1 U12272 ( .A1(n15802), .A2(n15803), .ZN(n15805) );
  AND2_X1 U12273 ( .A1(n15236), .A2(n10914), .ZN(n16436) );
  NAND2_X1 U12274 ( .A1(n10306), .A2(n10311), .ZN(n15600) );
  NAND2_X1 U12275 ( .A1(n15829), .A2(n10312), .ZN(n10306) );
  OR2_X1 U12276 ( .A1(n13052), .A2(n9894), .ZN(n13062) );
  INV_X1 U12277 ( .A(n10044), .ZN(n10344) );
  NAND2_X1 U12278 ( .A1(n11097), .A2(n11096), .ZN(n13826) );
  NAND2_X1 U12279 ( .A1(n13553), .A2(n11299), .ZN(n13470) );
  AND2_X1 U12280 ( .A1(n13470), .A2(n13469), .ZN(n13472) );
  XNOR2_X1 U12281 ( .A(n10845), .B(n13642), .ZN(n13640) );
  NAND2_X1 U12282 ( .A1(n13647), .A2(n13646), .ZN(n13645) );
  OR2_X1 U12283 ( .A1(n11076), .A2(n13642), .ZN(n13650) );
  NAND2_X1 U12284 ( .A1(n9920), .A2(n10295), .ZN(n13476) );
  NOR2_X1 U12285 ( .A1(n10291), .A2(n10294), .ZN(n10290) );
  NAND2_X1 U12286 ( .A1(n15835), .A2(n15836), .ZN(n15838) );
  INV_X2 U12287 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12923) );
  INV_X1 U12288 ( .A(n14491), .ZN(n19277) );
  NOR2_X2 U12289 ( .A1(n13098), .A2(n16486), .ZN(n19465) );
  NOR2_X2 U12290 ( .A1(n13097), .A2(n16486), .ZN(n19466) );
  INV_X1 U12291 ( .A(n19465), .ZN(n19456) );
  INV_X1 U12292 ( .A(n19466), .ZN(n19458) );
  NOR3_X1 U12293 ( .A1(n9810), .A2(n12150), .A3(n18889), .ZN(n18870) );
  OR2_X1 U12294 ( .A1(n16841), .A2(n17793), .ZN(n16839) );
  AND2_X1 U12295 ( .A1(n16873), .A2(n9807), .ZN(n16862) );
  OR2_X1 U12296 ( .A1(n16875), .A2(n17837), .ZN(n16873) );
  INV_X1 U12297 ( .A(n17143), .ZN(n17073) );
  NOR2_X1 U12298 ( .A1(n18870), .A2(n17683), .ZN(n17080) );
  INV_X1 U12299 ( .A(n17467), .ZN(n17462) );
  NOR2_X1 U12300 ( .A1(n17706), .A2(n10080), .ZN(n10079) );
  INV_X1 U12301 ( .A(n11461), .ZN(n17372) );
  NOR2_X1 U12302 ( .A1(n17683), .A2(n17645), .ZN(n17663) );
  NOR2_X1 U12303 ( .A1(n18929), .A2(n16750), .ZN(n17684) );
  NOR2_X1 U12304 ( .A1(n17786), .A2(n18114), .ZN(n18117) );
  NAND2_X1 U12305 ( .A1(n17950), .A2(n9824), .ZN(n17879) );
  NOR2_X1 U12306 ( .A1(n17934), .A2(n17933), .ZN(n17950) );
  AND3_X1 U12307 ( .A1(n17991), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17962) );
  AND2_X1 U12308 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17991) );
  INV_X1 U12309 ( .A(n17991), .ZN(n18005) );
  NAND2_X1 U12310 ( .A1(n17961), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17933) );
  NOR2_X1 U12311 ( .A1(n18048), .A2(n18049), .ZN(n17961) );
  INV_X1 U12312 ( .A(n17076), .ZN(n18061) );
  NOR2_X1 U12313 ( .A1(n16644), .A2(n9917), .ZN(n15883) );
  NAND2_X1 U12314 ( .A1(n10221), .A2(n10220), .ZN(n16642) );
  NAND2_X1 U12315 ( .A1(n16653), .A2(n10223), .ZN(n10220) );
  NAND2_X1 U12316 ( .A1(n11738), .A2(n10218), .ZN(n10221) );
  NAND2_X1 U12317 ( .A1(n17927), .A2(n10096), .ZN(n17786) );
  NOR3_X1 U12318 ( .A1(n11727), .A2(n18181), .A3(n10097), .ZN(n10096) );
  NAND2_X1 U12319 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10097) );
  NAND2_X1 U12320 ( .A1(n17897), .A2(n10216), .ZN(n18148) );
  AND4_X1 U12321 ( .A1(n10213), .A2(n10211), .A3(n10210), .A4(n10209), .ZN(
        n17796) );
  AOI22_X1 U12322 ( .A1(n11733), .A2(n10212), .B1(n17969), .B2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10211) );
  OR2_X1 U12323 ( .A1(n10318), .A2(n18002), .ZN(n10210) );
  OR2_X1 U12324 ( .A1(n17897), .A2(n10214), .ZN(n10213) );
  NOR2_X1 U12325 ( .A1(n10158), .A2(n18467), .ZN(n10156) );
  NAND2_X1 U12326 ( .A1(n17924), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18249) );
  INV_X1 U12327 ( .A(n10107), .ZN(n10106) );
  AOI21_X1 U12328 ( .B1(n9845), .B2(n18337), .A(n18287), .ZN(n10107) );
  INV_X1 U12329 ( .A(n17967), .ZN(n11699) );
  AND2_X1 U12330 ( .A1(n10108), .A2(n9845), .ZN(n18297) );
  OR2_X1 U12331 ( .A1(n18004), .A2(n18337), .ZN(n10108) );
  OAI22_X1 U12332 ( .A1(n18035), .A2(n10109), .B1(n11720), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18019) );
  AND2_X1 U12333 ( .A1(n11720), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10109) );
  XNOR2_X1 U12334 ( .A(n11681), .B(n10321), .ZN(n18051) );
  INV_X1 U12335 ( .A(n11680), .ZN(n10321) );
  NAND2_X1 U12336 ( .A1(n18057), .A2(n18058), .ZN(n18056) );
  XNOR2_X1 U12337 ( .A(n11676), .B(n11675), .ZN(n18070) );
  NAND2_X1 U12338 ( .A1(n18070), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18069) );
  NAND2_X1 U12339 ( .A1(n18081), .A2(n18080), .ZN(n18079) );
  NOR2_X1 U12340 ( .A1(n10322), .A2(n11670), .ZN(n18102) );
  NAND2_X1 U12341 ( .A1(n10155), .A2(n13951), .ZN(n18891) );
  NAND2_X1 U12342 ( .A1(n11577), .A2(n10156), .ZN(n10155) );
  NAND2_X1 U12343 ( .A1(n11577), .A2(n10157), .ZN(n18885) );
  INV_X1 U12344 ( .A(n10084), .ZN(n18889) );
  OAI211_X1 U12345 ( .C1(n17321), .C2(n17311), .A(n11506), .B(n11505), .ZN(
        n18441) );
  AOI211_X1 U12346 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n11504), .B(n11503), .ZN(n11505) );
  INV_X1 U12347 ( .A(n11601), .ZN(n18452) );
  NOR2_X1 U12348 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18440), .ZN(n18739) );
  NAND2_X1 U12349 ( .A1(n10148), .A2(n10147), .ZN(n18920) );
  NAND2_X1 U12350 ( .A1(n11603), .A2(n18872), .ZN(n10147) );
  NAND2_X1 U12351 ( .A1(n18867), .A2(n18868), .ZN(n10148) );
  INV_X1 U12352 ( .A(n13111), .ZN(n20089) );
  INV_X1 U12353 ( .A(n13348), .ZN(n20900) );
  NAND2_X1 U12354 ( .A1(n16027), .A2(n10060), .ZN(n14694) );
  AND2_X1 U12355 ( .A1(n10061), .A2(n14606), .ZN(n10060) );
  AND2_X1 U12356 ( .A1(n16031), .A2(n14538), .ZN(n14766) );
  NAND2_X1 U12357 ( .A1(n16027), .A2(n15999), .ZN(n16012) );
  INV_X1 U12358 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16008) );
  NOR2_X1 U12359 ( .A1(n21200), .A2(n14602), .ZN(n16027) );
  NOR2_X1 U12360 ( .A1(n21048), .A2(n16039), .ZN(n14516) );
  NOR3_X1 U12361 ( .A1(n20131), .A2(n13944), .A3(n13790), .ZN(n20116) );
  NOR2_X1 U12362 ( .A1(n20146), .A2(n21162), .ZN(n13727) );
  INV_X1 U12363 ( .A(n20154), .ZN(n20138) );
  NAND2_X1 U12364 ( .A1(n13593), .A2(n13592), .ZN(n20146) );
  INV_X1 U12365 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13419) );
  INV_X1 U12366 ( .A(n20153), .ZN(n20136) );
  AND2_X1 U12367 ( .A1(n13595), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20153) );
  INV_X1 U12368 ( .A(n20162), .ZN(n20144) );
  AND2_X2 U12369 ( .A1(n12640), .A2(n13111), .ZN(n20185) );
  INV_X1 U12370 ( .A(n20181), .ZN(n20171) );
  INV_X1 U12371 ( .A(n14813), .ZN(n14861) );
  INV_X1 U12372 ( .A(n14827), .ZN(n14863) );
  OR2_X1 U12373 ( .A1(n13110), .A2(n13109), .ZN(n13112) );
  INV_X2 U12374 ( .A(n14873), .ZN(n14879) );
  OR2_X1 U12375 ( .A1(n14873), .A2(n13115), .ZN(n14878) );
  AND2_X1 U12376 ( .A1(n12584), .A2(n13365), .ZN(n20189) );
  AND2_X1 U12377 ( .A1(n12623), .A2(n12508), .ZN(n20225) );
  CLKBUF_X1 U12378 ( .A(n14728), .Z(n14729) );
  NAND2_X1 U12379 ( .A1(n13906), .A2(n13905), .ZN(n14051) );
  INV_X1 U12380 ( .A(n16110), .ZN(n16084) );
  INV_X1 U12381 ( .A(n16116), .ZN(n16099) );
  XNOR2_X1 U12382 ( .A(n10352), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15048) );
  NAND2_X1 U12383 ( .A1(n10355), .A2(n10353), .ZN(n10352) );
  AND2_X1 U12384 ( .A1(n14639), .A2(n14638), .ZN(n15073) );
  OR3_X1 U12385 ( .A1(n15110), .A2(n15041), .A3(n15029), .ZN(n15078) );
  INV_X1 U12386 ( .A(n10139), .ZN(n14911) );
  INV_X1 U12387 ( .A(n10356), .ZN(n14955) );
  NAND2_X1 U12388 ( .A1(n10361), .A2(n13616), .ZN(n13771) );
  NAND2_X1 U12389 ( .A1(n16108), .A2(n16109), .ZN(n10361) );
  AND2_X1 U12390 ( .A1(n13021), .A2(n13008), .ZN(n16268) );
  AND2_X1 U12391 ( .A1(n13013), .A2(n16129), .ZN(n13038) );
  AND2_X1 U12392 ( .A1(n16133), .A2(n16136), .ZN(n16201) );
  NAND2_X1 U12393 ( .A1(n12765), .A2(n14597), .ZN(n13022) );
  XNOR2_X1 U12394 ( .A(n10229), .B(n12764), .ZN(n12765) );
  AND2_X1 U12395 ( .A1(n13021), .A2(n13020), .ZN(n16263) );
  INV_X1 U12396 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20670) );
  INV_X1 U12397 ( .A(n10141), .ZN(n20881) );
  INV_X1 U12398 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20228) );
  OAI21_X1 U12399 ( .B1(n13210), .B2(n16277), .A(n20396), .ZN(n20892) );
  AND2_X1 U12400 ( .A1(n20360), .A2(n20307), .ZN(n20351) );
  OAI21_X1 U12401 ( .B1(n20412), .B2(n20397), .A(n20708), .ZN(n20415) );
  OAI211_X1 U12402 ( .C1(n20463), .C2(n20637), .A(n20708), .B(n20448), .ZN(
        n20465) );
  NOR2_X2 U12403 ( .A1(n20473), .A2(n20669), .ZN(n20464) );
  OAI211_X1 U12404 ( .C1(n20518), .C2(n20637), .A(n20559), .B(n20503), .ZN(
        n20521) );
  OAI211_X1 U12405 ( .C1(n20662), .C2(n20637), .A(n20708), .B(n20636), .ZN(
        n20664) );
  NOR2_X2 U12406 ( .A1(n20602), .A2(n20601), .ZN(n20663) );
  INV_X1 U12407 ( .A(n20676), .ZN(n20694) );
  OAI211_X1 U12408 ( .C1(n20733), .C2(n20709), .A(n20708), .B(n20707), .ZN(
        n20737) );
  INV_X1 U12409 ( .A(n20710), .ZN(n20736) );
  INV_X1 U12410 ( .A(n20553), .ZN(n20744) );
  INV_X1 U12411 ( .A(n20562), .ZN(n20757) );
  INV_X1 U12412 ( .A(n20566), .ZN(n20763) );
  INV_X1 U12413 ( .A(n20570), .ZN(n20769) );
  INV_X1 U12414 ( .A(n20574), .ZN(n20775) );
  INV_X1 U12415 ( .A(n20578), .ZN(n20780) );
  INV_X1 U12416 ( .A(n20583), .ZN(n20785) );
  OR2_X1 U12417 ( .A1(n20698), .A2(n20697), .ZN(n20801) );
  INV_X1 U12418 ( .A(n20790), .ZN(n20797) );
  NOR2_X1 U12419 ( .A1(n20637), .A2(n12997), .ZN(n15958) );
  INV_X1 U12420 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20637) );
  OR2_X1 U12421 ( .A1(n12175), .A2(n12897), .ZN(n19104) );
  NAND2_X1 U12422 ( .A1(n11028), .A2(n11027), .ZN(n20076) );
  INV_X1 U12423 ( .A(n19266), .ZN(n19288) );
  NOR2_X1 U12424 ( .A1(n14491), .A2(n19301), .ZN(n19199) );
  INV_X1 U12425 ( .A(n19293), .ZN(n19271) );
  OR2_X1 U12426 ( .A1(n11382), .A2(n11381), .ZN(n13394) );
  OR2_X1 U12427 ( .A1(n11343), .A2(n11342), .ZN(n13136) );
  NOR2_X1 U12428 ( .A1(n11330), .A2(n11329), .ZN(n12840) );
  OR2_X1 U12429 ( .A1(n11315), .A2(n11314), .ZN(n12837) );
  CLKBUF_X1 U12430 ( .A(n12835), .Z(n12836) );
  AND2_X1 U12431 ( .A1(n12712), .A2(n12715), .ZN(n19326) );
  INV_X1 U12432 ( .A(n15346), .ZN(n15359) );
  AND2_X1 U12433 ( .A1(n12111), .A2(n11443), .ZN(n16319) );
  INV_X1 U12434 ( .A(n9992), .ZN(n9991) );
  CLKBUF_X1 U12435 ( .A(n15300), .Z(n15301) );
  INV_X1 U12436 ( .A(n16381), .ZN(n15404) );
  INV_X1 U12437 ( .A(n19360), .ZN(n19334) );
  INV_X1 U12438 ( .A(n19333), .ZN(n19359) );
  NOR2_X2 U12439 ( .A1(n19359), .A2(n12079), .ZN(n19361) );
  NOR2_X1 U12440 ( .A1(n19369), .A2(n19400), .ZN(n19384) );
  CLKBUF_X1 U12442 ( .A(n19376), .Z(n19400) );
  NOR2_X1 U12443 ( .A1(n12626), .A2(n11259), .ZN(n12801) );
  OR2_X1 U12444 ( .A1(n15723), .A2(n15550), .ZN(n15584) );
  INV_X1 U12445 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16473) );
  AND2_X1 U12446 ( .A1(n10295), .A2(n10289), .ZN(n12697) );
  INV_X1 U12447 ( .A(n16498), .ZN(n16477) );
  INV_X1 U12448 ( .A(n16478), .ZN(n16493) );
  NAND2_X1 U12449 ( .A1(n15609), .A2(n10256), .ZN(n10255) );
  INV_X1 U12450 ( .A(n10257), .ZN(n10256) );
  OAI21_X1 U12451 ( .B1(n16295), .B2(n19411), .A(n10258), .ZN(n10257) );
  OR2_X1 U12452 ( .A1(n12112), .A2(n15297), .ZN(n16329) );
  OR2_X1 U12453 ( .A1(n15490), .A2(n15489), .ZN(n16512) );
  AND2_X1 U12454 ( .A1(n10349), .A2(n10347), .ZN(n15486) );
  NAND2_X1 U12455 ( .A1(n16396), .A2(n10983), .ZN(n15503) );
  NAND2_X1 U12456 ( .A1(n10059), .A2(n10972), .ZN(n15512) );
  NAND2_X1 U12457 ( .A1(n10054), .A2(n10053), .ZN(n10059) );
  XNOR2_X1 U12458 ( .A(n9966), .B(n9898), .ZN(n15685) );
  AOI21_X1 U12459 ( .B1(n15569), .B2(n15566), .A(n15561), .ZN(n9966) );
  NAND2_X1 U12460 ( .A1(n15564), .A2(n10317), .ZN(n15674) );
  OR2_X1 U12461 ( .A1(n15570), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10317) );
  NAND2_X1 U12462 ( .A1(n10054), .A2(n15776), .ZN(n15771) );
  NAND2_X1 U12463 ( .A1(n13830), .A2(n10883), .ZN(n15822) );
  NAND2_X1 U12464 ( .A1(n10841), .A2(n10130), .ZN(n13512) );
  NAND2_X1 U12465 ( .A1(n9960), .A2(n15249), .ZN(n13152) );
  OR2_X1 U12466 ( .A1(n15846), .A2(n12633), .ZN(n20069) );
  INV_X1 U12467 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20056) );
  NAND2_X1 U12468 ( .A1(n12398), .A2(n11282), .ZN(n13158) );
  INV_X1 U12469 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15986) );
  XNOR2_X1 U12470 ( .A(n12683), .B(n12682), .ZN(n20038) );
  XNOR2_X1 U12471 ( .A(n12597), .B(n12599), .ZN(n20051) );
  NAND2_X1 U12472 ( .A1(n12901), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20031) );
  NOR2_X1 U12473 ( .A1(n19666), .A2(n19597), .ZN(n19522) );
  INV_X1 U12474 ( .A(n19582), .ZN(n19574) );
  OR3_X1 U12475 ( .A1(n19628), .A2(n19888), .A3(n19627), .ZN(n19647) );
  INV_X1 U12476 ( .A(n19641), .ZN(n19646) );
  INV_X1 U12477 ( .A(n19723), .ZN(n19724) );
  OAI21_X1 U12478 ( .B1(n19827), .B2(n13298), .A(n19804), .ZN(n19829) );
  INV_X1 U12479 ( .A(n19897), .ZN(n19805) );
  INV_X1 U12480 ( .A(n19901), .ZN(n19853) );
  INV_X1 U12481 ( .A(n19906), .ZN(n19856) );
  INV_X1 U12482 ( .A(n19911), .ZN(n19860) );
  INV_X1 U12483 ( .A(n19916), .ZN(n19863) );
  OAI22_X1 U12484 ( .A1(n20235), .A2(n19458), .B1(n18442), .B2(n19456), .ZN(
        n19894) );
  OAI22_X1 U12485 ( .A1(n20259), .A2(n19458), .B1(n19438), .B2(n19456), .ZN(
        n19903) );
  OAI22_X1 U12486 ( .A1(n14815), .A2(n19458), .B1(n19450), .B2(n19456), .ZN(
        n19913) );
  INV_X1 U12487 ( .A(n19823), .ZN(n19917) );
  INV_X1 U12488 ( .A(n19826), .ZN(n19922) );
  NAND2_X1 U12489 ( .A1(n19760), .A2(n19892), .ZN(n19934) );
  OAI22_X1 U12490 ( .A1(n20293), .A2(n19458), .B1(n19457), .B2(n19456), .ZN(
        n19929) );
  AND2_X1 U12491 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11074), .ZN(n16570) );
  INV_X1 U12492 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20067) );
  INV_X2 U12493 ( .A(n11751), .ZN(n16562) );
  INV_X1 U12494 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n11751) );
  NOR2_X1 U12495 ( .A1(n9810), .A2(n13957), .ZN(n16752) );
  INV_X1 U12496 ( .A(n17684), .ZN(n17683) );
  AND2_X1 U12497 ( .A1(n16839), .A2(n9807), .ZN(n16828) );
  AND2_X1 U12498 ( .A1(n17096), .A2(n10268), .ZN(n16895) );
  NAND2_X1 U12499 ( .A1(n17817), .A2(n16914), .ZN(n10268) );
  NOR2_X1 U12500 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17007), .ZN(n17006) );
  INV_X1 U12501 ( .A(n17121), .ZN(n17132) );
  NOR2_X1 U12502 ( .A1(n18922), .A2(n12164), .ZN(n17121) );
  NAND3_X1 U12503 ( .A1(n17066), .A2(n19097), .A3(n18927), .ZN(n17143) );
  INV_X1 U12504 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17459) );
  AND3_X1 U12505 ( .A1(n11495), .A2(n10418), .A3(n11494), .ZN(n10430) );
  NOR4_X1 U12506 ( .A1(n19084), .A2(n17081), .A3(n15987), .A4(n18929), .ZN(
        n17485) );
  INV_X1 U12507 ( .A(n17485), .ZN(n17488) );
  INV_X1 U12508 ( .A(n17482), .ZN(n17491) );
  NOR2_X1 U12509 ( .A1(n17488), .A2(n10430), .ZN(n17489) );
  INV_X1 U12510 ( .A(n17502), .ZN(n17498) );
  NAND2_X1 U12511 ( .A1(n17520), .A2(n9842), .ZN(n17511) );
  INV_X1 U12512 ( .A(n17526), .ZN(n17520) );
  NAND2_X1 U12513 ( .A1(n17520), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17519) );
  NOR2_X1 U12514 ( .A1(n17568), .A2(n10093), .ZN(n17530) );
  INV_X1 U12515 ( .A(n17541), .ZN(n10094) );
  NAND2_X1 U12516 ( .A1(n17530), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17529) );
  NOR2_X1 U12517 ( .A1(n17535), .A2(n17562), .ZN(n17551) );
  INV_X1 U12518 ( .A(n17572), .ZN(n17555) );
  NOR2_X1 U12519 ( .A1(n17750), .A2(n17575), .ZN(n17569) );
  NAND2_X1 U12520 ( .A1(n17569), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17568) );
  NOR2_X2 U12521 ( .A1(n18467), .A2(n17641), .ZN(n17567) );
  NOR2_X1 U12522 ( .A1(n17738), .A2(n17597), .ZN(n17590) );
  NOR2_X1 U12523 ( .A1(n17640), .A2(n17573), .ZN(n17608) );
  INV_X1 U12524 ( .A(n11704), .ZN(n17621) );
  INV_X1 U12525 ( .A(n11703), .ZN(n17628) );
  OR2_X1 U12526 ( .A1(n11634), .A2(n11633), .ZN(n10197) );
  AND2_X1 U12527 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11633) );
  INV_X1 U12528 ( .A(n17638), .ZN(n17633) );
  NOR2_X1 U12529 ( .A1(n11648), .A2(n11647), .ZN(n11649) );
  INV_X1 U12530 ( .A(n11645), .ZN(n10098) );
  AND2_X1 U12531 ( .A1(n11626), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11647) );
  NAND2_X1 U12532 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17642), .ZN(n17640) );
  INV_X2 U12533 ( .A(n17609), .ZN(n17641) );
  NOR2_X1 U12534 ( .A1(n17494), .A2(n17716), .ZN(n17642) );
  NOR2_X2 U12535 ( .A1(n18899), .A2(n17494), .ZN(n17638) );
  NOR2_X1 U12536 ( .A1(n15990), .A2(n17494), .ZN(n17639) );
  NOR2_X1 U12537 ( .A1(n19081), .A2(n17663), .ZN(n17660) );
  CLKBUF_X1 U12538 ( .A(n17660), .Z(n17679) );
  OAI211_X1 U12539 ( .C1(n19084), .C2(n19085), .A(n9810), .B(n17684), .ZN(
        n17744) );
  NAND2_X1 U12541 ( .A1(n10199), .A2(n10198), .ZN(n17765) );
  AND2_X1 U12542 ( .A1(n17885), .A2(n10159), .ZN(n17863) );
  NOR2_X1 U12543 ( .A1(n18181), .A2(n18221), .ZN(n10159) );
  AND2_X1 U12544 ( .A1(n17984), .A2(n10160), .ZN(n17885) );
  INV_X1 U12545 ( .A(n18213), .ZN(n10160) );
  INV_X1 U12546 ( .A(n17885), .ZN(n17899) );
  INV_X1 U12547 ( .A(n18815), .ZN(n18482) );
  NAND2_X1 U12548 ( .A1(n17950), .A2(n10426), .ZN(n17921) );
  OAI22_X1 U12549 ( .A1(n18297), .A2(n18108), .B1(n17943), .B2(n18295), .ZN(
        n17984) );
  INV_X1 U12550 ( .A(n17984), .ZN(n18000) );
  INV_X1 U12551 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18009) );
  INV_X1 U12552 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18023) );
  INV_X1 U12553 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18049) );
  NOR2_X2 U12554 ( .A1(n18488), .A2(n18599), .ZN(n18815) );
  NAND2_X1 U12555 ( .A1(n18103), .A2(n18060), .ZN(n18098) );
  INV_X1 U12556 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19042) );
  NAND2_X1 U12557 ( .A1(n18920), .A2(n10146), .ZN(n18107) );
  NOR2_X1 U12558 ( .A1(n19084), .A2(n18929), .ZN(n10146) );
  INV_X1 U12559 ( .A(n10222), .ZN(n17753) );
  AND2_X1 U12560 ( .A1(n18127), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10104) );
  OR2_X1 U12561 ( .A1(n18129), .A2(n18344), .ZN(n10101) );
  INV_X1 U12562 ( .A(n10217), .ZN(n17877) );
  NAND2_X1 U12563 ( .A1(n17896), .A2(n10318), .ZN(n17878) );
  NAND2_X1 U12564 ( .A1(n17613), .A2(n18423), .ZN(n18344) );
  INV_X1 U12565 ( .A(n18410), .ZN(n18404) );
  AOI21_X2 U12566 ( .B1(n15893), .B2(n15892), .A(n18929), .ZN(n18409) );
  AOI211_X1 U12567 ( .C1(n18872), .C2(n15889), .A(n15888), .B(n15887), .ZN(
        n15893) );
  NAND2_X1 U12568 ( .A1(n18426), .A2(n18427), .ZN(n18410) );
  INV_X1 U12569 ( .A(n18409), .ZN(n18427) );
  INV_X1 U12570 ( .A(n18385), .ZN(n18425) );
  NOR2_X1 U12571 ( .A1(n18427), .A2(n18873), .ZN(n18423) );
  INV_X1 U12572 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18905) );
  INV_X1 U12573 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18910) );
  OAI211_X1 U12574 ( .C1(n18929), .C2(n18908), .A(n18439), .B(n15872), .ZN(
        n19062) );
  INV_X1 U12575 ( .A(n19062), .ZN(n19065) );
  AND2_X1 U12576 ( .A1(n12144), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20230)
         );
  CLKBUF_X1 U12577 ( .A(n16733), .Z(n16739) );
  AOI211_X1 U12578 ( .C1(n14609), .C2(P1_REIP_REG_31__SCAN_IN), .A(n10076), 
        .B(n10235), .ZN(n10075) );
  NAND2_X1 U12579 ( .A1(n14536), .A2(n20128), .ZN(n10077) );
  NAND2_X1 U12580 ( .A1(n10132), .A2(n16105), .ZN(n10131) );
  AND2_X1 U12581 ( .A1(n16304), .A2(n16305), .ZN(n10161) );
  OAI21_X1 U12582 ( .B1(n16295), .B2(n15352), .A(n12129), .ZN(n12130) );
  NAND2_X1 U12583 ( .A1(n9990), .A2(n9988), .ZN(P2_U2858) );
  INV_X1 U12584 ( .A(n9989), .ZN(n9988) );
  OAI21_X1 U12585 ( .B1(n16309), .B2(n15352), .A(n15286), .ZN(n9989) );
  AOI211_X1 U12586 ( .C1(n16491), .C2(n16291), .A(n15442), .B(n15441), .ZN(
        n15443) );
  AOI21_X1 U12587 ( .B1(n16521), .B2(n16494), .A(n10045), .ZN(n16393) );
  NAND2_X1 U12588 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  OAI21_X1 U12589 ( .B1(n15674), .B2(n16478), .A(n10315), .ZN(P2_U2995) );
  INV_X1 U12590 ( .A(n9965), .ZN(n10315) );
  OAI21_X1 U12591 ( .B1(n15685), .B2(n16480), .A(n10316), .ZN(n9965) );
  AOI21_X1 U12592 ( .B1(n19148), .B2(n16491), .A(n15565), .ZN(n10316) );
  NOR2_X1 U12593 ( .A1(n10422), .A2(n14489), .ZN(n14490) );
  OAI21_X1 U12594 ( .B1(n16309), .B2(n19411), .A(n11454), .ZN(n11455) );
  NAND2_X1 U12595 ( .A1(n12123), .A2(n10282), .ZN(P2_U3018) );
  AND2_X1 U12596 ( .A1(n10286), .A2(n9877), .ZN(n10282) );
  OR2_X1 U12597 ( .A1(n15468), .A2(n19411), .ZN(n10286) );
  AOI21_X1 U12598 ( .B1(n16787), .B2(n17152), .A(n9861), .ZN(n10274) );
  OAI21_X1 U12599 ( .B1(n16616), .B2(n18015), .A(n9869), .ZN(P3_U2801) );
  OAI211_X1 U12600 ( .C1(n16620), .C2(n9831), .A(n10330), .B(n9872), .ZN(
        n10329) );
  NAND2_X1 U12601 ( .A1(n17820), .A2(n11741), .ZN(n17807) );
  NAND2_X1 U12602 ( .A1(n10102), .A2(n10099), .ZN(P3_U2836) );
  AND2_X1 U12603 ( .A1(n10101), .A2(n10100), .ZN(n10099) );
  OR2_X1 U12604 ( .A1(n10104), .A2(n10103), .ZN(n10102) );
  AOI21_X1 U12605 ( .B1(n18404), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n9934), .ZN(n10100) );
  AND3_X1 U12606 ( .A1(n9814), .A2(n17778), .A3(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9813) );
  INV_X1 U12607 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15250) );
  NAND2_X1 U12608 ( .A1(n10400), .A2(n10404), .ZN(n13764) );
  AND2_X1 U12609 ( .A1(n11741), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9814) );
  OR2_X1 U12610 ( .A1(n15349), .A2(n10301), .ZN(n9815) );
  OR2_X1 U12611 ( .A1(n14722), .A2(n10244), .ZN(n9816) );
  OR3_X1 U12612 ( .A1(n14797), .A2(n10237), .A3(n10236), .ZN(n9817) );
  OR2_X1 U12613 ( .A1(n14791), .A2(n10381), .ZN(n14764) );
  OR2_X1 U12614 ( .A1(n14717), .A2(n10370), .ZN(n14695) );
  INV_X1 U12615 ( .A(n12107), .ZN(n10127) );
  NAND2_X1 U12616 ( .A1(n9985), .A2(n9984), .ZN(n12712) );
  NAND2_X1 U12617 ( .A1(n9890), .A2(n10280), .ZN(n9818) );
  NAND2_X1 U12618 ( .A1(n19064), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11466) );
  AND2_X1 U12619 ( .A1(n10173), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9819) );
  AND2_X1 U12620 ( .A1(n10426), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9820) );
  OR3_X1 U12621 ( .A1(n15349), .A2(n15335), .A3(n10302), .ZN(n9821) );
  AND2_X1 U12622 ( .A1(n9855), .A2(n16237), .ZN(n9822) );
  AND4_X1 U12623 ( .A1(n11476), .A2(n11482), .A3(n10089), .A4(n9880), .ZN(
        n9823) );
  AND2_X1 U12624 ( .A1(n9820), .A2(n10270), .ZN(n9824) );
  AND3_X1 U12625 ( .A1(n12233), .A2(n12234), .A3(n10009), .ZN(n9825) );
  NAND2_X1 U12626 ( .A1(n9991), .A2(n15288), .ZN(n15294) );
  AND2_X1 U12627 ( .A1(n10398), .A2(n10397), .ZN(n15316) );
  INV_X1 U12628 ( .A(n10398), .ZN(n15328) );
  OAI21_X1 U12629 ( .B1(n16398), .B2(n10123), .A(n10120), .ZN(n11000) );
  AND2_X1 U12630 ( .A1(n11282), .A2(n9882), .ZN(n9826) );
  AND2_X1 U12631 ( .A1(n10358), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9827) );
  AND2_X1 U12632 ( .A1(n20233), .A2(n13431), .ZN(n9828) );
  INV_X2 U12633 ( .A(n11253), .ZN(n13682) );
  AND2_X1 U12634 ( .A1(n16644), .A2(n18002), .ZN(n9830) );
  AND2_X1 U12635 ( .A1(n16647), .A2(n16619), .ZN(n9831) );
  AND2_X1 U12636 ( .A1(n12688), .A2(n10292), .ZN(n9832) );
  AND3_X1 U12637 ( .A1(n9832), .A2(n12696), .A3(n10289), .ZN(n9833) );
  INV_X1 U12638 ( .A(n9911), .ZN(n14250) );
  NOR2_X1 U12639 ( .A1(n13745), .A2(n13747), .ZN(n13746) );
  INV_X1 U12640 ( .A(n13317), .ZN(n10171) );
  AND4_X1 U12641 ( .A1(n10171), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9834) );
  AND2_X1 U12642 ( .A1(n10177), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9835) );
  INV_X1 U12643 ( .A(n16652), .ZN(n10223) );
  AND2_X1 U12644 ( .A1(n10354), .A2(n9937), .ZN(n9836) );
  AND2_X1 U12645 ( .A1(n10738), .A2(n10683), .ZN(n9837) );
  OR2_X1 U12646 ( .A1(n10252), .A2(n13839), .ZN(n9838) );
  AND2_X1 U12647 ( .A1(n11782), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9839) );
  NAND2_X1 U12648 ( .A1(n11156), .A2(n11155), .ZN(n10295) );
  OR2_X1 U12649 ( .A1(n12835), .A2(n10410), .ZN(n13135) );
  NAND2_X1 U12650 ( .A1(n9858), .A2(n9823), .ZN(n18448) );
  AND2_X1 U12651 ( .A1(n10181), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9840) );
  AND2_X1 U12652 ( .A1(n15648), .A2(n10314), .ZN(n9841) );
  AND2_X1 U12653 ( .A1(n10079), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9842) );
  OR2_X1 U12654 ( .A1(n12096), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9843) );
  INV_X1 U12655 ( .A(n10384), .ZN(n12928) );
  OR2_X1 U12656 ( .A1(n11722), .A2(n11725), .ZN(n9845) );
  AND2_X2 U12657 ( .A1(n12064), .A2(n12883), .ZN(n10775) );
  OR2_X1 U12658 ( .A1(n11466), .A2(n11460), .ZN(n9847) );
  NAND2_X1 U12659 ( .A1(n16027), .A2(n10061), .ZN(n9848) );
  AND2_X1 U12660 ( .A1(n16078), .A2(n16075), .ZN(n9849) );
  NAND2_X1 U12661 ( .A1(n13830), .A2(n10344), .ZN(n15594) );
  OR2_X1 U12662 ( .A1(n15327), .A2(n15329), .ZN(n10398) );
  AND2_X1 U12663 ( .A1(n10614), .A2(n16562), .ZN(n10630) );
  OR2_X1 U12664 ( .A1(n14791), .A2(n14869), .ZN(n14782) );
  NOR2_X1 U12665 ( .A1(n14717), .A2(n10369), .ZN(n14682) );
  NOR2_X1 U12666 ( .A1(n14791), .A2(n10033), .ZN(n9850) );
  OR2_X1 U12667 ( .A1(n10985), .A2(n10192), .ZN(n9851) );
  INV_X1 U12668 ( .A(n10365), .ZN(n12420) );
  AND2_X1 U12669 ( .A1(n17520), .A2(n10079), .ZN(n9852) );
  OR2_X1 U12670 ( .A1(n16068), .A2(n14052), .ZN(n9853) );
  INV_X1 U12671 ( .A(n16068), .ZN(n10354) );
  INV_X1 U12672 ( .A(n12648), .ZN(n14261) );
  AND2_X1 U12673 ( .A1(n14505), .A2(n14104), .ZN(n14790) );
  AND2_X1 U12674 ( .A1(n13905), .A2(n9853), .ZN(n9854) );
  AND2_X1 U12676 ( .A1(n10424), .A2(n10241), .ZN(n9855) );
  INV_X1 U12677 ( .A(n14451), .ZN(n10114) );
  NAND2_X1 U12678 ( .A1(n10027), .A2(n12673), .ZN(n12720) );
  NOR3_X1 U12679 ( .A1(n14456), .A2(n10807), .A3(n14455), .ZN(n9856) );
  AND2_X1 U12680 ( .A1(n16109), .A2(n13770), .ZN(n9857) );
  AND4_X1 U12681 ( .A1(n11481), .A2(n11480), .A3(n11479), .A4(n11478), .ZN(
        n9858) );
  INV_X1 U12682 ( .A(n12150), .ZN(n13951) );
  NAND2_X1 U12683 ( .A1(n15300), .A2(n15303), .ZN(n15302) );
  AND2_X1 U12684 ( .A1(n15288), .A2(n9993), .ZN(n15293) );
  AND3_X1 U12685 ( .A1(n12235), .A2(n10011), .A3(n10010), .ZN(n9859) );
  OR3_X1 U12686 ( .A1(n10985), .A2(n10984), .A3(n10195), .ZN(n9860) );
  OR3_X1 U12687 ( .A1(n16777), .A2(n10276), .A3(n10275), .ZN(n9861) );
  NOR2_X1 U12688 ( .A1(n17529), .A2(n18478), .ZN(n17525) );
  NOR2_X1 U12689 ( .A1(n15316), .A2(n15318), .ZN(n15317) );
  AND2_X1 U12690 ( .A1(n9854), .A2(n14054), .ZN(n9862) );
  NOR2_X1 U12691 ( .A1(n11732), .A2(n11730), .ZN(n9863) );
  AND2_X1 U12692 ( .A1(n20233), .A2(n10366), .ZN(n9864) );
  OR2_X1 U12693 ( .A1(n16090), .A2(n15133), .ZN(n9865) );
  INV_X1 U12694 ( .A(n10158), .ZN(n10157) );
  AND2_X1 U12695 ( .A1(n10222), .A2(n11738), .ZN(n9866) );
  INV_X1 U12696 ( .A(n15510), .ZN(n10058) );
  OR2_X1 U12697 ( .A1(n13530), .A2(n12337), .ZN(n9867) );
  NAND2_X1 U12698 ( .A1(n9810), .A2(n18448), .ZN(n9868) );
  INV_X2 U12699 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n17094) );
  INV_X2 U12700 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12883) );
  NOR2_X1 U12701 ( .A1(n16617), .A2(n10329), .ZN(n9869) );
  NAND2_X1 U12702 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17892) );
  INV_X1 U12703 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17920) );
  NOR3_X1 U12704 ( .A1(n14791), .A2(n10033), .A3(n10036), .ZN(n9870) );
  INV_X1 U12705 ( .A(n10350), .ZN(n10126) );
  NOR2_X1 U12706 ( .A1(n15499), .A2(n10351), .ZN(n10350) );
  AND2_X1 U12707 ( .A1(n13772), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9871) );
  OR2_X1 U12708 ( .A1(n16614), .A2(n16615), .ZN(n9872) );
  AND2_X2 U12709 ( .A1(n12343), .A2(n12342), .ZN(n12997) );
  INV_X1 U12710 ( .A(n12997), .ZN(n10073) );
  OR2_X1 U12711 ( .A1(n12150), .A2(n11578), .ZN(n9873) );
  NOR2_X1 U12712 ( .A1(n15446), .A2(n10114), .ZN(n10335) );
  INV_X1 U12713 ( .A(n10023), .ZN(n10022) );
  NAND2_X1 U12714 ( .A1(n9854), .A2(n10024), .ZN(n10023) );
  INV_X1 U12715 ( .A(n10143), .ZN(n14069) );
  OAI21_X1 U12716 ( .B1(n10144), .B2(n14068), .A(n10354), .ZN(n10143) );
  OR2_X1 U12717 ( .A1(n10831), .A2(n11023), .ZN(n9874) );
  AND3_X1 U12718 ( .A1(n11530), .A2(n10153), .A3(n10149), .ZN(n9875) );
  AND3_X1 U12719 ( .A1(n11668), .A2(n10327), .A3(n10323), .ZN(n9876) );
  AND3_X1 U12720 ( .A1(n10285), .A2(n12122), .A3(n10283), .ZN(n9877) );
  AND3_X1 U12721 ( .A1(n10006), .A2(n10005), .A3(n10004), .ZN(n9878) );
  NOR2_X1 U12722 ( .A1(n15608), .A2(n10255), .ZN(n9879) );
  OR2_X1 U12723 ( .A1(n17415), .A2(n13990), .ZN(n9880) );
  AND2_X1 U12724 ( .A1(n9824), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9881) );
  AND2_X1 U12725 ( .A1(n10260), .A2(n19268), .ZN(n9882) );
  AND2_X1 U12726 ( .A1(n9822), .A2(n10242), .ZN(n9883) );
  INV_X1 U12727 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17004) );
  NAND2_X1 U12728 ( .A1(n14451), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9884) );
  BUF_X1 U12729 ( .A(n12660), .Z(n13263) );
  AOI21_X1 U12731 ( .B1(n10823), .B2(n11251), .A(n9976), .ZN(n10842) );
  NOR2_X1 U12732 ( .A1(n13654), .A2(n11785), .ZN(n9885) );
  NAND2_X1 U12733 ( .A1(n13588), .A2(n13589), .ZN(n13724) );
  NAND2_X1 U12734 ( .A1(n10262), .A2(n10263), .ZN(n15411) );
  NOR2_X1 U12735 ( .A1(n13890), .A2(n15345), .ZN(n15342) );
  AND2_X1 U12736 ( .A1(n10400), .A2(n10401), .ZN(n9886) );
  OR2_X1 U12737 ( .A1(n15349), .A2(n15192), .ZN(n9887) );
  OR2_X1 U12738 ( .A1(n13840), .A2(n9838), .ZN(n13855) );
  AND2_X1 U12739 ( .A1(n15181), .A2(n10173), .ZN(n9888) );
  AND2_X1 U12740 ( .A1(n10288), .A2(n13602), .ZN(n9889) );
  AND2_X1 U12741 ( .A1(n10281), .A2(n13143), .ZN(n9890) );
  NOR2_X1 U12742 ( .A1(n13226), .A2(n13227), .ZN(n13228) );
  OR2_X1 U12743 ( .A1(n13358), .A2(n14442), .ZN(n14774) );
  INV_X1 U12744 ( .A(n14774), .ZN(n20128) );
  NOR2_X1 U12745 ( .A1(n15753), .A2(n15206), .ZN(n13753) );
  AND2_X1 U12746 ( .A1(n12712), .A2(n11778), .ZN(n12686) );
  AND2_X1 U12747 ( .A1(n10783), .A2(n13682), .ZN(n9891) );
  OR2_X1 U12748 ( .A1(n9815), .A2(n15312), .ZN(n9892) );
  AND2_X1 U12749 ( .A1(n15249), .A2(n11137), .ZN(n9893) );
  OR2_X1 U12750 ( .A1(n10251), .A2(n13053), .ZN(n9894) );
  AND2_X1 U12751 ( .A1(n9889), .A2(n10287), .ZN(n9895) );
  NOR2_X1 U12752 ( .A1(n10829), .A2(n10828), .ZN(n9896) );
  NOR2_X1 U12753 ( .A1(n13840), .A2(n13839), .ZN(n9897) );
  AND2_X1 U12754 ( .A1(n15560), .A2(n15559), .ZN(n9898) );
  XNOR2_X1 U12755 ( .A(n11897), .B(n11924), .ZN(n15327) );
  XNOR2_X1 U12756 ( .A(n11952), .B(n11949), .ZN(n15309) );
  AND3_X1 U12757 ( .A1(n10187), .A2(n9799), .A3(n10826), .ZN(n9899) );
  AND2_X1 U12758 ( .A1(n10380), .A2(n10379), .ZN(n9900) );
  AND2_X1 U12759 ( .A1(n13445), .A2(n13444), .ZN(n9901) );
  INV_X1 U12760 ( .A(n10243), .ZN(n14687) );
  NOR3_X1 U12761 ( .A1(n14722), .A2(n10245), .A3(n10247), .ZN(n10243) );
  OR2_X1 U12762 ( .A1(n9994), .A2(n11785), .ZN(n9902) );
  AND2_X1 U12763 ( .A1(n11784), .A2(n11783), .ZN(n9903) );
  INV_X2 U12764 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20237) );
  OR2_X1 U12765 ( .A1(n10749), .A2(n10748), .ZN(n11290) );
  NOR2_X1 U12766 ( .A1(n15787), .A2(n15595), .ZN(n9904) );
  OR2_X1 U12767 ( .A1(n14889), .A2(n9937), .ZN(n9905) );
  INV_X1 U12768 ( .A(n10250), .ZN(n10249) );
  NOR2_X1 U12769 ( .A1(n9894), .A2(n13055), .ZN(n10250) );
  OR2_X1 U12770 ( .A1(n17969), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9906) );
  AND2_X1 U12771 ( .A1(n10374), .A2(n10372), .ZN(n9907) );
  AND2_X1 U12772 ( .A1(n9895), .A2(n13850), .ZN(n9908) );
  AND2_X1 U12773 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9909) );
  AND2_X1 U12774 ( .A1(n9837), .A2(n11290), .ZN(n9910) );
  INV_X1 U12775 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16448) );
  INV_X1 U12776 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16499) );
  OR2_X1 U12777 ( .A1(n13113), .A2(n12749), .ZN(n9911) );
  NOR2_X1 U12778 ( .A1(n13139), .A2(n13144), .ZN(n9912) );
  INV_X1 U12779 ( .A(n10984), .ZN(n10194) );
  NOR2_X1 U12780 ( .A1(n12835), .A2(n10408), .ZN(n13382) );
  NAND2_X1 U12781 ( .A1(n10399), .A2(n11782), .ZN(n14521) );
  NOR2_X2 U12782 ( .A1(n20285), .A2(n12749), .ZN(n14128) );
  INV_X1 U12783 ( .A(n14128), .ZN(n10037) );
  AND2_X1 U12784 ( .A1(n15186), .A2(n10177), .ZN(n9913) );
  AND2_X1 U12785 ( .A1(n16282), .A2(n10181), .ZN(n9914) );
  NOR2_X1 U12786 ( .A1(n14525), .A2(n12832), .ZN(n12831) );
  NAND2_X1 U12787 ( .A1(n12483), .A2(n12482), .ZN(n20390) );
  INV_X1 U12788 ( .A(n20390), .ZN(n10142) );
  NAND2_X1 U12789 ( .A1(n11924), .A2(n11923), .ZN(n9915) );
  OR2_X1 U12790 ( .A1(n11251), .A2(n11194), .ZN(n9916) );
  INV_X1 U12791 ( .A(n13920), .ZN(n10040) );
  AND2_X1 U12792 ( .A1(n10399), .A2(n9839), .ZN(n12834) );
  INV_X1 U12793 ( .A(n10239), .ZN(n14787) );
  NOR3_X1 U12794 ( .A1(n14797), .A2(n10237), .A3(n10240), .ZN(n10239) );
  INV_X1 U12795 ( .A(n10140), .ZN(n20359) );
  OR2_X1 U12796 ( .A1(n17969), .A2(n16640), .ZN(n9917) );
  AND2_X1 U12797 ( .A1(n10401), .A2(n13892), .ZN(n9918) );
  OR2_X1 U12798 ( .A1(n12835), .A2(n10406), .ZN(n13654) );
  INV_X1 U12799 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10175) );
  NOR2_X1 U12800 ( .A1(n13052), .A2(n10249), .ZN(n9919) );
  INV_X1 U12801 ( .A(n15296), .ZN(n10297) );
  AND2_X1 U12802 ( .A1(n10289), .A2(n10290), .ZN(n9920) );
  OR2_X1 U12803 ( .A1(n17049), .A2(n16782), .ZN(n9921) );
  INV_X1 U12804 ( .A(n11154), .ZN(n10289) );
  NOR2_X1 U12805 ( .A1(n13052), .A2(n13053), .ZN(n9922) );
  AND2_X1 U12806 ( .A1(n11282), .A2(n10260), .ZN(n9923) );
  AND2_X1 U12807 ( .A1(n10263), .A2(n10261), .ZN(n9924) );
  OR2_X1 U12808 ( .A1(n9838), .A2(n13893), .ZN(n9925) );
  AND2_X1 U12809 ( .A1(n17820), .A2(n9814), .ZN(n9927) );
  INV_X1 U12810 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10179) );
  NOR2_X1 U12811 ( .A1(n18931), .A2(n18935), .ZN(n19079) );
  INV_X1 U12812 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10168) );
  AND2_X1 U12813 ( .A1(n10267), .A2(n12110), .ZN(n9928) );
  INV_X1 U12814 ( .A(n10998), .ZN(n10191) );
  AND2_X2 U12815 ( .A1(n13174), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13169) );
  AND2_X1 U12816 ( .A1(n11429), .A2(n11428), .ZN(n9929) );
  AND2_X1 U12817 ( .A1(n10165), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9930) );
  NAND2_X1 U12818 ( .A1(n10232), .A2(n10231), .ZN(n16252) );
  INV_X1 U12819 ( .A(n16252), .ZN(n13734) );
  AND2_X1 U12820 ( .A1(n14556), .A2(n14555), .ZN(n9931) );
  INV_X1 U12821 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10215) );
  AND2_X1 U12822 ( .A1(n10190), .A2(n14452), .ZN(n9932) );
  INV_X1 U12823 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10273) );
  NOR2_X1 U12824 ( .A1(n20699), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n9933) );
  AND2_X1 U12825 ( .A1(n18416), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n9934) );
  NAND2_X1 U12826 ( .A1(n17950), .A2(n9820), .ZN(n10271) );
  INV_X1 U12827 ( .A(n15746), .ZN(n10314) );
  AND2_X1 U12828 ( .A1(n10313), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9935) );
  NAND2_X1 U12829 ( .A1(n15132), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9936) );
  INV_X1 U12830 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n10080) );
  INV_X1 U12831 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n9973) );
  INV_X1 U12832 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n9971) );
  OR2_X1 U12833 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9937) );
  INV_X1 U12834 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10166) );
  INV_X1 U12835 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10200) );
  INV_X1 U12836 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10174) );
  NAND3_X2 U12837 ( .A1(n13960), .A2(n18931), .A3(n19060), .ZN(n18426) );
  OAI22_X2 U12838 ( .A1(n20259), .A2(n20292), .B1(n21124), .B2(n20291), .ZN(
        n20717) );
  INV_X1 U12839 ( .A(n20796), .ZN(n9938) );
  INV_X1 U12840 ( .A(n9938), .ZN(n9939) );
  INV_X1 U12841 ( .A(n20711), .ZN(n9940) );
  INV_X1 U12842 ( .A(n9940), .ZN(n9941) );
  INV_X1 U12843 ( .A(n20770), .ZN(n9942) );
  INV_X1 U12844 ( .A(n9942), .ZN(n9943) );
  INV_X1 U12845 ( .A(n20723), .ZN(n9944) );
  INV_X1 U12846 ( .A(n9944), .ZN(n9945) );
  INV_X1 U12847 ( .A(n20727), .ZN(n9946) );
  INV_X1 U12848 ( .A(n9946), .ZN(n9947) );
  NOR3_X2 U12849 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18933), .A3(
        n18621), .ZN(n18638) );
  OAI22_X2 U12850 ( .A1(n20293), .A2(n20292), .B1(n21002), .B2(n20291), .ZN(
        n20735) );
  INV_X1 U12851 ( .A(n15304), .ZN(n10300) );
  CLKBUF_X1 U12852 ( .A(n12824), .Z(n9948) );
  NOR3_X1 U12853 ( .A1(n12626), .A2(n13682), .A3(n19951), .ZN(n12824) );
  CLKBUF_X1 U12854 ( .A(n20734), .Z(n9949) );
  AND2_X1 U12855 ( .A1(n16318), .A2(n14462), .ZN(n12107) );
  NOR2_X2 U12856 ( .A1(n15492), .A2(n14484), .ZN(n15451) );
  NAND2_X1 U12857 ( .A1(n10259), .A2(n9879), .ZN(n10254) );
  OAI21_X1 U12858 ( .B1(n15611), .B2(n19436), .A(n10253), .ZN(P2_U3016) );
  NAND3_X2 U12859 ( .A1(n15476), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15449) );
  AOI21_X1 U12860 ( .B1(n16296), .B2(n19420), .A(n10254), .ZN(n10253) );
  NAND2_X1 U12861 ( .A1(n15610), .A2(n19429), .ZN(n10259) );
  INV_X1 U12862 ( .A(n10660), .ZN(n9950) );
  NAND2_X1 U12863 ( .A1(n9951), .A2(n9953), .ZN(n13696) );
  NAND2_X1 U12864 ( .A1(n9952), .A2(n9953), .ZN(n19500) );
  AND4_X2 U12865 ( .A1(n11121), .A2(n10558), .A3(n10548), .A4(n12096), .ZN(
        n9955) );
  NAND4_X1 U12866 ( .A1(n10479), .A2(n10477), .A3(n10478), .A4(n10476), .ZN(
        n9957) );
  NAND4_X1 U12867 ( .A1(n10473), .A2(n10475), .A3(n10474), .A4(n10472), .ZN(
        n9959) );
  NAND3_X1 U12868 ( .A1(n10130), .A2(n10129), .A3(n10841), .ZN(n13514) );
  NAND3_X1 U12869 ( .A1(n10187), .A2(n10184), .A3(n9799), .ZN(n9975) );
  XNOR2_X2 U12870 ( .A(n10635), .B(n10634), .ZN(n10641) );
  NAND2_X1 U12871 ( .A1(n11779), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12687) );
  INV_X1 U12872 ( .A(n12714), .ZN(n9984) );
  INV_X1 U12873 ( .A(n12713), .ZN(n9985) );
  NAND2_X1 U12874 ( .A1(n11897), .A2(n10395), .ZN(n9987) );
  NAND3_X1 U12875 ( .A1(n15283), .A2(n15361), .A3(n15346), .ZN(n9990) );
  NAND2_X2 U12876 ( .A1(n9992), .A2(n15288), .ZN(n12025) );
  NOR2_X2 U12877 ( .A1(n13654), .A2(n9902), .ZN(n10403) );
  INV_X1 U12878 ( .A(n10403), .ZN(n13745) );
  NAND2_X1 U12879 ( .A1(n9995), .A2(n10359), .ZN(n16103) );
  NAND2_X1 U12880 ( .A1(n16108), .A2(n9857), .ZN(n9995) );
  NAND2_X1 U12881 ( .A1(n13607), .A2(n13606), .ZN(n9996) );
  OR2_X4 U12882 ( .A1(n9997), .A2(n10000), .ZN(n10136) );
  NAND4_X1 U12883 ( .A1(n9998), .A2(n9999), .A3(n12253), .A4(n10008), .ZN(
        n9997) );
  NAND4_X1 U12884 ( .A1(n9878), .A2(n10003), .A3(n10002), .A4(n10001), .ZN(
        n10000) );
  NAND3_X1 U12885 ( .A1(n12237), .A2(n10016), .A3(n10015), .ZN(n10014) );
  NAND2_X1 U12886 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10016) );
  NAND2_X2 U12887 ( .A1(n10143), .A2(n10017), .ZN(n14948) );
  OR2_X2 U12888 ( .A1(n14912), .A2(n14920), .ZN(n10139) );
  XNOR2_X2 U12889 ( .A(n12490), .B(n12489), .ZN(n12646) );
  NAND2_X1 U12890 ( .A1(n12646), .A2(n20237), .ZN(n10027) );
  AND2_X2 U12891 ( .A1(n13239), .A2(n13238), .ZN(n13253) );
  OR3_X2 U12892 ( .A1(n14791), .A2(n10033), .A3(n10032), .ZN(n14728) );
  INV_X1 U12893 ( .A(n14728), .ZN(n14218) );
  INV_X1 U12894 ( .A(n14753), .ZN(n10036) );
  NOR2_X2 U12895 ( .A1(n13540), .A2(n13542), .ZN(n13588) );
  AND2_X2 U12896 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13174) );
  OR2_X2 U12897 ( .A1(n14717), .A2(n10367), .ZN(n14671) );
  NAND2_X1 U12898 ( .A1(n10644), .A2(n10042), .ZN(n10623) );
  NAND2_X1 U12899 ( .A1(n10638), .A2(n10042), .ZN(n10384) );
  OAI211_X2 U12900 ( .C1(n10613), .C2(n10042), .A(n10612), .B(n10041), .ZN(
        n10635) );
  NAND3_X1 U12901 ( .A1(n10042), .A2(n10624), .A3(n10611), .ZN(n10041) );
  XNOR2_X1 U12902 ( .A(n10644), .B(n10042), .ZN(n19425) );
  XNOR2_X2 U12903 ( .A(n11150), .B(n11155), .ZN(n12716) );
  NAND3_X1 U12904 ( .A1(n10684), .A2(n10739), .A3(n9837), .ZN(n11088) );
  NAND3_X1 U12905 ( .A1(n10077), .A2(n10075), .A3(n10074), .ZN(P1_U2809) );
  NAND4_X1 U12906 ( .A1(n14633), .A2(n21285), .A3(P1_REIP_REG_30__SCAN_IN), 
        .A4(P1_REIP_REG_29__SCAN_IN), .ZN(n10074) );
  INV_X4 U12907 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19050) );
  INV_X1 U12908 ( .A(n17416), .ZN(n11637) );
  NAND3_X1 U12909 ( .A1(n10094), .A2(P3_EAX_REG_22__SCAN_IN), .A3(
        P3_EAX_REG_17__SCAN_IN), .ZN(n10093) );
  INV_X1 U12910 ( .A(n10108), .ZN(n18003) );
  AND2_X4 U12911 ( .A1(n11055), .A2(n12923), .ZN(n12066) );
  OAI21_X1 U12912 ( .B1(n11000), .B2(n9884), .A(n10110), .ZN(n15448) );
  OAI211_X1 U12913 ( .C1(n16398), .C2(n10126), .A(n10346), .B(n10124), .ZN(
        n10128) );
  NAND2_X1 U12914 ( .A1(n10346), .A2(n10122), .ZN(n10121) );
  NAND2_X1 U12915 ( .A1(n16398), .A2(n16397), .ZN(n16396) );
  NAND2_X1 U12916 ( .A1(n14887), .A2(n10131), .ZN(P1_U2969) );
  INV_X1 U12917 ( .A(n12388), .ZN(n10134) );
  AND2_X2 U12918 ( .A1(n12993), .A2(n10136), .ZN(n12297) );
  NAND2_X1 U12919 ( .A1(n13364), .A2(n10136), .ZN(n12983) );
  NOR2_X1 U12920 ( .A1(n13364), .A2(n10136), .ZN(n10135) );
  NAND2_X1 U12921 ( .A1(n12387), .A2(n10136), .ZN(n12259) );
  NAND2_X1 U12922 ( .A1(n13114), .A2(n10136), .ZN(n12456) );
  NAND2_X1 U12923 ( .A1(n20286), .A2(n10136), .ZN(n20570) );
  AOI21_X2 U12924 ( .B1(n14933), .B2(n14899), .A(n16068), .ZN(n14920) );
  XNOR2_X2 U12925 ( .A(n13166), .B(n20390), .ZN(n10141) );
  NAND2_X1 U12926 ( .A1(n10141), .A2(n13167), .ZN(n13184) );
  AND2_X1 U12927 ( .A1(n13189), .A2(n10141), .ZN(n20596) );
  NOR2_X1 U12928 ( .A1(n20241), .A2(n10141), .ZN(n10140) );
  NAND2_X1 U12929 ( .A1(n20151), .A2(n10141), .ZN(n13422) );
  NAND3_X1 U12930 ( .A1(n13617), .A2(n13781), .A3(n13618), .ZN(n13624) );
  INV_X2 U12931 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19057) );
  NAND4_X1 U12932 ( .A1(n10154), .A2(n11531), .A3(n11533), .A4(n9875), .ZN(
        n11534) );
  NOR2_X1 U12933 ( .A1(n11576), .A2(n11578), .ZN(n10158) );
  NAND3_X1 U12934 ( .A1(n16302), .A2(n16303), .A3(n10161), .ZN(P2_U2825) );
  NAND2_X1 U12935 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10170) );
  NAND3_X1 U12936 ( .A1(n10171), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13466) );
  INV_X1 U12937 ( .A(n10828), .ZN(n10187) );
  NAND4_X1 U12938 ( .A1(n10338), .A2(n10333), .A3(n10189), .A4(n10188), .ZN(
        n14465) );
  AND2_X1 U12939 ( .A1(n14457), .A2(n10190), .ZN(n14453) );
  NAND2_X1 U12940 ( .A1(n14457), .A2(n9932), .ZN(n14458) );
  NOR2_X1 U12941 ( .A1(n10985), .A2(n10984), .ZN(n10987) );
  NOR2_X2 U12942 ( .A1(n11635), .A2(n10197), .ZN(n17632) );
  NAND3_X1 U12943 ( .A1(n10199), .A2(n10198), .A3(n10200), .ZN(n17763) );
  INV_X1 U12944 ( .A(n11734), .ZN(n17776) );
  NAND2_X2 U12945 ( .A1(n10201), .A2(n17795), .ZN(n11734) );
  OAI21_X1 U12946 ( .B1(n17447), .B2(n17278), .A(n10205), .ZN(n10204) );
  NAND2_X1 U12947 ( .A1(n10202), .A2(n11627), .ZN(n10207) );
  INV_X2 U12948 ( .A(n17258), .ZN(n11626) );
  AND2_X2 U12949 ( .A1(n10217), .A2(n17969), .ZN(n17848) );
  NAND3_X1 U12950 ( .A1(n17896), .A2(n10318), .A3(n10215), .ZN(n10217) );
  INV_X1 U12951 ( .A(n18148), .ZN(n17794) );
  NAND2_X1 U12952 ( .A1(n11738), .A2(n16644), .ZN(n17754) );
  NOR2_X4 U12953 ( .A1(n10225), .A2(n10226), .ZN(n14366) );
  NAND2_X1 U12954 ( .A1(n10227), .A2(n10229), .ZN(n13028) );
  OR2_X1 U12955 ( .A1(n9804), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n10228) );
  XNOR2_X2 U12956 ( .A(n14601), .B(n14600), .ZN(n15024) );
  INV_X1 U12957 ( .A(n16003), .ZN(n10240) );
  NAND2_X1 U12958 ( .A1(n13734), .A2(n9883), .ZN(n13939) );
  OR2_X2 U12959 ( .A1(n13840), .A2(n9925), .ZN(n15428) );
  NAND2_X1 U12960 ( .A1(n12398), .A2(n9826), .ZN(n13551) );
  NAND2_X2 U12961 ( .A1(n12397), .A2(n12396), .ZN(n12398) );
  NAND2_X1 U12962 ( .A1(n10262), .A2(n9924), .ZN(n16370) );
  INV_X1 U12963 ( .A(n10271), .ZN(n17889) );
  OAI21_X1 U12964 ( .B1(n16781), .B2(n9921), .A(n10274), .ZN(P3_U2640) );
  INV_X1 U12965 ( .A(n13138), .ZN(n10277) );
  NAND2_X1 U12966 ( .A1(n10277), .A2(n10278), .ZN(n13659) );
  NAND2_X1 U12967 ( .A1(n13658), .A2(n9908), .ZN(n13849) );
  INV_X1 U12968 ( .A(n12688), .ZN(n10291) );
  INV_X1 U12969 ( .A(n12696), .ZN(n10294) );
  XNOR2_X2 U12970 ( .A(n10305), .B(n10304), .ZN(n13154) );
  NAND2_X1 U12971 ( .A1(n10739), .A2(n10738), .ZN(n10304) );
  NAND2_X1 U12972 ( .A1(n10684), .A2(n10683), .ZN(n10305) );
  NAND2_X2 U12973 ( .A1(n11737), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16644) );
  AND2_X2 U12974 ( .A1(n17763), .A2(n11736), .ZN(n11737) );
  NAND4_X1 U12975 ( .A1(n10328), .A2(n9876), .A3(n11671), .A4(n11669), .ZN(
        n10322) );
  INV_X1 U12976 ( .A(n10335), .ZN(n10334) );
  INV_X1 U12977 ( .A(n12104), .ZN(n10340) );
  NOR2_X2 U12978 ( .A1(n10546), .A2(n10538), .ZN(n10556) );
  NAND2_X4 U12979 ( .A1(n10342), .A2(n10341), .ZN(n19451) );
  NAND2_X1 U12980 ( .A1(n10466), .A2(n12883), .ZN(n10341) );
  NAND2_X1 U12981 ( .A1(n10471), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10342) );
  NAND2_X1 U12982 ( .A1(n14892), .A2(n14071), .ZN(n10353) );
  NAND2_X1 U12983 ( .A1(n14882), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10355) );
  INV_X2 U12984 ( .A(n13868), .ZN(n14241) );
  NAND2_X2 U12985 ( .A1(n12198), .A2(n13192), .ZN(n13868) );
  NOR2_X4 U12986 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15173) );
  NAND2_X1 U12987 ( .A1(n12420), .A2(n10364), .ZN(n12497) );
  NAND3_X1 U12988 ( .A1(n12297), .A2(n12420), .A3(n10364), .ZN(n12388) );
  NAND2_X1 U12989 ( .A1(n12418), .A2(n12659), .ZN(n10364) );
  NAND2_X1 U12990 ( .A1(n12296), .A2(n13113), .ZN(n10365) );
  NOR2_X1 U12991 ( .A1(n14717), .A2(n14719), .ZN(n14706) );
  INV_X1 U12992 ( .A(n14719), .ZN(n10371) );
  NAND2_X1 U12993 ( .A1(n14659), .A2(n10374), .ZN(n14623) );
  NAND2_X1 U12994 ( .A1(n14659), .A2(n14660), .ZN(n14646) );
  AND2_X2 U12995 ( .A1(n14659), .A2(n9907), .ZN(n14610) );
  AND3_X2 U12996 ( .A1(n13588), .A2(n13589), .A3(n9900), .ZN(n13918) );
  NAND3_X1 U12997 ( .A1(n13588), .A2(n13589), .A3(n10380), .ZN(n13822) );
  NAND2_X1 U12998 ( .A1(n12025), .A2(n10392), .ZN(n15283) );
  NAND2_X1 U12999 ( .A1(n12025), .A2(n15290), .ZN(n15284) );
  INV_X1 U13000 ( .A(n10386), .ZN(n10385) );
  OAI22_X1 U13001 ( .A1(n10392), .A2(n10390), .B1(n12052), .B2(n10391), .ZN(
        n10386) );
  CLKBUF_X1 U13002 ( .A(n10403), .Z(n10400) );
  NOR2_X1 U13003 ( .A1(n12835), .A2(n12840), .ZN(n13134) );
  INV_X1 U13004 ( .A(n12840), .ZN(n10411) );
  NAND3_X1 U13005 ( .A1(n12076), .A2(n10577), .A3(n16562), .ZN(n10595) );
  OAI21_X1 U13006 ( .B1(n15489), .B2(n12105), .A(n12104), .ZN(n12103) );
  CLKBUF_X1 U13007 ( .A(n12716), .Z(n15253) );
  NAND2_X1 U13008 ( .A1(n12716), .A2(n12888), .ZN(n10652) );
  NAND2_X1 U13009 ( .A1(n12716), .A2(n15261), .ZN(n10660) );
  OR2_X2 U13010 ( .A1(n12716), .A2(n15261), .ZN(n10649) );
  INV_X1 U13011 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12644) );
  NAND2_X1 U13012 ( .A1(n14072), .A2(n10040), .ZN(n13921) );
  INV_X1 U13013 ( .A(n13074), .ZN(n13070) );
  NAND2_X1 U13014 ( .A1(n10610), .A2(n10609), .ZN(n10612) );
  INV_X1 U13015 ( .A(n11759), .ZN(n12597) );
  INV_X1 U13016 ( .A(n12973), .ZN(n12748) );
  XNOR2_X1 U13017 ( .A(n13617), .B(n13580), .ZN(n13773) );
  CLKBUF_X1 U13018 ( .A(n13918), .Z(n13879) );
  OAI21_X1 U13019 ( .B1(n10627), .B2(n10605), .A(n10604), .ZN(n10607) );
  OR2_X2 U13020 ( .A1(n17126), .A2(n11465), .ZN(n10412) );
  INV_X1 U13021 ( .A(n19411), .ZN(n14475) );
  OR2_X1 U13022 ( .A1(n15440), .A2(n19419), .ZN(n10413) );
  AND3_X1 U13023 ( .A1(n18268), .A2(n18294), .A3(n11730), .ZN(n10414) );
  OR2_X1 U13024 ( .A1(n11697), .A2(n18333), .ZN(n10415) );
  OR2_X1 U13025 ( .A1(n10354), .A2(n15035), .ZN(n10417) );
  AND2_X1 U13026 ( .A1(n11490), .A2(n11489), .ZN(n10418) );
  OR3_X1 U13027 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16638), .A3(
        n17770), .ZN(n10419) );
  NOR2_X1 U13028 ( .A1(n13068), .A2(n13067), .ZN(n10420) );
  AND2_X1 U13029 ( .A1(n15445), .A2(n14451), .ZN(n10421) );
  AND2_X1 U13030 ( .A1(n16291), .A2(n14475), .ZN(n10422) );
  NAND2_X1 U13031 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11781) );
  AND2_X1 U13032 ( .A1(n16249), .A2(n16248), .ZN(n10424) );
  AND4_X1 U13033 ( .A1(n12728), .A2(n12727), .A3(n12726), .A4(n12725), .ZN(
        n10425) );
  NAND2_X2 U13034 ( .A1(n14879), .A2(n13115), .ZN(n14881) );
  AND2_X1 U13035 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10426) );
  INV_X2 U13036 ( .A(n17489), .ZN(n17468) );
  OR3_X1 U13037 ( .A1(n17847), .A2(n17756), .A3(n16640), .ZN(n10427) );
  NOR2_X1 U13038 ( .A1(n11369), .A2(n11368), .ZN(n13383) );
  INV_X1 U13039 ( .A(n13383), .ZN(n11784) );
  AND3_X1 U13040 ( .A1(n12100), .A2(n12099), .A3(n12098), .ZN(n10428) );
  INV_X1 U13041 ( .A(n11254), .ZN(n11319) );
  OR2_X1 U13042 ( .A1(n11356), .A2(n11355), .ZN(n11783) );
  AND3_X1 U13043 ( .A1(n10490), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10489), .ZN(n10429) );
  INV_X1 U13044 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20064) );
  INV_X1 U13045 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20112) );
  INV_X1 U13046 ( .A(n14061), .ZN(n15001) );
  NOR2_X1 U13047 ( .A1(n15376), .A2(n15375), .ZN(n10431) );
  INV_X1 U13048 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n14497) );
  INV_X1 U13049 ( .A(n12255), .ZN(n12724) );
  INV_X1 U13050 ( .A(n12267), .ZN(n12300) );
  INV_X1 U13051 ( .A(n9847), .ZN(n17436) );
  OR2_X1 U13052 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14363) );
  NAND2_X2 U13053 ( .A1(n10460), .A2(n10459), .ZN(n11752) );
  AND3_X1 U13054 ( .A1(n10957), .A2(n14459), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n10432) );
  AND2_X1 U13055 ( .A1(n15485), .A2(n11005), .ZN(n12104) );
  AND3_X1 U13056 ( .A1(n10598), .A2(n10597), .A3(n10596), .ZN(n10433) );
  NAND2_X1 U13057 ( .A1(n10582), .A2(n10581), .ZN(n10620) );
  INV_X1 U13058 ( .A(n20285), .ZN(n12458) );
  OR2_X1 U13059 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n12471), .ZN(
        n12277) );
  OR3_X1 U13060 ( .A1(n12331), .A2(n12330), .A3(n12329), .ZN(n12332) );
  NOR2_X1 U13061 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12198) );
  NAND2_X1 U13062 ( .A1(n10576), .A2(n19445), .ZN(n10498) );
  AND2_X1 U13063 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20064), .ZN(
        n10808) );
  NAND2_X1 U13064 ( .A1(n13113), .A2(n13002), .ZN(n12258) );
  INV_X1 U13065 ( .A(n13431), .ZN(n13432) );
  OR2_X1 U13066 ( .A1(n13443), .A2(n13442), .ZN(n13619) );
  AOI22_X1 U13067 ( .A1(n12647), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12195) );
  OR2_X1 U13069 ( .A1(n10877), .A2(n10876), .ZN(n11298) );
  NAND2_X1 U13070 ( .A1(n10819), .A2(n10818), .ZN(n10825) );
  OAI22_X1 U13071 ( .A1(n10654), .A2(n19701), .B1(n19881), .B2(n10653), .ZN(
        n10655) );
  AOI21_X1 U13072 ( .B1(n11062), .B2(n10809), .A(n10808), .ZN(n10817) );
  INV_X1 U13073 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11730) );
  NAND2_X1 U13074 ( .A1(n14446), .A2(n12258), .ZN(n12298) );
  NOR2_X1 U13075 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12644), .ZN(
        n12192) );
  INV_X1 U13076 ( .A(n13573), .ZN(n13574) );
  OR2_X1 U13077 ( .A1(n16090), .A2(n14060), .ZN(n14057) );
  AOI21_X1 U13078 ( .B1(n12287), .B2(n12286), .A(n12280), .ZN(n12293) );
  AOI22_X1 U13079 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12230) );
  NAND2_X1 U13080 ( .A1(n12659), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12966) );
  OR3_X1 U13081 ( .A1(n11026), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n15986), .ZN(n11023) );
  OR2_X1 U13082 ( .A1(n11168), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10604) );
  OR2_X1 U13083 ( .A1(n10782), .A2(n10781), .ZN(n11293) );
  NAND2_X1 U13084 ( .A1(n10488), .A2(n12883), .ZN(n10494) );
  INV_X1 U13086 ( .A(n14730), .ZN(n14217) );
  OR2_X1 U13087 ( .A1(n14323), .A2(n14929), .ZN(n14341) );
  NAND2_X1 U13088 ( .A1(n14061), .A2(n9849), .ZN(n14063) );
  AND2_X1 U13089 ( .A1(n13532), .A2(n13531), .ZN(n13573) );
  INV_X1 U13090 ( .A(n14999), .ZN(n16046) );
  OR2_X1 U13091 ( .A1(n11026), .A2(n11025), .ZN(n11028) );
  AND2_X1 U13092 ( .A1(n16328), .A2(n14462), .ZN(n12105) );
  NOR2_X1 U13093 ( .A1(n19451), .A2(n19460), .ZN(n10570) );
  AOI22_X1 U13094 ( .A1(n14468), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10617) );
  OAI21_X1 U13095 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n19050), .A(
        n11580), .ZN(n11581) );
  NAND2_X1 U13096 ( .A1(n11566), .A2(n11601), .ZN(n11578) );
  AND2_X1 U13097 ( .A1(n12294), .A2(n12337), .ZN(n12416) );
  AND2_X1 U13098 ( .A1(n13352), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14436) );
  OR2_X1 U13099 ( .A1(n14341), .A2(n14340), .ZN(n14344) );
  NAND2_X1 U13100 ( .A1(n14180), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14196) );
  INV_X1 U13101 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13535) );
  AND2_X1 U13102 ( .A1(n12749), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14439) );
  AND2_X1 U13103 ( .A1(n12390), .A2(n14597), .ZN(n13172) );
  NOR2_X1 U13104 ( .A1(n12426), .A2(n12275), .ZN(n12415) );
  INV_X1 U13105 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12471) );
  AND3_X1 U13106 ( .A1(n11359), .A2(n11358), .A3(n11357), .ZN(n15223) );
  OR2_X1 U13107 ( .A1(n11452), .A2(n15458), .ZN(n11453) );
  INV_X1 U13108 ( .A(n15805), .ZN(n16439) );
  OR2_X1 U13109 ( .A1(n10714), .A2(n10713), .ZN(n11252) );
  OR2_X1 U13110 ( .A1(n12373), .A2(n20076), .ZN(n11031) );
  INV_X1 U13111 ( .A(n11600), .ZN(n11569) );
  INV_X1 U13112 ( .A(n11493), .ZN(n11494) );
  NOR2_X1 U13114 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11459) );
  NAND2_X1 U13115 ( .A1(n19096), .A2(n13965), .ZN(n18393) );
  NOR2_X1 U13116 ( .A1(n17969), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11732) );
  INV_X1 U13117 ( .A(n18034), .ZN(n18036) );
  INV_X1 U13118 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16024) );
  OR2_X1 U13119 ( .A1(n13358), .A2(n13357), .ZN(n20140) );
  AND2_X1 U13120 ( .A1(n13883), .A2(n13882), .ZN(n13888) );
  INV_X1 U13121 ( .A(n13911), .ZN(n14089) );
  AND2_X1 U13122 ( .A1(n13723), .A2(n13722), .ZN(n13726) );
  AND2_X1 U13123 ( .A1(n13001), .A2(n13111), .ZN(n13021) );
  OAI21_X1 U13124 ( .B1(n20906), .B2(n16276), .A(n20875), .ZN(n20236) );
  INV_X1 U13125 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20594) );
  INV_X1 U13126 ( .A(n20329), .ZN(n20234) );
  NAND2_X1 U13127 ( .A1(n16105), .A2(n20230), .ZN(n20292) );
  INV_X1 U13128 ( .A(n19286), .ZN(n19256) );
  OR2_X1 U13129 ( .A1(n12001), .A2(n11780), .ZN(n12693) );
  NAND2_X1 U13130 ( .A1(n12928), .A2(n12349), .ZN(n11761) );
  AND3_X1 U13131 ( .A1(n11413), .A2(n11412), .A3(n11411), .ZN(n15206) );
  INV_X1 U13132 ( .A(n12900), .ZN(n12075) );
  AND2_X1 U13133 ( .A1(n13832), .A2(n11140), .ZN(n15795) );
  AND2_X1 U13134 ( .A1(n11304), .A2(n11303), .ZN(n13053) );
  INV_X1 U13135 ( .A(n19420), .ZN(n16551) );
  INV_X1 U13136 ( .A(n10807), .ZN(n14462) );
  NAND2_X1 U13137 ( .A1(n15701), .A2(n12408), .ZN(n19427) );
  NAND2_X1 U13138 ( .A1(n11032), .A2(n11031), .ZN(n12901) );
  INV_X1 U13139 ( .A(n19666), .ZN(n19699) );
  INV_X1 U13140 ( .A(n11121), .ZN(n19445) );
  INV_X1 U13141 ( .A(n18393), .ZN(n18890) );
  NOR2_X1 U13142 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16972), .ZN(n16958) );
  NOR2_X1 U13143 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17044), .ZN(n17015) );
  NAND2_X1 U13144 ( .A1(n17080), .A2(n18441), .ZN(n12164) );
  NOR4_X1 U13145 ( .A1(n17291), .A2(n17462), .A3(n13967), .A4(n17290), .ZN(
        n17272) );
  INV_X1 U13146 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17233) );
  NOR3_X1 U13147 ( .A1(n15987), .A2(n18441), .A3(n18448), .ZN(n15988) );
  NOR2_X1 U13148 ( .A1(n18114), .A2(n17785), .ZN(n18116) );
  INV_X1 U13149 ( .A(n18374), .ZN(n18394) );
  INV_X1 U13150 ( .A(n17925), .ZN(n18277) );
  INV_X1 U13151 ( .A(n18296), .ZN(n18276) );
  INV_X1 U13152 ( .A(n11677), .ZN(n11675) );
  NAND2_X1 U13153 ( .A1(n13595), .A2(n14540), .ZN(n20133) );
  INV_X1 U13154 ( .A(n20185), .ZN(n14801) );
  AND2_X1 U13155 ( .A1(n20185), .A2(n20294), .ZN(n20181) );
  AND2_X1 U13156 ( .A1(n14258), .A2(n14257), .ZN(n14707) );
  AND2_X1 U13157 ( .A1(n14448), .A2(n20229), .ZN(n14864) );
  NAND2_X1 U13158 ( .A1(n13112), .A2(n13111), .ZN(n14873) );
  INV_X1 U13159 ( .A(n12624), .ZN(n12619) );
  NAND2_X1 U13160 ( .A1(n13912), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13911) );
  AND2_X1 U13161 ( .A1(n13875), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13912) );
  AND2_X1 U13162 ( .A1(n13581), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13720) );
  OR2_X1 U13163 ( .A1(n16058), .A2(n16057), .ZN(n16175) );
  INV_X1 U13164 ( .A(n13038), .ZN(n16202) );
  NOR2_X1 U13165 ( .A1(n15025), .A2(n16266), .ZN(n16211) );
  INV_X1 U13166 ( .A(n16130), .ZN(n16205) );
  INV_X1 U13167 ( .A(n15958), .ZN(n20875) );
  NOR2_X1 U13168 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15169) );
  AND2_X1 U13169 ( .A1(n20232), .A2(n20883), .ZN(n20360) );
  OAI211_X1 U13170 ( .C1(n20335), .C2(n20334), .A(n20559), .B(n20333), .ZN(
        n20352) );
  AND2_X1 U13171 ( .A1(n20360), .A2(n20548), .ZN(n20384) );
  NOR2_X2 U13172 ( .A1(n20363), .A2(n20601), .ZN(n20414) );
  OR2_X1 U13173 ( .A1(n9811), .A2(n20234), .ZN(n20627) );
  NOR2_X2 U13174 ( .A1(n20473), .A2(n20697), .ZN(n20492) );
  NAND2_X1 U13175 ( .A1(n13069), .A2(n20389), .ZN(n20473) );
  INV_X1 U13176 ( .A(n20627), .ZN(n20496) );
  NOR2_X2 U13177 ( .A1(n20602), .A2(n20669), .ZN(n20588) );
  AND2_X1 U13178 ( .A1(n9811), .A2(n20329), .ZN(n20548) );
  OR2_X1 U13179 ( .A1(n9811), .A2(n20329), .ZN(n20669) );
  NOR2_X1 U13180 ( .A1(n20396), .A2(n20244), .ZN(n20743) );
  NOR2_X1 U13181 ( .A1(n20396), .A2(n20269), .ZN(n20768) );
  NOR2_X1 U13182 ( .A1(n20396), .A2(n20287), .ZN(n20784) );
  OR4_X1 U13183 ( .A1(n15948), .A2(n15947), .A3(n15946), .A4(n15945), .ZN(
        n15955) );
  INV_X1 U13184 ( .A(n19290), .ZN(n19203) );
  AND2_X1 U13185 ( .A1(n19104), .A2(n13482), .ZN(n19286) );
  INV_X1 U13186 ( .A(n19295), .ZN(n19243) );
  INV_X1 U13187 ( .A(n15556), .ZN(n19136) );
  OR2_X1 U13188 ( .A1(n11409), .A2(n11408), .ZN(n13601) );
  INV_X1 U13189 ( .A(n11783), .ZN(n13384) );
  INV_X1 U13190 ( .A(n12831), .ZN(n12842) );
  INV_X1 U13191 ( .A(n16570), .ZN(n14501) );
  INV_X1 U13192 ( .A(n20069), .ZN(n19364) );
  INV_X1 U13193 ( .A(n12829), .ZN(n16287) );
  CLKBUF_X1 U13194 ( .A(n12804), .Z(n12826) );
  AND2_X1 U13195 ( .A1(n16498), .A2(n12367), .ZN(n16488) );
  INV_X1 U13196 ( .A(n16480), .ZN(n16494) );
  INV_X1 U13197 ( .A(n15686), .ZN(n15731) );
  INV_X1 U13198 ( .A(n19419), .ZN(n19429) );
  NOR2_X2 U13199 ( .A1(n19666), .A2(n19557), .ZN(n19496) );
  OR2_X1 U13200 ( .A1(n19509), .A2(n19888), .ZN(n19527) );
  INV_X1 U13201 ( .A(n19541), .ZN(n19547) );
  OAI21_X1 U13202 ( .B1(n19577), .B2(n13298), .A(n19561), .ZN(n19579) );
  INV_X1 U13203 ( .A(n19601), .ZN(n19616) );
  INV_X1 U13204 ( .A(n19892), .ZN(n20041) );
  OR2_X1 U13205 ( .A1(n20051), .A2(n20060), .ZN(n19666) );
  AND2_X1 U13206 ( .A1(n19760), .A2(n19699), .ZN(n19751) );
  INV_X1 U13207 ( .A(n19832), .ZN(n19800) );
  INV_X1 U13208 ( .A(n20034), .ZN(n19771) );
  AND2_X1 U13209 ( .A1(n13124), .A2(n13123), .ZN(n13129) );
  INV_X1 U13210 ( .A(n19935), .ZN(n19875) );
  AOI21_X1 U13211 ( .B1(n11596), .B2(n11598), .A(n11595), .ZN(n18871) );
  INV_X1 U13212 ( .A(n17110), .ZN(n17139) );
  OR2_X1 U13213 ( .A1(n16849), .A2(P3_EBX_REG_23__SCAN_IN), .ZN(n16850) );
  NOR2_X1 U13214 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16943), .ZN(n16928) );
  NOR2_X1 U13215 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16999), .ZN(n16983) );
  NOR2_X2 U13216 ( .A1(n19034), .A2(n17073), .ZN(n17092) );
  NOR3_X1 U13217 ( .A1(n17288), .A2(n17488), .A3(n17472), .ZN(n17467) );
  AOI22_X1 U13218 ( .A1(n13965), .A2(n18868), .B1(n13964), .B2(n13963), .ZN(
        n15987) );
  NOR3_X1 U13219 ( .A1(n18478), .A2(n17689), .A3(n17568), .ZN(n17557) );
  AND2_X1 U13220 ( .A1(n18308), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n16639) );
  INV_X1 U13221 ( .A(n18344), .ZN(n18325) );
  NOR2_X1 U13222 ( .A1(n18211), .A2(n18347), .ZN(n18265) );
  INV_X1 U13223 ( .A(n18426), .ZN(n18416) );
  INV_X1 U13224 ( .A(n18739), .ZN(n18488) );
  NOR2_X1 U13225 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19034), .ZN(
        n19058) );
  AND2_X1 U13226 ( .A1(n19026), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18963) );
  NAND2_X1 U13227 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n13727), .ZN(n20131) );
  INV_X1 U13228 ( .A(n20165), .ZN(n13570) );
  OAI21_X1 U13229 ( .B1(n14505), .B2(n14506), .A(n14795), .ZN(n16082) );
  INV_X1 U13230 ( .A(n20189), .ZN(n20212) );
  NOR2_X1 U13231 ( .A1(n12583), .A2(n12507), .ZN(n12623) );
  NAND2_X1 U13232 ( .A1(n16116), .A2(n12852), .ZN(n16110) );
  INV_X1 U13233 ( .A(n16268), .ZN(n16215) );
  INV_X1 U13234 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13205) );
  NAND2_X1 U13235 ( .A1(n20360), .A2(n20496), .ZN(n20327) );
  AOI22_X1 U13236 ( .A1(n20331), .A2(n20334), .B1(n9933), .B2(n20552), .ZN(
        n20355) );
  AOI22_X1 U13237 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20364), .B1(n20367), 
        .B2(n20362), .ZN(n20388) );
  OR2_X1 U13238 ( .A1(n20473), .A2(n20627), .ZN(n20441) );
  AOI22_X1 U13239 ( .A1(n20447), .A2(n20444), .B1(n20630), .B2(n9933), .ZN(
        n20468) );
  OR2_X1 U13240 ( .A1(n20473), .A2(n20601), .ZN(n20499) );
  NAND2_X1 U13241 ( .A1(n20886), .A2(n20496), .ZN(n20547) );
  AOI22_X1 U13242 ( .A1(n20557), .A2(n20555), .B1(n20552), .B2(n20551), .ZN(
        n20593) );
  NAND2_X1 U13243 ( .A1(n20886), .A2(n20548), .ZN(n20624) );
  AOI22_X1 U13244 ( .A1(n20635), .A2(n20632), .B1(n20630), .B2(n20629), .ZN(
        n20668) );
  OR2_X1 U13245 ( .A1(n20698), .A2(n20669), .ZN(n20710) );
  OR2_X1 U13246 ( .A1(n20698), .A2(n20601), .ZN(n20790) );
  INV_X1 U13247 ( .A(n20863), .ZN(n20805) );
  AND2_X1 U13248 ( .A1(n20809), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20912) );
  OR2_X1 U13249 ( .A1(n12175), .A2(n12172), .ZN(n12626) );
  NAND2_X1 U13250 ( .A1(n16287), .A2(n13474), .ZN(n19290) );
  INV_X1 U13251 ( .A(n19326), .ZN(n20039) );
  INV_X1 U13252 ( .A(n12130), .ZN(n12131) );
  INV_X1 U13253 ( .A(n19361), .ZN(n15425) );
  AOI21_X2 U13254 ( .B1(n12860), .B2(n12078), .A(n14501), .ZN(n19333) );
  AND2_X1 U13255 ( .A1(n15404), .A2(n13054), .ZN(n19367) );
  NAND2_X1 U13256 ( .A1(n19369), .A2(n10553), .ZN(n12570) );
  INV_X1 U13257 ( .A(n19369), .ZN(n19402) );
  INV_X1 U13258 ( .A(n12801), .ZN(n12829) );
  INV_X1 U13259 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19197) );
  INV_X1 U13260 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16465) );
  OR2_X1 U13261 ( .A1(n12357), .A2(n12907), .ZN(n16480) );
  NAND2_X1 U13262 ( .A1(n11450), .A2(n20079), .ZN(n19419) );
  INV_X1 U13263 ( .A(n10641), .ZN(n15261) );
  INV_X1 U13264 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20048) );
  INV_X1 U13265 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15882) );
  AOI21_X1 U13266 ( .B1(n13673), .B2(n13672), .A(n13671), .ZN(n19471) );
  INV_X1 U13267 ( .A(n19522), .ZN(n19530) );
  OR2_X1 U13268 ( .A1(n19557), .A2(n20034), .ZN(n19541) );
  OR2_X1 U13269 ( .A1(n19597), .A2(n20034), .ZN(n19582) );
  INV_X1 U13270 ( .A(n19612), .ZN(n19619) );
  OR2_X1 U13271 ( .A1(n19597), .A2(n19596), .ZN(n19641) );
  INV_X1 U13272 ( .A(n19658), .ZN(n19665) );
  OR2_X1 U13273 ( .A1(n19597), .A2(n20041), .ZN(n19697) );
  OR2_X1 U13274 ( .A1(n19733), .A2(n19666), .ZN(n19723) );
  INV_X1 U13275 ( .A(n19751), .ZN(n19759) );
  INV_X1 U13276 ( .A(n19783), .ZN(n19793) );
  INV_X1 U13277 ( .A(n19913), .ZN(n19820) );
  INV_X1 U13278 ( .A(n19929), .ZN(n19833) );
  AOI211_X2 U13279 ( .C1(n13702), .C2(n13701), .A(n19888), .B(n13700), .ZN(
        n19880) );
  INV_X1 U13280 ( .A(n19867), .ZN(n19920) );
  INV_X1 U13281 ( .A(n19019), .ZN(n19093) );
  INV_X1 U13282 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17974) );
  INV_X1 U13283 ( .A(n17136), .ZN(n17140) );
  NOR2_X1 U13284 ( .A1(n16836), .A2(n17196), .ZN(n17200) );
  NOR2_X1 U13285 ( .A1(n17206), .A2(n17146), .ZN(n17211) );
  AND2_X1 U13286 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17359), .ZN(n17376) );
  INV_X1 U13287 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17476) );
  NOR2_X1 U13288 ( .A1(n10430), .A2(n17494), .ZN(n17609) );
  OR2_X1 U13289 ( .A1(n17579), .A2(n17602), .ZN(n17597) );
  NOR3_X1 U13290 ( .A1(n18478), .A2(n17640), .A3(n17573), .ZN(n17616) );
  INV_X1 U13291 ( .A(n17639), .ZN(n17636) );
  INV_X1 U13292 ( .A(n17663), .ZN(n17682) );
  INV_X1 U13293 ( .A(n17952), .ZN(n17938) );
  INV_X1 U13294 ( .A(n17997), .ZN(n18015) );
  OAI21_X1 U13295 ( .B1(n18265), .B2(n18212), .A(n18409), .ZN(n18329) );
  INV_X1 U13296 ( .A(n18423), .ZN(n18420) );
  INV_X1 U13297 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18903) );
  INV_X1 U13298 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18914) );
  INV_X1 U13299 ( .A(n19079), .ZN(n18929) );
  INV_X1 U13300 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19034) );
  INV_X1 U13301 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19066) );
  INV_X1 U13302 ( .A(n19093), .ZN(n19026) );
  NOR2_X1 U13303 ( .A1(n18944), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19019) );
  INV_X1 U13304 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10639) );
  NOR2_X4 U13305 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12889) );
  AND2_X4 U13306 ( .A1(n12889), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10670) );
  AND2_X4 U13307 ( .A1(n12889), .A2(n12923), .ZN(n10530) );
  AOI22_X1 U13308 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10440) );
  AND2_X4 U13309 ( .A1(n11055), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10671) );
  AOI22_X1 U13310 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10439) );
  AND2_X4 U13311 ( .A1(n10435), .A2(n12923), .ZN(n11867) );
  AND2_X4 U13312 ( .A1(n10435), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10529) );
  AOI22_X1 U13313 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10438) );
  AND2_X4 U13314 ( .A1(n12872), .A2(n12873), .ZN(n11868) );
  AND2_X4 U13315 ( .A1(n10436), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10669) );
  AOI22_X1 U13316 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10437) );
  NAND4_X1 U13317 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10441) );
  NAND2_X1 U13318 ( .A1(n10441), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10448) );
  AOI22_X1 U13319 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13320 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10444) );
  AOI22_X1 U13321 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U13322 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10442) );
  NAND4_X1 U13323 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n10446) );
  NAND2_X1 U13324 ( .A1(n10446), .A2(n12883), .ZN(n10447) );
  AOI22_X1 U13325 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13326 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13327 ( .A1(n10529), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11868), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U13328 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10449) );
  NAND4_X1 U13329 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10453) );
  NAND2_X1 U13330 ( .A1(n10453), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10460) );
  AOI22_X1 U13331 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U13332 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13333 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U13334 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10454) );
  NAND4_X1 U13335 ( .A1(n10457), .A2(n10456), .A3(n10455), .A4(n10454), .ZN(
        n10458) );
  NAND2_X1 U13336 ( .A1(n10458), .A2(n12883), .ZN(n10459) );
  INV_X1 U13337 ( .A(n11752), .ZN(n10461) );
  AOI22_X1 U13338 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13339 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13340 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13341 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13342 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13343 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U13344 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10467) );
  INV_X1 U13345 ( .A(n19451), .ZN(n10480) );
  AOI22_X1 U13346 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10475) );
  AOI22_X1 U13347 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11868), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10474) );
  AOI22_X1 U13348 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10529), .B1(
        n11867), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13349 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13350 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10479) );
  AOI22_X1 U13351 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10478) );
  AOI22_X1 U13352 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10477) );
  AOI21_X1 U13353 ( .B1(n10567), .B2(n10480), .A(n19460), .ZN(n10483) );
  INV_X1 U13354 ( .A(n11752), .ZN(n10560) );
  NAND2_X1 U13355 ( .A1(n10548), .A2(n10560), .ZN(n10566) );
  NAND2_X1 U13356 ( .A1(n10566), .A2(n10539), .ZN(n11044) );
  INV_X1 U13357 ( .A(n11044), .ZN(n10481) );
  NAND2_X1 U13358 ( .A1(n10481), .A2(n19451), .ZN(n10482) );
  NAND2_X1 U13359 ( .A1(n10483), .A2(n10482), .ZN(n11118) );
  AOI22_X1 U13360 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10487) );
  AOI22_X1 U13361 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13362 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13363 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13364 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13365 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13366 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12063), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13367 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10491) );
  NAND3_X1 U13368 ( .A1(n10429), .A2(n10492), .A3(n10491), .ZN(n10493) );
  NAND2_X1 U13369 ( .A1(n11118), .A2(n11121), .ZN(n10499) );
  AOI22_X1 U13370 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13371 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13372 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10501) );
  AOI22_X1 U13373 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10500) );
  NAND4_X1 U13374 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10504) );
  AOI22_X1 U13375 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13376 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U13377 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13378 ( .A1(n10529), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11868), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10505) );
  NAND4_X1 U13379 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10509) );
  AOI22_X1 U13380 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U13381 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10514) );
  AOI22_X1 U13382 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10513) );
  AOI22_X1 U13383 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10512) );
  NAND4_X1 U13384 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10516) );
  AOI22_X1 U13385 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10520) );
  AOI22_X1 U13386 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13387 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10518) );
  AOI22_X1 U13388 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10517) );
  NAND4_X1 U13389 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .ZN(
        n10521) );
  NAND2_X1 U13390 ( .A1(n10521), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10522) );
  AOI22_X1 U13391 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10527) );
  AOI22_X1 U13392 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13393 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13394 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10524) );
  NAND4_X1 U13395 ( .A1(n10527), .A2(n10526), .A3(n10525), .A4(n10524), .ZN(
        n10528) );
  NAND2_X1 U13396 ( .A1(n10528), .A2(n12883), .ZN(n10537) );
  AOI22_X1 U13397 ( .A1(n11867), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13398 ( .A1(n10670), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10530), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13399 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10671), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13400 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10669), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10531) );
  NAND4_X1 U13401 ( .A1(n10534), .A2(n10533), .A3(n10532), .A4(n10531), .ZN(
        n10535) );
  NAND2_X1 U13402 ( .A1(n10535), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10536) );
  NAND2_X1 U13403 ( .A1(n10557), .A2(n11048), .ZN(n10538) );
  INV_X1 U13404 ( .A(n10556), .ZN(n10544) );
  NAND2_X1 U13405 ( .A1(n10567), .A2(n11121), .ZN(n10541) );
  NOR2_X1 U13406 ( .A1(n19460), .A2(n10550), .ZN(n10540) );
  NAND3_X1 U13407 ( .A1(n10542), .A2(n10541), .A3(n10540), .ZN(n10543) );
  NAND3_X1 U13408 ( .A1(n10544), .A2(n13118), .A3(n10543), .ZN(n11124) );
  NAND2_X1 U13409 ( .A1(n12907), .A2(n12079), .ZN(n10587) );
  NAND2_X1 U13410 ( .A1(n10587), .A2(n13118), .ZN(n10545) );
  NAND2_X1 U13411 ( .A1(n11124), .A2(n10545), .ZN(n10589) );
  AOI21_X2 U13412 ( .B1(n10588), .B2(n11014), .A(n10589), .ZN(n10555) );
  INV_X1 U13413 ( .A(n10546), .ZN(n10547) );
  NAND3_X1 U13414 ( .A1(n12910), .A2(n19439), .A3(n11253), .ZN(n10552) );
  INV_X1 U13415 ( .A(n11049), .ZN(n10551) );
  NAND2_X1 U13416 ( .A1(n10552), .A2(n10551), .ZN(n11446) );
  INV_X1 U13417 ( .A(n11446), .ZN(n10554) );
  INV_X1 U13418 ( .A(n12373), .ZN(n10553) );
  OAI21_X2 U13419 ( .B1(n10555), .B2(n11751), .A(n10598), .ZN(n10627) );
  NAND2_X1 U13420 ( .A1(n10627), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10565) );
  NAND2_X1 U13421 ( .A1(n12909), .A2(n12172), .ZN(n11447) );
  INV_X1 U13422 ( .A(n10569), .ZN(n10559) );
  INV_X1 U13423 ( .A(n11258), .ZN(n12083) );
  NOR2_X1 U13424 ( .A1(n12083), .A2(n10560), .ZN(n10561) );
  NAND2_X1 U13425 ( .A1(n12077), .A2(n10561), .ZN(n10573) );
  INV_X1 U13426 ( .A(n10573), .ZN(n10562) );
  OR2_X2 U13427 ( .A1(n11447), .A2(n10562), .ZN(n12925) );
  AOI21_X2 U13428 ( .B1(n12925), .B2(n16562), .A(n10563), .ZN(n10564) );
  NAND2_X2 U13429 ( .A1(n10565), .A2(n10564), .ZN(n10621) );
  INV_X1 U13430 ( .A(n10621), .ZN(n10584) );
  NOR2_X1 U13431 ( .A1(n10566), .A2(n11253), .ZN(n10568) );
  INV_X1 U13432 ( .A(n10567), .ZN(n11255) );
  MUX2_X1 U13433 ( .A(n10568), .B(n11255), .S(n11121), .Z(n10571) );
  AND3_X2 U13434 ( .A1(n10571), .A2(n10570), .A3(n11116), .ZN(n12916) );
  INV_X1 U13435 ( .A(n11129), .ZN(n10602) );
  NAND2_X1 U13436 ( .A1(n12907), .A2(n12181), .ZN(n11060) );
  INV_X1 U13437 ( .A(n11060), .ZN(n10572) );
  NAND2_X1 U13438 ( .A1(n11049), .A2(n10572), .ZN(n12943) );
  INV_X1 U13439 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19422) );
  AND2_X1 U13440 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16562), .ZN(
        n10575) );
  NAND2_X1 U13441 ( .A1(n10614), .A2(n10575), .ZN(n10582) );
  NOR2_X1 U13442 ( .A1(n10602), .A2(n13477), .ZN(n10577) );
  INV_X1 U13443 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n15278) );
  NAND2_X1 U13444 ( .A1(n10616), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10579) );
  NAND2_X1 U13445 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10578) );
  OAI211_X1 U13446 ( .C1(n10595), .C2(n15278), .A(n10579), .B(n10578), .ZN(
        n10580) );
  INV_X1 U13447 ( .A(n10580), .ZN(n10581) );
  INV_X1 U13448 ( .A(n10620), .ZN(n10583) );
  NAND2_X1 U13449 ( .A1(n10627), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10586) );
  AOI21_X1 U13450 ( .B1(n11751), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10585) );
  INV_X1 U13451 ( .A(n10624), .ZN(n10608) );
  NAND2_X1 U13452 ( .A1(n10622), .A2(n10608), .ZN(n10613) );
  NAND2_X1 U13453 ( .A1(n10630), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10600) );
  NAND2_X1 U13454 ( .A1(n10588), .A2(n10587), .ZN(n11117) );
  AOI21_X1 U13455 ( .B1(n11117), .B2(n10590), .A(n11751), .ZN(n10591) );
  INV_X1 U13456 ( .A(n10591), .ZN(n10599) );
  INV_X1 U13457 ( .A(n12184), .ZN(n10593) );
  NAND2_X1 U13458 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U13459 ( .A1(n10593), .A2(n10592), .ZN(n10594) );
  AOI21_X1 U13460 ( .B1(n10616), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10594), .ZN(
        n10597) );
  INV_X1 U13461 ( .A(n10601), .ZN(n10603) );
  NOR2_X1 U13462 ( .A1(n10603), .A2(n10602), .ZN(n10605) );
  NAND2_X1 U13463 ( .A1(n10607), .A2(n10606), .ZN(n10637) );
  NAND2_X1 U13464 ( .A1(n10622), .A2(n10624), .ZN(n10610) );
  NAND2_X1 U13465 ( .A1(n10621), .A2(n10620), .ZN(n10611) );
  NAND2_X1 U13466 ( .A1(n10611), .A2(n10608), .ZN(n10609) );
  INV_X1 U13467 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10619) );
  NAND2_X1 U13468 ( .A1(n10614), .A2(n16562), .ZN(n10615) );
  INV_X1 U13469 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12410) );
  XNOR2_X2 U13470 ( .A(n10621), .B(n10583), .ZN(n10644) );
  NAND2_X1 U13471 ( .A1(n10623), .A2(n10622), .ZN(n10625) );
  NAND2_X1 U13472 ( .A1(n10625), .A2(n10624), .ZN(n10626) );
  OAI21_X2 U13473 ( .B1(n10635), .B2(n10634), .A(n10626), .ZN(n11150) );
  NAND2_X1 U13474 ( .A1(n10627), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10629) );
  NAND2_X1 U13475 ( .A1(n12184), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10628) );
  INV_X1 U13476 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10814) );
  NAND2_X1 U13477 ( .A1(n14468), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10632) );
  NAND2_X1 U13478 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10631) );
  OAI211_X1 U13479 ( .C1(n11206), .C2(n10814), .A(n10632), .B(n10631), .ZN(
        n10633) );
  OR2_X1 U13480 ( .A1(n10637), .A2(n10636), .ZN(n10638) );
  NAND2_X1 U13481 ( .A1(n12928), .A2(n10644), .ZN(n10657) );
  NOR2_X2 U13482 ( .A1(n10649), .A2(n10657), .ZN(n13094) );
  INV_X1 U13483 ( .A(n13094), .ZN(n10857) );
  OR2_X2 U13484 ( .A1(n10660), .A2(n10657), .ZN(n19763) );
  INV_X1 U13485 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11966) );
  OAI22_X1 U13486 ( .A1(n10639), .A2(n10857), .B1(n19763), .B2(n11966), .ZN(
        n10643) );
  INV_X1 U13487 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11956) );
  INV_X1 U13488 ( .A(n10644), .ZN(n10640) );
  NAND2_X1 U13489 ( .A1(n12928), .A2(n10640), .ZN(n10651) );
  INV_X1 U13490 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11965) );
  OAI22_X1 U13491 ( .A1(n11956), .A2(n19592), .B1(n13124), .B2(n11965), .ZN(
        n10642) );
  NOR2_X1 U13492 ( .A1(n10643), .A2(n10642), .ZN(n10667) );
  INV_X1 U13493 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11964) );
  INV_X1 U13494 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10645) );
  OAI22_X1 U13495 ( .A1(n11964), .A2(n19795), .B1(n13696), .B2(n10645), .ZN(
        n10648) );
  INV_X1 U13496 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10646) );
  INV_X1 U13497 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11967) );
  OAI22_X1 U13498 ( .A1(n10646), .A2(n19622), .B1(n19736), .B2(n11967), .ZN(
        n10647) );
  NOR2_X1 U13499 ( .A1(n10648), .A2(n10647), .ZN(n10666) );
  INV_X1 U13500 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11955) );
  OR2_X2 U13501 ( .A1(n10649), .A2(n10659), .ZN(n19554) );
  OR2_X2 U13502 ( .A1(n12716), .A2(n12888), .ZN(n10658) );
  INV_X1 U13503 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10650) );
  OAI22_X1 U13504 ( .A1(n11955), .A2(n19554), .B1(n19472), .B2(n10650), .ZN(
        n10656) );
  INV_X1 U13505 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10654) );
  OR2_X2 U13506 ( .A1(n10660), .A2(n10651), .ZN(n19701) );
  OR2_X2 U13507 ( .A1(n10652), .A2(n10657), .ZN(n19881) );
  INV_X1 U13508 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10653) );
  NOR2_X1 U13509 ( .A1(n10656), .A2(n10655), .ZN(n10665) );
  INV_X1 U13510 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11958) );
  OR2_X2 U13511 ( .A1(n10658), .A2(n10657), .ZN(n10762) );
  INV_X1 U13512 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11957) );
  OAI22_X1 U13513 ( .A1(n11958), .A2(n19500), .B1(n10762), .B2(n11957), .ZN(
        n10663) );
  INV_X1 U13514 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10661) );
  INV_X1 U13515 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11819) );
  OAI22_X1 U13516 ( .A1(n10661), .A2(n13669), .B1(n19668), .B2(n11819), .ZN(
        n10662) );
  NOR2_X1 U13517 ( .A1(n10663), .A2(n10662), .ZN(n10664) );
  NAND4_X1 U13518 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10684) );
  BUF_X1 U13519 ( .A(n11867), .Z(n10668) );
  AND2_X2 U13520 ( .A1(n9801), .A2(n12883), .ZN(n11305) );
  AND2_X2 U13521 ( .A1(n9801), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11883) );
  AOI22_X1 U13522 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11305), .B1(
        n11883), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10675) );
  AND2_X2 U13523 ( .A1(n12059), .A2(n12883), .ZN(n11884) );
  AND2_X2 U13524 ( .A1(n12059), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11816) );
  AOI22_X1 U13525 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11884), .B1(
        n11816), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10674) );
  BUF_X1 U13526 ( .A(n11868), .Z(n10676) );
  AND2_X2 U13527 ( .A1(n10676), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11889) );
  AOI22_X1 U13528 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10673) );
  AND2_X2 U13529 ( .A1(n12065), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12869) );
  AND2_X1 U13530 ( .A1(n12066), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10730) );
  AOI22_X1 U13531 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12869), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10672) );
  NAND4_X1 U13532 ( .A1(n10675), .A2(n10674), .A3(n10673), .A4(n10672), .ZN(
        n10682) );
  AND2_X2 U13533 ( .A1(n12064), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10729) );
  AOI22_X1 U13534 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10729), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10680) );
  NOR4_X2 U13535 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U13536 ( .A1(n11818), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n11882), .ZN(n10679) );
  AOI22_X1 U13537 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10776), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10678) );
  AND2_X2 U13538 ( .A1(n12058), .A2(n12883), .ZN(n11832) );
  AND2_X2 U13539 ( .A1(n10676), .A2(n12883), .ZN(n10704) );
  AOI22_X1 U13540 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10677) );
  NAND4_X1 U13541 ( .A1(n10680), .A2(n10679), .A3(n10678), .A4(n10677), .ZN(
        n10681) );
  NOR2_X1 U13542 ( .A1(n10682), .A2(n10681), .ZN(n11285) );
  NAND2_X1 U13543 ( .A1(n11285), .A2(n13682), .ZN(n10683) );
  INV_X1 U13544 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11901) );
  NAND2_X1 U13545 ( .A1(n13094), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10685) );
  OAI211_X1 U13546 ( .C1(n11901), .C2(n19500), .A(n10685), .B(n11259), .ZN(
        n10689) );
  INV_X1 U13547 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10687) );
  INV_X1 U13548 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10686) );
  NOR2_X1 U13549 ( .A1(n10689), .A2(n10688), .ZN(n10703) );
  INV_X1 U13550 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10691) );
  INV_X1 U13551 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10690) );
  OAI22_X1 U13552 ( .A1(n10691), .A2(n19472), .B1(n19622), .B2(n10690), .ZN(
        n10693) );
  INV_X1 U13553 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11898) );
  INV_X1 U13554 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11909) );
  OAI22_X1 U13555 ( .A1(n11898), .A2(n19554), .B1(n19763), .B2(n11909), .ZN(
        n10692) );
  NOR2_X1 U13556 ( .A1(n10693), .A2(n10692), .ZN(n10702) );
  INV_X1 U13557 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11899) );
  INV_X1 U13558 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11762) );
  OAI22_X1 U13559 ( .A1(n11899), .A2(n19592), .B1(n13669), .B2(n11762), .ZN(
        n10695) );
  INV_X1 U13560 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11900) );
  INV_X1 U13561 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11910) );
  OAI22_X1 U13562 ( .A1(n11900), .A2(n10762), .B1(n19736), .B2(n11910), .ZN(
        n10694) );
  NOR2_X1 U13563 ( .A1(n10695), .A2(n10694), .ZN(n10701) );
  INV_X1 U13564 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11908) );
  INV_X1 U13565 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10696) );
  INV_X1 U13566 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11907) );
  INV_X1 U13567 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10697) );
  OAI22_X1 U13568 ( .A1(n11907), .A2(n19795), .B1(n19701), .B2(n10697), .ZN(
        n10698) );
  NOR2_X1 U13569 ( .A1(n10699), .A2(n10698), .ZN(n10700) );
  AOI22_X1 U13570 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U13571 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11882), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13572 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11884), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13573 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10705) );
  NAND4_X1 U13574 ( .A1(n10708), .A2(n10707), .A3(n10706), .A4(n10705), .ZN(
        n10714) );
  AOI22_X1 U13575 ( .A1(n10729), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13576 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13577 ( .A1(n10798), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13578 ( .A1(n12869), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10709) );
  NAND4_X1 U13579 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10709), .ZN(
        n10713) );
  AND2_X1 U13580 ( .A1(n13682), .A2(n11252), .ZN(n12363) );
  AOI22_X1 U13581 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11832), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10718) );
  AOI22_X1 U13582 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n11882), .ZN(n10717) );
  AOI22_X1 U13583 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n11884), .ZN(n10716) );
  AOI22_X1 U13584 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10715) );
  NAND4_X1 U13585 ( .A1(n10718), .A2(n10717), .A3(n10716), .A4(n10715), .ZN(
        n10724) );
  AOI22_X1 U13586 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10775), .B1(
        n10729), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U13587 ( .A1(n10774), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13588 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10776), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U13589 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12869), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10719) );
  NAND4_X1 U13590 ( .A1(n10722), .A2(n10721), .A3(n10720), .A4(n10719), .ZN(
        n10723) );
  AND2_X1 U13591 ( .A1(n12363), .A2(n11077), .ZN(n11081) );
  INV_X1 U13592 ( .A(n11081), .ZN(n10737) );
  AOI22_X1 U13593 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n11882), .ZN(n10728) );
  AOI22_X1 U13594 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n11884), .ZN(n10727) );
  AOI22_X1 U13595 ( .A1(n11818), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n11816), .ZN(n10726) );
  AOI22_X1 U13596 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10725) );
  NAND4_X1 U13597 ( .A1(n10728), .A2(n10727), .A3(n10726), .A4(n10725), .ZN(
        n10736) );
  AOI22_X1 U13598 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10729), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13599 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U13600 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12869), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13601 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10776), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10731) );
  NAND4_X1 U13602 ( .A1(n10734), .A2(n10733), .A3(n10732), .A4(n10731), .ZN(
        n10735) );
  INV_X1 U13603 ( .A(n11273), .ZN(n11082) );
  NAND2_X1 U13604 ( .A1(n10737), .A2(n11082), .ZN(n10738) );
  INV_X1 U13605 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U13606 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11832), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13607 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n11882), .ZN(n10742) );
  AOI22_X1 U13608 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n11884), .ZN(n10741) );
  AOI22_X1 U13609 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10740) );
  NAND4_X1 U13610 ( .A1(n10743), .A2(n10742), .A3(n10741), .A4(n10740), .ZN(
        n10749) );
  AOI22_X1 U13611 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10729), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13612 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13613 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10798), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13614 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12869), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10744) );
  NAND4_X1 U13615 ( .A1(n10747), .A2(n10746), .A3(n10745), .A4(n10744), .ZN(
        n10748) );
  INV_X1 U13616 ( .A(n11290), .ZN(n11087) );
  INV_X1 U13617 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10750) );
  INV_X1 U13618 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12016) );
  OAI22_X1 U13619 ( .A1(n10750), .A2(n19472), .B1(n19763), .B2(n12016), .ZN(
        n10753) );
  INV_X1 U13620 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12006) );
  INV_X1 U13621 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10751) );
  OAI22_X1 U13622 ( .A1(n12006), .A2(n19554), .B1(n19701), .B2(n10751), .ZN(
        n10752) );
  NOR2_X1 U13623 ( .A1(n10753), .A2(n10752), .ZN(n10769) );
  INV_X1 U13624 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10755) );
  INV_X1 U13625 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10754) );
  OAI22_X1 U13626 ( .A1(n10755), .A2(n19881), .B1(n13696), .B2(n10754), .ZN(
        n10757) );
  INV_X1 U13627 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12014) );
  INV_X1 U13628 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12017) );
  OAI22_X1 U13629 ( .A1(n12014), .A2(n19795), .B1(n19736), .B2(n12017), .ZN(
        n10756) );
  NOR2_X1 U13630 ( .A1(n10757), .A2(n10756), .ZN(n10768) );
  INV_X1 U13631 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10759) );
  INV_X1 U13632 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10758) );
  OAI22_X1 U13633 ( .A1(n10759), .A2(n10857), .B1(n19622), .B2(n10758), .ZN(
        n10761) );
  INV_X1 U13634 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12007) );
  INV_X1 U13635 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12015) );
  OAI22_X1 U13636 ( .A1(n12007), .A2(n19592), .B1(n13124), .B2(n12015), .ZN(
        n10760) );
  NOR2_X1 U13637 ( .A1(n10761), .A2(n10760), .ZN(n10767) );
  INV_X1 U13638 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12008) );
  INV_X1 U13639 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13316) );
  OAI22_X1 U13640 ( .A1(n12008), .A2(n19500), .B1(n10762), .B2(n13316), .ZN(
        n10765) );
  INV_X1 U13641 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14529) );
  INV_X1 U13642 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10763) );
  OAI22_X1 U13643 ( .A1(n14529), .A2(n13669), .B1(n19668), .B2(n10763), .ZN(
        n10764) );
  NOR2_X1 U13644 ( .A1(n10765), .A2(n10764), .ZN(n10766) );
  AOI22_X1 U13645 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13646 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11882), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13647 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11884), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10771) );
  AOI22_X1 U13648 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10770) );
  NAND4_X1 U13649 ( .A1(n10773), .A2(n10772), .A3(n10771), .A4(n10770), .ZN(
        n10782) );
  AOI22_X1 U13650 ( .A1(n10729), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U13651 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10779) );
  AOI22_X1 U13652 ( .A1(n10798), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U13653 ( .A1(n12869), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10777) );
  NAND4_X1 U13654 ( .A1(n10780), .A2(n10779), .A3(n10778), .A4(n10777), .ZN(
        n10781) );
  INV_X1 U13655 ( .A(n11293), .ZN(n10783) );
  AOI22_X1 U13656 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n11882), .ZN(n10789) );
  INV_X1 U13657 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n19879) );
  NAND2_X1 U13658 ( .A1(n11818), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10788) );
  NAND2_X1 U13659 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10787) );
  AND3_X1 U13660 ( .A1(n10789), .A2(n10788), .A3(n10787), .ZN(n10806) );
  NAND2_X1 U13661 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10793) );
  NAND2_X1 U13662 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10792) );
  NAND2_X1 U13663 ( .A1(n11884), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10791) );
  NAND2_X1 U13664 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10790) );
  NAND2_X1 U13665 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10797) );
  NAND2_X1 U13666 ( .A1(n10774), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10796) );
  NAND2_X1 U13667 ( .A1(n10729), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10795) );
  NAND2_X1 U13668 ( .A1(n11889), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10794) );
  NAND2_X1 U13669 ( .A1(n10798), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10802) );
  NAND2_X1 U13670 ( .A1(n10730), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10801) );
  NAND2_X1 U13671 ( .A1(n10776), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10800) );
  NAND2_X1 U13672 ( .A1(n12869), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10799) );
  NAND4_X1 U13673 ( .A1(n10806), .A2(n10805), .A3(n10804), .A4(n10803), .ZN(
        n11302) );
  INV_X1 U13674 ( .A(n11302), .ZN(n10807) );
  MUX2_X1 U13675 ( .A(n20064), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11062) );
  INV_X1 U13676 ( .A(n11011), .ZN(n10809) );
  NAND2_X1 U13677 ( .A1(n12873), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10818) );
  NAND2_X1 U13678 ( .A1(n20056), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10816) );
  NAND2_X1 U13679 ( .A1(n10818), .A2(n10816), .ZN(n10810) );
  XNOR2_X1 U13680 ( .A(n10817), .B(n10810), .ZN(n11035) );
  INV_X1 U13681 ( .A(n11035), .ZN(n10811) );
  MUX2_X1 U13682 ( .A(n11273), .B(n10811), .S(n13477), .Z(n11061) );
  MUX2_X1 U13683 ( .A(n11061), .B(n10619), .S(n14459), .Z(n10839) );
  INV_X1 U13684 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U13685 ( .A1(n10812), .A2(n15278), .ZN(n10813) );
  NAND2_X1 U13686 ( .A1(n11077), .A2(n11251), .ZN(n11270) );
  OAI21_X1 U13687 ( .B1(n11251), .B2(n10813), .A(n11270), .ZN(n10838) );
  NAND2_X1 U13688 ( .A1(n10839), .A2(n10838), .ZN(n10829) );
  NAND2_X1 U13689 ( .A1(n11014), .A2(n11285), .ZN(n10815) );
  MUX2_X1 U13690 ( .A(n10815), .B(n10814), .S(n10990), .Z(n10822) );
  NAND2_X1 U13691 ( .A1(n13477), .A2(n11251), .ZN(n10831) );
  NAND2_X1 U13692 ( .A1(n10817), .A2(n10816), .ZN(n10819) );
  MUX2_X1 U13693 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n20048), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10824) );
  INV_X1 U13694 ( .A(n10824), .ZN(n10820) );
  XNOR2_X1 U13695 ( .A(n10825), .B(n10820), .ZN(n11022) );
  OR2_X1 U13696 ( .A1(n10831), .A2(n11022), .ZN(n10821) );
  NAND2_X1 U13697 ( .A1(n10822), .A2(n10821), .ZN(n10828) );
  NOR2_X1 U13698 ( .A1(n13477), .A2(n11290), .ZN(n10823) );
  INV_X1 U13699 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n11163) );
  MUX2_X1 U13700 ( .A(n11163), .B(n11293), .S(n11251), .Z(n10826) );
  OAI21_X1 U13701 ( .B1(n10827), .B2(n10826), .A(n10891), .ZN(n13554) );
  INV_X1 U13702 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13642) );
  XNOR2_X1 U13703 ( .A(n10829), .B(n10828), .ZN(n15249) );
  NAND2_X1 U13704 ( .A1(n11014), .A2(n11252), .ZN(n10830) );
  MUX2_X1 U13705 ( .A(n10830), .B(n10812), .S(n14459), .Z(n10833) );
  OAI21_X1 U13706 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20074), .A(
        n11011), .ZN(n11016) );
  OR2_X1 U13707 ( .A1(n10831), .A2(n11016), .ZN(n10832) );
  NAND2_X1 U13708 ( .A1(n10833), .A2(n10832), .ZN(n19287) );
  INV_X1 U13709 ( .A(n19287), .ZN(n10834) );
  INV_X1 U13710 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12364) );
  NOR2_X1 U13711 ( .A1(n10834), .A2(n12364), .ZN(n12573) );
  NAND2_X1 U13712 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10835) );
  NOR2_X1 U13713 ( .A1(n11251), .A2(n10835), .ZN(n10836) );
  OR2_X1 U13714 ( .A1(n10838), .A2(n10836), .ZN(n15274) );
  INV_X1 U13715 ( .A(n15274), .ZN(n12572) );
  NAND2_X1 U13716 ( .A1(n12573), .A2(n12572), .ZN(n12571) );
  NOR2_X1 U13717 ( .A1(n12573), .A2(n12572), .ZN(n10837) );
  AOI21_X1 U13718 ( .B1(n19422), .B2(n12571), .A(n10837), .ZN(n12347) );
  XNOR2_X1 U13719 ( .A(n10839), .B(n10838), .ZN(n15257) );
  XNOR2_X1 U13720 ( .A(n15257), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12346) );
  NOR2_X1 U13721 ( .A1(n15257), .A2(n12410), .ZN(n10840) );
  AOI21_X1 U13722 ( .B1(n12347), .B2(n12346), .A(n10840), .ZN(n13150) );
  XNOR2_X1 U13723 ( .A(n9896), .B(n9799), .ZN(n19265) );
  INV_X1 U13724 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19407) );
  XNOR2_X1 U13725 ( .A(n19265), .B(n19407), .ZN(n13511) );
  INV_X1 U13726 ( .A(n19265), .ZN(n10843) );
  NAND2_X1 U13727 ( .A1(n10843), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10844) );
  NAND2_X1 U13728 ( .A1(n13514), .A2(n10844), .ZN(n13639) );
  NAND2_X1 U13729 ( .A1(n13640), .A2(n13639), .ZN(n13638) );
  NAND2_X1 U13730 ( .A1(n10845), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10846) );
  INV_X1 U13731 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12038) );
  INV_X1 U13732 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12040) );
  OAI22_X1 U13733 ( .A1(n12038), .A2(n13124), .B1(n19763), .B2(n12040), .ZN(
        n10850) );
  INV_X1 U13734 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10848) );
  INV_X1 U13735 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10847) );
  OAI22_X1 U13736 ( .A1(n10848), .A2(n19472), .B1(n19701), .B2(n10847), .ZN(
        n10849) );
  NOR2_X1 U13737 ( .A1(n10850), .A2(n10849), .ZN(n10867) );
  INV_X1 U13738 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12036) );
  INV_X1 U13739 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10851) );
  OAI22_X1 U13740 ( .A1(n12036), .A2(n19795), .B1(n13696), .B2(n10851), .ZN(
        n10855) );
  INV_X1 U13741 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10853) );
  INV_X1 U13742 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10852) );
  OAI22_X1 U13743 ( .A1(n10853), .A2(n19622), .B1(n19668), .B2(n10852), .ZN(
        n10854) );
  NOR2_X1 U13744 ( .A1(n10855), .A2(n10854), .ZN(n10866) );
  INV_X1 U13745 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13104) );
  INV_X1 U13746 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10856) );
  OAI22_X1 U13747 ( .A1(n13104), .A2(n10857), .B1(n19592), .B2(n10856), .ZN(
        n10860) );
  INV_X1 U13748 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12028) );
  INV_X1 U13749 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10858) );
  OAI22_X1 U13750 ( .A1(n12028), .A2(n19554), .B1(n19881), .B2(n10858), .ZN(
        n10859) );
  NOR2_X1 U13751 ( .A1(n10860), .A2(n10859), .ZN(n10865) );
  INV_X1 U13752 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12029) );
  INV_X1 U13753 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12030) );
  OAI22_X1 U13754 ( .A1(n12029), .A2(n10762), .B1(n19500), .B2(n12030), .ZN(
        n10863) );
  INV_X1 U13755 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10861) );
  INV_X1 U13756 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12041) );
  OAI22_X1 U13757 ( .A1(n10861), .A2(n13669), .B1(n19736), .B2(n12041), .ZN(
        n10862) );
  NOR2_X1 U13758 ( .A1(n10863), .A2(n10862), .ZN(n10864) );
  NAND4_X1 U13759 ( .A1(n10867), .A2(n10866), .A3(n10865), .A4(n10864), .ZN(
        n10880) );
  AOI22_X1 U13760 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11832), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13761 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n11882), .ZN(n10870) );
  AOI22_X1 U13762 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11884), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13763 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10868) );
  NAND4_X1 U13764 ( .A1(n10871), .A2(n10870), .A3(n10869), .A4(n10868), .ZN(
        n10877) );
  AOI22_X1 U13765 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10729), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U13766 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10874) );
  AOI22_X1 U13767 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10798), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U13768 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10776), .B1(
        n12869), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10872) );
  NAND4_X1 U13769 ( .A1(n10875), .A2(n10874), .A3(n10873), .A4(n10872), .ZN(
        n10876) );
  INV_X1 U13770 ( .A(n11298), .ZN(n10878) );
  NAND2_X1 U13771 ( .A1(n10878), .A2(n13682), .ZN(n10879) );
  NAND2_X1 U13772 ( .A1(n11098), .A2(n10807), .ZN(n10881) );
  INV_X1 U13773 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n14535) );
  MUX2_X1 U13774 ( .A(n14535), .B(n11298), .S(n11251), .Z(n10889) );
  INV_X1 U13775 ( .A(n10889), .ZN(n10884) );
  XNOR2_X1 U13776 ( .A(n10891), .B(n10884), .ZN(n13493) );
  NAND2_X1 U13777 ( .A1(n10881), .A2(n13493), .ZN(n10882) );
  INV_X1 U13778 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11112) );
  XNOR2_X1 U13779 ( .A(n10882), .B(n11112), .ZN(n13827) );
  NAND2_X1 U13780 ( .A1(n10882), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10883) );
  NOR2_X1 U13781 ( .A1(n10891), .A2(n10884), .ZN(n10887) );
  INV_X1 U13782 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10885) );
  MUX2_X1 U13783 ( .A(n10885), .B(n11302), .S(n11251), .Z(n10888) );
  INV_X1 U13784 ( .A(n10888), .ZN(n10886) );
  XNOR2_X1 U13785 ( .A(n10887), .B(n10886), .ZN(n19253) );
  AND2_X1 U13786 ( .A1(n19253), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15819) );
  NAND2_X1 U13787 ( .A1(n10889), .A2(n10888), .ZN(n10890) );
  NAND2_X1 U13788 ( .A1(n14459), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10893) );
  INV_X1 U13789 ( .A(n10893), .ZN(n10892) );
  XNOR2_X1 U13790 ( .A(n10895), .B(n10892), .ZN(n19236) );
  NAND2_X1 U13791 ( .A1(n19236), .A2(n14462), .ZN(n15787) );
  INV_X1 U13792 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15595) );
  NAND2_X1 U13793 ( .A1(n10990), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10894) );
  INV_X1 U13794 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10898) );
  MUX2_X1 U13795 ( .A(n10894), .B(P2_EBX_REG_10__SCAN_IN), .S(n10902), .Z(
        n10896) );
  NAND2_X1 U13796 ( .A1(n10896), .A2(n10995), .ZN(n19225) );
  OR2_X1 U13797 ( .A1(n19225), .A2(n10807), .ZN(n10897) );
  INV_X1 U13798 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15797) );
  NAND2_X1 U13799 ( .A1(n10897), .A2(n15797), .ZN(n16438) );
  NOR2_X1 U13800 ( .A1(n11251), .A2(n10898), .ZN(n10899) );
  XNOR2_X1 U13801 ( .A(n10900), .B(n10899), .ZN(n15236) );
  NAND2_X1 U13802 ( .A1(n15236), .A2(n14462), .ZN(n10901) );
  INV_X1 U13803 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15814) );
  NAND2_X1 U13804 ( .A1(n10901), .A2(n15814), .ZN(n15790) );
  NAND2_X1 U13805 ( .A1(n15787), .A2(n15595), .ZN(n10909) );
  INV_X1 U13806 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13146) );
  INV_X1 U13807 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13142) );
  NAND2_X1 U13808 ( .A1(n13146), .A2(n10903), .ZN(n10919) );
  INV_X1 U13809 ( .A(n10903), .ZN(n10904) );
  NAND2_X1 U13810 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n10904), .ZN(n10905) );
  NOR2_X1 U13811 ( .A1(n11251), .A2(n10905), .ZN(n10906) );
  OR2_X1 U13812 ( .A1(n10918), .A2(n10906), .ZN(n15233) );
  OR2_X1 U13813 ( .A1(n15233), .A2(n10807), .ZN(n10912) );
  INV_X1 U13814 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10907) );
  NAND2_X1 U13815 ( .A1(n10912), .A2(n10907), .ZN(n16434) );
  INV_X1 U13816 ( .A(n19253), .ZN(n10908) );
  INV_X1 U13817 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15826) );
  NAND2_X1 U13818 ( .A1(n10908), .A2(n15826), .ZN(n15818) );
  AND4_X1 U13819 ( .A1(n15790), .A2(n10909), .A3(n16434), .A4(n15818), .ZN(
        n10910) );
  AND2_X1 U13820 ( .A1(n16438), .A2(n10910), .ZN(n10911) );
  INV_X1 U13821 ( .A(n10912), .ZN(n10913) );
  NAND2_X1 U13822 ( .A1(n10913), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16435) );
  AND2_X1 U13823 ( .A1(n14462), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10914) );
  NAND2_X1 U13824 ( .A1(n14462), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10915) );
  NOR2_X1 U13825 ( .A1(n19225), .A2(n10915), .ZN(n16437) );
  NOR2_X1 U13826 ( .A1(n16436), .A2(n16437), .ZN(n10916) );
  AND2_X1 U13827 ( .A1(n16435), .A2(n10916), .ZN(n15524) );
  NAND2_X1 U13828 ( .A1(n14459), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10917) );
  NAND3_X1 U13829 ( .A1(n14459), .A2(n10919), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n10920) );
  NAND2_X1 U13830 ( .A1(n10954), .A2(n10920), .ZN(n19213) );
  INV_X1 U13831 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15774) );
  OR3_X1 U13832 ( .A1(n19213), .A2(n10807), .A3(n15774), .ZN(n15775) );
  OR2_X1 U13833 ( .A1(n19213), .A2(n10807), .ZN(n10921) );
  NAND2_X1 U13834 ( .A1(n10921), .A2(n15774), .ZN(n15776) );
  INV_X1 U13835 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11194) );
  NOR2_X1 U13836 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n10922) );
  NOR2_X1 U13837 ( .A1(n11251), .A2(n10922), .ZN(n10923) );
  NOR2_X1 U13838 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n10924) );
  NOR2_X1 U13839 ( .A1(n11251), .A2(n10924), .ZN(n10925) );
  INV_X1 U13840 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11207) );
  NOR2_X1 U13841 ( .A1(n10940), .A2(n11207), .ZN(n10926) );
  MUX2_X1 U13842 ( .A(n10940), .B(n10926), .S(n14459), .Z(n10927) );
  INV_X1 U13843 ( .A(n10927), .ZN(n10928) );
  NAND2_X1 U13844 ( .A1(n10940), .A2(n11207), .ZN(n10930) );
  NAND2_X1 U13845 ( .A1(n10928), .A2(n10930), .ZN(n19152) );
  OR2_X1 U13846 ( .A1(n19152), .A2(n10807), .ZN(n10929) );
  NAND2_X1 U13847 ( .A1(n10929), .A2(n15689), .ZN(n15567) );
  NAND3_X1 U13848 ( .A1(n10930), .A2(n14459), .A3(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n10932) );
  OAI21_X1 U13849 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(P2_EBX_REG_18__SCAN_IN), 
        .A(n14459), .ZN(n10931) );
  NAND2_X1 U13850 ( .A1(n10932), .A2(n10956), .ZN(n19144) );
  OR2_X1 U13851 ( .A1(n19144), .A2(n10807), .ZN(n10963) );
  INV_X1 U13852 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15680) );
  NAND2_X1 U13853 ( .A1(n10963), .A2(n15680), .ZN(n15559) );
  NAND2_X1 U13854 ( .A1(n15567), .A2(n15559), .ZN(n15543) );
  NAND2_X1 U13855 ( .A1(n14459), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10933) );
  XNOR2_X1 U13856 ( .A(n10956), .B(n10933), .ZN(n19132) );
  NAND2_X1 U13857 ( .A1(n19132), .A2(n14462), .ZN(n10970) );
  INV_X1 U13858 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15669) );
  AND2_X1 U13859 ( .A1(n10970), .A2(n15669), .ZN(n15546) );
  NOR2_X1 U13860 ( .A1(n15543), .A2(n15546), .ZN(n15532) );
  INV_X1 U13861 ( .A(n10952), .ZN(n10934) );
  INV_X1 U13862 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10935) );
  NAND2_X1 U13863 ( .A1(n10934), .A2(n10935), .ZN(n10941) );
  NOR2_X1 U13864 ( .A1(n11251), .A2(n10935), .ZN(n10937) );
  INV_X1 U13865 ( .A(n10995), .ZN(n10936) );
  AOI21_X1 U13866 ( .B1(n10952), .B2(n10937), .A(n10936), .ZN(n10938) );
  NAND2_X1 U13867 ( .A1(n10941), .A2(n10938), .ZN(n19177) );
  OR2_X1 U13868 ( .A1(n19177), .A2(n10807), .ZN(n10939) );
  XNOR2_X1 U13869 ( .A(n10939), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15589) );
  INV_X1 U13870 ( .A(n10940), .ZN(n10943) );
  NAND3_X1 U13871 ( .A1(n10941), .A2(n10990), .A3(P2_EBX_REG_17__SCAN_IN), 
        .ZN(n10942) );
  NAND2_X1 U13872 ( .A1(n10943), .A2(n10942), .ZN(n19167) );
  OR2_X1 U13873 ( .A1(n19167), .A2(n10807), .ZN(n10944) );
  INV_X1 U13874 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11108) );
  NAND2_X1 U13875 ( .A1(n10944), .A2(n11108), .ZN(n15579) );
  NAND2_X1 U13876 ( .A1(n10946), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10945) );
  MUX2_X1 U13877 ( .A(n10946), .B(n10945), .S(n14459), .Z(n10947) );
  OR2_X1 U13878 ( .A1(n10946), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10951) );
  NAND2_X1 U13879 ( .A1(n19187), .A2(n14462), .ZN(n10948) );
  INV_X1 U13880 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15750) );
  NAND2_X1 U13881 ( .A1(n10948), .A2(n15750), .ZN(n15743) );
  INV_X1 U13882 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10949) );
  NOR2_X1 U13883 ( .A1(n11251), .A2(n10949), .ZN(n10950) );
  NAND2_X1 U13884 ( .A1(n10951), .A2(n10950), .ZN(n10953) );
  NAND2_X1 U13885 ( .A1(n10953), .A2(n10952), .ZN(n10968) );
  INV_X1 U13886 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15725) );
  OAI21_X1 U13887 ( .B1(n10968), .B2(n10807), .A(n15725), .ZN(n15735) );
  XNOR2_X1 U13888 ( .A(n10954), .B(n9916), .ZN(n19200) );
  NAND2_X1 U13889 ( .A1(n19200), .A2(n14462), .ZN(n10955) );
  INV_X1 U13890 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15764) );
  NAND2_X1 U13891 ( .A1(n10955), .A2(n15764), .ZN(n15768) );
  AND4_X1 U13892 ( .A1(n15579), .A2(n15743), .A3(n15735), .A4(n15768), .ZN(
        n10959) );
  NOR2_X1 U13893 ( .A1(n10973), .A2(n10432), .ZN(n15194) );
  NAND2_X1 U13894 ( .A1(n15194), .A2(n14462), .ZN(n10958) );
  INV_X1 U13895 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15655) );
  NAND2_X1 U13896 ( .A1(n10958), .A2(n15655), .ZN(n15535) );
  NAND4_X1 U13897 ( .A1(n15532), .A2(n15589), .A3(n10959), .A4(n15535), .ZN(
        n10960) );
  AND2_X1 U13898 ( .A1(n14462), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10961) );
  NAND2_X1 U13899 ( .A1(n15194), .A2(n10961), .ZN(n15534) );
  NAND2_X1 U13900 ( .A1(n14462), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10962) );
  OR2_X1 U13901 ( .A1(n19152), .A2(n10962), .ZN(n15566) );
  OR2_X1 U13902 ( .A1(n10963), .A2(n15680), .ZN(n15560) );
  AND2_X1 U13903 ( .A1(n15566), .A2(n15560), .ZN(n15531) );
  NAND2_X1 U13904 ( .A1(n14462), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10964) );
  OR2_X1 U13905 ( .A1(n19167), .A2(n10964), .ZN(n15578) );
  NAND2_X1 U13906 ( .A1(n14462), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10965) );
  OR2_X1 U13907 ( .A1(n19177), .A2(n10965), .ZN(n15575) );
  NAND2_X1 U13908 ( .A1(n15578), .A2(n15575), .ZN(n15530) );
  AND2_X1 U13909 ( .A1(n14462), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10966) );
  AND2_X1 U13910 ( .A1(n19200), .A2(n10966), .ZN(n15523) );
  AND2_X1 U13911 ( .A1(n14462), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10967) );
  NAND2_X1 U13912 ( .A1(n19187), .A2(n10967), .ZN(n15742) );
  INV_X1 U13913 ( .A(n10968), .ZN(n15217) );
  AND2_X1 U13914 ( .A1(n14462), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10969) );
  NAND2_X1 U13915 ( .A1(n15217), .A2(n10969), .ZN(n15734) );
  NAND2_X1 U13916 ( .A1(n15742), .A2(n15734), .ZN(n15528) );
  NOR3_X1 U13917 ( .A1(n15530), .A2(n15523), .A3(n15528), .ZN(n10971) );
  OR2_X1 U13918 ( .A1(n10970), .A2(n15669), .ZN(n15545) );
  AND4_X1 U13919 ( .A1(n15534), .A2(n15531), .A3(n10971), .A4(n15545), .ZN(
        n10972) );
  NAND2_X1 U13920 ( .A1(n14459), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10974) );
  INV_X1 U13921 ( .A(n10974), .ZN(n10975) );
  NAND2_X1 U13922 ( .A1(n10976), .A2(n10975), .ZN(n10977) );
  AND2_X1 U13923 ( .A1(n10985), .A2(n10977), .ZN(n15921) );
  NAND2_X1 U13924 ( .A1(n15921), .A2(n14462), .ZN(n10978) );
  INV_X1 U13925 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15639) );
  NAND2_X1 U13926 ( .A1(n10978), .A2(n15639), .ZN(n15510) );
  INV_X1 U13927 ( .A(n10978), .ZN(n10979) );
  NAND2_X1 U13928 ( .A1(n10979), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15511) );
  INV_X1 U13929 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10980) );
  NOR2_X1 U13930 ( .A1(n11251), .A2(n10980), .ZN(n10984) );
  XNOR2_X1 U13931 ( .A(n10985), .B(n10194), .ZN(n16369) );
  NAND2_X1 U13932 ( .A1(n16369), .A2(n14462), .ZN(n10981) );
  XNOR2_X1 U13933 ( .A(n10981), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16397) );
  INV_X1 U13934 ( .A(n10981), .ZN(n10982) );
  NAND2_X1 U13935 ( .A1(n10982), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10983) );
  INV_X1 U13936 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16357) );
  NAND2_X1 U13937 ( .A1(n14459), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10986) );
  OAI21_X1 U13938 ( .B1(n10987), .B2(n10986), .A(n10995), .ZN(n10988) );
  AND2_X1 U13939 ( .A1(n10989), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15499) );
  INV_X1 U13940 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15626) );
  NAND2_X1 U13941 ( .A1(n10990), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10991) );
  MUX2_X1 U13942 ( .A(n10991), .B(P2_EBX_REG_25__SCAN_IN), .S(n10994), .Z(
        n10992) );
  AND2_X1 U13943 ( .A1(n10992), .A2(n10995), .ZN(n16347) );
  AOI21_X1 U13944 ( .B1(n16347), .B2(n14462), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16390) );
  INV_X1 U13945 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10993) );
  NAND2_X1 U13946 ( .A1(n10995), .A2(n9851), .ZN(n14457) );
  NAND2_X1 U13947 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n9860), .ZN(n10996) );
  NOR2_X1 U13948 ( .A1(n11251), .A2(n10996), .ZN(n10997) );
  NOR2_X1 U13949 ( .A1(n14457), .A2(n10997), .ZN(n16338) );
  NAND2_X1 U13950 ( .A1(n16338), .A2(n14462), .ZN(n11003) );
  XNOR2_X1 U13951 ( .A(n11003), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15487) );
  NAND2_X1 U13952 ( .A1(n14459), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10998) );
  NAND2_X1 U13953 ( .A1(n10191), .A2(n9851), .ZN(n10999) );
  AND2_X1 U13954 ( .A1(n11008), .A2(n10999), .ZN(n16328) );
  NAND2_X1 U13955 ( .A1(n14459), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11006) );
  XNOR2_X1 U13956 ( .A(n11008), .B(n11006), .ZN(n16318) );
  INV_X1 U13957 ( .A(n11000), .ZN(n11001) );
  AND2_X1 U13958 ( .A1(n14462), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11002) );
  NAND2_X1 U13959 ( .A1(n16347), .A2(n11002), .ZN(n15485) );
  INV_X1 U13960 ( .A(n11003), .ZN(n11004) );
  NAND2_X1 U13961 ( .A1(n11004), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11005) );
  INV_X1 U13962 ( .A(n11006), .ZN(n11007) );
  NAND2_X1 U13963 ( .A1(n14459), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14452) );
  XNOR2_X1 U13964 ( .A(n14453), .B(n14452), .ZN(n11009) );
  INV_X1 U13965 ( .A(n11009), .ZN(n16306) );
  NAND3_X1 U13966 ( .A1(n16306), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14462), .ZN(n15445) );
  INV_X1 U13967 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11145) );
  OAI21_X1 U13968 ( .B1(n11009), .B2(n10807), .A(n11145), .ZN(n14451) );
  INV_X1 U13969 ( .A(n11016), .ZN(n11063) );
  XNOR2_X1 U13970 ( .A(n11062), .B(n11011), .ZN(n11036) );
  OAI21_X1 U13971 ( .B1(n11259), .B2(n11063), .A(n11036), .ZN(n11012) );
  OAI21_X1 U13972 ( .B1(n11035), .B2(n11259), .A(n11012), .ZN(n11013) );
  NAND2_X1 U13973 ( .A1(n11013), .A2(n13118), .ZN(n11018) );
  INV_X1 U13974 ( .A(n11062), .ZN(n11015) );
  OAI21_X1 U13975 ( .B1(n11016), .B2(n11015), .A(n11014), .ZN(n11017) );
  NAND2_X1 U13976 ( .A1(n11018), .A2(n11017), .ZN(n11021) );
  NAND2_X1 U13977 ( .A1(n12373), .A2(n11259), .ZN(n11019) );
  MUX2_X1 U13978 ( .A(n13477), .B(n11019), .S(n11035), .Z(n11020) );
  NAND2_X1 U13979 ( .A1(n11021), .A2(n11020), .ZN(n11024) );
  MUX2_X1 U13980 ( .A(n13477), .B(n11024), .S(n11066), .Z(n11029) );
  AND2_X1 U13981 ( .A1(n15986), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11025) );
  NAND2_X1 U13982 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15882), .ZN(
        n11027) );
  NAND2_X1 U13983 ( .A1(n11029), .A2(n20076), .ZN(n11030) );
  MUX2_X1 U13984 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11030), .S(
        n16562), .Z(n11032) );
  NAND2_X1 U13985 ( .A1(n12901), .A2(n11259), .ZN(n12863) );
  NOR2_X1 U13986 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19948) );
  AOI211_X1 U13987 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19948), .ZN(n12371) );
  INV_X1 U13988 ( .A(n12371), .ZN(n19943) );
  NAND2_X1 U13989 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19937) );
  INV_X1 U13990 ( .A(n19937), .ZN(n19951) );
  NOR2_X1 U13991 ( .A1(n19943), .A2(n19951), .ZN(n13473) );
  INV_X1 U13992 ( .A(n13473), .ZN(n12862) );
  OR3_X1 U13993 ( .A1(n12863), .A2(n19439), .A3(n12862), .ZN(n11073) );
  AOI21_X1 U13994 ( .B1(n11032), .B2(n13118), .A(n19451), .ZN(n11033) );
  NAND2_X1 U13995 ( .A1(n12863), .A2(n11033), .ZN(n11072) );
  INV_X1 U13996 ( .A(n11066), .ZN(n11034) );
  NOR2_X1 U13997 ( .A1(n11035), .A2(n11034), .ZN(n11052) );
  NAND2_X1 U13998 ( .A1(n11052), .A2(n11036), .ZN(n11037) );
  AND2_X1 U13999 ( .A1(n11049), .A2(n13473), .ZN(n11047) );
  NAND2_X1 U14000 ( .A1(n12079), .A2(n10480), .ZN(n11038) );
  NAND2_X1 U14001 ( .A1(n11038), .A2(n19439), .ZN(n11039) );
  NAND2_X1 U14002 ( .A1(n12909), .A2(n11039), .ZN(n11043) );
  NAND2_X1 U14003 ( .A1(n13682), .A2(n10480), .ZN(n11113) );
  NAND2_X1 U14004 ( .A1(n11113), .A2(n13118), .ZN(n11040) );
  NAND2_X1 U14005 ( .A1(n11040), .A2(n12096), .ZN(n11041) );
  AOI21_X1 U14006 ( .B1(n11041), .B2(n19439), .A(n11129), .ZN(n11042) );
  NAND2_X1 U14007 ( .A1(n11043), .A2(n11042), .ZN(n11114) );
  AOI21_X1 U14008 ( .B1(n11044), .B2(n12096), .A(n11060), .ZN(n11119) );
  NOR2_X1 U14009 ( .A1(n11044), .A2(n10480), .ZN(n11045) );
  OR3_X1 U14010 ( .A1(n11114), .A2(n11119), .A3(n11045), .ZN(n11046) );
  AOI21_X1 U14011 ( .B1(n12896), .B2(n11047), .A(n11046), .ZN(n12859) );
  MUX2_X1 U14012 ( .A(n11049), .B(n11048), .S(n13682), .Z(n11050) );
  NAND3_X1 U14013 ( .A1(n12896), .A2(n19937), .A3(n11050), .ZN(n11051) );
  NAND2_X1 U14014 ( .A1(n12859), .A2(n11051), .ZN(n11070) );
  NAND2_X1 U14015 ( .A1(n11052), .A2(n11063), .ZN(n11054) );
  AND2_X1 U14016 ( .A1(n12896), .A2(n14497), .ZN(n11053) );
  NAND2_X1 U14017 ( .A1(n11054), .A2(n11053), .ZN(n11058) );
  NAND2_X1 U14018 ( .A1(n11055), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11056) );
  NAND2_X1 U14019 ( .A1(n11056), .A2(n15882), .ZN(n12906) );
  INV_X1 U14020 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12905) );
  OAI21_X1 U14021 ( .B1(n11818), .B2(n12906), .A(n12905), .ZN(n11057) );
  NAND2_X1 U14022 ( .A1(n11057), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20066) );
  NAND2_X1 U14023 ( .A1(n11058), .A2(n20066), .ZN(n16560) );
  NOR2_X1 U14024 ( .A1(n12910), .A2(n13682), .ZN(n11059) );
  NAND2_X1 U14025 ( .A1(n16560), .A2(n11059), .ZN(n11069) );
  NOR2_X1 U14026 ( .A1(n12910), .A2(n11060), .ZN(n20079) );
  INV_X1 U14027 ( .A(n11061), .ZN(n11065) );
  NAND2_X1 U14028 ( .A1(n11063), .A2(n11062), .ZN(n11064) );
  NAND2_X1 U14029 ( .A1(n11065), .A2(n11064), .ZN(n11067) );
  NAND2_X1 U14030 ( .A1(n11067), .A2(n11066), .ZN(n20077) );
  NAND3_X1 U14031 ( .A1(n20079), .A2(n20076), .A3(n20077), .ZN(n11068) );
  NAND2_X1 U14032 ( .A1(n11069), .A2(n11068), .ZN(n12183) );
  NOR2_X1 U14033 ( .A1(n11070), .A2(n12183), .ZN(n11071) );
  NAND3_X1 U14034 ( .A1(n11073), .A2(n11072), .A3(n11071), .ZN(n11075) );
  NAND2_X1 U14035 ( .A1(n16562), .A2(n14497), .ZN(n13480) );
  INV_X1 U14036 ( .A(n13480), .ZN(n11074) );
  NOR2_X1 U14037 ( .A1(n12910), .A2(n13477), .ZN(n20080) );
  NAND2_X1 U14038 ( .A1(n11098), .A2(n13650), .ZN(n11093) );
  NAND2_X1 U14039 ( .A1(n11076), .A2(n13642), .ZN(n13647) );
  NOR2_X1 U14040 ( .A1(n12363), .A2(n12364), .ZN(n12362) );
  XNOR2_X1 U14041 ( .A(n11252), .B(n11077), .ZN(n11079) );
  INV_X1 U14042 ( .A(n11079), .ZN(n11078) );
  NAND2_X1 U14043 ( .A1(n12362), .A2(n11078), .ZN(n11080) );
  XNOR2_X1 U14044 ( .A(n12362), .B(n11079), .ZN(n12575) );
  NAND2_X1 U14045 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12575), .ZN(
        n12576) );
  NAND2_X1 U14046 ( .A1(n11080), .A2(n12576), .ZN(n11083) );
  XOR2_X1 U14047 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11083), .Z(
        n12356) );
  XOR2_X1 U14048 ( .A(n11082), .B(n11081), .Z(n12355) );
  NAND2_X1 U14049 ( .A1(n12356), .A2(n12355), .ZN(n12354) );
  NAND2_X1 U14050 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11083), .ZN(
        n11084) );
  NAND2_X1 U14051 ( .A1(n12354), .A2(n11084), .ZN(n11085) );
  XNOR2_X1 U14052 ( .A(n11085), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13153) );
  NAND2_X1 U14053 ( .A1(n11085), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11086) );
  XNOR2_X1 U14054 ( .A(n11088), .B(n11087), .ZN(n13508) );
  NAND2_X1 U14055 ( .A1(n13508), .A2(n19407), .ZN(n11089) );
  NAND2_X1 U14056 ( .A1(n13509), .A2(n11089), .ZN(n11092) );
  INV_X1 U14057 ( .A(n13508), .ZN(n11090) );
  NAND2_X1 U14058 ( .A1(n11090), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11091) );
  NAND2_X1 U14059 ( .A1(n11092), .A2(n11091), .ZN(n13646) );
  MUX2_X1 U14060 ( .A(n11098), .B(n11093), .S(n13645), .Z(n11097) );
  INV_X1 U14061 ( .A(n13650), .ZN(n11095) );
  NAND2_X1 U14062 ( .A1(n11095), .A2(n11101), .ZN(n11096) );
  NAND2_X1 U14063 ( .A1(n13826), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13825) );
  NAND2_X1 U14064 ( .A1(n13645), .A2(n13650), .ZN(n11099) );
  NAND2_X1 U14065 ( .A1(n11099), .A2(n11098), .ZN(n11100) );
  NAND2_X2 U14066 ( .A1(n13825), .A2(n11100), .ZN(n15829) );
  NAND2_X1 U14067 ( .A1(n11103), .A2(n10807), .ZN(n11104) );
  NAND2_X1 U14068 ( .A1(n11105), .A2(n11104), .ZN(n15827) );
  INV_X1 U14069 ( .A(n11105), .ZN(n11106) );
  NAND2_X1 U14070 ( .A1(n11106), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11107) );
  NAND2_X2 U14071 ( .A1(n15598), .A2(n11107), .ZN(n15813) );
  NAND2_X1 U14072 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15651) );
  INV_X1 U14073 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15719) );
  NOR3_X1 U14074 ( .A1(n15725), .A2(n15719), .A3(n11108), .ZN(n15687) );
  NAND2_X1 U14075 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15687), .ZN(
        n15663) );
  NOR2_X1 U14076 ( .A1(n15651), .A2(n15663), .ZN(n15520) );
  NAND2_X1 U14077 ( .A1(n15520), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11111) );
  NAND2_X1 U14078 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15746) );
  NAND2_X1 U14079 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11109) );
  NOR2_X1 U14080 ( .A1(n15746), .A2(n11109), .ZN(n11110) );
  NAND2_X1 U14081 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16541) );
  INV_X1 U14082 ( .A(n16541), .ZN(n15648) );
  NAND2_X1 U14083 ( .A1(n11110), .A2(n15648), .ZN(n15635) );
  OR2_X1 U14084 ( .A1(n11111), .A2(n15635), .ZN(n11133) );
  INV_X1 U14085 ( .A(n11133), .ZN(n11142) );
  NAND2_X2 U14086 ( .A1(n15813), .A2(n11142), .ZN(n15521) );
  NAND2_X1 U14087 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16530) );
  AND2_X2 U14088 ( .A1(n16400), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16388) );
  INV_X1 U14089 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16516) );
  INV_X1 U14090 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16502) );
  NOR2_X1 U14091 ( .A1(n16516), .A2(n16502), .ZN(n16500) );
  NAND2_X1 U14092 ( .A1(n16388), .A2(n16500), .ZN(n15492) );
  XNOR2_X1 U14093 ( .A(n15449), .B(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15464) );
  INV_X1 U14094 ( .A(n16530), .ZN(n11141) );
  NOR2_X1 U14095 ( .A1(n15826), .A2(n15595), .ZN(n11139) );
  NAND2_X1 U14096 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13831) );
  OR2_X1 U14097 ( .A1(n11112), .A2(n13831), .ZN(n11134) );
  NOR2_X1 U14098 ( .A1(n19422), .A2(n12364), .ZN(n12409) );
  INV_X1 U14099 ( .A(n12409), .ZN(n19426) );
  NAND2_X1 U14100 ( .A1(n11450), .A2(n12075), .ZN(n15701) );
  NOR2_X1 U14101 ( .A1(n12410), .A2(n19426), .ZN(n11136) );
  INV_X1 U14102 ( .A(n11136), .ZN(n11115) );
  AOI22_X1 U14103 ( .A1(n12410), .A2(n19426), .B1(n15701), .B2(n11115), .ZN(
        n13155) );
  NAND2_X1 U14104 ( .A1(n11117), .A2(n11116), .ZN(n11130) );
  NAND2_X1 U14105 ( .A1(n11118), .A2(n11259), .ZN(n12918) );
  INV_X1 U14106 ( .A(n11119), .ZN(n11120) );
  NAND2_X1 U14107 ( .A1(n12918), .A2(n11120), .ZN(n11122) );
  NAND2_X1 U14108 ( .A1(n11122), .A2(n11121), .ZN(n11127) );
  OAI22_X1 U14109 ( .A1(n11116), .A2(n19451), .B1(n13118), .B2(n19439), .ZN(
        n11123) );
  INV_X1 U14110 ( .A(n11123), .ZN(n11125) );
  AND2_X1 U14111 ( .A1(n11125), .A2(n11124), .ZN(n11126) );
  NAND2_X1 U14112 ( .A1(n11127), .A2(n11126), .ZN(n11128) );
  AOI21_X1 U14113 ( .B1(n11130), .B2(n11129), .A(n11128), .ZN(n12866) );
  INV_X1 U14114 ( .A(n12867), .ZN(n11131) );
  NAND2_X1 U14115 ( .A1(n12866), .A2(n11131), .ZN(n11132) );
  NAND2_X1 U14116 ( .A1(n11450), .A2(n11132), .ZN(n12408) );
  NAND3_X1 U14117 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13155), .A3(
        n19427), .ZN(n19408) );
  NOR2_X1 U14118 ( .A1(n11134), .A2(n19408), .ZN(n16548) );
  NAND2_X1 U14119 ( .A1(n11139), .A2(n16548), .ZN(n15794) );
  NOR2_X1 U14120 ( .A1(n11133), .A2(n15794), .ZN(n16531) );
  NAND2_X1 U14121 ( .A1(n11141), .A2(n16531), .ZN(n15623) );
  NOR2_X1 U14122 ( .A1(n15626), .A2(n15623), .ZN(n16513) );
  NAND2_X1 U14123 ( .A1(n16500), .A2(n16513), .ZN(n15613) );
  INV_X1 U14124 ( .A(n15613), .ZN(n12116) );
  NAND2_X1 U14125 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11451) );
  INV_X1 U14126 ( .A(n16500), .ZN(n11144) );
  INV_X1 U14127 ( .A(n19427), .ZN(n15834) );
  NAND2_X1 U14128 ( .A1(n19427), .A2(n11134), .ZN(n11138) );
  INV_X1 U14129 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11137) );
  INV_X1 U14130 ( .A(n15701), .ZN(n12407) );
  NAND3_X1 U14131 ( .A1(n12407), .A2(n19426), .A3(n12410), .ZN(n12400) );
  INV_X1 U14132 ( .A(n11450), .ZN(n11135) );
  NOR2_X2 U14133 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20037) );
  AND2_X2 U14134 ( .A1(n20037), .A2(n12184), .ZN(n19404) );
  INV_X2 U14135 ( .A(n19404), .ZN(n19254) );
  NAND2_X1 U14136 ( .A1(n11135), .A2(n19254), .ZN(n19423) );
  OAI211_X1 U14137 ( .C1(n11136), .C2(n12408), .A(n12400), .B(n19423), .ZN(
        n13156) );
  AOI21_X1 U14138 ( .B1(n11137), .B2(n19427), .A(n13156), .ZN(n19406) );
  AND2_X1 U14139 ( .A1(n11138), .A2(n19406), .ZN(n13832) );
  INV_X1 U14140 ( .A(n11139), .ZN(n16547) );
  NAND2_X1 U14141 ( .A1(n19427), .A2(n16547), .ZN(n11140) );
  OAI221_X1 U14142 ( .B1(n15834), .B2(n11142), .C1(n15834), .C2(n11141), .A(
        n15795), .ZN(n15631) );
  AOI21_X1 U14143 ( .B1(n15626), .B2(n19427), .A(n15631), .ZN(n16515) );
  INV_X1 U14144 ( .A(n16515), .ZN(n11143) );
  AOI21_X1 U14145 ( .B1(n11144), .B2(n19427), .A(n11143), .ZN(n14485) );
  INV_X1 U14146 ( .A(n14485), .ZN(n15618) );
  AOI21_X1 U14147 ( .B1(n12116), .B2(n11451), .A(n15618), .ZN(n12118) );
  NOR2_X1 U14148 ( .A1(n12118), .A2(n11145), .ZN(n11456) );
  NAND2_X1 U14149 ( .A1(n12128), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11149) );
  AOI22_X1 U14150 ( .A1(n14468), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11147) );
  NAND2_X1 U14151 ( .A1(n11169), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11146) );
  AND2_X1 U14152 ( .A1(n11147), .A2(n11146), .ZN(n11148) );
  NAND2_X1 U14153 ( .A1(n11149), .A2(n11148), .ZN(n13602) );
  INV_X1 U14154 ( .A(n11151), .ZN(n11152) );
  NOR2_X1 U14155 ( .A1(n11153), .A2(n11152), .ZN(n11154) );
  NAND2_X1 U14156 ( .A1(n12128), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11160) );
  AOI22_X1 U14157 ( .A1(n14468), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11158) );
  NAND2_X1 U14158 ( .A1(n11169), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11157) );
  AND2_X1 U14159 ( .A1(n11158), .A2(n11157), .ZN(n11159) );
  NAND2_X1 U14160 ( .A1(n11160), .A2(n11159), .ZN(n12696) );
  NAND2_X1 U14161 ( .A1(n12128), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11162) );
  AOI22_X1 U14162 ( .A1(n14468), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11161) );
  OAI211_X1 U14163 ( .C1(n11163), .C2(n11206), .A(n11162), .B(n11161), .ZN(
        n12688) );
  INV_X1 U14164 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11166) );
  NAND2_X1 U14165 ( .A1(n11169), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11165) );
  NAND2_X1 U14166 ( .A1(n14468), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11164) );
  OAI211_X1 U14167 ( .C1(n14497), .C2(n11166), .A(n11165), .B(n11164), .ZN(
        n11167) );
  AOI21_X1 U14168 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11167), .ZN(n13475) );
  NAND2_X1 U14169 ( .A1(n12128), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11173) );
  AOI22_X1 U14170 ( .A1(n14468), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11171) );
  NAND2_X1 U14171 ( .A1(n11169), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11170) );
  AND2_X1 U14172 ( .A1(n11171), .A2(n11170), .ZN(n11172) );
  NAND2_X1 U14173 ( .A1(n11173), .A2(n11172), .ZN(n14523) );
  NAND2_X1 U14174 ( .A1(n14522), .A2(n14523), .ZN(n14525) );
  AOI22_X1 U14175 ( .A1(n14468), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11175) );
  NAND2_X1 U14176 ( .A1(n11169), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11174) );
  NAND2_X1 U14177 ( .A1(n11175), .A2(n11174), .ZN(n11176) );
  AOI21_X1 U14178 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11176), .ZN(n12832) );
  AOI22_X1 U14179 ( .A1(n14468), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11178) );
  NAND2_X1 U14180 ( .A1(n11169), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11177) );
  NAND2_X1 U14181 ( .A1(n11178), .A2(n11177), .ZN(n11179) );
  AOI21_X1 U14182 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11179), .ZN(n12841) );
  NAND2_X1 U14183 ( .A1(n12831), .A2(n11180), .ZN(n13138) );
  NAND2_X1 U14184 ( .A1(n11169), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11182) );
  NAND2_X1 U14185 ( .A1(n14468), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11181) );
  OAI211_X1 U14186 ( .C1(n14497), .C2(n10175), .A(n11182), .B(n11181), .ZN(
        n11183) );
  AOI21_X1 U14187 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11183), .ZN(n13137) );
  NAND2_X1 U14188 ( .A1(n12128), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11187) );
  AOI22_X1 U14189 ( .A1(n14468), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11185) );
  NAND2_X1 U14190 ( .A1(n11169), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11184) );
  AND2_X1 U14191 ( .A1(n11185), .A2(n11184), .ZN(n11186) );
  NAND2_X1 U14192 ( .A1(n11187), .A2(n11186), .ZN(n13143) );
  INV_X1 U14193 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11190) );
  NAND2_X1 U14194 ( .A1(n11169), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11189) );
  NAND2_X1 U14195 ( .A1(n14468), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11188) );
  OAI211_X1 U14196 ( .C1(n14497), .C2(n11190), .A(n11189), .B(n11188), .ZN(
        n11191) );
  AOI21_X1 U14197 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11191), .ZN(n13388) );
  NAND2_X1 U14198 ( .A1(n12128), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11193) );
  AOI22_X1 U14199 ( .A1(n14468), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11192) );
  OAI211_X1 U14200 ( .C1(n11194), .C2(n11206), .A(n11193), .B(n11192), .ZN(
        n13396) );
  INV_X1 U14201 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U14202 ( .A1(n14468), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11195) );
  OAI21_X1 U14203 ( .B1(n11206), .B2(n13663), .A(n11195), .ZN(n11196) );
  AOI21_X1 U14204 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11196), .ZN(n13660) );
  NAND2_X1 U14205 ( .A1(n11169), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11198) );
  NAND2_X1 U14206 ( .A1(n14468), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11197) );
  OAI211_X1 U14207 ( .C1(n14497), .C2(n10179), .A(n11198), .B(n11197), .ZN(
        n11199) );
  AOI21_X1 U14208 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11199), .ZN(n13748) );
  INV_X1 U14209 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11202) );
  NAND2_X1 U14210 ( .A1(n11169), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11201) );
  NAND2_X1 U14211 ( .A1(n14468), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11200) );
  OAI211_X1 U14212 ( .C1(n14497), .C2(n11202), .A(n11201), .B(n11200), .ZN(
        n11203) );
  AOI21_X1 U14213 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11203), .ZN(n13767) );
  NAND2_X1 U14214 ( .A1(n12128), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11205) );
  AOI22_X1 U14215 ( .A1(n14468), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11204) );
  OAI211_X1 U14216 ( .C1(n11207), .C2(n11206), .A(n11205), .B(n11204), .ZN(
        n13850) );
  INV_X1 U14217 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15563) );
  NAND2_X1 U14218 ( .A1(n11169), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11209) );
  NAND2_X1 U14219 ( .A1(n14468), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11208) );
  OAI211_X1 U14220 ( .C1(n14497), .C2(n15563), .A(n11209), .B(n11208), .ZN(
        n11210) );
  AOI21_X1 U14221 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11210), .ZN(n15353) );
  AOI22_X1 U14222 ( .A1(n14468), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11212) );
  NAND2_X1 U14223 ( .A1(n11169), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11211) );
  NAND2_X1 U14224 ( .A1(n11212), .A2(n11211), .ZN(n11213) );
  AOI21_X1 U14225 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11213), .ZN(n15347) );
  INV_X1 U14226 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15538) );
  NAND2_X1 U14227 ( .A1(n11169), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U14228 ( .A1(n14468), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11214) );
  OAI211_X1 U14229 ( .C1(n14497), .C2(n15538), .A(n11215), .B(n11214), .ZN(
        n11216) );
  AOI21_X1 U14230 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11216), .ZN(n15192) );
  AOI22_X1 U14231 ( .A1(n14468), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11218) );
  NAND2_X1 U14232 ( .A1(n11169), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11217) );
  NAND2_X1 U14233 ( .A1(n11218), .A2(n11217), .ZN(n11219) );
  AOI21_X1 U14234 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11219), .ZN(n15335) );
  NAND2_X1 U14235 ( .A1(n12128), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11223) );
  AOI22_X1 U14236 ( .A1(n14468), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11221) );
  NAND2_X1 U14237 ( .A1(n11169), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11220) );
  AND2_X1 U14238 ( .A1(n11221), .A2(n11220), .ZN(n11222) );
  NAND2_X1 U14239 ( .A1(n11223), .A2(n11222), .ZN(n15325) );
  AOI22_X1 U14240 ( .A1(n14468), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11225) );
  NAND2_X1 U14241 ( .A1(n11169), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11224) );
  NAND2_X1 U14242 ( .A1(n11225), .A2(n11224), .ZN(n11226) );
  AOI21_X1 U14243 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11226), .ZN(n15321) );
  INV_X1 U14244 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11229) );
  NAND2_X1 U14245 ( .A1(n11169), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11228) );
  NAND2_X1 U14246 ( .A1(n14468), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11227) );
  OAI211_X1 U14247 ( .C1(n14497), .C2(n11229), .A(n11228), .B(n11227), .ZN(
        n11230) );
  AOI21_X1 U14248 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11230), .ZN(n15312) );
  AOI22_X1 U14249 ( .A1(n14468), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11232) );
  NAND2_X1 U14250 ( .A1(n11169), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11231) );
  NAND2_X1 U14251 ( .A1(n11232), .A2(n11231), .ZN(n11233) );
  AOI21_X1 U14252 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11233), .ZN(n15304) );
  NAND2_X1 U14253 ( .A1(n12128), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11237) );
  AOI22_X1 U14254 ( .A1(n14468), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11235) );
  NAND2_X1 U14255 ( .A1(n11169), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11234) );
  AND2_X1 U14256 ( .A1(n11235), .A2(n11234), .ZN(n11236) );
  NAND2_X1 U14257 ( .A1(n11237), .A2(n11236), .ZN(n15296) );
  NAND2_X1 U14258 ( .A1(n12128), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11241) );
  AOI22_X1 U14259 ( .A1(n14468), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11239) );
  NAND2_X1 U14260 ( .A1(n11169), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11238) );
  AND2_X1 U14261 ( .A1(n11239), .A2(n11238), .ZN(n11240) );
  NAND2_X1 U14262 ( .A1(n11241), .A2(n11240), .ZN(n12115) );
  NAND2_X1 U14263 ( .A1(n12128), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11245) );
  AOI22_X1 U14264 ( .A1(n14468), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11243) );
  NAND2_X1 U14265 ( .A1(n11169), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11242) );
  AND2_X1 U14266 ( .A1(n11243), .A2(n11242), .ZN(n11244) );
  NAND2_X1 U14267 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  OR2_X1 U14268 ( .A1(n12113), .A2(n11246), .ZN(n11247) );
  NAND2_X1 U14269 ( .A1(n14467), .A2(n11247), .ZN(n16309) );
  NAND2_X1 U14270 ( .A1(n12925), .A2(n12907), .ZN(n11248) );
  NAND2_X1 U14271 ( .A1(n11249), .A2(n11248), .ZN(n11250) );
  NAND2_X1 U14272 ( .A1(n11450), .A2(n11250), .ZN(n19411) );
  NAND2_X1 U14273 ( .A1(n11410), .A2(n11252), .ZN(n11257) );
  AND2_X1 U14274 ( .A1(n11253), .A2(n13298), .ZN(n11254) );
  NAND2_X1 U14275 ( .A1(n11255), .A2(n11254), .ZN(n11274) );
  NAND2_X1 U14276 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11256) );
  NAND4_X1 U14277 ( .A1(n11257), .A2(n9843), .A3(n11274), .A4(n11256), .ZN(
        n15835) );
  AND2_X2 U14278 ( .A1(n11258), .A2(n12631), .ZN(n11276) );
  NAND2_X1 U14279 ( .A1(n11276), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11264) );
  INV_X1 U14280 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n11261) );
  NAND2_X1 U14281 ( .A1(n11259), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11260) );
  OAI211_X1 U14282 ( .C1(n12096), .C2(n11261), .A(n11260), .B(n13298), .ZN(
        n11262) );
  INV_X1 U14283 ( .A(n11262), .ZN(n11263) );
  NAND2_X1 U14284 ( .A1(n11264), .A2(n11263), .ZN(n15836) );
  NAND2_X1 U14285 ( .A1(n11276), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11266) );
  INV_X2 U14286 ( .A(n9843), .ZN(n11440) );
  AOI22_X1 U14287 ( .A1(n11440), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11254), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11265) );
  XNOR2_X1 U14288 ( .A(n15838), .B(n11271), .ZN(n15270) );
  INV_X1 U14289 ( .A(n12631), .ZN(n11269) );
  NAND2_X1 U14290 ( .A1(n12079), .A2(n12096), .ZN(n11267) );
  MUX2_X1 U14291 ( .A(n11267), .B(n20064), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11268) );
  OAI21_X1 U14292 ( .B1(n11270), .B2(n11269), .A(n11268), .ZN(n15269) );
  NAND2_X1 U14293 ( .A1(n11271), .A2(n15838), .ZN(n11272) );
  NAND2_X1 U14294 ( .A1(n15272), .A2(n11272), .ZN(n11280) );
  NAND2_X1 U14295 ( .A1(n11410), .A2(n11273), .ZN(n11275) );
  OAI211_X1 U14296 ( .C1(n13298), .C2(n20056), .A(n11275), .B(n11274), .ZN(
        n11279) );
  XNOR2_X1 U14297 ( .A(n11280), .B(n11279), .ZN(n12397) );
  NAND2_X1 U14298 ( .A1(n11276), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11278) );
  AOI22_X1 U14299 ( .A1(n11440), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12080), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11277) );
  AND2_X1 U14300 ( .A1(n11278), .A2(n11277), .ZN(n12396) );
  INV_X1 U14301 ( .A(n11279), .ZN(n11281) );
  NAND2_X1 U14302 ( .A1(n11281), .A2(n11280), .ZN(n11282) );
  NAND2_X1 U14303 ( .A1(n11276), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U14304 ( .A1(n12080), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_3__SCAN_IN), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n11284) );
  NAND2_X1 U14305 ( .A1(n11440), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11283) );
  AND2_X1 U14306 ( .A1(n11284), .A2(n11283), .ZN(n11288) );
  INV_X1 U14307 ( .A(n11285), .ZN(n11286) );
  NAND2_X1 U14308 ( .A1(n11410), .A2(n11286), .ZN(n11287) );
  AOI22_X1 U14309 ( .A1(n11276), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n11410), 
        .B2(n11290), .ZN(n11292) );
  AOI22_X1 U14310 ( .A1(n11440), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12080), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11291) );
  NAND2_X1 U14311 ( .A1(n11292), .A2(n11291), .ZN(n19268) );
  INV_X1 U14312 ( .A(n13551), .ZN(n11297) );
  NAND2_X1 U14313 ( .A1(n11276), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11296) );
  NAND2_X1 U14314 ( .A1(n11410), .A2(n11293), .ZN(n11295) );
  AOI22_X1 U14315 ( .A1(n11440), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12080), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11294) );
  NAND3_X1 U14316 ( .A1(n11296), .A2(n11295), .A3(n11294), .ZN(n13549) );
  NAND2_X1 U14317 ( .A1(n11297), .A2(n13549), .ZN(n13553) );
  NAND2_X1 U14318 ( .A1(n11410), .A2(n11298), .ZN(n11299) );
  NAND2_X1 U14319 ( .A1(n11276), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11301) );
  INV_X2 U14320 ( .A(n11319), .ZN(n12080) );
  AOI22_X1 U14321 ( .A1(n11440), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12080), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11300) );
  NAND2_X1 U14322 ( .A1(n11301), .A2(n11300), .ZN(n13469) );
  AOI21_X1 U14323 ( .B1(n11410), .B2(n11302), .A(n13472), .ZN(n13052) );
  NAND2_X1 U14324 ( .A1(n11276), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14325 ( .A1(n11440), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12080), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11303) );
  NAND2_X1 U14326 ( .A1(n11276), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11318) );
  AOI22_X1 U14327 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14328 ( .A1(n11818), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11882), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14329 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11884), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14330 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11306) );
  NAND4_X1 U14331 ( .A1(n11309), .A2(n11308), .A3(n11307), .A4(n11306), .ZN(
        n11315) );
  AOI22_X1 U14332 ( .A1(n10729), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14333 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14334 ( .A1(n10798), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14335 ( .A1(n12869), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11310) );
  NAND4_X1 U14336 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n11314) );
  NAND2_X1 U14337 ( .A1(n11410), .A2(n12837), .ZN(n11317) );
  AOI22_X1 U14338 ( .A1(n11440), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12080), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11316) );
  NAND3_X1 U14339 ( .A1(n11318), .A2(n11317), .A3(n11316), .ZN(n13061) );
  INV_X1 U14340 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n11320) );
  OAI22_X1 U14341 ( .A1(n9843), .A2(n11320), .B1(n11319), .B2(n15814), .ZN(
        n11333) );
  INV_X1 U14342 ( .A(n11410), .ZN(n11331) );
  AOI22_X1 U14343 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11832), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14344 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n11882), .ZN(n11323) );
  AOI22_X1 U14345 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n11884), .ZN(n11322) );
  AOI22_X1 U14346 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11321) );
  NAND4_X1 U14347 ( .A1(n11324), .A2(n11323), .A3(n11322), .A4(n11321), .ZN(
        n11330) );
  AOI22_X1 U14348 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10774), .B1(
        n10729), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14349 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14350 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10730), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14351 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12869), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11325) );
  NAND4_X1 U14352 ( .A1(n11328), .A2(n11327), .A3(n11326), .A4(n11325), .ZN(
        n11329) );
  NOR2_X1 U14353 ( .A1(n11331), .A2(n12840), .ZN(n11332) );
  AOI211_X1 U14354 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n11276), .A(n11333), .B(
        n11332), .ZN(n13055) );
  NAND2_X1 U14355 ( .A1(n11276), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14356 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11832), .B1(
        n11305), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14357 ( .A1(n11818), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n11882), .ZN(n11336) );
  AOI22_X1 U14358 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11884), .B1(
        n11816), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14359 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11334) );
  NAND4_X1 U14360 ( .A1(n11337), .A2(n11336), .A3(n11335), .A4(n11334), .ZN(
        n11343) );
  AOI22_X1 U14361 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10774), .B1(
        n10729), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14362 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14363 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12869), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14364 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10798), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11338) );
  NAND4_X1 U14365 ( .A1(n11341), .A2(n11340), .A3(n11339), .A4(n11338), .ZN(
        n11342) );
  NAND2_X1 U14366 ( .A1(n11410), .A2(n13136), .ZN(n11345) );
  AOI22_X1 U14367 ( .A1(n11440), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11344) );
  NAND3_X1 U14368 ( .A1(n11346), .A2(n11345), .A3(n11344), .ZN(n13058) );
  NAND2_X1 U14369 ( .A1(n11276), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14370 ( .A1(n11440), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14371 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11832), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14372 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n11399), .ZN(n11349) );
  AOI22_X1 U14373 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__3__SCAN_IN), .B2(n11884), .ZN(n11348) );
  AOI22_X1 U14374 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11347) );
  NAND4_X1 U14375 ( .A1(n11350), .A2(n11349), .A3(n11348), .A4(n11347), .ZN(
        n11356) );
  AOI22_X1 U14376 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10774), .B1(
        n10729), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14377 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14378 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n10798), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14379 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12869), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11351) );
  NAND4_X1 U14380 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11355) );
  NAND2_X1 U14381 ( .A1(n11410), .A2(n11783), .ZN(n11357) );
  NAND2_X1 U14382 ( .A1(n11276), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14383 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11832), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14384 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n11399), .ZN(n11362) );
  AOI22_X1 U14385 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__4__SCAN_IN), .B2(n11884), .ZN(n11361) );
  AOI22_X1 U14386 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11360) );
  NAND4_X1 U14387 ( .A1(n11363), .A2(n11362), .A3(n11361), .A4(n11360), .ZN(
        n11369) );
  AOI22_X1 U14388 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10774), .B1(
        n10729), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14389 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14390 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10730), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14391 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12869), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11364) );
  NAND4_X1 U14392 ( .A1(n11367), .A2(n11366), .A3(n11365), .A4(n11364), .ZN(
        n11368) );
  NAND2_X1 U14393 ( .A1(n11410), .A2(n11784), .ZN(n11371) );
  AOI22_X1 U14394 ( .A1(n11440), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11370) );
  NAND3_X1 U14395 ( .A1(n11372), .A2(n11371), .A3(n11370), .ZN(n13080) );
  NAND2_X1 U14396 ( .A1(n15224), .A2(n13080), .ZN(n13226) );
  NAND2_X1 U14397 ( .A1(n11276), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14398 ( .A1(n11440), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14399 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14400 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11882), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14401 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11884), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11374) );
  AOI22_X1 U14402 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11373) );
  NAND4_X1 U14403 ( .A1(n11376), .A2(n11375), .A3(n11374), .A4(n11373), .ZN(
        n11382) );
  AOI22_X1 U14404 ( .A1(n10729), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14405 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14406 ( .A1(n10798), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14407 ( .A1(n12869), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11377) );
  NAND4_X1 U14408 ( .A1(n11380), .A2(n11379), .A3(n11378), .A4(n11377), .ZN(
        n11381) );
  NAND2_X1 U14409 ( .A1(n11410), .A2(n13394), .ZN(n11383) );
  NAND2_X1 U14410 ( .A1(n11276), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14411 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11305), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14412 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n11399), .ZN(n11388) );
  AOI22_X1 U14413 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n11816), .ZN(n11387) );
  AOI22_X1 U14414 ( .A1(n10704), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11884), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11386) );
  NAND4_X1 U14415 ( .A1(n11389), .A2(n11388), .A3(n11387), .A4(n11386), .ZN(
        n11395) );
  AOI22_X1 U14416 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10774), .B1(
        n10729), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14417 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14418 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10776), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14419 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12869), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11390) );
  NAND4_X1 U14420 ( .A1(n11393), .A2(n11392), .A3(n11391), .A4(n11390), .ZN(
        n11394) );
  NOR2_X1 U14421 ( .A1(n11395), .A2(n11394), .ZN(n11785) );
  INV_X1 U14422 ( .A(n11785), .ZN(n13656) );
  NAND2_X1 U14423 ( .A1(n11410), .A2(n13656), .ZN(n11397) );
  AOI22_X1 U14424 ( .A1(n11440), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11396) );
  NAND3_X1 U14425 ( .A1(n11398), .A2(n11397), .A3(n11396), .ZN(n15752) );
  NAND2_X1 U14426 ( .A1(n13228), .A2(n15752), .ZN(n15753) );
  NAND2_X1 U14427 ( .A1(n11276), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14428 ( .A1(n11440), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14429 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11832), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U14430 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n11399), .ZN(n11402) );
  AOI22_X1 U14431 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n11884), .ZN(n11401) );
  AOI22_X1 U14432 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11400) );
  NAND4_X1 U14433 ( .A1(n11403), .A2(n11402), .A3(n11401), .A4(n11400), .ZN(
        n11409) );
  AOI22_X1 U14434 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10774), .B1(
        n10729), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14435 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11406) );
  INV_X1 U14436 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19470) );
  AOI22_X1 U14437 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10798), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14438 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12869), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11404) );
  NAND4_X1 U14439 ( .A1(n11407), .A2(n11406), .A3(n11405), .A4(n11404), .ZN(
        n11408) );
  NAND2_X1 U14440 ( .A1(n11410), .A2(n13601), .ZN(n11411) );
  NAND2_X1 U14441 ( .A1(n11276), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11415) );
  AOI22_X1 U14442 ( .A1(n11440), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11414) );
  NAND2_X1 U14443 ( .A1(n11415), .A2(n11414), .ZN(n13754) );
  NAND2_X1 U14444 ( .A1(n13753), .A2(n13754), .ZN(n13840) );
  NAND2_X1 U14445 ( .A1(n11276), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14446 ( .A1(n11440), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11416) );
  NAND2_X1 U14447 ( .A1(n11276), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14448 ( .A1(n11440), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11418) );
  NAND2_X1 U14449 ( .A1(n11419), .A2(n11418), .ZN(n13856) );
  NAND2_X1 U14450 ( .A1(n11276), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14451 ( .A1(n11440), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11420) );
  AND2_X1 U14452 ( .A1(n11421), .A2(n11420), .ZN(n13893) );
  NAND2_X1 U14453 ( .A1(n11276), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14454 ( .A1(n11440), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11422) );
  AND2_X1 U14455 ( .A1(n11423), .A2(n11422), .ZN(n15427) );
  OR2_X2 U14456 ( .A1(n15428), .A2(n15427), .ZN(n15430) );
  NAND2_X1 U14457 ( .A1(n11276), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14458 ( .A1(n11440), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11424) );
  AND2_X1 U14459 ( .A1(n11425), .A2(n11424), .ZN(n15195) );
  NAND2_X1 U14460 ( .A1(n11276), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14461 ( .A1(n11440), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11426) );
  NAND2_X1 U14462 ( .A1(n11427), .A2(n11426), .ZN(n15409) );
  NAND2_X1 U14463 ( .A1(n11276), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14464 ( .A1(n11440), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11428) );
  NAND2_X1 U14465 ( .A1(n11276), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14466 ( .A1(n11440), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11430) );
  AND2_X1 U14467 ( .A1(n11431), .A2(n11430), .ZN(n15399) );
  OR2_X2 U14468 ( .A1(n16370), .A2(n15399), .ZN(n15401) );
  NAND2_X1 U14469 ( .A1(n11276), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14470 ( .A1(n11440), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11432) );
  AND2_X1 U14471 ( .A1(n11433), .A2(n11432), .ZN(n15391) );
  NOR2_X2 U14472 ( .A1(n15401), .A2(n15391), .ZN(n15392) );
  NAND2_X1 U14473 ( .A1(n11276), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14474 ( .A1(n11440), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11434) );
  NAND2_X1 U14475 ( .A1(n11435), .A2(n11434), .ZN(n15382) );
  NAND2_X1 U14476 ( .A1(n11276), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14477 ( .A1(n11440), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11436) );
  NAND2_X1 U14478 ( .A1(n11437), .A2(n11436), .ZN(n15374) );
  NAND2_X1 U14479 ( .A1(n11276), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14480 ( .A1(n11440), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11438) );
  NAND2_X1 U14481 ( .A1(n11439), .A2(n11438), .ZN(n12110) );
  NAND2_X1 U14482 ( .A1(n11276), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U14483 ( .A1(n11440), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11441) );
  AND2_X1 U14484 ( .A1(n11442), .A2(n11441), .ZN(n11444) );
  NAND2_X1 U14485 ( .A1(n11443), .A2(n11444), .ZN(n11445) );
  NAND2_X1 U14486 ( .A1(n12916), .A2(n11446), .ZN(n12898) );
  NAND2_X1 U14487 ( .A1(n11447), .A2(n11259), .ZN(n11448) );
  NAND2_X1 U14488 ( .A1(n12898), .A2(n11448), .ZN(n11449) );
  NOR3_X1 U14489 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n11451), .A3(
        n15613), .ZN(n11452) );
  INV_X1 U14490 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20014) );
  NOR2_X1 U14491 ( .A1(n19254), .A2(n20014), .ZN(n15458) );
  AOI211_X1 U14492 ( .C1(n15464), .C2(n19429), .A(n11456), .B(n11455), .ZN(
        n11457) );
  OAI21_X1 U14493 ( .B1(n15466), .B2(n19436), .A(n11457), .ZN(P2_U3017) );
  INV_X1 U14494 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17327) );
  NOR2_X4 U14495 ( .A1(n17094), .A2(n11467), .ZN(n17438) );
  AOI22_X1 U14496 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11475) );
  NAND3_X2 U14497 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n18887), .ZN(n11517) );
  INV_X4 U14498 ( .A(n9803), .ZN(n17447) );
  INV_X1 U14499 ( .A(n17126), .ZN(n11458) );
  AOI22_X1 U14500 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14501 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11462) );
  OAI211_X1 U14502 ( .C1(n17447), .C2(n17459), .A(n11463), .B(n11462), .ZN(
        n11473) );
  INV_X1 U14503 ( .A(n11466), .ZN(n11464) );
  AOI22_X1 U14504 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14505 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11470) );
  INV_X1 U14506 ( .A(n11625), .ZN(n11491) );
  INV_X2 U14507 ( .A(n11491), .ZN(n17165) );
  AOI22_X1 U14508 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11469) );
  NAND2_X1 U14509 ( .A1(n11665), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11468) );
  NAND4_X1 U14510 ( .A1(n11471), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(
        n11472) );
  AOI211_X1 U14511 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n11473), .B(n11472), .ZN(n11474) );
  OAI211_X1 U14512 ( .C1(n10412), .C2(n17327), .A(n11475), .B(n11474), .ZN(
        n17613) );
  INV_X1 U14513 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17414) );
  INV_X2 U14514 ( .A(n9847), .ZN(n17394) );
  INV_X2 U14515 ( .A(n11496), .ZN(n17410) );
  AOI22_X1 U14516 ( .A1(n17410), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11476) );
  AOI22_X1 U14517 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11626), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14518 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11480) );
  INV_X4 U14519 ( .A(n10416), .ZN(n17396) );
  AOI22_X1 U14520 ( .A1(n11629), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11479) );
  NAND2_X1 U14521 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11478) );
  INV_X1 U14522 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17326) );
  AOI22_X1 U14523 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11665), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11483) );
  OAI21_X1 U14524 ( .B1(n10412), .B2(n17326), .A(n11483), .ZN(n11487) );
  INV_X1 U14525 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U14526 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14527 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11484) );
  OAI211_X1 U14528 ( .C1(n11517), .C2(n17328), .A(n11485), .B(n11484), .ZN(
        n11486) );
  AOI211_X1 U14529 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n11487), .B(n11486), .ZN(n11495) );
  AOI22_X1 U14530 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11490) );
  INV_X1 U14531 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U14532 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11492) );
  OAI21_X1 U14533 ( .B1(n17453), .B2(n17325), .A(n11492), .ZN(n11493) );
  AOI22_X1 U14534 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11506) );
  INV_X1 U14535 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17446) );
  AOI22_X1 U14536 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14537 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11497) );
  OAI211_X1 U14538 ( .C1(n17441), .C2(n17446), .A(n11498), .B(n11497), .ZN(
        n11504) );
  AOI22_X1 U14539 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14540 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14541 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11500) );
  NAND2_X1 U14542 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11499) );
  NAND4_X1 U14543 ( .A1(n11502), .A2(n11501), .A3(n11500), .A4(n11499), .ZN(
        n11503) );
  INV_X1 U14544 ( .A(n11565), .ZN(n11547) );
  INV_X1 U14545 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17361) );
  AOI22_X1 U14546 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11516) );
  INV_X1 U14547 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17363) );
  AOI22_X1 U14548 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14549 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11507) );
  OAI211_X1 U14550 ( .C1(n17447), .C2(n17363), .A(n11508), .B(n11507), .ZN(
        n11514) );
  AOI22_X1 U14551 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14552 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14553 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11510) );
  NAND2_X1 U14554 ( .A1(n11665), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11509) );
  NAND4_X1 U14555 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11513) );
  AOI211_X1 U14556 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n11514), .B(n11513), .ZN(n11515) );
  AOI22_X1 U14557 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14558 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14559 ( .A1(n11629), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11665), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11525) );
  INV_X1 U14560 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17260) );
  OAI22_X1 U14561 ( .A1(n17258), .A2(n17476), .B1(n17416), .B2(n17260), .ZN(
        n11523) );
  AOI22_X1 U14562 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14563 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14564 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11519) );
  NAND2_X1 U14565 ( .A1(n9803), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11518) );
  NAND4_X1 U14566 ( .A1(n11521), .A2(n11520), .A3(n11519), .A4(n11518), .ZN(
        n11522) );
  AOI211_X1 U14567 ( .C1(n17438), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n11523), .B(n11522), .ZN(n11524) );
  NAND4_X1 U14568 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(
        n18457) );
  NOR2_X1 U14569 ( .A1(n18462), .A2(n18457), .ZN(n13964) );
  AOI22_X1 U14570 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11528) );
  INV_X1 U14571 ( .A(n11528), .ZN(n11535) );
  INV_X1 U14572 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17355) );
  AOI22_X1 U14573 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11533) );
  INV_X1 U14574 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U14575 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11529) );
  OAI21_X1 U14576 ( .B1(n17453), .B2(n17214), .A(n11529), .ZN(n11532) );
  AOI22_X1 U14577 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14578 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14579 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11536) );
  OAI21_X1 U14580 ( .B1(n17453), .B2(n17233), .A(n11536), .ZN(n11546) );
  INV_X1 U14581 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U14582 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11544) );
  INV_X1 U14583 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14584 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11537) );
  OAI21_X1 U14585 ( .B1(n17426), .B2(n11538), .A(n11537), .ZN(n11542) );
  INV_X1 U14586 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15859) );
  AOI22_X1 U14587 ( .A1(n17396), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U14588 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11626), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11539) );
  OAI211_X1 U14589 ( .C1(n17447), .C2(n15859), .A(n11540), .B(n11539), .ZN(
        n11541) );
  AOI211_X1 U14590 ( .C1(n11665), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n11542), .B(n11541), .ZN(n11543) );
  OAI211_X1 U14591 ( .C1(n10412), .C2(n17229), .A(n11544), .B(n11543), .ZN(
        n11545) );
  NAND3_X1 U14592 ( .A1(n11547), .A2(n13964), .A3(n11563), .ZN(n11568) );
  INV_X1 U14593 ( .A(n18462), .ZN(n11560) );
  INV_X1 U14594 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14595 ( .A1(n14033), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14596 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11548) );
  OAI211_X1 U14597 ( .C1(n17426), .C2(n11550), .A(n11549), .B(n11548), .ZN(
        n11558) );
  INV_X1 U14598 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14024) );
  AOI22_X1 U14599 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11556) );
  INV_X1 U14600 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17278) );
  AOI22_X1 U14601 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11551) );
  OAI21_X1 U14602 ( .B1(n17258), .B2(n17278), .A(n11551), .ZN(n11554) );
  INV_X1 U14603 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17405) );
  AOI22_X1 U14604 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11552) );
  OAI21_X1 U14605 ( .B1(n17447), .B2(n17405), .A(n11552), .ZN(n11553) );
  AOI211_X1 U14606 ( .C1(n11667), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n11554), .B(n11553), .ZN(n11555) );
  OAI211_X1 U14607 ( .C1(n17415), .C2(n14024), .A(n11556), .B(n11555), .ZN(
        n11557) );
  AOI211_X4 U14608 ( .C1(n11665), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n11558), .B(n11557), .ZN(n11601) );
  NAND2_X1 U14609 ( .A1(n18467), .A2(n11601), .ZN(n15886) );
  NAND2_X1 U14610 ( .A1(n11567), .A2(n15886), .ZN(n11574) );
  NOR2_X1 U14611 ( .A1(n17081), .A2(n18448), .ZN(n11572) );
  NAND2_X1 U14612 ( .A1(n13962), .A2(n18467), .ZN(n18899) );
  NAND2_X1 U14613 ( .A1(n18478), .A2(n18899), .ZN(n15990) );
  NAND2_X1 U14614 ( .A1(n11572), .A2(n15990), .ZN(n13954) );
  NAND2_X1 U14615 ( .A1(n11601), .A2(n11563), .ZN(n15890) );
  AOI21_X1 U14616 ( .B1(n11567), .B2(n15890), .A(n18441), .ZN(n11564) );
  NOR2_X2 U14617 ( .A1(n19084), .A2(n18441), .ZN(n11600) );
  AOI211_X1 U14618 ( .C1(n11560), .C2(n18467), .A(n11600), .B(n18452), .ZN(
        n11562) );
  OAI21_X1 U14619 ( .B1(n11563), .B2(n10430), .A(n18462), .ZN(n11561) );
  NAND2_X1 U14620 ( .A1(n13962), .A2(n18462), .ZN(n11576) );
  NOR2_X1 U14621 ( .A1(n11601), .A2(n11568), .ZN(n13957) );
  NOR2_X1 U14622 ( .A1(n16752), .A2(n11569), .ZN(n12150) );
  NOR2_X1 U14623 ( .A1(n19084), .A2(n12150), .ZN(n11571) );
  AOI21_X1 U14624 ( .B1(n11571), .B2(n11573), .A(n11570), .ZN(n11577) );
  INV_X2 U14625 ( .A(n18900), .ZN(n18878) );
  NOR2_X1 U14626 ( .A1(n11600), .A2(n11572), .ZN(n19096) );
  INV_X1 U14627 ( .A(n11573), .ZN(n11575) );
  NAND2_X1 U14628 ( .A1(n11575), .A2(n11574), .ZN(n11599) );
  NAND2_X1 U14629 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18903), .ZN(
        n11593) );
  OAI22_X1 U14630 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18914), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11581), .ZN(n11586) );
  NOR2_X1 U14631 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18914), .ZN(
        n11582) );
  NAND2_X1 U14632 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11581), .ZN(
        n11587) );
  AOI22_X1 U14633 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11586), .B1(
        n11582), .B2(n11587), .ZN(n11591) );
  OAI21_X1 U14634 ( .B1(n18903), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11593), .ZN(n11592) );
  NOR2_X1 U14635 ( .A1(n11594), .A2(n11592), .ZN(n11590) );
  OAI21_X1 U14636 ( .B1(n11585), .B2(n11584), .A(n11591), .ZN(n11583) );
  AOI21_X1 U14637 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11587), .A(
        n11586), .ZN(n11588) );
  AOI21_X1 U14638 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18914), .A(
        n11588), .ZN(n11589) );
  INV_X1 U14639 ( .A(n11589), .ZN(n11595) );
  INV_X1 U14640 ( .A(n11592), .ZN(n11597) );
  XOR2_X1 U14641 ( .A(n11594), .B(n11593), .Z(n11596) );
  AOI21_X1 U14642 ( .B1(n11598), .B2(n11597), .A(n16750), .ZN(n18872) );
  INV_X1 U14643 ( .A(n13962), .ZN(n18473) );
  AOI211_X1 U14644 ( .C1(n18473), .C2(n18462), .A(n11600), .B(n11599), .ZN(
        n13956) );
  NAND2_X1 U14645 ( .A1(n11601), .A2(n18448), .ZN(n11602) );
  NOR2_X1 U14646 ( .A1(n13962), .A2(n11602), .ZN(n15889) );
  NAND2_X1 U14647 ( .A1(n13956), .A2(n15889), .ZN(n18873) );
  INV_X1 U14648 ( .A(n18873), .ZN(n11603) );
  INV_X1 U14649 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18931) );
  NAND2_X1 U14650 ( .A1(n19042), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18935) );
  NOR2_X2 U14651 ( .A1(n18448), .A2(n16753), .ZN(n18040) );
  NOR2_X1 U14652 ( .A1(n18012), .A2(n18040), .ZN(n17847) );
  INV_X1 U14653 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18109) );
  NAND2_X1 U14654 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18114) );
  INV_X1 U14655 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18221) );
  INV_X1 U14656 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18185) );
  NAND2_X1 U14657 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18184) );
  NOR3_X1 U14658 ( .A1(n18221), .A2(n18185), .A3(n18184), .ZN(n18171) );
  NAND2_X1 U14659 ( .A1(n18171), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16637) );
  INV_X1 U14660 ( .A(n16637), .ZN(n17801) );
  NAND2_X1 U14661 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17801), .ZN(
        n11727) );
  NAND2_X1 U14662 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18181) );
  INV_X1 U14663 ( .A(n18181), .ZN(n18218) );
  INV_X1 U14664 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18268) );
  NAND2_X1 U14665 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18303) );
  INV_X1 U14666 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18307) );
  NOR2_X1 U14667 ( .A1(n18303), .A2(n18307), .ZN(n17947) );
  NAND2_X1 U14668 ( .A1(n17947), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18287) );
  INV_X1 U14669 ( .A(n18287), .ZN(n17907) );
  NAND2_X1 U14670 ( .A1(n17907), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18263) );
  NOR2_X1 U14671 ( .A1(n18268), .A2(n18263), .ZN(n18248) );
  INV_X1 U14672 ( .A(n18248), .ZN(n18239) );
  INV_X1 U14673 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U14674 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11613) );
  INV_X1 U14675 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17469) );
  AOI22_X1 U14676 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14677 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11604) );
  OAI211_X1 U14678 ( .C1(n17447), .C2(n17469), .A(n11605), .B(n11604), .ZN(
        n11611) );
  AOI22_X1 U14679 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14680 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14681 ( .A1(n11665), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11607) );
  NAND2_X1 U14682 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11606) );
  NAND4_X1 U14683 ( .A1(n11609), .A2(n11608), .A3(n11607), .A4(n11606), .ZN(
        n11610) );
  AOI211_X1 U14684 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n11611), .B(n11610), .ZN(n11612) );
  OAI211_X1 U14685 ( .C1(n17453), .C2(n17227), .A(n11613), .B(n11612), .ZN(
        n11704) );
  AOI22_X1 U14686 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11623) );
  INV_X1 U14687 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17388) );
  AOI22_X1 U14688 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14689 ( .A1(n14033), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11614) );
  OAI211_X1 U14690 ( .C1(n17426), .C2(n17388), .A(n11615), .B(n11614), .ZN(
        n11621) );
  AOI22_X1 U14691 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11626), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14692 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14693 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11617) );
  NAND2_X1 U14694 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11616) );
  NAND4_X1 U14695 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n11620) );
  AOI211_X1 U14696 ( .C1(n11665), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n11621), .B(n11620), .ZN(n11622) );
  OAI211_X1 U14697 ( .C1(n17447), .C2(n17476), .A(n11623), .B(n11622), .ZN(
        n11703) );
  INV_X1 U14698 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17393) );
  AOI22_X1 U14699 ( .A1(n14033), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11631) );
  INV_X1 U14700 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U14701 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11624) );
  OAI21_X1 U14702 ( .B1(n17441), .B2(n17281), .A(n11624), .ZN(n11628) );
  AOI22_X1 U14703 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11625), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11627) );
  OAI211_X1 U14704 ( .C1(n17415), .C2(n17393), .A(n11631), .B(n11630), .ZN(
        n11635) );
  INV_X1 U14705 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14021) );
  AOI22_X1 U14706 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11632) );
  OAI21_X1 U14707 ( .B1(n10416), .B2(n14021), .A(n11632), .ZN(n11634) );
  INV_X1 U14708 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14709 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17410), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11643) );
  INV_X1 U14710 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U14711 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11636) );
  OAI21_X1 U14712 ( .B1(n17484), .B2(n11517), .A(n11636), .ZN(n11641) );
  INV_X1 U14713 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17412) );
  AOI22_X1 U14714 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n11637), .ZN(n11639) );
  AOI22_X1 U14715 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11461), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11638) );
  OAI211_X1 U14716 ( .C1(n17426), .C2(n17412), .A(n11639), .B(n11638), .ZN(
        n11640) );
  AOI211_X1 U14717 ( .C1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(n11665), .A(
        n11641), .B(n11640), .ZN(n11642) );
  OAI211_X1 U14718 ( .C1(n10412), .C2(n11644), .A(n11643), .B(n11642), .ZN(
        n11645) );
  AOI22_X1 U14719 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17394), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17396), .ZN(n11646) );
  OAI21_X1 U14720 ( .B1(n13990), .B2(n17453), .A(n11646), .ZN(n11648) );
  INV_X1 U14721 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14045) );
  AOI22_X1 U14722 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11650) );
  OAI21_X1 U14723 ( .B1(n10416), .B2(n14045), .A(n11650), .ZN(n11659) );
  INV_X1 U14724 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17371) );
  AOI22_X1 U14725 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11657) );
  INV_X1 U14726 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17246) );
  AOI22_X1 U14727 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11651) );
  OAI21_X1 U14728 ( .B1(n17441), .B2(n17246), .A(n11651), .ZN(n11655) );
  INV_X1 U14729 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17473) );
  AOI22_X1 U14730 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14731 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11652) );
  OAI211_X1 U14732 ( .C1(n17447), .C2(n17473), .A(n11653), .B(n11652), .ZN(
        n11654) );
  AOI211_X1 U14733 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n11655), .B(n11654), .ZN(n11656) );
  OAI211_X1 U14734 ( .C1(n10412), .C2(n17371), .A(n11657), .B(n11656), .ZN(
        n11658) );
  INV_X1 U14735 ( .A(n17625), .ZN(n11660) );
  XOR2_X1 U14736 ( .A(n17621), .B(n11683), .Z(n11680) );
  XNOR2_X1 U14737 ( .A(n17625), .B(n11661), .ZN(n11662) );
  NAND2_X1 U14738 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11662), .ZN(
        n11679) );
  XOR2_X1 U14739 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11662), .Z(
        n18058) );
  NAND2_X1 U14740 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11663), .ZN(
        n11674) );
  NAND2_X1 U14741 ( .A1(n11702), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11673) );
  INV_X1 U14742 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19044) );
  INV_X1 U14743 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17320) );
  AOI22_X1 U14744 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11664) );
  OAI21_X1 U14745 ( .B1(n10416), .B2(n17320), .A(n11664), .ZN(n11672) );
  INV_X1 U14746 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17435) );
  AOI22_X1 U14747 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11671) );
  INV_X1 U14748 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U14749 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11665), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11666) );
  OAI21_X1 U14750 ( .B1(n17415), .B2(n17452), .A(n11666), .ZN(n11670) );
  INV_X1 U14751 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14001) );
  AOI22_X1 U14752 ( .A1(n14033), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14753 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11668) );
  INV_X1 U14754 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19061) );
  NOR2_X1 U14755 ( .A1(n18102), .A2(n19061), .ZN(n18101) );
  NAND2_X1 U14756 ( .A1(n11674), .A2(n18079), .ZN(n11676) );
  XOR2_X1 U14757 ( .A(n17628), .B(n11712), .Z(n11677) );
  NAND2_X1 U14758 ( .A1(n11677), .A2(n11676), .ZN(n11678) );
  NAND2_X1 U14759 ( .A1(n11680), .A2(n11681), .ZN(n11682) );
  NAND2_X1 U14760 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18051), .ZN(
        n18050) );
  NAND2_X1 U14761 ( .A1(n11682), .A2(n18050), .ZN(n18030) );
  INV_X1 U14762 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18333) );
  INV_X1 U14763 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14764 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11685) );
  OAI21_X1 U14765 ( .B1(n11496), .B2(n11686), .A(n11685), .ZN(n11696) );
  INV_X1 U14766 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17464) );
  AOI22_X1 U14767 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11694) );
  INV_X1 U14768 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U14769 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11687) );
  OAI21_X1 U14770 ( .B1(n17258), .B2(n17164), .A(n11687), .ZN(n11692) );
  INV_X1 U14771 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14772 ( .A1(n17396), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14773 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11688) );
  OAI211_X1 U14774 ( .C1(n17426), .C2(n11690), .A(n11689), .B(n11688), .ZN(
        n11691) );
  AOI211_X1 U14775 ( .C1(n11665), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n11692), .B(n11691), .ZN(n11693) );
  OAI211_X1 U14776 ( .C1(n11517), .C2(n17464), .A(n11694), .B(n11693), .ZN(
        n11695) );
  XNOR2_X1 U14777 ( .A(n18333), .B(n11705), .ZN(n18038) );
  XOR2_X1 U14778 ( .A(n11698), .B(n18038), .Z(n18031) );
  NAND2_X1 U14779 ( .A1(n18030), .A2(n18031), .ZN(n18029) );
  XNOR2_X1 U14780 ( .A(n11705), .B(n11698), .ZN(n11697) );
  AND2_X2 U14781 ( .A1(n18029), .A2(n10415), .ZN(n17967) );
  NAND2_X1 U14782 ( .A1(n11700), .A2(n11699), .ZN(n11701) );
  NAND2_X1 U14783 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17794), .ZN(
        n17785) );
  NAND2_X1 U14784 ( .A1(n11711), .A2(n11703), .ZN(n11708) );
  NOR2_X1 U14785 ( .A1(n17625), .A2(n11708), .ZN(n11706) );
  NAND2_X1 U14786 ( .A1(n11706), .A2(n11704), .ZN(n18034) );
  NAND2_X1 U14787 ( .A1(n11705), .A2(n18036), .ZN(n11721) );
  NOR2_X1 U14788 ( .A1(n11721), .A2(n11739), .ZN(n11726) );
  INV_X1 U14789 ( .A(n11726), .ZN(n11722) );
  XOR2_X1 U14790 ( .A(n18036), .B(n11705), .Z(n11720) );
  XNOR2_X1 U14791 ( .A(n11706), .B(n17621), .ZN(n11707) );
  NAND2_X1 U14792 ( .A1(n11707), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11719) );
  XOR2_X1 U14793 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11707), .Z(
        n18046) );
  XOR2_X1 U14794 ( .A(n11708), .B(n17625), .Z(n11709) );
  NAND2_X1 U14795 ( .A1(n11709), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11718) );
  XOR2_X1 U14796 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11709), .Z(
        n18064) );
  XNOR2_X1 U14797 ( .A(n11711), .B(n17628), .ZN(n11710) );
  NAND2_X1 U14798 ( .A1(n11710), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11717) );
  INV_X1 U14799 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15894) );
  XNOR2_X1 U14800 ( .A(n15894), .B(n11710), .ZN(n18073) );
  OAI21_X1 U14801 ( .B1(n18102), .B2(n11712), .A(n11711), .ZN(n11715) );
  NAND2_X1 U14802 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11715), .ZN(
        n11716) );
  INV_X1 U14803 ( .A(n18102), .ZN(n18092) );
  AOI21_X1 U14804 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17637), .A(
        n18092), .ZN(n11714) );
  NOR2_X1 U14805 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17637), .ZN(
        n11713) );
  AOI221_X1 U14806 ( .B1(n18092), .B2(n17637), .C1(n11714), .C2(n19061), .A(
        n11713), .ZN(n18085) );
  XOR2_X1 U14807 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11715), .Z(
        n18084) );
  NAND2_X1 U14808 ( .A1(n18085), .A2(n18084), .ZN(n18083) );
  NAND2_X1 U14809 ( .A1(n11716), .A2(n18083), .ZN(n18072) );
  NAND2_X1 U14810 ( .A1(n18073), .A2(n18072), .ZN(n18071) );
  NAND2_X1 U14811 ( .A1(n11717), .A2(n18071), .ZN(n18063) );
  NAND2_X1 U14812 ( .A1(n18064), .A2(n18063), .ZN(n18062) );
  XNOR2_X1 U14813 ( .A(n11739), .B(n11721), .ZN(n18020) );
  NAND2_X1 U14814 ( .A1(n18019), .A2(n18020), .ZN(n18018) );
  NAND2_X1 U14815 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18018), .ZN(
        n11725) );
  NOR2_X1 U14816 ( .A1(n18019), .A2(n18020), .ZN(n11724) );
  NOR2_X1 U14817 ( .A1(n11726), .A2(n11725), .ZN(n11723) );
  AOI211_X1 U14818 ( .C1(n11726), .C2(n11725), .A(n11724), .B(n11723), .ZN(
        n18004) );
  INV_X1 U14819 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18337) );
  NOR2_X2 U14820 ( .A1(n18268), .A2(n17928), .ZN(n17927) );
  OAI22_X1 U14821 ( .A1(n18116), .A2(n17943), .B1(n18117), .B2(n18108), .ZN(
        n17771) );
  NOR2_X1 U14822 ( .A1(n18109), .A2(n17771), .ZN(n17756) );
  INV_X1 U14823 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16640) );
  INV_X1 U14824 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17811) );
  INV_X1 U14825 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18151) );
  INV_X1 U14826 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18135) );
  NOR3_X1 U14827 ( .A1(n17811), .A2(n18151), .A3(n18135), .ZN(n18130) );
  NAND2_X1 U14828 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18130), .ZN(
        n18110) );
  NOR2_X1 U14829 ( .A1(n18109), .A2(n18110), .ZN(n16603) );
  INV_X1 U14830 ( .A(n16603), .ZN(n16638) );
  NAND2_X1 U14831 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18248), .ZN(
        n18213) );
  NOR2_X1 U14832 ( .A1(n18181), .A2(n18213), .ZN(n17797) );
  INV_X1 U14833 ( .A(n17797), .ZN(n15898) );
  NOR2_X1 U14834 ( .A1(n16637), .A2(n15898), .ZN(n15905) );
  NAND2_X1 U14835 ( .A1(n15905), .A2(n17984), .ZN(n17770) );
  INV_X1 U14836 ( .A(n11727), .ZN(n18144) );
  NAND2_X1 U14837 ( .A1(n18221), .A2(n17969), .ZN(n17867) );
  NOR2_X1 U14838 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17867), .ZN(
        n11728) );
  INV_X1 U14839 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18201) );
  NAND2_X1 U14840 ( .A1(n11728), .A2(n18201), .ZN(n17831) );
  NOR2_X1 U14841 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17831), .ZN(
        n17815) );
  INV_X1 U14842 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18173) );
  NAND3_X1 U14843 ( .A1(n17815), .A2(n17811), .A3(n18173), .ZN(n11733) );
  NOR2_X2 U14844 ( .A1(n11729), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17968) );
  INV_X1 U14845 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18328) );
  INV_X1 U14846 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18315) );
  NAND2_X1 U14847 ( .A1(n18328), .A2(n18315), .ZN(n17982) );
  INV_X1 U14848 ( .A(n17982), .ZN(n17970) );
  NAND3_X1 U14849 ( .A1(n17968), .A2(n17970), .A3(n18307), .ZN(n17931) );
  NOR2_X2 U14850 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17931), .ZN(
        n17908) );
  INV_X1 U14851 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18294) );
  NAND2_X1 U14852 ( .A1(n17908), .A2(n10414), .ZN(n11731) );
  NAND2_X2 U14853 ( .A1(n11731), .A2(n17969), .ZN(n17896) );
  INV_X1 U14854 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18233) );
  NAND2_X1 U14855 ( .A1(n17796), .A2(n18151), .ZN(n17795) );
  NAND2_X1 U14856 ( .A1(n17969), .A2(n17795), .ZN(n17775) );
  NOR2_X4 U14857 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11737), .ZN(
        n16653) );
  INV_X1 U14858 ( .A(n16653), .ZN(n11738) );
  AOI22_X1 U14859 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17969), .B1(
        n18002), .B2(n16640), .ZN(n16652) );
  AOI211_X1 U14860 ( .C1(n9866), .C2(n16652), .A(n16642), .B(n18015), .ZN(
        n11740) );
  INV_X1 U14861 ( .A(n11740), .ZN(n11750) );
  OAI21_X1 U14862 ( .B1(n19042), .B2(n18931), .A(n19034), .ZN(n19078) );
  INV_X1 U14863 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19083) );
  NOR2_X1 U14864 ( .A1(n19042), .A2(n19083), .ZN(n17935) );
  INV_X1 U14865 ( .A(n17935), .ZN(n18060) );
  INV_X1 U14866 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16812) );
  INV_X1 U14867 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18097) );
  NAND2_X1 U14868 ( .A1(n17962), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17934) );
  NAND2_X1 U14869 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17076) );
  NAND2_X1 U14870 ( .A1(n18061), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18048) );
  INV_X1 U14871 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16927) );
  NAND3_X1 U14872 ( .A1(n17857), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17842) );
  INV_X1 U14873 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17841) );
  NOR2_X2 U14874 ( .A1(n17842), .A2(n17841), .ZN(n17820) );
  INV_X1 U14875 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17780) );
  NAND2_X1 U14876 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11743) );
  INV_X1 U14877 ( .A(n11743), .ZN(n17778) );
  INV_X1 U14878 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17758) );
  OR3_X1 U14879 ( .A1(n18097), .A2(n12155), .A3(n17758), .ZN(n16771) );
  INV_X1 U14880 ( .A(n16584), .ZN(n16612) );
  AOI21_X1 U14881 ( .B1(n16812), .B2(n16771), .A(n16587), .ZN(n16806) );
  INV_X1 U14882 ( .A(n16806), .ZN(n11747) );
  INV_X1 U14883 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n13960) );
  NAND2_X1 U14884 ( .A1(n13960), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18104) );
  INV_X1 U14885 ( .A(n17819), .ZN(n16585) );
  NAND2_X1 U14886 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17820), .ZN(
        n12159) );
  NOR2_X1 U14887 ( .A1(n17821), .A2(n12159), .ZN(n17779) );
  NAND2_X1 U14888 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17779), .ZN(
        n12162) );
  NOR2_X1 U14889 ( .A1(n11743), .A2(n12162), .ZN(n12154) );
  OAI21_X1 U14890 ( .B1(n12154), .B2(n18104), .A(n18103), .ZN(n11742) );
  AOI21_X1 U14891 ( .B1(n17935), .B2(n12155), .A(n11742), .ZN(n17766) );
  OAI21_X1 U14892 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n16585), .A(
        n17766), .ZN(n17751) );
  AOI221_X1 U14893 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19042), .C1(n18931), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n19058), .ZN(n18440) );
  NAND3_X1 U14894 ( .A1(n19034), .A2(n18931), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18599) );
  AOI21_X1 U14895 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17819), .A(
        n18815), .ZN(n17891) );
  INV_X1 U14896 ( .A(n17891), .ZN(n17949) );
  NAND2_X1 U14897 ( .A1(n9927), .A2(n17949), .ZN(n17791) );
  NOR3_X1 U14898 ( .A1(n11743), .A2(n10273), .A3(n17791), .ZN(n17759) );
  XOR2_X1 U14899 ( .A(n16812), .B(n17758), .Z(n11744) );
  AOI22_X1 U14900 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17751), .B1(
        n17759), .B2(n11744), .ZN(n11746) );
  NOR2_X1 U14901 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19060) );
  INV_X2 U14902 ( .A(n18426), .ZN(n18308) );
  NAND2_X1 U14903 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18308), .ZN(n11745) );
  OAI211_X1 U14904 ( .C1(n17938), .C2(n11747), .A(n11746), .B(n11745), .ZN(
        n11748) );
  INV_X1 U14905 ( .A(n11748), .ZN(n11749) );
  NAND4_X1 U14906 ( .A1(n10427), .A2(n10419), .A3(n11750), .A4(n11749), .ZN(
        P3_U2802) );
  NAND2_X1 U14907 ( .A1(n10495), .A2(n16562), .ZN(n11753) );
  INV_X1 U14908 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n13298) );
  NAND2_X1 U14909 ( .A1(n11753), .A2(n13298), .ZN(n11774) );
  INV_X1 U14910 ( .A(n20037), .ZN(n20042) );
  NAND2_X1 U14911 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13300) );
  NAND2_X1 U14912 ( .A1(n13300), .A2(n20056), .ZN(n11754) );
  NOR2_X1 U14913 ( .A1(n20056), .A2(n20064), .ZN(n13695) );
  NAND2_X1 U14914 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13695), .ZN(
        n11770) );
  NAND2_X1 U14915 ( .A1(n11754), .A2(n11770), .ZN(n19553) );
  NOR2_X1 U14916 ( .A1(n20042), .A2(n19553), .ZN(n11755) );
  AOI21_X1 U14917 ( .B1(n11774), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11755), .ZN(n11756) );
  NOR2_X1 U14918 ( .A1(n10495), .A2(n11751), .ZN(n12629) );
  OAI21_X1 U14919 ( .B1(n11758), .B2(n11757), .A(n11768), .ZN(n11759) );
  AOI22_X1 U14920 ( .A1(n11774), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20037), .B2(n20074), .ZN(n11760) );
  NAND2_X1 U14921 ( .A1(n11774), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11763) );
  NAND2_X1 U14922 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20074), .ZN(
        n19729) );
  NAND2_X1 U14923 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20064), .ZN(
        n19698) );
  NAND2_X1 U14924 ( .A1(n19729), .A2(n19698), .ZN(n19552) );
  NAND2_X1 U14925 ( .A1(n20037), .A2(n19552), .ZN(n19732) );
  NAND2_X1 U14926 ( .A1(n11763), .A2(n19732), .ZN(n11764) );
  INV_X1 U14927 ( .A(n11765), .ZN(n11766) );
  NOR2_X1 U14928 ( .A1(n15846), .A2(n11766), .ZN(n11767) );
  INV_X1 U14929 ( .A(n11768), .ZN(n11769) );
  AOI21_X1 U14930 ( .B1(n12597), .B2(n12598), .A(n11769), .ZN(n12713) );
  INV_X1 U14931 ( .A(n11770), .ZN(n11771) );
  NAND2_X1 U14932 ( .A1(n11771), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19889) );
  OAI211_X1 U14933 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n11771), .A(
        n19889), .B(n20037), .ZN(n11772) );
  INV_X1 U14934 ( .A(n11772), .ZN(n11773) );
  AOI21_X1 U14935 ( .B1(n11774), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11773), .ZN(n11775) );
  NAND2_X1 U14936 ( .A1(n11776), .A2(n11775), .ZN(n11779) );
  AND2_X1 U14937 ( .A1(n11947), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11777) );
  NAND2_X1 U14938 ( .A1(n11779), .A2(n11777), .ZN(n12694) );
  OAI21_X1 U14939 ( .B1(n11779), .B2(n11777), .A(n12694), .ZN(n12714) );
  NAND2_X1 U14940 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10495), .ZN(
        n11778) );
  INV_X1 U14941 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11780) );
  NAND2_X1 U14942 ( .A1(n12834), .A2(n12837), .ZN(n12835) );
  AOI22_X1 U14943 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U14944 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11882), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U14945 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11884), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14946 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11786) );
  NAND4_X1 U14947 ( .A1(n11789), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n11795) );
  AOI22_X1 U14948 ( .A1(n10729), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14949 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14950 ( .A1(n10798), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U14951 ( .A1(n12869), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11790) );
  NAND4_X1 U14952 ( .A1(n11793), .A2(n11792), .A3(n11791), .A4(n11790), .ZN(
        n11794) );
  NOR2_X1 U14953 ( .A1(n11795), .A2(n11794), .ZN(n13747) );
  AOI22_X1 U14954 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11818), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14955 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n11882), .ZN(n11798) );
  AOI22_X1 U14956 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n11884), .ZN(n11797) );
  AOI22_X1 U14957 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11796) );
  NAND4_X1 U14958 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11805) );
  AOI22_X1 U14959 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10729), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U14960 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U14961 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10730), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U14962 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12869), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11800) );
  NAND4_X1 U14963 ( .A1(n11803), .A2(n11802), .A3(n11801), .A4(n11800), .ZN(
        n11804) );
  AOI22_X1 U14964 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n11818), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U14965 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n11882), .ZN(n11808) );
  AOI22_X1 U14966 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__2__SCAN_IN), .B2(n11884), .ZN(n11807) );
  AOI22_X1 U14967 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11806) );
  NAND4_X1 U14968 ( .A1(n11809), .A2(n11808), .A3(n11807), .A4(n11806), .ZN(
        n11815) );
  AOI22_X1 U14969 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10729), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U14970 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U14971 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10730), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U14972 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12869), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11810) );
  NAND4_X1 U14973 ( .A1(n11813), .A2(n11812), .A3(n11811), .A4(n11810), .ZN(
        n11814) );
  NOR2_X1 U14974 ( .A1(n11815), .A2(n11814), .ZN(n13848) );
  INV_X1 U14975 ( .A(n11816), .ZN(n11817) );
  NOR2_X1 U14976 ( .A1(n11817), .A2(n11965), .ZN(n11823) );
  INV_X1 U14977 ( .A(n11818), .ZN(n11821) );
  INV_X1 U14978 ( .A(n11832), .ZN(n11820) );
  OAI22_X1 U14979 ( .A1(n10661), .A2(n11821), .B1(n11820), .B2(n11819), .ZN(
        n11822) );
  AOI211_X1 U14980 ( .C1(n11882), .C2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n11823), .B(n11822), .ZN(n11831) );
  AOI22_X1 U14981 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__3__SCAN_IN), .B2(n11884), .ZN(n11830) );
  AOI22_X1 U14982 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14983 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10729), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U14984 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U14985 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10730), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14986 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12869), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11824) );
  AND4_X1 U14987 ( .A1(n11827), .A2(n11826), .A3(n11825), .A4(n11824), .ZN(
        n11828) );
  NAND4_X1 U14988 ( .A1(n11831), .A2(n11830), .A3(n11829), .A4(n11828), .ZN(
        n13892) );
  AOI22_X1 U14989 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11818), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U14990 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n11882), .ZN(n11835) );
  AOI22_X1 U14991 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__4__SCAN_IN), .B2(n11884), .ZN(n11834) );
  AOI22_X1 U14992 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11833) );
  NAND4_X1 U14993 ( .A1(n11836), .A2(n11835), .A3(n11834), .A4(n11833), .ZN(
        n11842) );
  AOI22_X1 U14994 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10729), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U14995 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U14996 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10730), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14997 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12869), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11837) );
  NAND4_X1 U14998 ( .A1(n11840), .A2(n11839), .A3(n11838), .A4(n11837), .ZN(
        n11841) );
  NOR2_X1 U14999 ( .A1(n11842), .A2(n11841), .ZN(n15345) );
  AOI22_X1 U15000 ( .A1(n11832), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11818), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U15001 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11882), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U15002 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11884), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U15003 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11843) );
  NAND4_X1 U15004 ( .A1(n11846), .A2(n11845), .A3(n11844), .A4(n11843), .ZN(
        n11852) );
  AOI22_X1 U15005 ( .A1(n10729), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U15006 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U15007 ( .A1(n10798), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10730), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U15008 ( .A1(n12869), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11847) );
  NAND4_X1 U15009 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11851) );
  OR2_X1 U15010 ( .A1(n11852), .A2(n11851), .ZN(n15343) );
  NAND2_X1 U15011 ( .A1(n15342), .A2(n15343), .ZN(n15332) );
  AOI22_X1 U15012 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n11818), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U15013 ( .A1(n11816), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n11882), .ZN(n11855) );
  AOI22_X1 U15014 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11884), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U15015 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10704), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11853) );
  NAND4_X1 U15016 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(
        n11862) );
  AOI22_X1 U15017 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10729), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U15018 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U15019 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10730), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U15020 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12869), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11857) );
  NAND4_X1 U15021 ( .A1(n11860), .A2(n11859), .A3(n11858), .A4(n11857), .ZN(
        n11861) );
  NOR2_X1 U15022 ( .A1(n11862), .A2(n11861), .ZN(n15334) );
  INV_X1 U15023 ( .A(n12064), .ZN(n12039) );
  INV_X1 U15024 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n19600) );
  INV_X1 U15025 ( .A(n12063), .ZN(n12037) );
  INV_X1 U15026 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11863) );
  OAI22_X1 U15027 ( .A1(n12039), .A2(n19600), .B1(n12037), .B2(n11863), .ZN(
        n11866) );
  INV_X1 U15028 ( .A(n12066), .ZN(n12042) );
  INV_X1 U15029 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11864) );
  INV_X1 U15030 ( .A(n12065), .ZN(n12887) );
  INV_X1 U15031 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n19533) );
  OAI22_X1 U15032 ( .A1(n12042), .A2(n11864), .B1(n12887), .B2(n19533), .ZN(
        n11865) );
  NOR2_X1 U15033 ( .A1(n11866), .A2(n11865), .ZN(n11871) );
  AOI22_X1 U15034 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U15035 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11869) );
  XNOR2_X1 U15036 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12055) );
  NAND4_X1 U15037 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n12055), .ZN(
        n11881) );
  INV_X1 U15038 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13133) );
  INV_X1 U15039 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11872) );
  OAI22_X1 U15040 ( .A1(n12039), .A2(n13133), .B1(n12037), .B2(n11872), .ZN(
        n11876) );
  INV_X1 U15041 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11874) );
  INV_X1 U15042 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11873) );
  OAI22_X1 U15043 ( .A1(n12042), .A2(n11874), .B1(n12887), .B2(n11873), .ZN(
        n11875) );
  NOR2_X1 U15044 ( .A1(n11876), .A2(n11875), .ZN(n11879) );
  INV_X1 U15045 ( .A(n12055), .ZN(n12061) );
  AOI22_X1 U15046 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U15047 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11877) );
  NAND4_X1 U15048 ( .A1(n11879), .A2(n12061), .A3(n11878), .A4(n11877), .ZN(
        n11880) );
  AND2_X1 U15049 ( .A1(n11881), .A2(n11880), .ZN(n11921) );
  NAND2_X1 U15050 ( .A1(n11259), .A2(n11921), .ZN(n11896) );
  AOI22_X1 U15051 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11818), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U15052 ( .A1(n11883), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n11882), .ZN(n11887) );
  AOI22_X1 U15053 ( .A1(n11305), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n11816), .ZN(n11886) );
  AOI22_X1 U15054 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10704), .B1(
        n11884), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11885) );
  NAND4_X1 U15055 ( .A1(n11888), .A2(n11887), .A3(n11886), .A4(n11885), .ZN(
        n11895) );
  AOI22_X1 U15056 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10729), .B1(
        n10774), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U15057 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11889), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U15058 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12869), .B1(
        n10798), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U15059 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10730), .B1(
        n10776), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11890) );
  NAND4_X1 U15060 ( .A1(n11893), .A2(n11892), .A3(n11891), .A4(n11890), .ZN(
        n11894) );
  OR2_X1 U15061 ( .A1(n11895), .A2(n11894), .ZN(n11918) );
  XNOR2_X1 U15062 ( .A(n11896), .B(n11918), .ZN(n11924) );
  NAND2_X1 U15063 ( .A1(n13682), .A2(n11921), .ZN(n15329) );
  OAI22_X1 U15064 ( .A1(n12039), .A2(n11899), .B1(n12037), .B2(n11898), .ZN(
        n11903) );
  OAI22_X1 U15065 ( .A1(n12042), .A2(n11901), .B1(n12887), .B2(n11900), .ZN(
        n11902) );
  NOR2_X1 U15066 ( .A1(n11903), .A2(n11902), .ZN(n11906) );
  AOI22_X1 U15067 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U15068 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11904) );
  NAND4_X1 U15069 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n12055), .ZN(
        n11917) );
  OAI22_X1 U15070 ( .A1(n12039), .A2(n11908), .B1(n12037), .B2(n11907), .ZN(
        n11912) );
  OAI22_X1 U15071 ( .A1(n12042), .A2(n11910), .B1(n12887), .B2(n11909), .ZN(
        n11911) );
  NOR2_X1 U15072 ( .A1(n11912), .A2(n11911), .ZN(n11915) );
  AOI22_X1 U15073 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U15074 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11913) );
  NAND4_X1 U15075 ( .A1(n11915), .A2(n12061), .A3(n11914), .A4(n11913), .ZN(
        n11916) );
  NAND2_X1 U15076 ( .A1(n11917), .A2(n11916), .ZN(n11925) );
  NAND2_X1 U15077 ( .A1(n11918), .A2(n11921), .ZN(n11926) );
  XOR2_X1 U15078 ( .A(n11925), .B(n11926), .Z(n11919) );
  NAND2_X1 U15079 ( .A1(n11919), .A2(n11947), .ZN(n15318) );
  INV_X1 U15080 ( .A(n11925), .ZN(n11920) );
  NAND2_X1 U15081 ( .A1(n13682), .A2(n11920), .ZN(n15320) );
  INV_X1 U15082 ( .A(n11921), .ZN(n11922) );
  NOR2_X1 U15083 ( .A1(n15320), .A2(n11922), .ZN(n11923) );
  NOR2_X1 U15084 ( .A1(n11926), .A2(n11925), .ZN(n11948) );
  INV_X1 U15085 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11928) );
  INV_X1 U15086 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11927) );
  OAI22_X1 U15087 ( .A1(n12039), .A2(n11928), .B1(n12037), .B2(n11927), .ZN(
        n11932) );
  INV_X1 U15088 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11930) );
  INV_X1 U15089 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11929) );
  OAI22_X1 U15090 ( .A1(n12042), .A2(n11930), .B1(n12887), .B2(n11929), .ZN(
        n11931) );
  NOR2_X1 U15091 ( .A1(n11932), .A2(n11931), .ZN(n11935) );
  AOI22_X1 U15092 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U15093 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11933) );
  NAND4_X1 U15094 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n12055), .ZN(
        n11946) );
  INV_X1 U15095 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11937) );
  INV_X1 U15096 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11936) );
  OAI22_X1 U15097 ( .A1(n12039), .A2(n11937), .B1(n12037), .B2(n11936), .ZN(
        n11941) );
  INV_X1 U15098 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11939) );
  INV_X1 U15099 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11938) );
  OAI22_X1 U15100 ( .A1(n12042), .A2(n11939), .B1(n12887), .B2(n11938), .ZN(
        n11940) );
  NOR2_X1 U15101 ( .A1(n11941), .A2(n11940), .ZN(n11944) );
  AOI22_X1 U15102 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11943) );
  AOI22_X1 U15103 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11942) );
  NAND4_X1 U15104 ( .A1(n11944), .A2(n12061), .A3(n11943), .A4(n11942), .ZN(
        n11945) );
  AND2_X1 U15105 ( .A1(n11946), .A2(n11945), .ZN(n11950) );
  NAND2_X1 U15106 ( .A1(n11948), .A2(n11950), .ZN(n11975) );
  OAI211_X1 U15107 ( .C1(n11948), .C2(n11950), .A(n11975), .B(n11947), .ZN(
        n11953) );
  INV_X1 U15108 ( .A(n11953), .ZN(n11949) );
  INV_X1 U15109 ( .A(n11950), .ZN(n11951) );
  NOR2_X1 U15110 ( .A1(n11259), .A2(n11951), .ZN(n15311) );
  OAI22_X1 U15111 ( .A1(n12039), .A2(n11956), .B1(n12037), .B2(n11955), .ZN(
        n11960) );
  OAI22_X1 U15112 ( .A1(n12042), .A2(n11958), .B1(n12887), .B2(n11957), .ZN(
        n11959) );
  NOR2_X1 U15113 ( .A1(n11960), .A2(n11959), .ZN(n11963) );
  AOI22_X1 U15114 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15115 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11961) );
  NAND4_X1 U15116 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n12055), .ZN(
        n11974) );
  OAI22_X1 U15117 ( .A1(n12039), .A2(n11965), .B1(n12037), .B2(n11964), .ZN(
        n11969) );
  OAI22_X1 U15118 ( .A1(n12042), .A2(n11967), .B1(n12887), .B2(n11966), .ZN(
        n11968) );
  NOR2_X1 U15119 ( .A1(n11969), .A2(n11968), .ZN(n11972) );
  AOI22_X1 U15120 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11971) );
  AOI22_X1 U15121 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11970) );
  NAND4_X1 U15122 ( .A1(n11972), .A2(n12061), .A3(n11971), .A4(n11970), .ZN(
        n11973) );
  NAND2_X1 U15123 ( .A1(n11974), .A2(n11973), .ZN(n11977) );
  AOI21_X1 U15124 ( .B1(n11975), .B2(n11977), .A(n12001), .ZN(n11976) );
  OR2_X1 U15125 ( .A1(n11975), .A2(n11977), .ZN(n12002) );
  NAND2_X1 U15126 ( .A1(n11976), .A2(n12002), .ZN(n11979) );
  NOR2_X1 U15127 ( .A1(n11259), .A2(n11977), .ZN(n15303) );
  INV_X1 U15128 ( .A(n11978), .ZN(n11980) );
  INV_X1 U15129 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11982) );
  INV_X1 U15130 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11981) );
  OAI22_X1 U15131 ( .A1(n12039), .A2(n11982), .B1(n12037), .B2(n11981), .ZN(
        n11986) );
  INV_X1 U15132 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11984) );
  INV_X1 U15133 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11983) );
  OAI22_X1 U15134 ( .A1(n12042), .A2(n11984), .B1(n12887), .B2(n11983), .ZN(
        n11985) );
  NOR2_X1 U15135 ( .A1(n11986), .A2(n11985), .ZN(n11989) );
  AOI22_X1 U15136 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15137 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11987) );
  NAND4_X1 U15138 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n12055), .ZN(
        n12000) );
  INV_X1 U15139 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11991) );
  INV_X1 U15140 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11990) );
  OAI22_X1 U15141 ( .A1(n12039), .A2(n11991), .B1(n12037), .B2(n11990), .ZN(
        n11995) );
  INV_X1 U15142 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11993) );
  INV_X1 U15143 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11992) );
  OAI22_X1 U15144 ( .A1(n12042), .A2(n11993), .B1(n12887), .B2(n11992), .ZN(
        n11994) );
  NOR2_X1 U15145 ( .A1(n11995), .A2(n11994), .ZN(n11998) );
  AOI22_X1 U15146 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U15147 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11996) );
  NAND4_X1 U15148 ( .A1(n11998), .A2(n12061), .A3(n11997), .A4(n11996), .ZN(
        n11999) );
  NAND2_X1 U15149 ( .A1(n12000), .A2(n11999), .ZN(n12005) );
  NOR2_X1 U15150 ( .A1(n12002), .A2(n12005), .ZN(n12026) );
  NOR2_X1 U15151 ( .A1(n11259), .A2(n12005), .ZN(n15295) );
  OAI22_X1 U15152 ( .A1(n12039), .A2(n12007), .B1(n12037), .B2(n12006), .ZN(
        n12010) );
  OAI22_X1 U15153 ( .A1(n12042), .A2(n12008), .B1(n12887), .B2(n13316), .ZN(
        n12009) );
  NOR2_X1 U15154 ( .A1(n12010), .A2(n12009), .ZN(n12013) );
  AOI22_X1 U15155 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15156 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12011) );
  NAND4_X1 U15157 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n12055), .ZN(
        n12024) );
  OAI22_X1 U15158 ( .A1(n12039), .A2(n12015), .B1(n12037), .B2(n12014), .ZN(
        n12019) );
  OAI22_X1 U15159 ( .A1(n12042), .A2(n12017), .B1(n12887), .B2(n12016), .ZN(
        n12018) );
  NOR2_X1 U15160 ( .A1(n12019), .A2(n12018), .ZN(n12022) );
  AOI22_X1 U15161 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15162 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12020) );
  NAND4_X1 U15163 ( .A1(n12022), .A2(n12061), .A3(n12021), .A4(n12020), .ZN(
        n12023) );
  INV_X1 U15164 ( .A(n12026), .ZN(n15287) );
  NAND2_X1 U15165 ( .A1(n11259), .A2(n15290), .ZN(n12027) );
  NOR2_X1 U15166 ( .A1(n15287), .A2(n12027), .ZN(n12051) );
  OAI22_X1 U15167 ( .A1(n10856), .A2(n12039), .B1(n12037), .B2(n12028), .ZN(
        n12032) );
  OAI22_X1 U15168 ( .A1(n12042), .A2(n12030), .B1(n12887), .B2(n12029), .ZN(
        n12031) );
  NOR2_X1 U15169 ( .A1(n12032), .A2(n12031), .ZN(n12035) );
  AOI22_X1 U15170 ( .A1(n12058), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15171 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10676), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12033) );
  NAND4_X1 U15172 ( .A1(n12035), .A2(n12034), .A3(n12033), .A4(n12055), .ZN(
        n12049) );
  OAI22_X1 U15173 ( .A1(n12039), .A2(n12038), .B1(n12037), .B2(n12036), .ZN(
        n12044) );
  OAI22_X1 U15174 ( .A1(n12042), .A2(n12041), .B1(n12887), .B2(n12040), .ZN(
        n12043) );
  NOR2_X1 U15175 ( .A1(n12044), .A2(n12043), .ZN(n12047) );
  AOI22_X1 U15176 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15177 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12045) );
  NAND4_X1 U15178 ( .A1(n12047), .A2(n12061), .A3(n12046), .A4(n12045), .ZN(
        n12048) );
  AND2_X1 U15179 ( .A1(n12049), .A2(n12048), .ZN(n12050) );
  NAND2_X1 U15180 ( .A1(n12051), .A2(n12050), .ZN(n12052) );
  OAI21_X1 U15181 ( .B1(n12051), .B2(n12050), .A(n12052), .ZN(n15285) );
  AOI22_X1 U15182 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12063), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15183 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12053) );
  NAND2_X1 U15184 ( .A1(n12054), .A2(n12053), .ZN(n12072) );
  AOI22_X1 U15185 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15186 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12056) );
  NAND3_X1 U15187 ( .A1(n12057), .A2(n12056), .A3(n12055), .ZN(n12071) );
  AOI22_X1 U15188 ( .A1(n9802), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12058), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15189 ( .A1(n11868), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12059), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12060) );
  NAND3_X1 U15190 ( .A1(n12062), .A2(n12061), .A3(n12060), .ZN(n12070) );
  AOI22_X1 U15191 ( .A1(n12064), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12063), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15192 ( .A1(n12066), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12065), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12067) );
  NAND2_X1 U15193 ( .A1(n12068), .A2(n12067), .ZN(n12069) );
  OAI22_X1 U15194 ( .A1(n12072), .A2(n12071), .B1(n12070), .B2(n12069), .ZN(
        n12073) );
  AND2_X1 U15195 ( .A1(n11116), .A2(n19937), .ZN(n12178) );
  AND2_X1 U15196 ( .A1(n11447), .A2(n12178), .ZN(n12074) );
  NAND2_X1 U15197 ( .A1(n12077), .A2(n12076), .ZN(n12078) );
  NAND2_X1 U15198 ( .A1(n12124), .A2(n19361), .ZN(n12101) );
  NAND2_X1 U15199 ( .A1(n11276), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15200 ( .A1(n11440), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12080), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12081) );
  NAND2_X1 U15201 ( .A1(n12082), .A2(n12081), .ZN(n14477) );
  XNOR2_X1 U15202 ( .A(n14476), .B(n14477), .ZN(n16296) );
  NOR2_X2 U15203 ( .A1(n19359), .A2(n12096), .ZN(n19360) );
  AOI22_X1 U15204 ( .A1(n16296), .A2(n19360), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19359), .ZN(n12100) );
  NOR2_X2 U15205 ( .A1(n19359), .A2(n12083), .ZN(n16381) );
  NOR4_X1 U15206 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12087) );
  NOR4_X1 U15207 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12086) );
  NOR4_X1 U15208 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12085) );
  NOR4_X1 U15209 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12084) );
  NAND4_X1 U15210 ( .A1(n12087), .A2(n12086), .A3(n12085), .A4(n12084), .ZN(
        n12092) );
  NOR4_X1 U15211 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12090) );
  NOR4_X1 U15212 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12089) );
  NOR4_X1 U15213 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12088) );
  INV_X1 U15214 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19962) );
  NAND4_X1 U15215 ( .A1(n12090), .A2(n12089), .A3(n12088), .A4(n19962), .ZN(
        n12091) );
  OAI21_X1 U15216 ( .B1(n12092), .B2(n12091), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12093) );
  INV_X1 U15217 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16677) );
  OR2_X1 U15218 ( .A1(n13097), .A2(n16677), .ZN(n12095) );
  NAND2_X1 U15219 ( .A1(n13097), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12094) );
  NAND2_X1 U15220 ( .A1(n12095), .A2(n12094), .ZN(n19310) );
  NAND2_X1 U15221 ( .A1(n16381), .A2(n19310), .ZN(n12099) );
  AND2_X1 U15222 ( .A1(n12096), .A2(n10495), .ZN(n12097) );
  NAND2_X1 U15223 ( .A1(n19333), .A2(n12097), .ZN(n13054) );
  NOR2_X2 U15224 ( .A1(n13054), .A2(n13098), .ZN(n19302) );
  NOR2_X2 U15225 ( .A1(n13054), .A2(n13097), .ZN(n19304) );
  AOI22_X1 U15226 ( .A1(n19302), .A2(BUF2_REG_30__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12098) );
  NAND2_X1 U15227 ( .A1(n12101), .A2(n10428), .ZN(P2_U2889) );
  NAND2_X1 U15228 ( .A1(n15477), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15478) );
  OAI21_X1 U15229 ( .B1(n15489), .B2(n10340), .A(n12105), .ZN(n12106) );
  NAND2_X1 U15230 ( .A1(n15478), .A2(n12106), .ZN(n12109) );
  XNOR2_X1 U15231 ( .A(n12107), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12108) );
  XNOR2_X1 U15232 ( .A(n12109), .B(n12108), .ZN(n15467) );
  NAND2_X1 U15233 ( .A1(n15467), .A2(n19414), .ZN(n12123) );
  OR2_X1 U15234 ( .A1(n15376), .A2(n12110), .ZN(n12111) );
  INV_X1 U15235 ( .A(n12113), .ZN(n12114) );
  NAND2_X1 U15236 ( .A1(n19404), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15471) );
  AOI21_X1 U15237 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n12116), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12117) );
  NOR2_X1 U15238 ( .A1(n12118), .A2(n12117), .ZN(n12119) );
  INV_X1 U15239 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12120) );
  NOR2_X1 U15240 ( .A1(n15492), .A2(n12120), .ZN(n12121) );
  OAI21_X1 U15241 ( .B1(n12121), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15449), .ZN(n15475) );
  NOR2_X1 U15242 ( .A1(n12901), .A2(n12898), .ZN(n12858) );
  NAND2_X1 U15243 ( .A1(n12124), .A2(n15346), .ZN(n12132) );
  INV_X1 U15244 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15453) );
  NAND2_X1 U15245 ( .A1(n11169), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12126) );
  NAND2_X1 U15246 ( .A1(n14468), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12125) );
  OAI211_X1 U15247 ( .C1(n14497), .C2(n15453), .A(n12126), .B(n12125), .ZN(
        n12127) );
  AOI21_X1 U15248 ( .B1(n12128), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12127), .ZN(n14466) );
  NAND2_X1 U15249 ( .A1(n15352), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12129) );
  NAND2_X1 U15250 ( .A1(n12132), .A2(n12131), .ZN(P2_U2857) );
  NOR2_X1 U15251 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12134) );
  NOR4_X1 U15252 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12133) );
  NAND4_X1 U15253 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12134), .A4(n12133), .ZN(n12147) );
  NOR2_X1 U15254 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12147), .ZN(n16733)
         );
  NOR4_X1 U15255 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12138) );
  NOR4_X1 U15256 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12137) );
  NOR4_X1 U15257 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12136) );
  NOR4_X1 U15258 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12135) );
  AND4_X1 U15259 ( .A1(n12138), .A2(n12137), .A3(n12136), .A4(n12135), .ZN(
        n12143) );
  NOR4_X1 U15260 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12141) );
  NOR4_X1 U15261 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12140) );
  NOR4_X1 U15262 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12139) );
  INV_X1 U15263 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20824) );
  AND4_X1 U15264 ( .A1(n12141), .A2(n12140), .A3(n12139), .A4(n20824), .ZN(
        n12142) );
  NAND2_X1 U15265 ( .A1(n12143), .A2(n12142), .ZN(n12144) );
  INV_X1 U15266 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21282) );
  INV_X1 U15267 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21178) );
  NOR4_X1 U15268 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        n21282), .A4(n21178), .ZN(n12146) );
  NOR4_X1 U15269 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12145)
         );
  NAND3_X1 U15270 ( .A1(n20230), .A2(n12146), .A3(n12145), .ZN(U214) );
  NOR2_X1 U15271 ( .A1(n13097), .A2(n12147), .ZN(n16659) );
  NAND2_X1 U15272 ( .A1(n16659), .A2(U214), .ZN(U212) );
  NOR3_X1 U15273 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17125) );
  INV_X1 U15274 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17100) );
  NAND2_X1 U15275 ( .A1(n17125), .A2(n17100), .ZN(n17099) );
  NOR2_X1 U15276 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17099), .ZN(n17085) );
  INV_X1 U15277 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17463) );
  NAND2_X1 U15278 ( .A1(n17085), .A2(n17463), .ZN(n17070) );
  NOR2_X1 U15279 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17070), .ZN(n17053) );
  INV_X1 U15280 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17047) );
  NAND2_X1 U15281 ( .A1(n17053), .A2(n17047), .ZN(n17044) );
  INV_X1 U15282 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17430) );
  NAND2_X1 U15283 ( .A1(n17015), .A2(n17430), .ZN(n17007) );
  INV_X1 U15284 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17000) );
  NAND2_X1 U15285 ( .A1(n17006), .A2(n17000), .ZN(n16999) );
  INV_X1 U15286 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16973) );
  NAND2_X1 U15287 ( .A1(n16983), .A2(n16973), .ZN(n16972) );
  INV_X1 U15288 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16947) );
  NAND2_X1 U15289 ( .A1(n16958), .A2(n16947), .ZN(n16943) );
  INV_X1 U15290 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16924) );
  NAND2_X1 U15291 ( .A1(n16928), .A2(n16924), .ZN(n16923) );
  NOR2_X1 U15292 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16923), .ZN(n16905) );
  INV_X1 U15293 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17273) );
  NAND2_X1 U15294 ( .A1(n16905), .A2(n17273), .ZN(n16902) );
  NOR2_X1 U15295 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16902), .ZN(n16881) );
  INV_X1 U15296 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17241) );
  NAND2_X1 U15297 ( .A1(n16881), .A2(n17241), .ZN(n16871) );
  NOR2_X1 U15298 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16871), .ZN(n16863) );
  INV_X1 U15299 ( .A(n16863), .ZN(n16849) );
  NOR2_X1 U15300 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16850), .ZN(n16842) );
  INV_X1 U15301 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16836) );
  NAND2_X1 U15302 ( .A1(n16842), .A2(n16836), .ZN(n16835) );
  NOR2_X1 U15303 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16835), .ZN(n16822) );
  NAND2_X1 U15304 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19085) );
  INV_X1 U15305 ( .A(n12148), .ZN(n12149) );
  NAND2_X1 U15306 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18448), .ZN(n12151) );
  AOI211_X4 U15307 ( .C1(n19085), .C2(n19083), .A(n12164), .B(n12151), .ZN(
        n17110) );
  AOI211_X1 U15308 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16835), .A(n16822), .B(
        n17139), .ZN(n12169) );
  INV_X1 U15309 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19010) );
  INV_X1 U15310 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18944) );
  NOR2_X1 U15311 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18945) );
  NOR3_X1 U15312 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18963), .A3(n18945), 
        .ZN(n13953) );
  INV_X1 U15313 ( .A(n13953), .ZN(n19082) );
  INV_X1 U15314 ( .A(n19085), .ZN(n18932) );
  AOI211_X1 U15315 ( .C1(n19082), .C2(n19084), .A(n18932), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n12165) );
  INV_X1 U15316 ( .A(n12165), .ZN(n18922) );
  INV_X1 U15317 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19008) );
  INV_X1 U15318 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19004) );
  INV_X1 U15319 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18987) );
  INV_X1 U15320 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18982) );
  INV_X1 U15321 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18975) );
  INV_X1 U15322 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18972) );
  INV_X1 U15323 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18968) );
  INV_X1 U15324 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18964) );
  INV_X1 U15325 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18961) );
  NOR2_X1 U15326 ( .A1(n19066), .A2(n18961), .ZN(n17107) );
  INV_X1 U15327 ( .A(n17107), .ZN(n17120) );
  NOR2_X1 U15328 ( .A1(n18964), .A2(n17120), .ZN(n17086) );
  NAND2_X1 U15329 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17086), .ZN(n17060) );
  NOR2_X1 U15330 ( .A1(n18968), .A2(n17060), .ZN(n17055) );
  NAND2_X1 U15331 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17055), .ZN(n17031) );
  NOR3_X1 U15332 ( .A1(n18975), .A2(n18972), .A3(n17031), .ZN(n17010) );
  NAND4_X1 U15333 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n17010), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16969) );
  NOR2_X1 U15334 ( .A1(n18982), .A2(n16969), .ZN(n16968) );
  NAND2_X1 U15335 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16968), .ZN(n16956) );
  NOR2_X1 U15336 ( .A1(n18987), .A2(n16956), .ZN(n16889) );
  INV_X1 U15337 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18996) );
  INV_X1 U15338 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18992) );
  NAND2_X1 U15339 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16937) );
  NOR2_X1 U15340 ( .A1(n18992), .A2(n16937), .ZN(n16891) );
  NAND2_X1 U15341 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16891), .ZN(n16892) );
  NOR2_X1 U15342 ( .A1(n18996), .A2(n16892), .ZN(n16886) );
  NAND3_X1 U15343 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16889), .A3(n16886), 
        .ZN(n16866) );
  NAND2_X1 U15344 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n16854) );
  NOR3_X1 U15345 ( .A1(n19004), .A2(n16866), .A3(n16854), .ZN(n16845) );
  NAND2_X1 U15346 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16845), .ZN(n16831) );
  NOR2_X1 U15347 ( .A1(n19008), .A2(n16831), .ZN(n12152) );
  NAND2_X1 U15348 ( .A1(n17121), .A2(n12152), .ZN(n16769) );
  NAND3_X1 U15349 ( .A1(n13960), .A2(n18931), .A3(n19083), .ZN(n18940) );
  NOR2_X2 U15350 ( .A1(n19042), .A2(n18940), .ZN(n17084) );
  NOR2_X1 U15351 ( .A1(n18308), .A2(n17084), .ZN(n17066) );
  INV_X1 U15352 ( .A(n17080), .ZN(n19097) );
  NAND2_X1 U15353 ( .A1(n18931), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18809) );
  OR2_X1 U15354 ( .A1(n18935), .A2(n18809), .ZN(n18927) );
  OAI221_X1 U15355 ( .B1(n17132), .B2(P3_REIP_REG_26__SCAN_IN), .C1(n17132), 
        .C2(n12152), .A(n17143), .ZN(n16819) );
  INV_X1 U15356 ( .A(n16819), .ZN(n12153) );
  AOI21_X1 U15357 ( .B1(n19010), .B2(n16769), .A(n12153), .ZN(n12168) );
  INV_X1 U15358 ( .A(n12154), .ZN(n12156) );
  NOR2_X1 U15359 ( .A1(n18097), .A2(n12155), .ZN(n16772) );
  AOI21_X1 U15360 ( .B1(n10273), .B2(n12156), .A(n16772), .ZN(n17769) );
  INV_X1 U15361 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17790) );
  NOR2_X1 U15362 ( .A1(n17790), .A2(n12162), .ZN(n12161) );
  OAI21_X1 U15363 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n12161), .A(
        n12156), .ZN(n17781) );
  INV_X1 U15364 ( .A(n17781), .ZN(n16829) );
  OAI21_X1 U15365 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17779), .A(
        n12162), .ZN(n12157) );
  INV_X1 U15366 ( .A(n12157), .ZN(n17804) );
  INV_X1 U15367 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17825) );
  INV_X1 U15368 ( .A(n12159), .ZN(n12160) );
  NAND2_X1 U15369 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12160), .ZN(
        n12158) );
  AOI21_X1 U15370 ( .B1(n17825), .B2(n12158), .A(n17779), .ZN(n17823) );
  NOR2_X1 U15371 ( .A1(n18097), .A2(n17842), .ZN(n17817) );
  INV_X1 U15372 ( .A(n17817), .ZN(n16893) );
  AOI21_X1 U15373 ( .B1(n17841), .B2(n16893), .A(n12160), .ZN(n17846) );
  NAND2_X1 U15374 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17889), .ZN(
        n16942) );
  INV_X1 U15375 ( .A(n16942), .ZN(n17890) );
  NAND2_X1 U15376 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17890), .ZN(
        n16941) );
  NOR2_X1 U15377 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16941), .ZN(
        n16914) );
  INV_X1 U15378 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16779) );
  INV_X1 U15379 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16794) );
  INV_X1 U15380 ( .A(n16587), .ZN(n16608) );
  NOR2_X1 U15381 ( .A1(n17846), .A2(n16895), .ZN(n16882) );
  NOR2_X1 U15382 ( .A1(n16882), .A2(n17116), .ZN(n16875) );
  INV_X1 U15383 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17834) );
  AOI22_X1 U15384 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12160), .B1(
        n12159), .B2(n17834), .ZN(n17837) );
  NOR2_X1 U15385 ( .A1(n17823), .A2(n16862), .ZN(n16861) );
  NOR2_X1 U15386 ( .A1(n16861), .A2(n17116), .ZN(n16853) );
  NOR2_X1 U15387 ( .A1(n17804), .A2(n16853), .ZN(n16852) );
  NOR2_X1 U15388 ( .A1(n16852), .A2(n17116), .ZN(n16841) );
  AOI21_X1 U15389 ( .B1(n17790), .B2(n12162), .A(n12161), .ZN(n17793) );
  NOR2_X1 U15390 ( .A1(n16829), .A2(n16828), .ZN(n16827) );
  NOR2_X1 U15391 ( .A1(n16827), .A2(n17116), .ZN(n12163) );
  NOR2_X1 U15392 ( .A1(n17769), .A2(n12163), .ZN(n16773) );
  INV_X1 U15393 ( .A(n17084), .ZN(n18938) );
  AOI211_X1 U15394 ( .C1(n17769), .C2(n12163), .A(n16773), .B(n18938), .ZN(
        n12167) );
  AOI211_X4 U15395 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18448), .A(n12165), .B(
        n12164), .ZN(n17136) );
  INV_X1 U15396 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17195) );
  OAI22_X1 U15397 ( .A1(n10273), .A2(n17127), .B1(n17140), .B2(n17195), .ZN(
        n12166) );
  OR4_X1 U15398 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        P3_U2645) );
  NAND2_X1 U15399 ( .A1(n12896), .A2(n16570), .ZN(n12175) );
  INV_X1 U15400 ( .A(n12175), .ZN(n12171) );
  INV_X1 U15401 ( .A(n12909), .ZN(n12170) );
  AND2_X1 U15402 ( .A1(n12171), .A2(n12170), .ZN(n19297) );
  INV_X1 U15403 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12174) );
  AND2_X1 U15404 ( .A1(n20037), .A2(n14497), .ZN(n12176) );
  INV_X1 U15405 ( .A(n12176), .ZN(n12173) );
  OAI211_X1 U15406 ( .C1(n19297), .C2(n12174), .A(n12173), .B(n12626), .ZN(
        P2_U2814) );
  INV_X1 U15407 ( .A(n11116), .ZN(n12188) );
  INV_X1 U15408 ( .A(n11447), .ZN(n12897) );
  OAI21_X1 U15409 ( .B1(n12176), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19104), 
        .ZN(n12177) );
  OAI21_X1 U15410 ( .B1(n12188), .B2(n19104), .A(n12177), .ZN(P2_U3612) );
  NOR2_X1 U15411 ( .A1(n12178), .A2(n13473), .ZN(n12179) );
  AND2_X1 U15412 ( .A1(n11447), .A2(n12179), .ZN(n12180) );
  AND2_X1 U15413 ( .A1(n12896), .A2(n12180), .ZN(n12913) );
  NOR2_X1 U15414 ( .A1(n12913), .A2(n14501), .ZN(n20084) );
  AND2_X1 U15415 ( .A1(n12181), .A2(n16570), .ZN(n12182) );
  NAND2_X1 U15416 ( .A1(n12183), .A2(n12182), .ZN(n12357) );
  OAI21_X1 U15417 ( .B1(n20084), .B2(n12905), .A(n12357), .ZN(P2_U2819) );
  NAND2_X1 U15418 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12944) );
  NOR2_X1 U15419 ( .A1(n16562), .A2(n12944), .ZN(n19376) );
  NOR2_X1 U15420 ( .A1(n12184), .A2(n20067), .ZN(n12941) );
  OAI21_X1 U15421 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n12941), .A(n19104), 
        .ZN(n12185) );
  AOI21_X1 U15422 ( .B1(n19400), .B2(n19937), .A(n12185), .ZN(n12191) );
  INV_X1 U15423 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19947) );
  AOI21_X1 U15424 ( .B1(n20067), .B2(n14497), .A(n16562), .ZN(n16565) );
  AOI21_X1 U15425 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19937), .A(n16565), 
        .ZN(n12186) );
  NOR2_X1 U15426 ( .A1(n12191), .A2(n12186), .ZN(n12190) );
  OAI21_X1 U15427 ( .B1(n11259), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n12371), 
        .ZN(n12187) );
  NAND3_X1 U15428 ( .A1(n12188), .A2(n16562), .A3(n12187), .ZN(n12189) );
  AOI22_X1 U15429 ( .A1(n12191), .A2(n19947), .B1(n12190), .B2(n12189), .ZN(
        P2_U3610) );
  AND2_X4 U15430 ( .A1(n13169), .A2(n13332), .ZN(n12660) );
  AOI22_X1 U15431 ( .A1(n14389), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15432 ( .A1(n14418), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12196) );
  NOR2_X1 U15434 ( .A1(n13175), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12193) );
  AOI22_X1 U15435 ( .A1(n14394), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12648), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12194) );
  NAND4_X1 U15436 ( .A1(n12197), .A2(n12196), .A3(n12195), .A4(n12194), .ZN(
        n12211) );
  AOI22_X1 U15437 ( .A1(n12252), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12209) );
  AND2_X4 U15438 ( .A1(n13176), .A2(n12199), .ZN(n14422) );
  AND2_X2 U15439 ( .A1(n13176), .A2(n12200), .ZN(n12255) );
  AOI22_X1 U15440 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12208) );
  AND2_X2 U15441 ( .A1(n15173), .A2(n12205), .ZN(n12665) );
  INV_X1 U15442 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12202) );
  INV_X1 U15443 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12201) );
  NOR2_X1 U15444 ( .A1(n12202), .A2(n12201), .ZN(n12203) );
  AND2_X2 U15445 ( .A1(n15173), .A2(n12203), .ZN(n12256) );
  AOI22_X1 U15446 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12207) );
  INV_X1 U15447 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12454) );
  AND2_X2 U15448 ( .A1(n12205), .A2(n13174), .ZN(n12236) );
  AOI22_X1 U15449 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12236), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12206) );
  NAND4_X1 U15450 ( .A1(n12209), .A2(n12208), .A3(n12207), .A4(n12206), .ZN(
        n12210) );
  OR2_X2 U15451 ( .A1(n12211), .A2(n12210), .ZN(n12250) );
  AOI22_X1 U15452 ( .A1(n12252), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12236), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15453 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15454 ( .A1(n12647), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15455 ( .A1(n14418), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15456 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15457 ( .A1(n14394), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12648), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15458 ( .A1(n12255), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12665), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15459 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12216) );
  NAND2_X2 U15460 ( .A1(n12221), .A2(n12220), .ZN(n20285) );
  NAND2_X1 U15461 ( .A1(n20280), .A2(n20285), .ZN(n12239) );
  AOI22_X1 U15462 ( .A1(n12647), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15463 ( .A1(n12252), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14420), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12224) );
  NAND2_X1 U15464 ( .A1(n14418), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12223) );
  NAND2_X1 U15465 ( .A1(n14366), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12222) );
  AOI22_X1 U15466 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15467 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15468 ( .A1(n14394), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12648), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15469 ( .A1(n12236), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12226) );
  INV_X2 U15470 ( .A(n12250), .ZN(n12846) );
  NOR2_X1 U15471 ( .A1(n13002), .A2(n12846), .ZN(n12261) );
  AOI22_X1 U15472 ( .A1(n14418), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15473 ( .A1(n12647), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15474 ( .A1(n12252), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14394), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12233) );
  BUF_X4 U15475 ( .A(n12256), .Z(n14421) );
  AOI22_X1 U15476 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U15477 ( .A1(n12648), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12237) );
  MUX2_X1 U15478 ( .A(n12239), .B(n12261), .S(n20260), .Z(n12260) );
  AOI22_X1 U15479 ( .A1(n9809), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15480 ( .A1(n14418), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15481 ( .A1(n12647), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15482 ( .A1(n14394), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12648), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12240) );
  NAND4_X1 U15483 ( .A1(n12243), .A2(n12242), .A3(n12241), .A4(n12240), .ZN(
        n12249) );
  AOI22_X1 U15484 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15485 ( .A1(n12252), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15486 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15487 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12236), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12244) );
  NAND4_X1 U15488 ( .A1(n12247), .A2(n12246), .A3(n12245), .A4(n12244), .ZN(
        n12248) );
  INV_X1 U15489 ( .A(n12258), .ZN(n12251) );
  NOR2_X2 U15490 ( .A1(n20285), .A2(n12846), .ZN(n12418) );
  NAND2_X1 U15491 ( .A1(n12251), .A2(n12418), .ZN(n12387) );
  AOI22_X1 U15492 ( .A1(n12647), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15493 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12648), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15494 ( .A1(n14394), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12257) );
  NAND3_X1 U15495 ( .A1(n12260), .A2(n12259), .A3(n12298), .ZN(n12426) );
  AOI22_X1 U15496 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15497 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15498 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15499 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12236), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15500 ( .A1(n14389), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15501 ( .A1(n14394), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12648), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12271) );
  BUF_X4 U15502 ( .A(n14418), .Z(n14367) );
  AND3_X4 U15503 ( .A1(n12274), .A2(n12273), .A3(n12272), .ZN(n13364) );
  NAND2_X1 U15504 ( .A1(n12492), .A2(n13364), .ZN(n12275) );
  MUX2_X1 U15505 ( .A(n20631), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12290) );
  NAND2_X1 U15506 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20670), .ZN(
        n12314) );
  INV_X1 U15507 ( .A(n12314), .ZN(n12289) );
  NAND2_X1 U15508 ( .A1(n12290), .A2(n12289), .ZN(n12288) );
  NAND2_X1 U15509 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20631), .ZN(
        n12276) );
  NAND2_X1 U15510 ( .A1(n12288), .A2(n12276), .ZN(n12285) );
  NAND2_X1 U15511 ( .A1(n12285), .A2(n12277), .ZN(n12279) );
  NAND2_X1 U15512 ( .A1(n12471), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12278) );
  NAND2_X1 U15513 ( .A1(n12279), .A2(n12278), .ZN(n12287) );
  MUX2_X1 U15514 ( .A(n20594), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12286) );
  NOR2_X1 U15515 ( .A1(n13332), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12280) );
  NAND2_X1 U15516 ( .A1(n20228), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12281) );
  NAND2_X1 U15517 ( .A1(n12293), .A2(n12281), .ZN(n12283) );
  NAND2_X1 U15518 ( .A1(n13205), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12282) );
  MUX2_X1 U15519 ( .A(n12471), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12284) );
  XNOR2_X1 U15520 ( .A(n12285), .B(n12284), .ZN(n12329) );
  XNOR2_X1 U15521 ( .A(n12287), .B(n12286), .ZN(n12335) );
  OAI21_X1 U15522 ( .B1(n12290), .B2(n12289), .A(n12288), .ZN(n12322) );
  NOR3_X1 U15523 ( .A1(n12329), .A2(n12335), .A3(n12322), .ZN(n12291) );
  OR2_X1 U15524 ( .A1(n12311), .A2(n12291), .ZN(n12294) );
  NOR2_X1 U15525 ( .A1(n20228), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12292) );
  NAND2_X1 U15526 ( .A1(n12293), .A2(n12292), .ZN(n12337) );
  NOR2_X1 U15527 ( .A1(n12416), .A2(n20089), .ZN(n12295) );
  NAND2_X1 U15528 ( .A1(n12424), .A2(n12295), .ZN(n12381) );
  INV_X1 U15529 ( .A(n12381), .ZN(n12344) );
  INV_X1 U15530 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21225) );
  INV_X1 U15531 ( .A(n20625), .ZN(n20747) );
  NOR2_X1 U15532 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20747), .ZN(n13594) );
  INV_X1 U15533 ( .A(n13594), .ZN(n20092) );
  NAND2_X1 U15534 ( .A1(n12846), .A2(n20285), .ZN(n12296) );
  INV_X2 U15535 ( .A(n13364), .ZN(n20238) );
  AOI22_X1 U15536 ( .A1(n14389), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15537 ( .A1(n14418), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U15538 ( .A1(n12647), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15539 ( .A1(n14394), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12648), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12301) );
  NAND4_X1 U15540 ( .A1(n12304), .A2(n12303), .A3(n12302), .A4(n12301), .ZN(
        n12310) );
  AOI22_X1 U15541 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15542 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15543 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15544 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12236), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12305) );
  NAND4_X1 U15545 ( .A1(n12308), .A2(n12307), .A3(n12306), .A4(n12305), .ZN(
        n12309) );
  OR2_X4 U15546 ( .A1(n12310), .A2(n12309), .ZN(n20254) );
  NAND2_X1 U15547 ( .A1(n20280), .A2(n20254), .ZN(n13258) );
  NAND2_X1 U15548 ( .A1(n12336), .A2(n12311), .ZN(n12343) );
  NAND2_X1 U15549 ( .A1(n13364), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12967) );
  NAND2_X1 U15550 ( .A1(n12311), .A2(n13576), .ZN(n12341) );
  NOR2_X1 U15551 ( .A1(n20280), .A2(n20237), .ZN(n12312) );
  AOI21_X1 U15552 ( .B1(n13576), .B2(n20254), .A(n12312), .ZN(n12324) );
  INV_X1 U15553 ( .A(n12324), .ZN(n12313) );
  NOR2_X1 U15554 ( .A1(n12322), .A2(n12313), .ZN(n12321) );
  INV_X1 U15555 ( .A(n13576), .ZN(n12331) );
  OAI21_X1 U15556 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20670), .A(
        n12314), .ZN(n12316) );
  NOR2_X1 U15557 ( .A1(n12331), .A2(n12316), .ZN(n12320) );
  INV_X1 U15558 ( .A(n12492), .ZN(n12318) );
  OR2_X1 U15559 ( .A1(n20280), .A2(n13364), .ZN(n12315) );
  NAND2_X1 U15560 ( .A1(n12315), .A2(n12508), .ZN(n12330) );
  INV_X1 U15561 ( .A(n12316), .ZN(n12317) );
  OAI211_X1 U15562 ( .C1(n13364), .C2(n12318), .A(n12330), .B(n12317), .ZN(
        n12319) );
  OAI21_X1 U15563 ( .B1(n12336), .B2(n12320), .A(n12319), .ZN(n12323) );
  NAND2_X1 U15564 ( .A1(n12321), .A2(n12323), .ZN(n12328) );
  NAND2_X1 U15565 ( .A1(n12324), .A2(n20254), .ZN(n12340) );
  OAI211_X1 U15566 ( .C1(n12324), .C2(n12323), .A(n12322), .B(n12340), .ZN(
        n12327) );
  NAND2_X1 U15567 ( .A1(n13530), .A2(n12329), .ZN(n12325) );
  OAI211_X1 U15568 ( .C1(n12331), .C2(n12329), .A(n12325), .B(n12330), .ZN(
        n12326) );
  NAND3_X1 U15569 ( .A1(n12328), .A2(n12327), .A3(n12326), .ZN(n12333) );
  AOI22_X1 U15570 ( .A1(n13579), .A2(n12335), .B1(n12333), .B2(n12332), .ZN(
        n12334) );
  INV_X1 U15571 ( .A(n12337), .ZN(n12338) );
  NAND2_X1 U15572 ( .A1(n13530), .A2(n12338), .ZN(n12339) );
  OAI211_X1 U15573 ( .C1(n12344), .C2(n21225), .A(n20092), .B(n12583), .ZN(
        P1_U2801) );
  NAND2_X1 U15574 ( .A1(n16565), .A2(n12944), .ZN(n12345) );
  XNOR2_X1 U15575 ( .A(n12347), .B(n12346), .ZN(n12403) );
  INV_X1 U15576 ( .A(n12403), .ZN(n12360) );
  NAND2_X1 U15577 ( .A1(n14497), .A2(n13298), .ZN(n20030) );
  INV_X1 U15578 ( .A(n20030), .ZN(n20035) );
  OR2_X1 U15579 ( .A1(n20037), .A2(n20035), .ZN(n20065) );
  NAND2_X1 U15580 ( .A1(n20065), .A2(n11751), .ZN(n12348) );
  INV_X1 U15581 ( .A(n12349), .ZN(n12352) );
  INV_X1 U15582 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n12350) );
  NAND2_X1 U15583 ( .A1(n12350), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12351) );
  NAND2_X1 U15584 ( .A1(n12352), .A2(n12351), .ZN(n12367) );
  OAI21_X1 U15585 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13317), .ZN(n15263) );
  NAND2_X1 U15586 ( .A1(n19404), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12401) );
  NAND2_X1 U15587 ( .A1(n16477), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12353) );
  OAI211_X1 U15588 ( .C1(n16475), .C2(n15263), .A(n12401), .B(n12353), .ZN(
        n12359) );
  OAI21_X1 U15589 ( .B1(n12356), .B2(n12355), .A(n12354), .ZN(n12402) );
  NOR2_X1 U15590 ( .A1(n12402), .A2(n16478), .ZN(n12358) );
  AOI211_X1 U15591 ( .C1(n16494), .C2(n12360), .A(n12359), .B(n12358), .ZN(
        n12361) );
  OAI21_X1 U15592 ( .B1(n15261), .B2(n16486), .A(n12361), .ZN(P2_U3012) );
  AOI21_X1 U15593 ( .B1(n12363), .B2(n12364), .A(n12362), .ZN(n15839) );
  XNOR2_X1 U15594 ( .A(n19287), .B(n12364), .ZN(n15842) );
  INV_X1 U15595 ( .A(n15842), .ZN(n12365) );
  INV_X1 U15596 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19120) );
  NAND2_X1 U15597 ( .A1(n19404), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n15840) );
  OAI21_X1 U15598 ( .B1(n16480), .B2(n12365), .A(n15840), .ZN(n12366) );
  AOI21_X1 U15599 ( .B1(n16493), .B2(n15839), .A(n12366), .ZN(n12369) );
  OAI21_X1 U15600 ( .B1(n16477), .B2(n12367), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12368) );
  OAI211_X1 U15601 ( .C1(n10384), .C2(n16486), .A(n12369), .B(n12368), .ZN(
        P2_U3014) );
  INV_X1 U15602 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12830) );
  OR3_X1 U15603 ( .A1(n12863), .A2(n12909), .A3(n14501), .ZN(n12370) );
  NAND2_X1 U15604 ( .A1(n12829), .A2(n12370), .ZN(n12372) );
  AOI22_X1 U15605 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n19384), .B1(n19376), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12374) );
  OAI21_X1 U15606 ( .B1(n12830), .B2(n12570), .A(n12374), .ZN(P2_U2921) );
  INV_X1 U15607 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15608 ( .A1(n19376), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19384), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12375) );
  OAI21_X1 U15609 ( .B1(n12376), .B2(n12570), .A(n12375), .ZN(P2_U2928) );
  INV_X1 U15610 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n12821) );
  AOI22_X1 U15611 ( .A1(n19376), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19384), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12377) );
  OAI21_X1 U15612 ( .B1(n12821), .B2(n12570), .A(n12377), .ZN(P2_U2926) );
  INV_X1 U15613 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15377) );
  AOI22_X1 U15614 ( .A1(n19376), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19384), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12378) );
  OAI21_X1 U15615 ( .B1(n15377), .B2(n12570), .A(n12378), .ZN(P2_U2924) );
  INV_X1 U15616 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15402) );
  AOI22_X1 U15617 ( .A1(n19376), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19384), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12379) );
  OAI21_X1 U15618 ( .B1(n15402), .B2(n12570), .A(n12379), .ZN(P2_U2927) );
  INV_X1 U15619 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U15620 ( .A1(n19376), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19384), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12380) );
  OAI21_X1 U15621 ( .B1(n12818), .B2(n12570), .A(n12380), .ZN(P2_U2922) );
  INV_X1 U15622 ( .A(n13355), .ZN(n13106) );
  OAI21_X1 U15623 ( .B1(n13594), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13348), 
        .ZN(n12382) );
  OAI21_X1 U15624 ( .B1(n12457), .B2(n13348), .A(n12382), .ZN(P1_U3487) );
  INV_X1 U15625 ( .A(n12416), .ZN(n12383) );
  NAND2_X1 U15626 ( .A1(n12424), .A2(n12383), .ZN(n12385) );
  AND2_X1 U15627 ( .A1(n12997), .A2(n13106), .ZN(n12384) );
  AOI21_X1 U15628 ( .B1(n12385), .B2(n12299), .A(n12384), .ZN(n20088) );
  NAND2_X1 U15629 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20813) );
  OAI21_X1 U15630 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20813), .ZN(n12438) );
  OR2_X1 U15631 ( .A1(n12438), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15979) );
  NAND2_X1 U15632 ( .A1(n20238), .A2(n20254), .ZN(n13735) );
  NAND3_X1 U15633 ( .A1(n13106), .A2(n15979), .A3(n14593), .ZN(n12386) );
  NAND2_X1 U15634 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20902) );
  NAND2_X1 U15635 ( .A1(n12386), .A2(n20902), .ZN(n20903) );
  AND2_X1 U15636 ( .A1(n20088), .A2(n20903), .ZN(n15941) );
  NOR2_X1 U15637 ( .A1(n15941), .A2(n20089), .ZN(n20096) );
  INV_X1 U15638 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21242) );
  NOR2_X1 U15639 ( .A1(n15164), .A2(n12847), .ZN(n12390) );
  AND2_X1 U15640 ( .A1(n15164), .A2(n13364), .ZN(n12389) );
  NOR2_X1 U15641 ( .A1(n12388), .A2(n12389), .ZN(n12423) );
  NAND2_X1 U15642 ( .A1(n12423), .A2(n12492), .ZN(n15942) );
  NAND2_X1 U15643 ( .A1(n12390), .A2(n13355), .ZN(n13171) );
  NAND3_X1 U15644 ( .A1(n12299), .A2(n15942), .A3(n13171), .ZN(n12391) );
  MUX2_X1 U15645 ( .A(n13172), .B(n12391), .S(n12997), .Z(n12393) );
  AND2_X1 U15646 ( .A1(n12424), .A2(n12416), .ZN(n12392) );
  NOR2_X1 U15647 ( .A1(n12393), .A2(n12392), .ZN(n15943) );
  INV_X1 U15648 ( .A(n15943), .ZN(n12394) );
  NAND2_X1 U15649 ( .A1(n20096), .A2(n12394), .ZN(n12395) );
  OAI21_X1 U15650 ( .B1(n20096), .B2(n21242), .A(n12395), .ZN(P1_U3484) );
  OR2_X1 U15651 ( .A1(n12397), .A2(n12396), .ZN(n12399) );
  NAND2_X1 U15652 ( .A1(n12399), .A2(n12398), .ZN(n20050) );
  OAI211_X1 U15653 ( .C1(n19419), .C2(n12402), .A(n12401), .B(n12400), .ZN(
        n12405) );
  NOR2_X1 U15654 ( .A1(n12403), .A2(n19436), .ZN(n12404) );
  AOI211_X1 U15655 ( .C1(n19420), .C2(n20050), .A(n12405), .B(n12404), .ZN(
        n12414) );
  OAI21_X1 U15656 ( .B1(n12409), .B2(n12408), .A(n19423), .ZN(n12406) );
  AOI21_X1 U15657 ( .B1(n12407), .B2(n12409), .A(n12406), .ZN(n12412) );
  INV_X1 U15658 ( .A(n12408), .ZN(n15703) );
  NAND2_X1 U15659 ( .A1(n15703), .A2(n12409), .ZN(n12411) );
  MUX2_X1 U15660 ( .A(n12412), .B(n12411), .S(n12410), .Z(n12413) );
  OAI211_X1 U15661 ( .C1(n15261), .C2(n19411), .A(n12414), .B(n12413), .ZN(
        P2_U3044) );
  NAND2_X2 U15662 ( .A1(n12415), .A2(n12508), .ZN(n13007) );
  INV_X1 U15663 ( .A(n20902), .ZN(n20811) );
  NOR2_X1 U15664 ( .A1(n20811), .A2(n12416), .ZN(n12988) );
  INV_X1 U15665 ( .A(n12988), .ZN(n12417) );
  OAI22_X1 U15666 ( .A1(n13007), .A2(n12417), .B1(n12997), .B2(n13171), .ZN(
        n13109) );
  INV_X1 U15667 ( .A(n13109), .ZN(n12435) );
  NAND2_X1 U15668 ( .A1(n13364), .A2(n20254), .ZN(n13378) );
  BUF_X1 U15669 ( .A(n12418), .Z(n12419) );
  AOI21_X1 U15670 ( .B1(n12419), .B2(n20254), .A(n13364), .ZN(n12422) );
  INV_X1 U15671 ( .A(n12419), .ZN(n13114) );
  NAND2_X1 U15672 ( .A1(n13114), .A2(n12659), .ZN(n12421) );
  OR2_X2 U15673 ( .A1(n12421), .A2(n10365), .ZN(n12443) );
  NAND2_X1 U15674 ( .A1(n12422), .A2(n12443), .ZN(n12495) );
  AND2_X1 U15675 ( .A1(n12423), .A2(n12495), .ZN(n12425) );
  OR2_X1 U15676 ( .A1(n12425), .A2(n12424), .ZN(n12999) );
  NAND2_X1 U15677 ( .A1(n13172), .A2(n12997), .ZN(n12639) );
  OAI211_X1 U15678 ( .C1(n13378), .C2(n20260), .A(n12999), .B(n12639), .ZN(
        n12433) );
  INV_X1 U15679 ( .A(n13378), .ZN(n12427) );
  NAND2_X1 U15680 ( .A1(n12427), .A2(n12492), .ZN(n12428) );
  NOR2_X1 U15681 ( .A1(n12455), .A2(n12428), .ZN(n15925) );
  INV_X1 U15682 ( .A(n15979), .ZN(n13365) );
  NAND2_X1 U15683 ( .A1(n15925), .A2(n13365), .ZN(n12431) );
  OAI21_X1 U15684 ( .B1(n13365), .B2(n14597), .A(n12429), .ZN(n12430) );
  AOI21_X1 U15685 ( .B1(n12431), .B2(n12430), .A(n13107), .ZN(n12432) );
  NOR2_X1 U15686 ( .A1(n12433), .A2(n12432), .ZN(n12434) );
  NAND2_X1 U15687 ( .A1(n12435), .A2(n12434), .ZN(n15928) );
  NOR2_X1 U15688 ( .A1(n12749), .A2(n16272), .ZN(n16276) );
  NAND2_X1 U15689 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16276), .ZN(n16277) );
  INV_X1 U15690 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21158) );
  NOR2_X1 U15691 ( .A1(n16277), .A2(n21158), .ZN(n12436) );
  AOI21_X1 U15692 ( .B1(n15928), .B2(n13111), .A(n12436), .ZN(n12485) );
  NAND2_X1 U15693 ( .A1(n20237), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n12437) );
  AND2_X1 U15694 ( .A1(n12485), .A2(n12437), .ZN(n20876) );
  INV_X1 U15695 ( .A(n20876), .ZN(n20878) );
  INV_X1 U15696 ( .A(n14446), .ZN(n12641) );
  NAND2_X1 U15697 ( .A1(n12492), .A2(n9846), .ZN(n13011) );
  NAND2_X1 U15698 ( .A1(n20238), .A2(n20260), .ZN(n12491) );
  OAI211_X1 U15699 ( .C1(n20905), .C2(n12659), .A(n13011), .B(n12491), .ZN(
        n12460) );
  INV_X1 U15700 ( .A(n13168), .ZN(n12441) );
  NAND2_X1 U15701 ( .A1(n12441), .A2(n13378), .ZN(n12442) );
  NOR2_X1 U15702 ( .A1(n12460), .A2(n12442), .ZN(n12445) );
  NAND2_X1 U15703 ( .A1(n12455), .A2(n13364), .ZN(n12444) );
  NAND3_X1 U15704 ( .A1(n12445), .A2(n12444), .A3(n12461), .ZN(n12446) );
  OAI21_X2 U15705 ( .B1(n12449), .B2(n12446), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12475) );
  NAND2_X1 U15706 ( .A1(n15169), .A2(n20237), .ZN(n12704) );
  NAND2_X1 U15707 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12473) );
  OAI21_X1 U15708 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n12473), .ZN(n20699) );
  NAND2_X1 U15709 ( .A1(n15952), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12467) );
  OAI21_X1 U15710 ( .B1(n12704), .B2(n20699), .A(n12467), .ZN(n12447) );
  INV_X1 U15711 ( .A(n12447), .ZN(n12448) );
  OAI21_X2 U15712 ( .B1(n12475), .B2(n15166), .A(n12448), .ZN(n12451) );
  XNOR2_X2 U15713 ( .A(n12451), .B(n12466), .ZN(n20356) );
  INV_X1 U15714 ( .A(n15952), .ZN(n12452) );
  MUX2_X1 U15715 ( .A(n12452), .B(n12704), .S(n20670), .Z(n12453) );
  OAI21_X2 U15716 ( .B1(n12475), .B2(n12454), .A(n12453), .ZN(n12490) );
  NAND2_X1 U15717 ( .A1(n12455), .A2(n13355), .ZN(n12500) );
  AOI22_X1 U15718 ( .A1(n12457), .A2(n12456), .B1(n13786), .B2(n10365), .ZN(
        n12465) );
  NAND2_X1 U15719 ( .A1(n13168), .A2(n12458), .ZN(n13009) );
  NAND4_X1 U15720 ( .A1(n13009), .A2(n15169), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .A4(n13378), .ZN(n12459) );
  NOR2_X1 U15721 ( .A1(n12460), .A2(n12459), .ZN(n12464) );
  INV_X1 U15722 ( .A(n12461), .ZN(n12462) );
  NAND2_X1 U15723 ( .A1(n12462), .A2(n20254), .ZN(n12463) );
  NAND4_X1 U15724 ( .A1(n12500), .A2(n12465), .A3(n12464), .A4(n12463), .ZN(
        n12488) );
  INV_X1 U15725 ( .A(n12466), .ZN(n12469) );
  NAND2_X1 U15726 ( .A1(n12467), .A2(n15166), .ZN(n12468) );
  NAND2_X1 U15727 ( .A1(n12469), .A2(n12468), .ZN(n12470) );
  INV_X1 U15728 ( .A(n12473), .ZN(n12472) );
  NAND2_X1 U15729 ( .A1(n12472), .A2(n12471), .ZN(n20595) );
  NAND2_X1 U15730 ( .A1(n12473), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12474) );
  OR2_X1 U15731 ( .A1(n12478), .A2(n13175), .ZN(n12477) );
  NAND2_X1 U15732 ( .A1(n15952), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12476) );
  NAND2_X2 U15733 ( .A1(n12954), .A2(n12953), .ZN(n13166) );
  OR2_X1 U15734 ( .A1(n12478), .A2(n13332), .ZN(n12483) );
  INV_X1 U15735 ( .A(n12704), .ZN(n12481) );
  NAND3_X1 U15736 ( .A1(n20594), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20471) );
  INV_X1 U15737 ( .A(n20471), .ZN(n20474) );
  NAND2_X1 U15738 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20474), .ZN(
        n20469) );
  NAND2_X1 U15739 ( .A1(n20594), .A2(n20469), .ZN(n12480) );
  NAND3_X1 U15740 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20748) );
  INV_X1 U15741 ( .A(n20748), .ZN(n12479) );
  NAND2_X1 U15742 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12479), .ZN(
        n20740) );
  AND2_X1 U15743 ( .A1(n12480), .A2(n20740), .ZN(n20497) );
  AOI22_X1 U15744 ( .A1(n12481), .A2(n20497), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15952), .ZN(n12482) );
  OR2_X1 U15745 ( .A1(n13166), .A2(n10142), .ZN(n12484) );
  XNOR2_X1 U15746 ( .A(n12484), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20152) );
  INV_X1 U15747 ( .A(n13007), .ZN(n13203) );
  INV_X1 U15748 ( .A(n12485), .ZN(n12486) );
  NAND4_X1 U15749 ( .A1(n20152), .A2(n13203), .A3(n15169), .A4(n12486), .ZN(
        n12487) );
  OAI21_X1 U15750 ( .B1(n20878), .B2(n13205), .A(n12487), .ZN(P1_U3468) );
  INV_X1 U15751 ( .A(n12488), .ZN(n12489) );
  OAI21_X1 U15752 ( .B1(n12492), .B2(n13378), .A(n12491), .ZN(n12493) );
  INV_X1 U15753 ( .A(n12493), .ZN(n12494) );
  OAI211_X1 U15754 ( .C1(n14567), .C2(n12297), .A(n12495), .B(n12494), .ZN(
        n12496) );
  INV_X1 U15755 ( .A(n12496), .ZN(n12499) );
  OAI21_X1 U15756 ( .B1(n12497), .B2(n13168), .A(n20254), .ZN(n12498) );
  AND3_X1 U15757 ( .A1(n12500), .A2(n12499), .A3(n12498), .ZN(n13010) );
  AND2_X1 U15758 ( .A1(n13011), .A2(n20280), .ZN(n12501) );
  NAND3_X1 U15759 ( .A1(n13007), .A2(n13010), .A3(n12501), .ZN(n13167) );
  NOR2_X1 U15760 ( .A1(n15164), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12502) );
  AOI21_X1 U15761 ( .B1(n12646), .B2(n13167), .A(n12502), .ZN(n15927) );
  INV_X1 U15762 ( .A(n15927), .ZN(n12504) );
  OAI22_X1 U15763 ( .A1(n16272), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20875), .ZN(n12503) );
  AOI21_X1 U15764 ( .B1(n12504), .B2(n15169), .A(n12503), .ZN(n12506) );
  AOI21_X1 U15765 ( .B1(n15925), .B2(n15169), .A(n20876), .ZN(n12505) );
  OAI22_X1 U15766 ( .A1(n12506), .A2(n20876), .B1(n12505), .B2(n12644), .ZN(
        P1_U3474) );
  AND2_X1 U15767 ( .A1(n20905), .A2(n20811), .ZN(n12507) );
  INV_X2 U15768 ( .A(n12623), .ZN(n20224) );
  AOI22_X1 U15769 ( .A1(n20225), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20224), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n12512) );
  NAND2_X1 U15770 ( .A1(n12623), .A2(n20254), .ZN(n12624) );
  INV_X1 U15771 ( .A(n20230), .ZN(n20229) );
  NAND2_X1 U15772 ( .A1(n20229), .A2(DATAI_1_), .ZN(n12510) );
  NAND2_X1 U15773 ( .A1(n20230), .A2(BUF1_REG_1__SCAN_IN), .ZN(n12509) );
  AND2_X1 U15774 ( .A1(n12510), .A2(n12509), .ZN(n20255) );
  INV_X1 U15775 ( .A(n20255), .ZN(n12511) );
  NAND2_X1 U15776 ( .A1(n12619), .A2(n12511), .ZN(n12533) );
  NAND2_X1 U15777 ( .A1(n12512), .A2(n12533), .ZN(P1_U2953) );
  AOI22_X1 U15778 ( .A1(n20225), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20224), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n12515) );
  INV_X1 U15779 ( .A(DATAI_7_), .ZN(n12513) );
  MUX2_X1 U15780 ( .A(n12513), .B(n16691), .S(n20230), .Z(n20297) );
  INV_X1 U15781 ( .A(n20297), .ZN(n12514) );
  NAND2_X1 U15782 ( .A1(n12619), .A2(n12514), .ZN(n12520) );
  NAND2_X1 U15783 ( .A1(n12515), .A2(n12520), .ZN(P1_U2959) );
  AOI22_X1 U15784 ( .A1(n20225), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20224), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n12519) );
  INV_X1 U15785 ( .A(DATAI_3_), .ZN(n12517) );
  INV_X1 U15786 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n12516) );
  MUX2_X1 U15787 ( .A(n12517), .B(n12516), .S(n20230), .Z(n20269) );
  INV_X1 U15788 ( .A(n20269), .ZN(n12518) );
  NAND2_X1 U15789 ( .A1(n12619), .A2(n12518), .ZN(n12552) );
  NAND2_X1 U15790 ( .A1(n12519), .A2(n12552), .ZN(P1_U2955) );
  AOI22_X1 U15791 ( .A1(n20225), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20224), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n12521) );
  NAND2_X1 U15792 ( .A1(n12521), .A2(n12520), .ZN(P1_U2944) );
  AOI22_X1 U15793 ( .A1(n20225), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20224), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n12525) );
  INV_X1 U15794 ( .A(DATAI_6_), .ZN(n12523) );
  INV_X1 U15795 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n12522) );
  MUX2_X1 U15796 ( .A(n12523), .B(n12522), .S(n20230), .Z(n20287) );
  INV_X1 U15797 ( .A(n20287), .ZN(n12524) );
  NAND2_X1 U15798 ( .A1(n12619), .A2(n12524), .ZN(n12546) );
  NAND2_X1 U15799 ( .A1(n12525), .A2(n12546), .ZN(P1_U2958) );
  AOI22_X1 U15800 ( .A1(n20225), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20224), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n12528) );
  INV_X1 U15801 ( .A(DATAI_2_), .ZN(n12526) );
  MUX2_X1 U15802 ( .A(n12526), .B(n16699), .S(n20230), .Z(n20262) );
  INV_X1 U15803 ( .A(n20262), .ZN(n12527) );
  NAND2_X1 U15804 ( .A1(n12619), .A2(n12527), .ZN(n12535) );
  NAND2_X1 U15805 ( .A1(n12528), .A2(n12535), .ZN(P1_U2939) );
  AOI22_X1 U15806 ( .A1(n20225), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20224), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n12532) );
  NAND2_X1 U15807 ( .A1(n20229), .A2(DATAI_0_), .ZN(n12530) );
  NAND2_X1 U15808 ( .A1(n20230), .A2(BUF1_REG_0__SCAN_IN), .ZN(n12529) );
  AND2_X1 U15809 ( .A1(n12530), .A2(n12529), .ZN(n20244) );
  INV_X1 U15810 ( .A(n20244), .ZN(n12531) );
  NAND2_X1 U15811 ( .A1(n12619), .A2(n12531), .ZN(n12541) );
  NAND2_X1 U15812 ( .A1(n12532), .A2(n12541), .ZN(P1_U2952) );
  AOI22_X1 U15813 ( .A1(n20225), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20224), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n12534) );
  NAND2_X1 U15814 ( .A1(n12534), .A2(n12533), .ZN(P1_U2938) );
  AOI22_X1 U15815 ( .A1(n20225), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20224), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n12536) );
  NAND2_X1 U15816 ( .A1(n12536), .A2(n12535), .ZN(P1_U2954) );
  AOI22_X1 U15817 ( .A1(n20225), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20224), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n12540) );
  INV_X1 U15818 ( .A(DATAI_5_), .ZN(n12538) );
  INV_X1 U15819 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n12537) );
  MUX2_X1 U15820 ( .A(n12538), .B(n12537), .S(n20230), .Z(n20281) );
  INV_X1 U15821 ( .A(n20281), .ZN(n12539) );
  NAND2_X1 U15822 ( .A1(n12619), .A2(n12539), .ZN(n12550) );
  NAND2_X1 U15823 ( .A1(n12540), .A2(n12550), .ZN(P1_U2957) );
  AOI22_X1 U15824 ( .A1(n20225), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20224), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n12542) );
  NAND2_X1 U15825 ( .A1(n12542), .A2(n12541), .ZN(P1_U2937) );
  AOI22_X1 U15826 ( .A1(n20225), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20224), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n12545) );
  INV_X1 U15827 ( .A(DATAI_4_), .ZN(n12543) );
  MUX2_X1 U15828 ( .A(n12543), .B(n16696), .S(n20230), .Z(n20274) );
  INV_X1 U15829 ( .A(n20274), .ZN(n12544) );
  NAND2_X1 U15830 ( .A1(n12619), .A2(n12544), .ZN(n12548) );
  NAND2_X1 U15831 ( .A1(n12545), .A2(n12548), .ZN(P1_U2956) );
  AOI22_X1 U15832 ( .A1(n20225), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20224), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U15833 ( .A1(n12547), .A2(n12546), .ZN(P1_U2943) );
  AOI22_X1 U15834 ( .A1(n20225), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20224), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n12549) );
  NAND2_X1 U15835 ( .A1(n12549), .A2(n12548), .ZN(P1_U2941) );
  AOI22_X1 U15836 ( .A1(n20225), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20224), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n12551) );
  NAND2_X1 U15837 ( .A1(n12551), .A2(n12550), .ZN(P1_U2942) );
  AOI22_X1 U15838 ( .A1(n20225), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20224), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n12553) );
  NAND2_X1 U15839 ( .A1(n12553), .A2(n12552), .ZN(P1_U2940) );
  INV_X1 U15840 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15841 ( .A1(n19400), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12554) );
  OAI21_X1 U15842 ( .B1(n12555), .B2(n12570), .A(n12554), .ZN(P2_U2931) );
  INV_X1 U15843 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15844 ( .A1(n19400), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12556) );
  OAI21_X1 U15845 ( .B1(n12557), .B2(n12570), .A(n12556), .ZN(P2_U2935) );
  INV_X1 U15846 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U15847 ( .A1(n19400), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12558) );
  OAI21_X1 U15848 ( .B1(n12559), .B2(n12570), .A(n12558), .ZN(P2_U2934) );
  INV_X1 U15849 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U15850 ( .A1(n19400), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12560) );
  OAI21_X1 U15851 ( .B1(n12561), .B2(n12570), .A(n12560), .ZN(P2_U2932) );
  INV_X1 U15852 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15853 ( .A1(n19400), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12562) );
  OAI21_X1 U15854 ( .B1(n12563), .B2(n12570), .A(n12562), .ZN(P2_U2933) );
  INV_X1 U15855 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n15385) );
  AOI22_X1 U15856 ( .A1(n19376), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12564) );
  OAI21_X1 U15857 ( .B1(n15385), .B2(n12570), .A(n12564), .ZN(P2_U2925) );
  INV_X1 U15858 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U15859 ( .A1(n19376), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12565) );
  OAI21_X1 U15860 ( .B1(n12566), .B2(n12570), .A(n12565), .ZN(P2_U2929) );
  INV_X1 U15861 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15862 ( .A1(n19376), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12567) );
  OAI21_X1 U15863 ( .B1(n12568), .B2(n12570), .A(n12567), .ZN(P2_U2930) );
  INV_X1 U15864 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15368) );
  AOI22_X1 U15865 ( .A1(n19376), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12569) );
  OAI21_X1 U15866 ( .B1(n15368), .B2(n12570), .A(n12569), .ZN(P2_U2923) );
  OAI21_X1 U15867 ( .B1(n12573), .B2(n12572), .A(n12571), .ZN(n12574) );
  XOR2_X1 U15868 ( .A(n12574), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n19437) );
  OR2_X1 U15869 ( .A1(n12575), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12577) );
  AND2_X1 U15870 ( .A1(n12577), .A2(n12576), .ZN(n19428) );
  NAND2_X1 U15871 ( .A1(n19404), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19434) );
  INV_X1 U15872 ( .A(n19434), .ZN(n12579) );
  MUX2_X1 U15873 ( .A(n16488), .B(n16477), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n12578) );
  AOI211_X1 U15874 ( .C1(n19428), .C2(n16493), .A(n12579), .B(n12578), .ZN(
        n12581) );
  NAND2_X1 U15875 ( .A1(n19425), .A2(n16491), .ZN(n12580) );
  OAI211_X1 U15876 ( .C1(n19437), .C2(n16480), .A(n12581), .B(n12580), .ZN(
        P2_U3013) );
  INV_X1 U15877 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n21149) );
  NAND3_X1 U15878 ( .A1(n15925), .A2(n13111), .A3(n10073), .ZN(n12582) );
  OAI21_X1 U15879 ( .B1(n12583), .B2(n20254), .A(n12582), .ZN(n12584) );
  NAND2_X1 U15880 ( .A1(n20189), .A2(n20238), .ZN(n13087) );
  NAND2_X1 U15881 ( .A1(n20237), .A2(n16276), .ZN(n20187) );
  INV_X2 U15882 ( .A(n20187), .ZN(n20210) );
  NOR2_X4 U15883 ( .A1(n20189), .A2(n20210), .ZN(n15982) );
  AOI22_X1 U15884 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12585) );
  OAI21_X1 U15885 ( .B1(n21149), .B2(n13087), .A(n12585), .ZN(P1_U2907) );
  INV_X1 U15886 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n21023) );
  AOI22_X1 U15887 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12586) );
  OAI21_X1 U15888 ( .B1(n21023), .B2(n13087), .A(n12586), .ZN(P1_U2909) );
  INV_X1 U15889 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12588) );
  AOI22_X1 U15890 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12587) );
  OAI21_X1 U15891 ( .B1(n12588), .B2(n13087), .A(n12587), .ZN(P1_U2917) );
  INV_X1 U15892 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U15893 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12589) );
  OAI21_X1 U15894 ( .B1(n12607), .B2(n13087), .A(n12589), .ZN(P1_U2912) );
  INV_X1 U15895 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15896 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12590) );
  OAI21_X1 U15897 ( .B1(n12591), .B2(n13087), .A(n12590), .ZN(P1_U2913) );
  INV_X1 U15898 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n21191) );
  AOI22_X1 U15899 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12592) );
  OAI21_X1 U15900 ( .B1(n21191), .B2(n13087), .A(n12592), .ZN(P1_U2914) );
  INV_X1 U15901 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21132) );
  AOI22_X1 U15902 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12593) );
  OAI21_X1 U15903 ( .B1(n21132), .B2(n13087), .A(n12593), .ZN(P1_U2915) );
  INV_X1 U15904 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21197) );
  AOI22_X1 U15905 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12594) );
  OAI21_X1 U15906 ( .B1(n21197), .B2(n13087), .A(n12594), .ZN(P1_U2911) );
  INV_X1 U15907 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n21068) );
  AOI22_X1 U15908 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12595) );
  OAI21_X1 U15909 ( .B1(n21068), .B2(n13087), .A(n12595), .ZN(P1_U2908) );
  INV_X1 U15910 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n21155) );
  AOI22_X1 U15911 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12596) );
  OAI21_X1 U15912 ( .B1(n21155), .B2(n13087), .A(n12596), .ZN(P1_U2916) );
  INV_X1 U15913 ( .A(n12598), .ZN(n12599) );
  NAND2_X1 U15914 ( .A1(n20051), .A2(n15346), .ZN(n12601) );
  INV_X2 U15915 ( .A(n15352), .ZN(n15356) );
  NAND2_X1 U15916 ( .A1(n12888), .A2(n15356), .ZN(n12600) );
  OAI211_X1 U15917 ( .C1(n15356), .C2(n10619), .A(n12601), .B(n12600), .ZN(
        P2_U2885) );
  INV_X1 U15918 ( .A(n20225), .ZN(n12625) );
  INV_X1 U15919 ( .A(DATAI_12_), .ZN(n12603) );
  NAND2_X1 U15920 ( .A1(n20230), .A2(BUF1_REG_12__SCAN_IN), .ZN(n12602) );
  OAI21_X1 U15921 ( .B1(n20230), .B2(n12603), .A(n12602), .ZN(n14812) );
  NAND2_X1 U15922 ( .A1(n12619), .A2(n14812), .ZN(n20220) );
  NAND2_X1 U15923 ( .A1(n20224), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n12604) );
  OAI211_X1 U15924 ( .C1(n12625), .C2(n21068), .A(n20220), .B(n12604), .ZN(
        P1_U2949) );
  NAND2_X1 U15925 ( .A1(n20224), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n12606) );
  INV_X1 U15926 ( .A(DATAI_8_), .ZN(n21194) );
  INV_X1 U15927 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16689) );
  MUX2_X1 U15928 ( .A(n21194), .B(n16689), .S(n20230), .Z(n14832) );
  INV_X1 U15929 ( .A(n14832), .ZN(n12605) );
  NAND2_X1 U15930 ( .A1(n12619), .A2(n12605), .ZN(n12608) );
  OAI211_X1 U15931 ( .C1(n12625), .C2(n12607), .A(n12606), .B(n12608), .ZN(
        P1_U2945) );
  INV_X1 U15932 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20199) );
  NAND2_X1 U15933 ( .A1(n20224), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n12609) );
  OAI211_X1 U15934 ( .C1(n12625), .C2(n20199), .A(n12609), .B(n12608), .ZN(
        P1_U2960) );
  INV_X1 U15935 ( .A(DATAI_11_), .ZN(n21243) );
  INV_X1 U15936 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16683) );
  MUX2_X1 U15937 ( .A(n21243), .B(n16683), .S(n20230), .Z(n14818) );
  INV_X1 U15938 ( .A(n14818), .ZN(n12610) );
  NAND2_X1 U15939 ( .A1(n12619), .A2(n12610), .ZN(n20218) );
  NAND2_X1 U15940 ( .A1(n20224), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n12611) );
  OAI211_X1 U15941 ( .C1(n12625), .C2(n21023), .A(n20218), .B(n12611), .ZN(
        P1_U2948) );
  INV_X1 U15942 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13079) );
  INV_X1 U15943 ( .A(DATAI_14_), .ZN(n20989) );
  NAND2_X1 U15944 ( .A1(n20230), .A2(BUF1_REG_14__SCAN_IN), .ZN(n12612) );
  OAI21_X1 U15945 ( .B1(n20230), .B2(n20989), .A(n12612), .ZN(n14874) );
  NAND2_X1 U15946 ( .A1(n12619), .A2(n14874), .ZN(n20226) );
  NAND2_X1 U15947 ( .A1(n20224), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n12613) );
  OAI211_X1 U15948 ( .C1(n12625), .C2(n13079), .A(n20226), .B(n12613), .ZN(
        P1_U2951) );
  INV_X1 U15949 ( .A(DATAI_9_), .ZN(n21196) );
  INV_X1 U15950 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16687) );
  MUX2_X1 U15951 ( .A(n21196), .B(n16687), .S(n20230), .Z(n14828) );
  INV_X1 U15952 ( .A(n14828), .ZN(n12614) );
  NAND2_X1 U15953 ( .A1(n12619), .A2(n12614), .ZN(n20214) );
  NAND2_X1 U15954 ( .A1(n20224), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n12615) );
  OAI211_X1 U15955 ( .C1(n12625), .C2(n21197), .A(n20214), .B(n12615), .ZN(
        P1_U2946) );
  INV_X1 U15956 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21206) );
  INV_X1 U15957 ( .A(DATAI_10_), .ZN(n21234) );
  INV_X1 U15958 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16685) );
  MUX2_X1 U15959 ( .A(n21234), .B(n16685), .S(n20230), .Z(n14823) );
  INV_X1 U15960 ( .A(n14823), .ZN(n12616) );
  NAND2_X1 U15961 ( .A1(n12619), .A2(n12616), .ZN(n20216) );
  NAND2_X1 U15962 ( .A1(n20224), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n12617) );
  OAI211_X1 U15963 ( .C1(n12625), .C2(n21206), .A(n20216), .B(n12617), .ZN(
        P1_U2947) );
  INV_X1 U15964 ( .A(DATAI_13_), .ZN(n21021) );
  INV_X1 U15965 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16679) );
  MUX2_X1 U15966 ( .A(n21021), .B(n16679), .S(n20230), .Z(n14877) );
  INV_X1 U15967 ( .A(n14877), .ZN(n12618) );
  NAND2_X1 U15968 ( .A1(n12619), .A2(n12618), .ZN(n20222) );
  NAND2_X1 U15969 ( .A1(n20224), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n12620) );
  OAI211_X1 U15970 ( .C1(n12625), .C2(n21149), .A(n20222), .B(n12620), .ZN(
        P1_U2950) );
  INV_X1 U15971 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14871) );
  INV_X1 U15972 ( .A(DATAI_15_), .ZN(n12622) );
  INV_X1 U15973 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12621) );
  MUX2_X1 U15974 ( .A(n12622), .B(n12621), .S(n20230), .Z(n14870) );
  INV_X1 U15975 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20188) );
  OAI222_X1 U15976 ( .A1(n12625), .A2(n14871), .B1(n12624), .B2(n14870), .C1(
        n12623), .C2(n20188), .ZN(P1_U2967) );
  INV_X1 U15977 ( .A(n9948), .ZN(n12628) );
  AOI22_X1 U15978 ( .A1(n13098), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13097), .ZN(n19309) );
  INV_X1 U15979 ( .A(n12626), .ZN(n13484) );
  OAI21_X1 U15980 ( .B1(n12907), .B2(n19937), .A(n13484), .ZN(n12804) );
  AOI22_X1 U15981 ( .A1(P2_LWORD_REG_15__SCAN_IN), .A2(n12826), .B1(n12801), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n12627) );
  OAI21_X1 U15982 ( .B1(n12628), .B2(n19309), .A(n12627), .ZN(P2_U2982) );
  NOR2_X1 U15983 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12630) );
  OAI21_X1 U15984 ( .B1(n12631), .B2(n12630), .A(n12629), .ZN(n12632) );
  INV_X1 U15985 ( .A(n12632), .ZN(n12633) );
  MUX2_X1 U15986 ( .A(n10384), .B(n10812), .S(n15323), .Z(n12634) );
  OAI21_X1 U15987 ( .B1(n20069), .B2(n15359), .A(n12634), .ZN(P2_U2887) );
  INV_X1 U15988 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15170) );
  NAND2_X1 U15989 ( .A1(n14567), .A2(n15170), .ZN(n12636) );
  NAND2_X1 U15990 ( .A1(n14591), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12635) );
  AND2_X1 U15991 ( .A1(n12636), .A2(n12764), .ZN(n13502) );
  INV_X1 U15992 ( .A(n13502), .ZN(n12680) );
  NOR2_X1 U15993 ( .A1(n12458), .A2(n13113), .ZN(n12637) );
  NAND4_X1 U15994 ( .A1(n13168), .A2(n12637), .A3(n12846), .A4(n12659), .ZN(
        n13105) );
  OR2_X1 U15995 ( .A1(n13105), .A2(n14593), .ZN(n12638) );
  NAND2_X1 U15996 ( .A1(n12639), .A2(n12638), .ZN(n12640) );
  INV_X1 U15997 ( .A(n13113), .ZN(n20294) );
  INV_X1 U15998 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n20997) );
  NAND2_X1 U15999 ( .A1(n12641), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13333) );
  NAND2_X1 U16000 ( .A1(n12749), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12643) );
  NAND2_X1 U16001 ( .A1(n14250), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12642) );
  OAI211_X1 U16002 ( .C1(n13333), .C2(n12644), .A(n12643), .B(n12642), .ZN(
        n12645) );
  AOI21_X1 U16003 ( .B1(n12646), .B2(n14128), .A(n12645), .ZN(n12754) );
  AOI22_X1 U16004 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U16005 ( .A1(n14418), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U16006 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12650) );
  INV_X1 U16007 ( .A(n14394), .ZN(n14263) );
  INV_X2 U16008 ( .A(n14263), .ZN(n14368) );
  AOI22_X1 U16009 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12648), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12649) );
  NAND4_X1 U16010 ( .A1(n12652), .A2(n12651), .A3(n12650), .A4(n12649), .ZN(
        n12658) );
  INV_X2 U16011 ( .A(n12724), .ZN(n14414) );
  AOI22_X1 U16012 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14414), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U16013 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U16014 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U16015 ( .A1(n14352), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12236), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12653) );
  NAND4_X1 U16016 ( .A1(n12656), .A2(n12655), .A3(n12654), .A4(n12653), .ZN(
        n12657) );
  NAND2_X1 U16017 ( .A1(n12659), .A2(n13784), .ZN(n12674) );
  NOR2_X1 U16018 ( .A1(n12966), .A2(n13784), .ZN(n12723) );
  AOI22_X1 U16019 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U16020 ( .A1(n14418), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U16021 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U16022 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12661) );
  NAND4_X1 U16023 ( .A1(n12664), .A2(n12663), .A3(n12662), .A4(n12661), .ZN(
        n12671) );
  AOI22_X1 U16024 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14422), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U16025 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12668) );
  AOI22_X1 U16026 ( .A1(n14352), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U16028 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12236), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12666) );
  NAND4_X1 U16029 ( .A1(n12669), .A2(n12668), .A3(n12667), .A4(n12666), .ZN(
        n12670) );
  MUX2_X1 U16030 ( .A(n13782), .B(n12723), .S(n12979), .Z(n12672) );
  INV_X1 U16031 ( .A(n12672), .ZN(n12673) );
  INV_X1 U16032 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12676) );
  AOI21_X1 U16033 ( .B1(n13364), .B2(n12979), .A(n20237), .ZN(n12675) );
  OAI211_X1 U16034 ( .C1(n13579), .C2(n12676), .A(n12675), .B(n12674), .ZN(
        n12719) );
  NAND2_X1 U16035 ( .A1(n20329), .A2(n12458), .ZN(n12677) );
  NAND2_X1 U16036 ( .A1(n12677), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12679) );
  OR2_X1 U16037 ( .A1(n12679), .A2(n12754), .ZN(n12757) );
  INV_X1 U16038 ( .A(n12757), .ZN(n12678) );
  AOI21_X1 U16039 ( .B1(n12754), .B2(n12679), .A(n12678), .ZN(n12710) );
  INV_X1 U16040 ( .A(n12710), .ZN(n13507) );
  NAND2_X2 U16041 ( .A1(n20185), .A2(n13113), .ZN(n14803) );
  OAI222_X1 U16042 ( .A1(n12680), .A2(n20171), .B1(n20997), .B2(n20185), .C1(
        n13507), .C2(n14803), .ZN(P1_U2872) );
  INV_X1 U16043 ( .A(n12681), .ZN(n12683) );
  NOR2_X1 U16044 ( .A1(n15356), .A2(n15278), .ZN(n12684) );
  AOI21_X1 U16045 ( .B1(n19425), .B2(n15356), .A(n12684), .ZN(n12685) );
  OAI21_X1 U16046 ( .B1(n20038), .B2(n15359), .A(n12685), .ZN(P2_U2886) );
  AOI21_X1 U16047 ( .B1(n12686), .B2(n12687), .A(n12693), .ZN(n14528) );
  XNOR2_X1 U16048 ( .A(n14528), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12692) );
  OR2_X1 U16049 ( .A1(n12699), .A2(n12688), .ZN(n12689) );
  AND2_X1 U16050 ( .A1(n12689), .A2(n13476), .ZN(n16490) );
  NOR2_X1 U16051 ( .A1(n15356), .A2(n11163), .ZN(n12690) );
  AOI21_X1 U16052 ( .B1(n16490), .B2(n15356), .A(n12690), .ZN(n12691) );
  OAI21_X1 U16053 ( .B1(n12692), .B2(n15359), .A(n12691), .ZN(P2_U2882) );
  AND3_X1 U16054 ( .A1(n12694), .A2(n12686), .A3(n12693), .ZN(n12695) );
  OR2_X1 U16055 ( .A1(n12695), .A2(n14528), .ZN(n19336) );
  INV_X1 U16056 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19270) );
  NOR2_X1 U16057 ( .A1(n12697), .A2(n12696), .ZN(n12698) );
  OR2_X1 U16058 ( .A1(n12699), .A2(n12698), .ZN(n19412) );
  MUX2_X1 U16059 ( .A(n19270), .B(n19412), .S(n15356), .Z(n12700) );
  OAI21_X1 U16060 ( .B1(n19336), .B2(n15359), .A(n12700), .ZN(P2_U2883) );
  AND2_X1 U16061 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20625), .ZN(n20885) );
  OAI21_X1 U16062 ( .B1(n20905), .B2(n12979), .A(n12983), .ZN(n12701) );
  INV_X1 U16063 ( .A(n12701), .ZN(n12702) );
  OAI21_X1 U16064 ( .B1(n20329), .B2(n13258), .A(n12702), .ZN(n12703) );
  NAND2_X1 U16065 ( .A1(n12703), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12950) );
  OAI21_X1 U16066 ( .B1(n12703), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12950), .ZN(n13044) );
  NAND2_X1 U16067 ( .A1(n16255), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13037) );
  NAND2_X1 U16068 ( .A1(n12704), .A2(n20747), .ZN(n20901) );
  NAND2_X1 U16069 ( .A1(n20901), .A2(n20237), .ZN(n12705) );
  NAND2_X1 U16070 ( .A1(n20237), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12707) );
  INV_X1 U16071 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20703) );
  NAND2_X1 U16072 ( .A1(n20703), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12706) );
  NAND2_X1 U16073 ( .A1(n12707), .A2(n12706), .ZN(n12852) );
  OAI21_X1 U16074 ( .B1(n16099), .B2(n12852), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12708) );
  OAI211_X1 U16075 ( .C1(n13044), .C2(n20095), .A(n13037), .B(n12708), .ZN(
        n12709) );
  AOI21_X1 U16076 ( .B1(n12710), .B2(n16105), .A(n12709), .ZN(n12711) );
  INV_X1 U16077 ( .A(n12711), .ZN(P1_U2999) );
  NAND2_X1 U16078 ( .A1(n12713), .A2(n12714), .ZN(n12715) );
  MUX2_X1 U16079 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n15253), .S(n15356), .Z(
        n12717) );
  AOI21_X1 U16080 ( .B1(n19326), .B2(n15346), .A(n12717), .ZN(n12718) );
  INV_X1 U16081 ( .A(n12718), .ZN(P2_U2884) );
  INV_X1 U16082 ( .A(n13782), .ZN(n12721) );
  INV_X1 U16083 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12738) );
  INV_X1 U16084 ( .A(n12723), .ZN(n12737) );
  AOI22_X1 U16085 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U16086 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U16087 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12726) );
  AOI22_X1 U16088 ( .A1(n14331), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U16089 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U16090 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12731) );
  NAND2_X1 U16091 ( .A1(n14198), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12730) );
  NAND2_X1 U16092 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12729) );
  AND4_X1 U16093 ( .A1(n12732), .A2(n12731), .A3(n12730), .A4(n12729), .ZN(
        n12735) );
  AOI22_X1 U16094 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12734) );
  OR2_X1 U16095 ( .A1(n12967), .A2(n12978), .ZN(n12736) );
  OAI211_X1 U16096 ( .C1(n13579), .C2(n12738), .A(n12737), .B(n12736), .ZN(
        n12974) );
  INV_X1 U16097 ( .A(n12974), .ZN(n12739) );
  INV_X1 U16098 ( .A(n20356), .ZN(n12742) );
  INV_X1 U16099 ( .A(n12740), .ZN(n12741) );
  NAND2_X1 U16100 ( .A1(n20302), .A2(n12743), .ZN(n13216) );
  INV_X1 U16101 ( .A(n13216), .ZN(n12744) );
  NAND2_X1 U16102 ( .A1(n12744), .A2(n20237), .ZN(n12746) );
  OR2_X1 U16103 ( .A1(n12966), .A2(n12978), .ZN(n12745) );
  INV_X1 U16104 ( .A(n12972), .ZN(n12747) );
  NAND2_X1 U16105 ( .A1(n13211), .A2(n14128), .ZN(n12753) );
  AOI22_X1 U16106 ( .A1(n14250), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n12749), .ZN(n12751) );
  INV_X1 U16107 ( .A(n13333), .ZN(n13401) );
  NAND2_X1 U16108 ( .A1(n13401), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12750) );
  AND2_X1 U16109 ( .A1(n12751), .A2(n12750), .ZN(n12752) );
  NAND2_X1 U16110 ( .A1(n12753), .A2(n12752), .ZN(n12759) );
  INV_X1 U16111 ( .A(n12754), .ZN(n12755) );
  OR2_X1 U16112 ( .A1(n12755), .A2(n14363), .ZN(n12756) );
  NAND2_X1 U16113 ( .A1(n12757), .A2(n12756), .ZN(n12758) );
  NAND2_X1 U16114 ( .A1(n12759), .A2(n12758), .ZN(n13073) );
  OAI21_X1 U16115 ( .B1(n12759), .B2(n12758), .A(n13073), .ZN(n13571) );
  INV_X1 U16116 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12760) );
  NAND2_X1 U16117 ( .A1(n14591), .A2(n12760), .ZN(n12761) );
  OAI211_X1 U16118 ( .C1(n13735), .C2(P1_EBX_REG_1__SCAN_IN), .A(n14614), .B(
        n12761), .ZN(n12763) );
  INV_X1 U16119 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n21128) );
  NAND2_X1 U16120 ( .A1(n9804), .A2(n21128), .ZN(n12762) );
  OAI21_X1 U16121 ( .B1(n12765), .B2(n14597), .A(n13022), .ZN(n13565) );
  AOI22_X1 U16122 ( .A1(n20181), .A2(n13565), .B1(n14801), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n12766) );
  OAI21_X1 U16123 ( .B1(n13571), .B2(n14803), .A(n12766), .ZN(P1_U2871) );
  AOI22_X1 U16124 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n12826), .B1(n12801), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U16125 ( .A1(n13098), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13097), .ZN(n19331) );
  INV_X1 U16126 ( .A(n19331), .ZN(n15419) );
  NAND2_X1 U16127 ( .A1(n9948), .A2(n15419), .ZN(n12799) );
  NAND2_X1 U16128 ( .A1(n12767), .A2(n12799), .ZN(P2_U2957) );
  AOI22_X1 U16129 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U16130 ( .A1(n13098), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13097), .ZN(n19368) );
  INV_X1 U16131 ( .A(n19368), .ZN(n13756) );
  NAND2_X1 U16132 ( .A1(n9948), .A2(n13756), .ZN(n12781) );
  NAND2_X1 U16133 ( .A1(n12768), .A2(n12781), .ZN(P2_U2952) );
  AOI22_X1 U16134 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U16135 ( .A1(n13098), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13097), .ZN(n19452) );
  INV_X1 U16136 ( .A(n19452), .ZN(n15431) );
  NAND2_X1 U16137 ( .A1(n9948), .A2(n15431), .ZN(n12802) );
  NAND2_X1 U16138 ( .A1(n12769), .A2(n12802), .ZN(P2_U2971) );
  AOI22_X1 U16139 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U16140 ( .A1(n13098), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13097), .ZN(n19446) );
  INV_X1 U16141 ( .A(n19446), .ZN(n13895) );
  NAND2_X1 U16142 ( .A1(n9948), .A2(n13895), .ZN(n12805) );
  NAND2_X1 U16143 ( .A1(n12770), .A2(n12805), .ZN(P2_U2970) );
  AOI22_X1 U16144 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n12804), .B1(n16287), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U16145 ( .A1(n13098), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13097), .ZN(n19440) );
  INV_X1 U16146 ( .A(n19440), .ZN(n13858) );
  NAND2_X1 U16147 ( .A1(n9948), .A2(n13858), .ZN(n12810) );
  NAND2_X1 U16148 ( .A1(n12771), .A2(n12810), .ZN(P2_U2954) );
  AOI22_X1 U16149 ( .A1(P2_LWORD_REG_12__SCAN_IN), .A2(n12804), .B1(n16287), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U16150 ( .A1(n13098), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n13097), .ZN(n15369) );
  INV_X1 U16151 ( .A(n15369), .ZN(n12772) );
  NAND2_X1 U16152 ( .A1(n9948), .A2(n12772), .ZN(n12791) );
  NAND2_X1 U16153 ( .A1(n12773), .A2(n12791), .ZN(P2_U2979) );
  AOI22_X1 U16154 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12777) );
  OR2_X1 U16155 ( .A1(n13097), .A2(n16683), .ZN(n12775) );
  NAND2_X1 U16156 ( .A1(n13097), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12774) );
  AND2_X1 U16157 ( .A1(n12775), .A2(n12774), .ZN(n19316) );
  INV_X1 U16158 ( .A(n19316), .ZN(n12776) );
  NAND2_X1 U16159 ( .A1(n9948), .A2(n12776), .ZN(n12787) );
  NAND2_X1 U16160 ( .A1(n12777), .A2(n12787), .ZN(P2_U2978) );
  AOI22_X1 U16161 ( .A1(P2_LWORD_REG_10__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n12780) );
  OR2_X1 U16162 ( .A1(n13097), .A2(n16685), .ZN(n12779) );
  NAND2_X1 U16163 ( .A1(n13097), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12778) );
  NAND2_X1 U16164 ( .A1(n12779), .A2(n12778), .ZN(n15387) );
  NAND2_X1 U16165 ( .A1(n9948), .A2(n15387), .ZN(n12789) );
  NAND2_X1 U16166 ( .A1(n12780), .A2(n12789), .ZN(P2_U2977) );
  AOI22_X1 U16167 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n12804), .B1(n16287), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n12782) );
  NAND2_X1 U16168 ( .A1(n12782), .A2(n12781), .ZN(P2_U2967) );
  AOI22_X1 U16169 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U16170 ( .A1(n13098), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n13097), .ZN(n15403) );
  INV_X1 U16171 ( .A(n15403), .ZN(n12783) );
  NAND2_X1 U16172 ( .A1(n9948), .A2(n12783), .ZN(n12793) );
  NAND2_X1 U16173 ( .A1(n12784), .A2(n12793), .ZN(P2_U2975) );
  AOI22_X1 U16174 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12785) );
  OAI22_X1 U16175 ( .A1(n13097), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13098), .ZN(n19463) );
  INV_X1 U16176 ( .A(n19463), .ZN(n16380) );
  NAND2_X1 U16177 ( .A1(n9948), .A2(n16380), .ZN(n12795) );
  NAND2_X1 U16178 ( .A1(n12785), .A2(n12795), .ZN(P2_U2974) );
  AOI22_X1 U16179 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U16180 ( .A1(n13098), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13097), .ZN(n19322) );
  INV_X1 U16181 ( .A(n19322), .ZN(n15413) );
  NAND2_X1 U16182 ( .A1(n9948), .A2(n15413), .ZN(n12797) );
  NAND2_X1 U16183 ( .A1(n12786), .A2(n12797), .ZN(P2_U2973) );
  AOI22_X1 U16184 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n12804), .B1(n12801), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12788) );
  NAND2_X1 U16185 ( .A1(n12788), .A2(n12787), .ZN(P2_U2963) );
  AOI22_X1 U16186 ( .A1(P2_UWORD_REG_10__SCAN_IN), .A2(n12804), .B1(n12801), 
        .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n12790) );
  NAND2_X1 U16187 ( .A1(n12790), .A2(n12789), .ZN(P2_U2962) );
  AOI22_X1 U16188 ( .A1(P2_UWORD_REG_12__SCAN_IN), .A2(n12804), .B1(n16287), 
        .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n12792) );
  NAND2_X1 U16189 ( .A1(n12792), .A2(n12791), .ZN(P2_U2964) );
  AOI22_X1 U16190 ( .A1(P2_UWORD_REG_8__SCAN_IN), .A2(n12804), .B1(n12801), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n12794) );
  NAND2_X1 U16191 ( .A1(n12794), .A2(n12793), .ZN(P2_U2960) );
  AOI22_X1 U16192 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n12804), .B1(n12801), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12796) );
  NAND2_X1 U16193 ( .A1(n12796), .A2(n12795), .ZN(P2_U2959) );
  AOI22_X1 U16194 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n12804), .B1(n12801), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n12798) );
  NAND2_X1 U16195 ( .A1(n12798), .A2(n12797), .ZN(P2_U2958) );
  AOI22_X1 U16196 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12800) );
  NAND2_X1 U16197 ( .A1(n12800), .A2(n12799), .ZN(P2_U2972) );
  AOI22_X1 U16198 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n12826), .B1(n12801), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12803) );
  NAND2_X1 U16199 ( .A1(n12803), .A2(n12802), .ZN(P2_U2956) );
  AOI22_X1 U16200 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n12804), .B1(n16287), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12806) );
  NAND2_X1 U16201 ( .A1(n12806), .A2(n12805), .ZN(P2_U2955) );
  AOI22_X1 U16202 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U16203 ( .A1(n13098), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13097), .ZN(n19358) );
  INV_X1 U16204 ( .A(n19358), .ZN(n13842) );
  NAND2_X1 U16205 ( .A1(n9948), .A2(n13842), .ZN(n12808) );
  NAND2_X1 U16206 ( .A1(n12807), .A2(n12808), .ZN(P2_U2968) );
  AOI22_X1 U16207 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12809) );
  NAND2_X1 U16208 ( .A1(n12809), .A2(n12808), .ZN(P2_U2953) );
  AOI22_X1 U16209 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n12826), .B1(n16287), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12811) );
  NAND2_X1 U16210 ( .A1(n12811), .A2(n12810), .ZN(P2_U2969) );
  OR2_X1 U16211 ( .A1(n13097), .A2(n16687), .ZN(n12813) );
  NAND2_X1 U16212 ( .A1(n13097), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12812) );
  NAND2_X1 U16213 ( .A1(n12813), .A2(n12812), .ZN(n15395) );
  NAND2_X1 U16214 ( .A1(n9948), .A2(n15395), .ZN(n12820) );
  NAND2_X1 U16215 ( .A1(n12826), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n12814) );
  OAI211_X1 U16216 ( .C1(n11320), .C2(n12829), .A(n12820), .B(n12814), .ZN(
        P2_U2976) );
  OR2_X1 U16217 ( .A1(n13097), .A2(n16679), .ZN(n12816) );
  NAND2_X1 U16218 ( .A1(n13097), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12815) );
  NAND2_X1 U16219 ( .A1(n12816), .A2(n12815), .ZN(n15362) );
  NAND2_X1 U16220 ( .A1(n9948), .A2(n15362), .ZN(n12823) );
  NAND2_X1 U16221 ( .A1(n12826), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n12817) );
  OAI211_X1 U16222 ( .C1(n12818), .C2(n12829), .A(n12823), .B(n12817), .ZN(
        P2_U2965) );
  NAND2_X1 U16223 ( .A1(n12826), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12819) );
  OAI211_X1 U16224 ( .C1(n12821), .C2(n12829), .A(n12820), .B(n12819), .ZN(
        P2_U2961) );
  INV_X1 U16225 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19375) );
  NAND2_X1 U16226 ( .A1(n12826), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n12822) );
  OAI211_X1 U16227 ( .C1(n19375), .C2(n12829), .A(n12823), .B(n12822), .ZN(
        P2_U2980) );
  INV_X1 U16228 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19373) );
  NAND2_X1 U16229 ( .A1(n9948), .A2(n19310), .ZN(n12828) );
  NAND2_X1 U16230 ( .A1(n12826), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12825) );
  OAI211_X1 U16231 ( .C1(n19373), .C2(n12829), .A(n12828), .B(n12825), .ZN(
        P2_U2981) );
  NAND2_X1 U16232 ( .A1(n12826), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12827) );
  OAI211_X1 U16233 ( .C1(n12830), .C2(n12829), .A(n12828), .B(n12827), .ZN(
        P2_U2966) );
  NAND2_X1 U16234 ( .A1(n14525), .A2(n12832), .ZN(n12833) );
  NAND2_X1 U16235 ( .A1(n12842), .A2(n12833), .ZN(n19242) );
  OAI211_X1 U16236 ( .C1(n12834), .C2(n12837), .A(n12836), .B(n15346), .ZN(
        n12839) );
  NAND2_X1 U16237 ( .A1(n15352), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12838) );
  OAI211_X1 U16238 ( .C1(n19242), .C2(n15352), .A(n12839), .B(n12838), .ZN(
        P2_U2879) );
  XNOR2_X1 U16239 ( .A(n12836), .B(n12840), .ZN(n12845) );
  NAND2_X1 U16240 ( .A1(n12842), .A2(n12841), .ZN(n12843) );
  AND2_X1 U16241 ( .A1(n13138), .A2(n12843), .ZN(n16458) );
  INV_X1 U16242 ( .A(n16458), .ZN(n15809) );
  MUX2_X1 U16243 ( .A(n15809), .B(n10898), .S(n15323), .Z(n12844) );
  OAI21_X1 U16244 ( .B1(n12845), .B2(n15359), .A(n12844), .ZN(P2_U2878) );
  NAND2_X1 U16245 ( .A1(n12972), .A2(n20254), .ZN(n12851) );
  XNOR2_X1 U16246 ( .A(n12978), .B(n12979), .ZN(n12849) );
  OR2_X1 U16247 ( .A1(n12847), .A2(n12846), .ZN(n12848) );
  AOI21_X1 U16248 ( .B1(n13786), .B2(n12849), .A(n12848), .ZN(n12850) );
  NAND2_X1 U16249 ( .A1(n12851), .A2(n12850), .ZN(n12948) );
  XNOR2_X1 U16250 ( .A(n12947), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13051) );
  INV_X1 U16251 ( .A(n13571), .ZN(n12856) );
  NAND2_X1 U16252 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12854) );
  INV_X1 U16253 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21013) );
  OR2_X1 U16254 ( .A1(n12853), .A2(n21013), .ZN(n13045) );
  OAI211_X1 U16255 ( .C1(n16110), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n12854), .B(n13045), .ZN(n12855) );
  AOI21_X1 U16256 ( .B1(n12856), .B2(n16105), .A(n12855), .ZN(n12857) );
  OAI21_X1 U16257 ( .B1(n13051), .B2(n20095), .A(n12857), .ZN(P1_U2998) );
  NAND2_X1 U16258 ( .A1(n12350), .A2(n13473), .ZN(n16286) );
  INV_X1 U16259 ( .A(n12858), .ZN(n12861) );
  NAND3_X1 U16260 ( .A1(n12861), .A2(n12860), .A3(n12859), .ZN(n12865) );
  NOR3_X1 U16261 ( .A1(n12863), .A2(n12862), .A3(n12909), .ZN(n12864) );
  NOR2_X1 U16262 ( .A1(n12865), .A2(n12864), .ZN(n14502) );
  INV_X1 U16263 ( .A(n14502), .ZN(n12940) );
  INV_X1 U16264 ( .A(n12866), .ZN(n12927) );
  NOR2_X1 U16265 ( .A1(n12868), .A2(n12867), .ZN(n12895) );
  NAND2_X1 U16266 ( .A1(n12895), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12871) );
  INV_X1 U16267 ( .A(n12869), .ZN(n12870) );
  NAND2_X1 U16268 ( .A1(n12871), .A2(n12870), .ZN(n12881) );
  INV_X1 U16269 ( .A(n11055), .ZN(n12876) );
  INV_X1 U16270 ( .A(n12872), .ZN(n12874) );
  NAND2_X1 U16271 ( .A1(n12874), .A2(n12873), .ZN(n12886) );
  INV_X1 U16272 ( .A(n12886), .ZN(n12875) );
  AOI21_X1 U16273 ( .B1(n12925), .B2(n12876), .A(n12875), .ZN(n12880) );
  NAND2_X1 U16274 ( .A1(n12887), .A2(n12883), .ZN(n12877) );
  AOI21_X1 U16275 ( .B1(n12925), .B2(n11055), .A(n12877), .ZN(n12879) );
  NAND2_X1 U16276 ( .A1(n12900), .A2(n12898), .ZN(n12891) );
  NAND2_X1 U16277 ( .A1(n12891), .A2(n12886), .ZN(n12878) );
  AOI22_X1 U16278 ( .A1(n12881), .A2(n12880), .B1(n12879), .B2(n12878), .ZN(
        n12882) );
  AOI21_X1 U16279 ( .B1(n15253), .B2(n12927), .A(n12882), .ZN(n20029) );
  NAND2_X1 U16280 ( .A1(n20029), .A2(n12940), .ZN(n12885) );
  NAND2_X1 U16281 ( .A1(n14502), .A2(n12883), .ZN(n12884) );
  NAND2_X1 U16282 ( .A1(n12885), .A2(n12884), .ZN(n12935) );
  NAND2_X1 U16283 ( .A1(n12887), .A2(n12886), .ZN(n12894) );
  NAND2_X1 U16284 ( .A1(n12888), .A2(n12927), .ZN(n12893) );
  NOR2_X1 U16285 ( .A1(n11055), .A2(n12889), .ZN(n12890) );
  AOI22_X1 U16286 ( .A1(n12891), .A2(n12894), .B1(n12890), .B2(n12925), .ZN(
        n12892) );
  OAI211_X1 U16287 ( .C1(n12895), .C2(n12894), .A(n12893), .B(n12892), .ZN(
        n14498) );
  MUX2_X1 U16288 ( .A(n14498), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n14502), .Z(n12931) );
  INV_X1 U16289 ( .A(n12931), .ZN(n12934) );
  INV_X1 U16290 ( .A(n12901), .ZN(n12899) );
  OAI22_X1 U16291 ( .A1(n12899), .A2(n12898), .B1(n12897), .B2(n12896), .ZN(
        n12903) );
  NOR2_X1 U16292 ( .A1(n12901), .A2(n12900), .ZN(n12902) );
  NOR2_X1 U16293 ( .A1(n12903), .A2(n12902), .ZN(n20083) );
  INV_X1 U16294 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n12904) );
  NAND2_X1 U16295 ( .A1(n12905), .A2(n12904), .ZN(n12912) );
  NAND2_X1 U16296 ( .A1(n12907), .A2(n12906), .ZN(n12908) );
  OR2_X1 U16297 ( .A1(n12909), .A2(n12908), .ZN(n15879) );
  OAI21_X1 U16298 ( .B1(n13118), .B2(n12910), .A(n15879), .ZN(n12911) );
  AOI21_X1 U16299 ( .B1(n12913), .B2(n12912), .A(n12911), .ZN(n12914) );
  OAI211_X1 U16300 ( .C1(n12935), .C2(n12934), .A(n20083), .B(n12914), .ZN(
        n12915) );
  INV_X1 U16301 ( .A(n12915), .ZN(n12939) );
  INV_X1 U16302 ( .A(n12925), .ZN(n12920) );
  INV_X1 U16303 ( .A(n12916), .ZN(n12917) );
  AND2_X1 U16304 ( .A1(n12918), .A2(n12917), .ZN(n12922) );
  XNOR2_X1 U16305 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12919) );
  OAI22_X1 U16306 ( .A1(n12920), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n12922), .B2(n12919), .ZN(n12921) );
  AOI21_X1 U16307 ( .B1(n19425), .B2(n12927), .A(n12921), .ZN(n15852) );
  INV_X1 U16308 ( .A(n15852), .ZN(n12930) );
  INV_X1 U16309 ( .A(n12922), .ZN(n12924) );
  MUX2_X1 U16310 ( .A(n12925), .B(n12924), .S(n12923), .Z(n12926) );
  AOI21_X1 U16311 ( .B1(n12928), .B2(n12927), .A(n12926), .ZN(n15847) );
  OAI211_X1 U16312 ( .C1(n15852), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15847), .ZN(n12929) );
  OAI211_X1 U16313 ( .C1(n12930), .C2(n20064), .A(n12929), .B(n12940), .ZN(
        n12933) );
  NOR2_X1 U16314 ( .A1(n12931), .A2(n20056), .ZN(n12932) );
  AOI211_X1 U16315 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n12935), .A(
        n12933), .B(n12932), .ZN(n12937) );
  NAND2_X1 U16316 ( .A1(n20048), .A2(n20056), .ZN(n19501) );
  OAI22_X1 U16317 ( .A1(n12935), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        n19501), .B2(n12934), .ZN(n12936) );
  OAI21_X1 U16318 ( .B1(n12937), .B2(n12936), .A(n15986), .ZN(n12938) );
  OAI211_X1 U16319 ( .C1(n12940), .C2(n15882), .A(n12939), .B(n12938), .ZN(
        n16569) );
  OAI21_X1 U16320 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n16569), .A(n16562), 
        .ZN(n12942) );
  OAI211_X1 U16321 ( .C1(n16286), .C2(n12943), .A(n12942), .B(n12941), .ZN(
        n16567) );
  INV_X1 U16322 ( .A(n16567), .ZN(n13036) );
  OAI21_X1 U16323 ( .B1(n13036), .B2(n11751), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12946) );
  NOR2_X1 U16324 ( .A1(n11751), .A2(n12944), .ZN(n16561) );
  INV_X1 U16325 ( .A(n16561), .ZN(n12945) );
  NAND2_X1 U16326 ( .A1(n12946), .A2(n12945), .ZN(P2_U3593) );
  NAND2_X1 U16327 ( .A1(n12947), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12952) );
  INV_X1 U16328 ( .A(n12948), .ZN(n12949) );
  OR2_X1 U16329 ( .A1(n12950), .A2(n12949), .ZN(n12951) );
  INV_X1 U16330 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13023) );
  NAND2_X1 U16332 ( .A1(n12955), .A2(n13166), .ZN(n13188) );
  AOI22_X1 U16333 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U16334 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12958) );
  INV_X2 U16335 ( .A(n12300), .ZN(n14199) );
  AOI22_X1 U16336 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U16337 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12956) );
  NAND4_X1 U16338 ( .A1(n12959), .A2(n12958), .A3(n12957), .A4(n12956), .ZN(
        n12965) );
  AOI22_X1 U16339 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14414), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U16340 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12962) );
  AOI22_X1 U16341 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12961) );
  AOI22_X1 U16342 ( .A1(n14352), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12960) );
  NAND4_X1 U16343 ( .A1(n12963), .A2(n12962), .A3(n12961), .A4(n12960), .ZN(
        n12964) );
  NOR2_X1 U16344 ( .A1(n12965), .A2(n12964), .ZN(n12982) );
  OAI22_X2 U16345 ( .A1(n13188), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12982), 
        .B2(n12966), .ZN(n12971) );
  INV_X1 U16346 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12968) );
  OAI22_X1 U16347 ( .A1(n12968), .A2(n13579), .B1(n12967), .B2(n12982), .ZN(
        n12969) );
  INV_X1 U16348 ( .A(n12969), .ZN(n12970) );
  XNOR2_X2 U16349 ( .A(n12971), .B(n12970), .ZN(n13238) );
  NAND2_X1 U16350 ( .A1(n12973), .A2(n12972), .ZN(n12977) );
  XNOR2_X2 U16351 ( .A(n13238), .B(n13237), .ZN(n13069) );
  INV_X1 U16352 ( .A(n13258), .ZN(n13781) );
  NAND2_X1 U16353 ( .A1(n13069), .A2(n13781), .ZN(n12987) );
  INV_X1 U16354 ( .A(n12978), .ZN(n12980) );
  NAND2_X1 U16355 ( .A1(n12980), .A2(n12979), .ZN(n12981) );
  NAND2_X1 U16356 ( .A1(n12981), .A2(n12982), .ZN(n13277) );
  OAI21_X1 U16357 ( .B1(n12982), .B2(n12981), .A(n13277), .ZN(n12985) );
  INV_X1 U16358 ( .A(n12983), .ZN(n12984) );
  AOI21_X1 U16359 ( .B1(n12985), .B2(n13786), .A(n12984), .ZN(n12986) );
  NAND2_X1 U16360 ( .A1(n12987), .A2(n12986), .ZN(n13232) );
  XNOR2_X1 U16361 ( .A(n13233), .B(n13232), .ZN(n13093) );
  NAND2_X1 U16362 ( .A1(n20254), .A2(n15979), .ZN(n12989) );
  NAND2_X1 U16363 ( .A1(n12989), .A2(n12988), .ZN(n12995) );
  AOI21_X1 U16364 ( .B1(n12429), .B2(n20902), .A(n13364), .ZN(n12991) );
  NOR2_X1 U16365 ( .A1(n20905), .A2(n13365), .ZN(n12990) );
  OAI21_X1 U16366 ( .B1(n12991), .B2(n12990), .A(n14446), .ZN(n12992) );
  NAND2_X1 U16367 ( .A1(n12992), .A2(n10073), .ZN(n12994) );
  MUX2_X1 U16368 ( .A(n12995), .B(n12994), .S(n12993), .Z(n13000) );
  INV_X1 U16369 ( .A(n15164), .ZN(n12996) );
  NAND3_X1 U16370 ( .A1(n12997), .A2(n12996), .A3(n20254), .ZN(n12998) );
  NAND3_X1 U16371 ( .A1(n13000), .A2(n12999), .A3(n12998), .ZN(n13001) );
  INV_X1 U16372 ( .A(n13019), .ZN(n13003) );
  NAND2_X1 U16373 ( .A1(n13003), .A2(n13002), .ZN(n13004) );
  AND2_X1 U16374 ( .A1(n13171), .A2(n13004), .ZN(n13006) );
  NAND4_X1 U16375 ( .A1(n13007), .A2(n13006), .A3(n13108), .A4(n15942), .ZN(
        n13008) );
  AOI21_X1 U16376 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13630) );
  NAND2_X1 U16377 ( .A1(n16205), .A2(n13630), .ZN(n13285) );
  NAND2_X1 U16378 ( .A1(n13021), .A2(n15925), .ZN(n16133) );
  OAI211_X1 U16379 ( .C1(n13011), .C2(n20238), .A(n13010), .B(n13009), .ZN(
        n13012) );
  NAND2_X1 U16380 ( .A1(n13021), .A2(n13012), .ZN(n16136) );
  OR2_X1 U16381 ( .A1(n16136), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13013) );
  OR2_X1 U16382 ( .A1(n13021), .A2(n16255), .ZN(n16129) );
  OAI21_X1 U16383 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n16201), .A(
        n13038), .ZN(n13032) );
  INV_X1 U16384 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13014) );
  OR2_X1 U16385 ( .A1(n12853), .A2(n13014), .ZN(n13018) );
  NAND4_X1 U16386 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A4(n16205), .ZN(n13017) );
  INV_X1 U16387 ( .A(n16133), .ZN(n13015) );
  NOR2_X1 U16388 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13015), .ZN(
        n13047) );
  OR3_X1 U16389 ( .A1(n12760), .A2(n16206), .A3(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13016) );
  NAND3_X1 U16390 ( .A1(n13018), .A2(n13017), .A3(n13016), .ZN(n13031) );
  OAI22_X1 U16391 ( .A1(n12299), .A2(n20254), .B1(n13002), .B2(n13019), .ZN(
        n13020) );
  NAND2_X1 U16392 ( .A1(n14591), .A2(n13023), .ZN(n13024) );
  OAI211_X1 U16393 ( .C1(n14593), .C2(P1_EBX_REG_2__SCAN_IN), .A(n14614), .B(
        n13024), .ZN(n13026) );
  INV_X1 U16394 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13075) );
  NAND2_X1 U16395 ( .A1(n9804), .A2(n13075), .ZN(n13025) );
  AND2_X1 U16396 ( .A1(n13026), .A2(n13025), .ZN(n13027) );
  NAND2_X1 U16397 ( .A1(n13028), .A2(n13027), .ZN(n13029) );
  NAND2_X1 U16398 ( .A1(n13411), .A2(n13029), .ZN(n13362) );
  NOR2_X1 U16399 ( .A1(n16242), .A2(n13362), .ZN(n13030) );
  AOI211_X1 U16400 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n13032), .A(
        n13031), .B(n13030), .ZN(n13033) );
  OAI211_X1 U16401 ( .C1(n13093), .C2(n16215), .A(n13285), .B(n13033), .ZN(
        P1_U3029) );
  NOR2_X1 U16402 ( .A1(n19951), .A2(n11751), .ZN(n15984) );
  AOI21_X1 U16403 ( .B1(n15984), .B2(n20035), .A(n16570), .ZN(n13035) );
  NOR2_X1 U16404 ( .A1(n11751), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19103) );
  OAI211_X1 U16405 ( .C1(n13036), .C2(n19103), .A(n19951), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n13034) );
  NAND4_X1 U16406 ( .A1(n20067), .A2(n11751), .A3(n12350), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19301) );
  OAI211_X1 U16407 ( .C1(n13036), .C2(n13035), .A(n13034), .B(n19301), .ZN(
        P2_U3177) );
  INV_X1 U16408 ( .A(n13037), .ZN(n13042) );
  AOI21_X1 U16409 ( .B1(n16205), .B2(n15170), .A(n16202), .ZN(n13046) );
  INV_X1 U16410 ( .A(n16136), .ZN(n13039) );
  NOR3_X1 U16411 ( .A1(n16205), .A2(n13039), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13040) );
  AOI21_X1 U16412 ( .B1(n13046), .B2(n16133), .A(n13040), .ZN(n13041) );
  AOI211_X1 U16413 ( .C1(n16263), .C2(n13502), .A(n13042), .B(n13041), .ZN(
        n13043) );
  OAI21_X1 U16414 ( .B1(n13044), .B2(n16215), .A(n13043), .ZN(P1_U3031) );
  OAI21_X1 U16415 ( .B1(n13046), .B2(n12760), .A(n13045), .ZN(n13049) );
  NAND2_X1 U16416 ( .A1(n16201), .A2(n16130), .ZN(n16161) );
  INV_X1 U16417 ( .A(n16161), .ZN(n15044) );
  NOR3_X1 U16418 ( .A1(n15044), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13047), .ZN(n13048) );
  AOI211_X1 U16419 ( .C1(n16263), .C2(n13565), .A(n13049), .B(n13048), .ZN(
        n13050) );
  OAI21_X1 U16420 ( .B1(n13051), .B2(n16215), .A(n13050), .ZN(P1_U3030) );
  XOR2_X1 U16421 ( .A(n13053), .B(n13052), .Z(n15825) );
  INV_X1 U16422 ( .A(n15825), .ZN(n19258) );
  OR2_X1 U16423 ( .A1(n19361), .A2(n19360), .ZN(n19324) );
  INV_X1 U16424 ( .A(n19324), .ZN(n19318) );
  INV_X1 U16425 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19388) );
  OAI222_X1 U16426 ( .A1(n19258), .A2(n19318), .B1(n19333), .B2(n19388), .C1(
        n19367), .C2(n19463), .ZN(P2_U2912) );
  AOI21_X1 U16427 ( .B1(n13055), .B2(n13062), .A(n9919), .ZN(n15806) );
  INV_X1 U16428 ( .A(n15806), .ZN(n13057) );
  INV_X1 U16429 ( .A(n15395), .ZN(n13056) );
  OAI222_X1 U16430 ( .A1(n13057), .A2(n19318), .B1(n13056), .B2(n19367), .C1(
        n11320), .C2(n19333), .ZN(P2_U2910) );
  OR2_X1 U16431 ( .A1(n13058), .A2(n9919), .ZN(n13059) );
  NAND2_X1 U16432 ( .A1(n13059), .A2(n15222), .ZN(n19235) );
  INV_X1 U16433 ( .A(n15387), .ZN(n13060) );
  INV_X1 U16434 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19382) );
  OAI222_X1 U16435 ( .A1(n19235), .A2(n19318), .B1(n13060), .B2(n19367), .C1(
        n19382), .C2(n19333), .ZN(P2_U2909) );
  OR2_X1 U16436 ( .A1(n13061), .A2(n9922), .ZN(n13063) );
  NAND2_X1 U16437 ( .A1(n13063), .A2(n13062), .ZN(n19249) );
  INV_X1 U16438 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19386) );
  OAI222_X1 U16439 ( .A1(n19249), .A2(n19318), .B1(n15403), .B2(n19367), .C1(
        n19386), .C2(n19333), .ZN(P2_U2911) );
  NAND2_X1 U16440 ( .A1(n14439), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13325) );
  INV_X1 U16441 ( .A(n13325), .ZN(n13068) );
  INV_X2 U16442 ( .A(n14363), .ZN(n14437) );
  XNOR2_X1 U16443 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13363) );
  AOI21_X1 U16444 ( .B1(n14437), .B2(n13363), .A(n14439), .ZN(n13065) );
  NAND2_X1 U16445 ( .A1(n14250), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n13064) );
  OAI211_X1 U16446 ( .C1(n13333), .C2(n13175), .A(n13065), .B(n13064), .ZN(
        n13066) );
  INV_X1 U16447 ( .A(n13066), .ZN(n13067) );
  INV_X1 U16448 ( .A(n13326), .ZN(n13072) );
  AOI21_X1 U16449 ( .B1(n13074), .B2(n13073), .A(n13072), .ZN(n13116) );
  INV_X1 U16450 ( .A(n14803), .ZN(n20182) );
  OAI22_X1 U16451 ( .A1(n20171), .A2(n13362), .B1(n13075), .B2(n20185), .ZN(
        n13076) );
  AOI21_X1 U16452 ( .B1(n13116), .B2(n20182), .A(n13076), .ZN(n13077) );
  INV_X1 U16453 ( .A(n13077), .ZN(P1_U2870) );
  AOI22_X1 U16454 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20210), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15982), .ZN(n13078) );
  OAI21_X1 U16455 ( .B1(n13079), .B2(n13087), .A(n13078), .ZN(P1_U2906) );
  OR2_X1 U16456 ( .A1(n13080), .A2(n15224), .ZN(n13081) );
  NAND2_X1 U16457 ( .A1(n13081), .A2(n13226), .ZN(n19224) );
  INV_X1 U16458 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19378) );
  OAI222_X1 U16459 ( .A1(n19224), .A2(n19318), .B1(n15369), .B2(n19367), .C1(
        n19378), .C2(n19333), .ZN(P2_U2907) );
  INV_X1 U16460 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U16461 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13082) );
  OAI21_X1 U16462 ( .B1(n13083), .B2(n13087), .A(n13082), .ZN(P1_U2919) );
  INV_X1 U16463 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14860) );
  AOI22_X1 U16464 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13084) );
  OAI21_X1 U16465 ( .B1(n14860), .B2(n13087), .A(n13084), .ZN(P1_U2920) );
  AOI22_X1 U16466 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13085) );
  OAI21_X1 U16467 ( .B1(n21206), .B2(n13087), .A(n13085), .ZN(P1_U2910) );
  INV_X1 U16468 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13088) );
  AOI22_X1 U16469 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13086) );
  OAI21_X1 U16470 ( .B1(n13088), .B2(n13087), .A(n13086), .ZN(P1_U2918) );
  NOR2_X1 U16471 ( .A1(n16110), .A2(n13363), .ZN(n13091) );
  INV_X1 U16472 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13089) );
  OAI22_X1 U16473 ( .A1(n16116), .A2(n13089), .B1(n12853), .B2(n13014), .ZN(
        n13090) );
  AOI211_X1 U16474 ( .C1(n13116), .C2(n16105), .A(n13091), .B(n13090), .ZN(
        n13092) );
  OAI21_X1 U16475 ( .B1(n20095), .B2(n13093), .A(n13092), .ZN(P1_U2997) );
  NOR2_X1 U16476 ( .A1(n19326), .A2(n12350), .ZN(n19585) );
  INV_X1 U16477 ( .A(n19585), .ZN(n20043) );
  NAND2_X1 U16478 ( .A1(n20048), .A2(n13695), .ZN(n19620) );
  OAI21_X1 U16479 ( .B1(n20043), .B2(n20041), .A(n19620), .ZN(n13096) );
  NOR2_X1 U16480 ( .A1(n20074), .A2(n19620), .ZN(n19673) );
  OR3_X1 U16481 ( .A1(n13094), .A2(n19673), .A3(n20067), .ZN(n13099) );
  INV_X1 U16482 ( .A(n19673), .ZN(n19670) );
  NAND2_X1 U16483 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19670), .ZN(n13095) );
  NAND4_X1 U16484 ( .A1(n13096), .A2(n19737), .A3(n13099), .A4(n13095), .ZN(
        n19662) );
  INV_X1 U16485 ( .A(n19662), .ZN(n13122) );
  INV_X1 U16486 ( .A(n19697), .ZN(n19689) );
  AOI22_X1 U16487 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19466), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19465), .ZN(n19925) );
  INV_X1 U16488 ( .A(n19925), .ZN(n19870) );
  NOR2_X2 U16489 ( .A1(n20041), .A2(n19557), .ZN(n19658) );
  AOI22_X1 U16490 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19466), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19465), .ZN(n19826) );
  AOI22_X1 U16491 ( .A1(n19689), .A2(n19870), .B1(n19658), .B2(n19922), .ZN(
        n13103) );
  NOR2_X1 U16492 ( .A1(n13298), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19474) );
  INV_X1 U16493 ( .A(n13099), .ZN(n13100) );
  AOI211_X2 U16494 ( .C1(n19620), .C2(n20067), .A(n19474), .B(n13100), .ZN(
        n19661) );
  NOR2_X2 U16495 ( .A1(n10560), .A2(n19459), .ZN(n19921) );
  AOI22_X1 U16496 ( .A1(n19661), .A2(n13101), .B1(n19673), .B2(n19921), .ZN(
        n13102) );
  OAI211_X1 U16497 ( .C1(n13122), .C2(n13104), .A(n13103), .B(n13102), .ZN(
        P2_U3110) );
  OAI22_X1 U16498 ( .A1(n13108), .A2(n13107), .B1(n13106), .B2(n13105), .ZN(
        n13110) );
  NAND2_X1 U16499 ( .A1(n13114), .A2(n13113), .ZN(n13115) );
  INV_X1 U16500 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20213) );
  OAI222_X1 U16501 ( .A1(n14881), .A2(n13507), .B1(n14879), .B2(n20213), .C1(
        n14878), .C2(n20244), .ZN(P1_U2904) );
  INV_X1 U16502 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20209) );
  OAI222_X1 U16503 ( .A1(n14881), .A2(n13571), .B1(n14879), .B2(n20209), .C1(
        n14878), .C2(n20255), .ZN(P1_U2903) );
  INV_X1 U16504 ( .A(n13116), .ZN(n13381) );
  INV_X1 U16505 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20207) );
  OAI222_X1 U16506 ( .A1(n14881), .A2(n13381), .B1(n14879), .B2(n20207), .C1(
        n14878), .C2(n20262), .ZN(P1_U2902) );
  INV_X1 U16507 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U16508 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19466), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19465), .ZN(n19897) );
  INV_X1 U16509 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20235) );
  INV_X1 U16510 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18442) );
  AOI22_X1 U16511 ( .A1(n19689), .A2(n19805), .B1(n19658), .B2(n19894), .ZN(
        n13120) );
  NOR2_X2 U16512 ( .A1(n13118), .A2(n19459), .ZN(n19885) );
  AOI22_X1 U16513 ( .A1(n19661), .A2(n13117), .B1(n19885), .B2(n19673), .ZN(
        n13119) );
  OAI211_X1 U16514 ( .C1(n13122), .C2(n13121), .A(n13120), .B(n13119), .ZN(
        P2_U3104) );
  INV_X1 U16515 ( .A(n19596), .ZN(n19584) );
  NOR3_X1 U16516 ( .A1(n20056), .A2(n20048), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19796) );
  AOI21_X1 U16517 ( .B1(n19891), .B2(n19584), .A(n19796), .ZN(n13126) );
  NAND2_X1 U16518 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19796), .ZN(
        n13130) );
  AND2_X1 U16519 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13130), .ZN(n13123) );
  AND2_X1 U16520 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n13130), .ZN(n13125) );
  NOR4_X2 U16521 ( .A1(n13126), .A2(n19888), .A3(n13129), .A4(n13125), .ZN(
        n19852) );
  INV_X1 U16522 ( .A(n19760), .ZN(n13127) );
  NOR2_X2 U16523 ( .A1(n13127), .A2(n19596), .ZN(n19874) );
  NOR2_X2 U16524 ( .A1(n19733), .A2(n19596), .ZN(n19848) );
  AOI22_X1 U16525 ( .A1(n19874), .A2(n19805), .B1(n19848), .B2(n19894), .ZN(
        n13132) );
  AOI21_X1 U16526 ( .B1(n13298), .B2(n19796), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13128) );
  NOR2_X1 U16527 ( .A1(n13129), .A2(n13128), .ZN(n19847) );
  INV_X1 U16528 ( .A(n13130), .ZN(n19846) );
  AOI22_X1 U16529 ( .A1(n19847), .A2(n13117), .B1(n19885), .B2(n19846), .ZN(
        n13131) );
  OAI211_X1 U16530 ( .C1(n19852), .C2(n13133), .A(n13132), .B(n13131), .ZN(
        P2_U3152) );
  OAI211_X1 U16531 ( .C1(n13134), .C2(n13136), .A(n13135), .B(n15346), .ZN(
        n13141) );
  AND2_X1 U16532 ( .A1(n13138), .A2(n13137), .ZN(n13139) );
  NAND2_X1 U16533 ( .A1(n9912), .A2(n15356), .ZN(n13140) );
  OAI211_X1 U16534 ( .C1(n15356), .C2(n13142), .A(n13141), .B(n13140), .ZN(
        P2_U2877) );
  XNOR2_X1 U16535 ( .A(n13135), .B(n13384), .ZN(n13149) );
  OR2_X1 U16536 ( .A1(n13144), .A2(n13143), .ZN(n13145) );
  AND2_X1 U16537 ( .A1(n13145), .A2(n13387), .ZN(n16539) );
  NOR2_X1 U16538 ( .A1(n15356), .A2(n13146), .ZN(n13147) );
  AOI21_X1 U16539 ( .B1(n16539), .B2(n15356), .A(n13147), .ZN(n13148) );
  OAI21_X1 U16540 ( .B1(n13149), .B2(n15359), .A(n13148), .ZN(P2_U2876) );
  XNOR2_X1 U16541 ( .A(n13150), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13151) );
  XNOR2_X1 U16542 ( .A(n13152), .B(n13151), .ZN(n13324) );
  XNOR2_X1 U16543 ( .A(n13154), .B(n13153), .ZN(n13320) );
  INV_X1 U16544 ( .A(n13320), .ZN(n13164) );
  AND2_X1 U16545 ( .A1(n13155), .A2(n19427), .ZN(n13157) );
  MUX2_X1 U16546 ( .A(n13157), .B(n13156), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13163) );
  INV_X1 U16547 ( .A(n15253), .ZN(n13161) );
  NAND2_X1 U16548 ( .A1(n19404), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n13318) );
  AOI21_X1 U16549 ( .B1(n13159), .B2(n13158), .A(n19269), .ZN(n20046) );
  NAND2_X1 U16550 ( .A1(n19420), .A2(n20046), .ZN(n13160) );
  OAI211_X1 U16551 ( .C1(n13161), .C2(n19411), .A(n13318), .B(n13160), .ZN(
        n13162) );
  AOI211_X1 U16552 ( .C1(n13164), .C2(n19429), .A(n13163), .B(n13162), .ZN(
        n13165) );
  OAI21_X1 U16553 ( .B1(n19436), .B2(n13324), .A(n13165), .ZN(P2_U3043) );
  INV_X1 U16554 ( .A(n13167), .ZN(n15160) );
  NAND2_X1 U16555 ( .A1(n15160), .A2(n13168), .ZN(n13197) );
  NOR2_X1 U16556 ( .A1(n13169), .A2(n13332), .ZN(n13170) );
  NOR2_X1 U16557 ( .A1(n12660), .A2(n13170), .ZN(n20865) );
  INV_X1 U16558 ( .A(n13171), .ZN(n13173) );
  OR2_X1 U16559 ( .A1(n13173), .A2(n13172), .ZN(n13195) );
  INV_X1 U16560 ( .A(n15172), .ZN(n15161) );
  NAND2_X1 U16561 ( .A1(n15161), .A2(n13175), .ZN(n13190) );
  NAND2_X1 U16562 ( .A1(n13190), .A2(n13332), .ZN(n13178) );
  INV_X1 U16563 ( .A(n13176), .ZN(n13177) );
  AOI22_X1 U16564 ( .A1(n13178), .A2(n13177), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n15172), .ZN(n13180) );
  XNOR2_X1 U16565 ( .A(n13192), .B(n13332), .ZN(n13179) );
  AOI22_X1 U16566 ( .A1(n13195), .A2(n13180), .B1(n15925), .B2(n13179), .ZN(
        n13181) );
  OAI21_X1 U16567 ( .B1(n13197), .B2(n20865), .A(n13181), .ZN(n13182) );
  INV_X1 U16568 ( .A(n13182), .ZN(n13183) );
  NAND2_X1 U16569 ( .A1(n13184), .A2(n13183), .ZN(n20864) );
  NAND2_X1 U16570 ( .A1(n20864), .A2(n15928), .ZN(n13187) );
  INV_X1 U16571 ( .A(n15928), .ZN(n13185) );
  NAND2_X1 U16572 ( .A1(n13185), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13186) );
  NAND2_X1 U16573 ( .A1(n13187), .A2(n13186), .ZN(n15936) );
  NAND2_X1 U16574 ( .A1(n15936), .A2(n16272), .ZN(n13202) );
  NOR2_X1 U16575 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16272), .ZN(n13207) );
  NAND2_X1 U16576 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13207), .ZN(
        n13201) );
  INV_X1 U16577 ( .A(n13169), .ZN(n13191) );
  NAND2_X1 U16578 ( .A1(n13191), .A2(n13190), .ZN(n20874) );
  NOR2_X1 U16579 ( .A1(n13193), .A2(n13192), .ZN(n13194) );
  AOI22_X1 U16580 ( .A1(n13195), .A2(n20874), .B1(n15925), .B2(n13194), .ZN(
        n13196) );
  OAI21_X1 U16581 ( .B1(n13197), .B2(n20874), .A(n13196), .ZN(n13198) );
  INV_X1 U16582 ( .A(n13198), .ZN(n13199) );
  OAI21_X1 U16583 ( .B1(n13189), .B2(n15160), .A(n13199), .ZN(n20869) );
  MUX2_X1 U16584 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n20869), .S(
        n15928), .Z(n15935) );
  AOI22_X1 U16585 ( .A1(n13207), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16272), .B2(n15935), .ZN(n13200) );
  AOI21_X1 U16586 ( .B1(n13202), .B2(n13201), .A(n13200), .ZN(n15947) );
  INV_X1 U16587 ( .A(n15173), .ZN(n15162) );
  AND2_X1 U16588 ( .A1(n15947), .A2(n15162), .ZN(n13222) );
  NAND2_X1 U16589 ( .A1(n20152), .A2(n13203), .ZN(n13204) );
  OAI21_X1 U16590 ( .B1(n15928), .B2(n13205), .A(n13204), .ZN(n13206) );
  NAND2_X1 U16591 ( .A1(n13206), .A2(n16272), .ZN(n13209) );
  NAND2_X1 U16592 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13207), .ZN(
        n13208) );
  NAND2_X1 U16593 ( .A1(n13209), .A2(n13208), .ZN(n15946) );
  NOR3_X1 U16594 ( .A1(n13222), .A2(n15946), .A3(P1_FLUSH_REG_SCAN_IN), .ZN(
        n13210) );
  NOR2_X1 U16595 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20906) );
  AND2_X1 U16596 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20637), .ZN(n20880) );
  NAND2_X1 U16597 ( .A1(n9811), .A2(n20885), .ZN(n20599) );
  OR2_X1 U16598 ( .A1(n9811), .A2(n20747), .ZN(n13212) );
  NAND2_X1 U16599 ( .A1(n20703), .A2(n20625), .ZN(n20882) );
  AND2_X1 U16600 ( .A1(n13212), .A2(n20882), .ZN(n20745) );
  MUX2_X1 U16601 ( .A(n20599), .B(n20745), .S(n13069), .Z(n13213) );
  OAI21_X1 U16602 ( .B1(n20880), .B2(n13189), .A(n13213), .ZN(n13214) );
  NAND2_X1 U16603 ( .A1(n20892), .A2(n13214), .ZN(n13215) );
  OAI21_X1 U16604 ( .B1(n20892), .B2(n12471), .A(n13215), .ZN(P1_U3476) );
  NOR2_X1 U16605 ( .A1(n20702), .A2(n20880), .ZN(n13219) );
  INV_X1 U16606 ( .A(n20882), .ZN(n13217) );
  MUX2_X1 U16607 ( .A(n20885), .B(n13217), .S(n9811), .Z(n13218) );
  OAI21_X1 U16608 ( .B1(n13219), .B2(n13218), .A(n20892), .ZN(n13220) );
  OAI21_X1 U16609 ( .B1(n20631), .B2(n20892), .A(n13220), .ZN(P1_U3477) );
  INV_X1 U16610 ( .A(n16276), .ZN(n13221) );
  NOR3_X1 U16611 ( .A1(n13222), .A2(n15946), .A3(n13221), .ZN(n15953) );
  INV_X1 U16612 ( .A(n12646), .ZN(n13223) );
  OAI22_X1 U16613 ( .A1(n20329), .A2(n20747), .B1(n13223), .B2(n20880), .ZN(
        n13224) );
  OAI21_X1 U16614 ( .B1(n15953), .B2(n13224), .A(n20892), .ZN(n13225) );
  OAI21_X1 U16615 ( .B1(n20892), .B2(n20670), .A(n13225), .ZN(P1_U3478) );
  NAND2_X1 U16616 ( .A1(n13227), .A2(n13226), .ZN(n13230) );
  INV_X1 U16617 ( .A(n13228), .ZN(n13229) );
  NAND2_X1 U16618 ( .A1(n13230), .A2(n13229), .ZN(n19201) );
  INV_X1 U16619 ( .A(n15362), .ZN(n13231) );
  OAI222_X1 U16620 ( .A1(n19201), .A2(n19318), .B1(n13231), .B2(n19367), .C1(
        n19375), .C2(n19333), .ZN(P2_U2906) );
  NAND2_X1 U16621 ( .A1(n13233), .A2(n13232), .ZN(n13236) );
  NAND2_X1 U16622 ( .A1(n13234), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13235) );
  NAND2_X1 U16623 ( .A1(n13236), .A2(n13235), .ZN(n13339) );
  INV_X1 U16624 ( .A(n13237), .ZN(n13239) );
  INV_X1 U16625 ( .A(n13253), .ZN(n13252) );
  AOI22_X1 U16626 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U16627 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16628 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13241) );
  AOI22_X1 U16629 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13240) );
  NAND4_X1 U16630 ( .A1(n13243), .A2(n13242), .A3(n13241), .A4(n13240), .ZN(
        n13249) );
  AOI22_X1 U16631 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14422), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U16632 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13246) );
  AOI22_X1 U16633 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13245) );
  AOI22_X1 U16634 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13244) );
  NAND4_X1 U16635 ( .A1(n13247), .A2(n13246), .A3(n13245), .A4(n13244), .ZN(
        n13248) );
  AOI22_X1 U16636 ( .A1(n13576), .A2(n13276), .B1(n13530), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13250) );
  INV_X1 U16637 ( .A(n20233), .ZN(n20389) );
  NAND2_X1 U16638 ( .A1(n13252), .A2(n20389), .ZN(n13254) );
  INV_X1 U16639 ( .A(n13276), .ZN(n13255) );
  XNOR2_X1 U16640 ( .A(n13277), .B(n13255), .ZN(n13256) );
  NAND2_X1 U16641 ( .A1(n13256), .A2(n13786), .ZN(n13257) );
  OAI21_X1 U16642 ( .B1(n20883), .B2(n13258), .A(n13257), .ZN(n13260) );
  INV_X1 U16643 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13259) );
  XNOR2_X1 U16644 ( .A(n13260), .B(n13259), .ZN(n13338) );
  NAND2_X1 U16645 ( .A1(n13339), .A2(n13338), .ZN(n13262) );
  NAND2_X1 U16646 ( .A1(n13260), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13261) );
  AOI22_X1 U16647 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13267) );
  AOI22_X1 U16648 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13266) );
  AOI22_X1 U16649 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13265) );
  AOI22_X1 U16650 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13264) );
  NAND4_X1 U16651 ( .A1(n13267), .A2(n13266), .A3(n13265), .A4(n13264), .ZN(
        n13273) );
  AOI22_X1 U16652 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14414), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13271) );
  AOI22_X1 U16653 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13270) );
  AOI22_X1 U16654 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13269) );
  AOI22_X1 U16655 ( .A1(n14352), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13268) );
  NAND4_X1 U16656 ( .A1(n13271), .A2(n13270), .A3(n13269), .A4(n13268), .ZN(
        n13272) );
  NAND2_X1 U16657 ( .A1(n13576), .A2(n13280), .ZN(n13275) );
  NAND2_X1 U16658 ( .A1(n13530), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13274) );
  NAND2_X1 U16659 ( .A1(n13275), .A2(n13274), .ZN(n13431) );
  XNOR2_X1 U16660 ( .A(n13433), .B(n13431), .ZN(n13409) );
  NAND2_X1 U16661 ( .A1(n13409), .A2(n13781), .ZN(n13283) );
  NAND2_X1 U16662 ( .A1(n13277), .A2(n13276), .ZN(n13279) );
  INV_X1 U16663 ( .A(n13279), .ZN(n13281) );
  INV_X1 U16664 ( .A(n13280), .ZN(n13278) );
  OR2_X1 U16665 ( .A1(n13279), .A2(n13278), .ZN(n13621) );
  OAI211_X1 U16666 ( .C1(n13281), .C2(n13280), .A(n13786), .B(n13621), .ZN(
        n13282) );
  NAND2_X1 U16667 ( .A1(n13283), .A2(n13282), .ZN(n13608) );
  INV_X1 U16668 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13284) );
  XNOR2_X1 U16669 ( .A(n13608), .B(n13284), .ZN(n13606) );
  XNOR2_X1 U16670 ( .A(n13607), .B(n13606), .ZN(n13429) );
  INV_X1 U16671 ( .A(n16201), .ZN(n15038) );
  NAND2_X1 U16672 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15026) );
  AOI21_X1 U16673 ( .B1(n15038), .B2(n15026), .A(n16202), .ZN(n16225) );
  NAND2_X1 U16674 ( .A1(n16225), .A2(n13285), .ZN(n15154) );
  INV_X1 U16675 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20823) );
  NOR2_X1 U16676 ( .A1(n12853), .A2(n20823), .ZN(n13424) );
  MUX2_X1 U16677 ( .A(n14586), .B(n9804), .S(P1_EBX_REG_3__SCAN_IN), .Z(n13286) );
  INV_X1 U16678 ( .A(n13286), .ZN(n13288) );
  NAND2_X1 U16679 ( .A1(n14567), .A2(n13259), .ZN(n13287) );
  NAND2_X1 U16680 ( .A1(n13288), .A2(n13287), .ZN(n13410) );
  MUX2_X1 U16681 ( .A(n9804), .B(n10135), .S(P1_EBX_REG_4__SCAN_IN), .Z(n13289) );
  INV_X1 U16682 ( .A(n13289), .ZN(n13291) );
  NAND2_X1 U16683 ( .A1(n14593), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13290) );
  NAND2_X1 U16684 ( .A1(n13291), .A2(n13290), .ZN(n13292) );
  OR2_X1 U16685 ( .A1(n13413), .A2(n13292), .ZN(n13293) );
  NAND2_X1 U16686 ( .A1(n13462), .A2(n13293), .ZN(n20163) );
  NOR2_X1 U16687 ( .A1(n16242), .A2(n20163), .ZN(n13294) );
  AOI211_X1 U16688 ( .C1(n15154), .C2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13424), .B(n13294), .ZN(n13296) );
  OAI22_X1 U16689 ( .A1(n13630), .A2(n16130), .B1(n15026), .B2(n16206), .ZN(
        n15153) );
  NAND2_X1 U16690 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13632) );
  OAI211_X1 U16691 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n15153), .B(n13632), .ZN(n13295) );
  OAI211_X1 U16692 ( .C1(n13429), .C2(n16215), .A(n13296), .B(n13295), .ZN(
        P1_U3027) );
  NAND2_X1 U16693 ( .A1(n19585), .A2(n19771), .ZN(n13297) );
  OR2_X1 U16694 ( .A1(n20064), .A2(n19501), .ZN(n13306) );
  NAND2_X1 U16695 ( .A1(n13297), .A2(n13306), .ZN(n13304) );
  NAND2_X1 U16696 ( .A1(n10762), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13299) );
  NAND2_X1 U16697 ( .A1(n13299), .A2(n13298), .ZN(n13302) );
  INV_X1 U16698 ( .A(n13300), .ZN(n19762) );
  INV_X1 U16699 ( .A(n19501), .ZN(n13301) );
  NAND2_X1 U16700 ( .A1(n19762), .A2(n13301), .ZN(n13308) );
  AOI21_X1 U16701 ( .B1(n13302), .B2(n13308), .A(n19888), .ZN(n13303) );
  NAND2_X1 U16702 ( .A1(n13304), .A2(n13303), .ZN(n19549) );
  INV_X1 U16703 ( .A(n19549), .ZN(n19534) );
  INV_X1 U16704 ( .A(n13306), .ZN(n13307) );
  NAND2_X1 U16705 ( .A1(n13307), .A2(n20037), .ZN(n13311) );
  INV_X1 U16706 ( .A(n10762), .ZN(n13309) );
  INV_X1 U16707 ( .A(n13308), .ZN(n19546) );
  OAI21_X1 U16708 ( .B1(n13309), .B2(n19546), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13310) );
  NAND2_X1 U16709 ( .A1(n13311), .A2(n13310), .ZN(n19548) );
  AOI22_X1 U16710 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19466), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19465), .ZN(n19823) );
  INV_X1 U16711 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20277) );
  INV_X1 U16712 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18470) );
  OAI22_X1 U16713 ( .A1(n20277), .A2(n19458), .B1(n18470), .B2(n19456), .ZN(
        n19867) );
  AOI22_X1 U16714 ( .A1(n19574), .A2(n19867), .B1(n13312), .B2(n19546), .ZN(
        n13313) );
  OAI21_X1 U16715 ( .B1(n19541), .B2(n19823), .A(n13313), .ZN(n13314) );
  AOI21_X1 U16716 ( .B1(n13305), .B2(n19548), .A(n13314), .ZN(n13315) );
  OAI21_X1 U16717 ( .B1(n19534), .B2(n13316), .A(n13315), .ZN(P2_U3077) );
  AOI21_X1 U16718 ( .B1(n15250), .B2(n13317), .A(n13467), .ZN(n15246) );
  NAND2_X1 U16719 ( .A1(n16488), .A2(n15246), .ZN(n13319) );
  OAI211_X1 U16720 ( .C1(n15250), .C2(n16498), .A(n13319), .B(n13318), .ZN(
        n13322) );
  NOR2_X1 U16721 ( .A1(n13320), .A2(n16478), .ZN(n13321) );
  AOI211_X1 U16722 ( .C1(n16491), .C2(n15253), .A(n13322), .B(n13321), .ZN(
        n13323) );
  OAI21_X1 U16723 ( .B1(n16480), .B2(n13324), .A(n13323), .ZN(P2_U3011) );
  INV_X1 U16724 ( .A(n16105), .ZN(n16111) );
  INV_X1 U16725 ( .A(n13327), .ZN(n13329) );
  INV_X1 U16726 ( .A(n13404), .ZN(n13328) );
  OAI21_X1 U16727 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13329), .A(
        n13328), .ZN(n13414) );
  AOI22_X1 U16728 ( .A1(n14437), .A2(n13414), .B1(n14439), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13331) );
  NAND2_X1 U16729 ( .A1(n14250), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n13330) );
  OAI211_X1 U16730 ( .C1(n13333), .C2(n13332), .A(n13331), .B(n13330), .ZN(
        n13334) );
  INV_X1 U16731 ( .A(n13334), .ZN(n13335) );
  NAND2_X1 U16732 ( .A1(n13336), .A2(n13337), .ZN(n13430) );
  OAI21_X1 U16733 ( .B1(n13337), .B2(n13336), .A(n13430), .ZN(n20179) );
  XOR2_X1 U16734 ( .A(n13339), .B(n13338), .Z(n15152) );
  INV_X1 U16735 ( .A(n20095), .ZN(n16113) );
  NAND2_X1 U16736 ( .A1(n15152), .A2(n16113), .ZN(n13342) );
  INV_X1 U16737 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13415) );
  NOR2_X1 U16738 ( .A1(n12853), .A2(n13415), .ZN(n15155) );
  NOR2_X1 U16739 ( .A1(n16110), .A2(n13414), .ZN(n13340) );
  AOI211_X1 U16740 ( .C1(n16099), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15155), .B(n13340), .ZN(n13341) );
  OAI211_X1 U16741 ( .C1(n16111), .C2(n20179), .A(n13342), .B(n13341), .ZN(
        P1_U2996) );
  INV_X1 U16742 ( .A(n20906), .ZN(n13343) );
  NOR2_X1 U16743 ( .A1(n20637), .A2(n13343), .ZN(n15956) );
  AOI21_X1 U16744 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n15956), .A(n16255), 
        .ZN(n13346) );
  AND2_X1 U16745 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20237), .ZN(n13344) );
  NAND2_X1 U16746 ( .A1(n14437), .A2(n13344), .ZN(n13345) );
  NAND2_X1 U16747 ( .A1(n13595), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13358) );
  INV_X1 U16748 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14743) );
  INV_X1 U16749 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14929) );
  INV_X1 U16750 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14340) );
  INV_X1 U16751 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U16752 ( .A1(n14382), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14404) );
  INV_X1 U16753 ( .A(n14404), .ZN(n13352) );
  NAND2_X1 U16754 ( .A1(n14436), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13354) );
  INV_X1 U16755 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13353) );
  XNOR2_X1 U16756 ( .A(n13354), .B(n13353), .ZN(n14442) );
  INV_X1 U16757 ( .A(n13377), .ZN(n13359) );
  NAND2_X1 U16758 ( .A1(n13355), .A2(n13359), .ZN(n13356) );
  NAND2_X1 U16759 ( .A1(n14774), .A2(n13356), .ZN(n20165) );
  INV_X1 U16760 ( .A(n14442), .ZN(n13357) );
  AND2_X1 U16761 ( .A1(n20902), .A2(n20703), .ZN(n15950) );
  INV_X1 U16762 ( .A(n15950), .ZN(n13360) );
  NAND3_X1 U16763 ( .A1(n13360), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n13359), 
        .ZN(n13361) );
  OAI22_X1 U16764 ( .A1(n20140), .A2(n13363), .B1(n20162), .B2(n13362), .ZN(
        n13376) );
  OR2_X1 U16765 ( .A1(n13364), .A2(n13377), .ZN(n13367) );
  OAI21_X1 U16766 ( .B1(n20254), .B2(n13365), .A(n15950), .ZN(n13368) );
  NAND2_X1 U16767 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13591) );
  NAND2_X1 U16768 ( .A1(n13593), .A2(n13591), .ZN(n13371) );
  NAND2_X1 U16769 ( .A1(n13595), .A2(n13371), .ZN(n13416) );
  AND2_X1 U16770 ( .A1(n20254), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13366) );
  NOR2_X1 U16771 ( .A1(n13367), .A2(n13366), .ZN(n13369) );
  AND2_X2 U16772 ( .A1(n13369), .A2(n13368), .ZN(n20110) );
  NAND2_X1 U16773 ( .A1(n20110), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13370) );
  OAI21_X1 U16774 ( .B1(n13371), .B2(n21013), .A(n13370), .ZN(n13372) );
  AOI21_X1 U16775 ( .B1(n13416), .B2(P1_REIP_REG_2__SCAN_IN), .A(n13372), .ZN(
        n13374) );
  NAND2_X1 U16776 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13373) );
  NAND2_X1 U16777 ( .A1(n13374), .A2(n13373), .ZN(n13375) );
  NOR2_X1 U16778 ( .A1(n13376), .A2(n13375), .ZN(n13380) );
  INV_X1 U16779 ( .A(n13189), .ZN(n20241) );
  NOR2_X1 U16780 ( .A1(n13378), .A2(n13377), .ZN(n20151) );
  NAND2_X1 U16781 ( .A1(n20241), .A2(n20151), .ZN(n13379) );
  OAI211_X1 U16782 ( .C1(n13381), .C2(n13570), .A(n13380), .B(n13379), .ZN(
        P1_U2838) );
  INV_X1 U16783 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13393) );
  INV_X1 U16784 ( .A(n13382), .ZN(n13386) );
  OAI21_X1 U16785 ( .B1(n13135), .B2(n13384), .A(n13383), .ZN(n13385) );
  NAND3_X1 U16786 ( .A1(n13386), .A2(n15346), .A3(n13385), .ZN(n13392) );
  NAND2_X1 U16787 ( .A1(n13388), .A2(n13387), .ZN(n13390) );
  INV_X1 U16788 ( .A(n13395), .ZN(n13389) );
  AND2_X1 U16789 ( .A1(n13390), .A2(n13389), .ZN(n19220) );
  NAND2_X1 U16790 ( .A1(n15356), .A2(n19220), .ZN(n13391) );
  OAI211_X1 U16791 ( .C1(n15356), .C2(n13393), .A(n13392), .B(n13391), .ZN(
        P2_U2875) );
  XNOR2_X1 U16792 ( .A(n13382), .B(n13394), .ZN(n13400) );
  OR2_X1 U16793 ( .A1(n13396), .A2(n13395), .ZN(n13397) );
  AND2_X1 U16794 ( .A1(n13397), .A2(n13659), .ZN(n19202) );
  NOR2_X1 U16795 ( .A1(n15356), .A2(n11194), .ZN(n13398) );
  AOI21_X1 U16796 ( .B1(n19202), .B2(n15356), .A(n13398), .ZN(n13399) );
  OAI21_X1 U16797 ( .B1(n13400), .B2(n15359), .A(n13399), .ZN(P2_U2874) );
  NAND2_X1 U16798 ( .A1(n13401), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13407) );
  INV_X1 U16799 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13402) );
  AOI21_X1 U16800 ( .B1(n13402), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13403) );
  AOI21_X1 U16801 ( .B1(n14250), .B2(P1_EAX_REG_4__SCAN_IN), .A(n13403), .ZN(
        n13406) );
  NOR2_X1 U16802 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n13404), .ZN(
        n13405) );
  NOR2_X1 U16803 ( .A1(n13446), .A2(n13405), .ZN(n20159) );
  AOI22_X1 U16804 ( .A1(n13407), .A2(n13406), .B1(n14437), .B2(n20159), .ZN(
        n13408) );
  NOR2_X1 U16805 ( .A1(n13430), .A2(n13452), .ZN(n13455) );
  AOI21_X1 U16806 ( .B1(n13452), .B2(n13430), .A(n13455), .ZN(n20166) );
  INV_X1 U16807 ( .A(n20166), .ZN(n13500) );
  INV_X1 U16808 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21221) );
  OAI222_X1 U16809 ( .A1(n13500), .A2(n14803), .B1(n20185), .B2(n21221), .C1(
        n20163), .C2(n20171), .ZN(P1_U2868) );
  AND2_X1 U16810 ( .A1(n13411), .A2(n13410), .ZN(n13412) );
  NOR2_X1 U16811 ( .A1(n13413), .A2(n13412), .ZN(n20180) );
  NOR2_X1 U16812 ( .A1(n20140), .A2(n13414), .ZN(n13421) );
  NOR2_X1 U16813 ( .A1(n14540), .A2(n13591), .ZN(n20150) );
  AOI22_X1 U16814 ( .A1(n20110), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n20150), .B2(
        n13415), .ZN(n13418) );
  NAND2_X1 U16815 ( .A1(n13416), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13417) );
  OAI211_X1 U16816 ( .C1(n20136), .C2(n13419), .A(n13418), .B(n13417), .ZN(
        n13420) );
  AOI211_X1 U16817 ( .C1(n20180), .C2(n20144), .A(n13421), .B(n13420), .ZN(
        n13423) );
  OAI211_X1 U16818 ( .C1(n20179), .C2(n13570), .A(n13423), .B(n13422), .ZN(
        P1_U2837) );
  INV_X1 U16819 ( .A(n20159), .ZN(n13426) );
  AOI21_X1 U16820 ( .B1(n16099), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13424), .ZN(n13425) );
  OAI21_X1 U16821 ( .B1(n13426), .B2(n16110), .A(n13425), .ZN(n13427) );
  AOI21_X1 U16822 ( .B1(n20166), .B2(n16105), .A(n13427), .ZN(n13428) );
  OAI21_X1 U16823 ( .B1(n20095), .B2(n13429), .A(n13428), .ZN(P1_U2995) );
  INV_X1 U16824 ( .A(n13430), .ZN(n13454) );
  AOI22_X1 U16825 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n9808), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13437) );
  AOI22_X1 U16826 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n14367), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13436) );
  AOI22_X1 U16827 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U16828 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13434) );
  NAND4_X1 U16829 ( .A1(n13437), .A2(n13436), .A3(n13435), .A4(n13434), .ZN(
        n13443) );
  AOI22_X1 U16830 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n14368), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13441) );
  AOI22_X1 U16831 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13440) );
  AOI22_X1 U16832 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13439) );
  AOI22_X1 U16833 ( .A1(n14331), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13438) );
  NAND4_X1 U16834 ( .A1(n13441), .A2(n13440), .A3(n13439), .A4(n13438), .ZN(
        n13442) );
  NAND2_X1 U16835 ( .A1(n13576), .A2(n13619), .ZN(n13445) );
  NAND2_X1 U16836 ( .A1(n13530), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13444) );
  NAND2_X1 U16837 ( .A1(n13610), .A2(n14128), .ZN(n13451) );
  INV_X1 U16838 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13448) );
  OAI21_X1 U16839 ( .B1(n13446), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n13533), .ZN(n20141) );
  AOI22_X1 U16840 ( .A1(n20141), .A2(n14437), .B1(n14439), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13447) );
  OAI21_X1 U16841 ( .B1(n9911), .B2(n13448), .A(n13447), .ZN(n13449) );
  INV_X1 U16842 ( .A(n13449), .ZN(n13450) );
  NAND2_X1 U16843 ( .A1(n13451), .A2(n13450), .ZN(n13456) );
  NAND3_X1 U16844 ( .A1(n13454), .A2(n13456), .A3(n13453), .ZN(n13540) );
  INV_X1 U16845 ( .A(n13455), .ZN(n13458) );
  INV_X1 U16846 ( .A(n13456), .ZN(n13457) );
  NAND2_X1 U16847 ( .A1(n13458), .A2(n13457), .ZN(n13459) );
  NAND2_X1 U16848 ( .A1(n13540), .A2(n13459), .ZN(n20134) );
  INV_X1 U16849 ( .A(n14586), .ZN(n14582) );
  NAND2_X1 U16850 ( .A1(n14614), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13460) );
  OAI211_X1 U16851 ( .C1(n14593), .C2(P1_EBX_REG_5__SCAN_IN), .A(n14591), .B(
        n13460), .ZN(n13461) );
  OAI21_X1 U16852 ( .B1(n14582), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13461), .ZN(
        n13463) );
  AOI21_X1 U16853 ( .B1(n13463), .B2(n13462), .A(n13734), .ZN(n20143) );
  AOI22_X1 U16854 ( .A1(n20143), .A2(n20181), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14801), .ZN(n13464) );
  OAI21_X1 U16855 ( .B1(n20134), .B2(n14803), .A(n13464), .ZN(P1_U2867) );
  INV_X1 U16856 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14471) );
  INV_X1 U16857 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15480) );
  INV_X1 U16858 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16405) );
  INV_X1 U16859 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16415) );
  AOI21_X1 U16860 ( .B1(n16499), .B2(n13466), .A(n9834), .ZN(n16487) );
  OAI22_X1 U16861 ( .A1(n11751), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16562), .ZN(n14495) );
  INV_X1 U16862 ( .A(n14495), .ZN(n19285) );
  AOI22_X1 U16863 ( .A1(n16562), .A2(n19422), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n11751), .ZN(n14492) );
  NOR2_X1 U16864 ( .A1(n19285), .A2(n14492), .ZN(n14493) );
  NAND2_X1 U16865 ( .A1(n14493), .A2(n15263), .ZN(n15244) );
  NOR2_X1 U16866 ( .A1(n15246), .A2(n15244), .ZN(n19276) );
  OAI21_X1 U16867 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13467), .A(
        n13466), .ZN(n19275) );
  NAND2_X1 U16868 ( .A1(n19276), .A2(n19275), .ZN(n13547) );
  NOR2_X1 U16869 ( .A1(n16487), .A2(n13547), .ZN(n15179) );
  NOR2_X1 U16870 ( .A1(n19277), .A2(n15179), .ZN(n13468) );
  OAI21_X1 U16871 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9834), .A(
        n15178), .ZN(n16474) );
  XNOR2_X1 U16872 ( .A(n13468), .B(n16474), .ZN(n13497) );
  NOR2_X1 U16873 ( .A1(n13470), .A2(n13469), .ZN(n13471) );
  OR2_X1 U16874 ( .A1(n13472), .A2(n13471), .ZN(n19319) );
  AND2_X1 U16875 ( .A1(n12350), .A2(n13473), .ZN(n13474) );
  XNOR2_X1 U16876 ( .A(n13476), .B(n13475), .ZN(n16485) );
  INV_X1 U16877 ( .A(n16485), .ZN(n14532) );
  NOR2_X1 U16878 ( .A1(n19104), .A2(n13477), .ZN(n13492) );
  AND2_X1 U16879 ( .A1(n19937), .A2(n12350), .ZN(n13478) );
  NAND2_X1 U16880 ( .A1(n13492), .A2(n13478), .ZN(n19295) );
  INV_X1 U16881 ( .A(n19474), .ZN(n13479) );
  NOR2_X1 U16882 ( .A1(n13480), .A2(n13479), .ZN(n16559) );
  OR2_X1 U16883 ( .A1(n19404), .A2(n19245), .ZN(n13481) );
  NOR2_X1 U16884 ( .A1(n16559), .A2(n13481), .ZN(n13482) );
  NAND2_X1 U16885 ( .A1(n19286), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n13488) );
  NAND2_X1 U16886 ( .A1(n19256), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19264) );
  INV_X2 U16887 ( .A(n19264), .ZN(n19298) );
  NAND2_X1 U16888 ( .A1(n16287), .A2(n16286), .ZN(n13486) );
  NAND2_X1 U16889 ( .A1(n19937), .A2(n12350), .ZN(n13490) );
  INV_X1 U16890 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13483) );
  NAND3_X1 U16891 ( .A1(n13484), .A2(n13490), .A3(n13483), .ZN(n13485) );
  AOI22_X1 U16892 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19298), .B1(
        P2_EBX_REG_6__SCAN_IN), .B2(n19293), .ZN(n13487) );
  NAND3_X1 U16893 ( .A1(n13488), .A2(n13487), .A3(n19254), .ZN(n13489) );
  AOI21_X1 U16894 ( .B1(n14532), .B2(n19243), .A(n13489), .ZN(n13495) );
  AND2_X1 U16895 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13490), .ZN(n13491) );
  NAND2_X1 U16896 ( .A1(n13492), .A2(n13491), .ZN(n19266) );
  OR2_X1 U16897 ( .A1(n19266), .A2(n13493), .ZN(n13494) );
  OAI211_X1 U16898 ( .C1(n19319), .C2(n19290), .A(n13495), .B(n13494), .ZN(
        n13496) );
  AOI21_X1 U16899 ( .B1(n13497), .B2(n19245), .A(n13496), .ZN(n13498) );
  INV_X1 U16900 ( .A(n13498), .ZN(P2_U2849) );
  OAI222_X1 U16901 ( .A1(n14881), .A2(n20134), .B1(n14879), .B2(n13448), .C1(
        n14878), .C2(n20281), .ZN(P1_U2899) );
  INV_X1 U16902 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13499) );
  OAI222_X1 U16903 ( .A1(n20179), .A2(n14881), .B1(n13499), .B2(n14879), .C1(
        n14878), .C2(n20269), .ZN(P1_U2901) );
  INV_X1 U16904 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20204) );
  OAI222_X1 U16905 ( .A1(n13500), .A2(n14881), .B1(n20204), .B2(n14879), .C1(
        n14878), .C2(n20274), .ZN(P1_U2900) );
  INV_X1 U16906 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21207) );
  NAND2_X1 U16907 ( .A1(n20136), .A2(n20140), .ZN(n13501) );
  NAND2_X1 U16908 ( .A1(n13501), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13504) );
  AOI22_X1 U16909 ( .A1(n13502), .A2(n20144), .B1(n20110), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13503) );
  OAI211_X1 U16910 ( .C1(n15998), .C2(n21207), .A(n13504), .B(n13503), .ZN(
        n13505) );
  AOI21_X1 U16911 ( .B1(n12646), .B2(n20151), .A(n13505), .ZN(n13506) );
  OAI21_X1 U16912 ( .B1(n13507), .B2(n13570), .A(n13506), .ZN(P1_U2840) );
  XNOR2_X1 U16913 ( .A(n13508), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13510) );
  XNOR2_X1 U16914 ( .A(n13510), .B(n13509), .ZN(n19418) );
  NAND2_X1 U16915 ( .A1(n13512), .A2(n13511), .ZN(n13513) );
  AND2_X1 U16916 ( .A1(n13514), .A2(n13513), .ZN(n19415) );
  INV_X1 U16917 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19964) );
  OAI22_X1 U16918 ( .A1(n19964), .A2(n19254), .B1(n16475), .B2(n19275), .ZN(
        n13516) );
  INV_X1 U16919 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19263) );
  NOR2_X1 U16920 ( .A1(n16498), .A2(n19263), .ZN(n13515) );
  NOR2_X1 U16921 ( .A1(n13516), .A2(n13515), .ZN(n13517) );
  OAI21_X1 U16922 ( .B1(n19412), .B2(n16486), .A(n13517), .ZN(n13518) );
  AOI21_X1 U16923 ( .B1(n19415), .B2(n16494), .A(n13518), .ZN(n13519) );
  OAI21_X1 U16924 ( .B1(n16478), .B2(n19418), .A(n13519), .ZN(P2_U3010) );
  AOI22_X1 U16925 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13523) );
  AOI22_X1 U16926 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13522) );
  AOI22_X1 U16927 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13521) );
  AOI22_X1 U16928 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13520) );
  NAND4_X1 U16929 ( .A1(n13523), .A2(n13522), .A3(n13521), .A4(n13520), .ZN(
        n13529) );
  AOI22_X1 U16930 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13527) );
  AOI22_X1 U16931 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13526) );
  AOI22_X1 U16932 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13525) );
  AOI22_X1 U16933 ( .A1(n14352), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13524) );
  NAND4_X1 U16934 ( .A1(n13527), .A2(n13526), .A3(n13525), .A4(n13524), .ZN(
        n13528) );
  NAND2_X1 U16935 ( .A1(n13576), .A2(n13785), .ZN(n13532) );
  NAND2_X1 U16936 ( .A1(n13530), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13531) );
  NAND2_X1 U16937 ( .A1(n13572), .A2(n13573), .ZN(n13618) );
  INV_X1 U16938 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13538) );
  AND2_X1 U16939 ( .A1(n13533), .A2(n13535), .ZN(n13534) );
  OR2_X1 U16940 ( .A1(n13534), .A2(n13581), .ZN(n13626) );
  INV_X1 U16941 ( .A(n14439), .ZN(n13914) );
  NOR2_X1 U16942 ( .A1(n13914), .A2(n13535), .ZN(n13536) );
  AOI21_X1 U16943 ( .B1(n13626), .B2(n14437), .A(n13536), .ZN(n13537) );
  OAI21_X1 U16944 ( .B1(n9911), .B2(n13538), .A(n13537), .ZN(n13539) );
  AOI21_X1 U16945 ( .B1(n13542), .B2(n13540), .A(n13541), .ZN(n13628) );
  INV_X1 U16946 ( .A(n13628), .ZN(n13600) );
  MUX2_X1 U16947 ( .A(n9804), .B(n10135), .S(P1_EBX_REG_6__SCAN_IN), .Z(n13543) );
  INV_X1 U16948 ( .A(n13543), .ZN(n13545) );
  NAND2_X1 U16949 ( .A1(n14593), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13544) );
  NAND2_X1 U16950 ( .A1(n13545), .A2(n13544), .ZN(n16248) );
  XNOR2_X1 U16951 ( .A(n16252), .B(n16248), .ZN(n13634) );
  AOI22_X1 U16952 ( .A1(n13634), .A2(n20181), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14801), .ZN(n13546) );
  OAI21_X1 U16953 ( .B1(n13600), .B2(n14803), .A(n13546), .ZN(P1_U2866) );
  NAND2_X1 U16954 ( .A1(n9797), .A2(n13547), .ZN(n13548) );
  XNOR2_X1 U16955 ( .A(n16487), .B(n13548), .ZN(n13561) );
  INV_X1 U16956 ( .A(n13549), .ZN(n13550) );
  NAND2_X1 U16957 ( .A1(n13551), .A2(n13550), .ZN(n13552) );
  NAND2_X1 U16958 ( .A1(n13553), .A2(n13552), .ZN(n19323) );
  INV_X1 U16959 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19966) );
  OAI22_X1 U16960 ( .A1(n19271), .A2(n11163), .B1(n13554), .B2(n19266), .ZN(
        n13555) );
  INV_X1 U16961 ( .A(n13555), .ZN(n13556) );
  OAI211_X1 U16962 ( .C1(n19966), .C2(n19256), .A(n13556), .B(n19254), .ZN(
        n13557) );
  AOI21_X1 U16963 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19298), .A(
        n13557), .ZN(n13559) );
  NAND2_X1 U16964 ( .A1(n16490), .A2(n19243), .ZN(n13558) );
  OAI211_X1 U16965 ( .C1(n19323), .C2(n19290), .A(n13559), .B(n13558), .ZN(
        n13560) );
  AOI21_X1 U16966 ( .B1(n13561), .B2(n19245), .A(n13560), .ZN(n13562) );
  INV_X1 U16967 ( .A(n13562), .ZN(P2_U2850) );
  OAI222_X1 U16968 ( .A1(n14881), .A2(n13600), .B1(n14879), .B2(n13538), .C1(
        n14878), .C2(n20287), .ZN(P1_U2898) );
  INV_X1 U16969 ( .A(n20702), .ZN(n20705) );
  INV_X1 U16970 ( .A(n20110), .ZN(n20156) );
  OAI22_X1 U16971 ( .A1(n20156), .A2(n21128), .B1(P1_REIP_REG_1__SCAN_IN), 
        .B2(n14540), .ZN(n13564) );
  NOR2_X1 U16972 ( .A1(n13595), .A2(n21013), .ZN(n13563) );
  AOI211_X1 U16973 ( .C1(n20144), .C2(n13565), .A(n13564), .B(n13563), .ZN(
        n13567) );
  NAND2_X1 U16974 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13566) );
  OAI211_X1 U16975 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20140), .A(
        n13567), .B(n13566), .ZN(n13568) );
  AOI21_X1 U16976 ( .B1(n20705), .B2(n20151), .A(n13568), .ZN(n13569) );
  OAI21_X1 U16977 ( .B1(n13571), .B2(n13570), .A(n13569), .ZN(P1_U2839) );
  NAND2_X1 U16978 ( .A1(n13575), .A2(n13574), .ZN(n13617) );
  INV_X1 U16979 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13578) );
  NAND2_X1 U16980 ( .A1(n13576), .A2(n13784), .ZN(n13577) );
  OAI21_X1 U16981 ( .B1(n13579), .B2(n13578), .A(n13577), .ZN(n13580) );
  NAND2_X1 U16982 ( .A1(n13773), .A2(n14128), .ZN(n13587) );
  INV_X1 U16983 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13590) );
  NOR2_X1 U16984 ( .A1(n13581), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13582) );
  OR2_X1 U16985 ( .A1(n13720), .A2(n13582), .ZN(n20125) );
  AOI22_X1 U16986 ( .A1(n20125), .A2(n14437), .B1(n14439), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13583) );
  INV_X1 U16987 ( .A(n13583), .ZN(n13584) );
  NAND2_X1 U16988 ( .A1(n13587), .A2(n13586), .ZN(n13589) );
  OAI21_X1 U16989 ( .B1(n13541), .B2(n13589), .A(n13724), .ZN(n16104) );
  OAI222_X1 U16990 ( .A1(n16104), .A2(n14881), .B1(n13590), .B2(n14879), .C1(
        n14878), .C2(n20297), .ZN(P1_U2897) );
  INV_X1 U16991 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21215) );
  INV_X1 U16992 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21162) );
  NOR3_X1 U16993 ( .A1(n20823), .A2(n13415), .A3(n13591), .ZN(n13592) );
  NAND2_X1 U16994 ( .A1(n13592), .A2(n13595), .ZN(n20132) );
  NOR3_X1 U16995 ( .A1(n21215), .A2(n21162), .A3(n20132), .ZN(n13728) );
  NOR2_X1 U16996 ( .A1(n15998), .A2(n13728), .ZN(n20127) );
  NAND2_X1 U16997 ( .A1(n13595), .A2(n13594), .ZN(n20154) );
  AOI21_X1 U16998 ( .B1(n20153), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20138), .ZN(n13597) );
  AOI22_X1 U16999 ( .A1(n13634), .A2(n20144), .B1(n20110), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n13596) );
  OAI211_X1 U17000 ( .C1(n13626), .C2(n20140), .A(n13597), .B(n13596), .ZN(
        n13598) );
  AOI221_X1 U17001 ( .B1(n20127), .B2(P1_REIP_REG_6__SCAN_IN), .C1(n13727), 
        .C2(n21215), .A(n13598), .ZN(n13599) );
  OAI21_X1 U17002 ( .B1(n13600), .B2(n14774), .A(n13599), .ZN(P1_U2834) );
  XNOR2_X1 U17003 ( .A(n9885), .B(n13601), .ZN(n13605) );
  OR2_X1 U17004 ( .A1(n13602), .A2(n13658), .ZN(n13603) );
  AND2_X1 U17005 ( .A1(n13749), .A2(n13603), .ZN(n16408) );
  INV_X1 U17006 ( .A(n16408), .ZN(n15729) );
  MUX2_X1 U17007 ( .A(n15729), .B(n10949), .S(n15323), .Z(n13604) );
  OAI21_X1 U17008 ( .B1(n13605), .B2(n15359), .A(n13604), .ZN(P2_U2872) );
  NAND2_X1 U17009 ( .A1(n13608), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13609) );
  NAND2_X1 U17010 ( .A1(n13610), .A2(n13781), .ZN(n13613) );
  XNOR2_X1 U17011 ( .A(n13621), .B(n13619), .ZN(n13611) );
  NAND2_X1 U17012 ( .A1(n13611), .A2(n13786), .ZN(n13612) );
  NAND2_X1 U17013 ( .A1(n13613), .A2(n13612), .ZN(n13615) );
  INV_X1 U17014 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13614) );
  XNOR2_X1 U17015 ( .A(n13615), .B(n13614), .ZN(n16109) );
  NAND2_X1 U17016 ( .A1(n13615), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13616) );
  INV_X1 U17017 ( .A(n13619), .ZN(n13620) );
  OR2_X1 U17018 ( .A1(n13621), .A2(n13620), .ZN(n13774) );
  XNOR2_X1 U17019 ( .A(n13774), .B(n13785), .ZN(n13622) );
  NAND2_X1 U17020 ( .A1(n13622), .A2(n13786), .ZN(n13623) );
  NAND2_X1 U17021 ( .A1(n13624), .A2(n13623), .ZN(n13772) );
  INV_X1 U17022 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13797) );
  XNOR2_X1 U17023 ( .A(n13772), .B(n13797), .ZN(n13770) );
  XNOR2_X1 U17024 ( .A(n13771), .B(n13770), .ZN(n13637) );
  NOR2_X1 U17025 ( .A1(n12853), .A2(n21215), .ZN(n13633) );
  AOI21_X1 U17026 ( .B1(n16099), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13633), .ZN(n13625) );
  OAI21_X1 U17027 ( .B1(n13626), .B2(n16110), .A(n13625), .ZN(n13627) );
  AOI21_X1 U17028 ( .B1(n13628), .B2(n16105), .A(n13627), .ZN(n13629) );
  OAI21_X1 U17029 ( .B1(n20095), .B2(n13637), .A(n13629), .ZN(P1_U2993) );
  OR2_X1 U17030 ( .A1(n13632), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16265) );
  OR2_X1 U17031 ( .A1(n13614), .A2(n13632), .ZN(n15025) );
  NOR2_X1 U17032 ( .A1(n13630), .A2(n15025), .ZN(n16226) );
  OAI21_X1 U17033 ( .B1(n16226), .B2(n16130), .A(n16225), .ZN(n13631) );
  AOI21_X1 U17034 ( .B1(n15038), .B2(n13632), .A(n13631), .ZN(n16271) );
  OAI21_X1 U17035 ( .B1(n16206), .B2(n16265), .A(n16271), .ZN(n13796) );
  INV_X1 U17036 ( .A(n15153), .ZN(n16266) );
  AOI22_X1 U17037 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13796), .B1(
        n16211), .B2(n13797), .ZN(n13636) );
  AOI21_X1 U17038 ( .B1(n13634), .B2(n16263), .A(n13633), .ZN(n13635) );
  OAI211_X1 U17039 ( .C1(n13637), .C2(n16215), .A(n13636), .B(n13635), .ZN(
        P1_U3025) );
  OAI21_X1 U17040 ( .B1(n13640), .B2(n13639), .A(n13638), .ZN(n16489) );
  OAI22_X1 U17041 ( .A1(n19323), .A2(n16551), .B1(n19966), .B2(n19254), .ZN(
        n13644) );
  OAI21_X1 U17042 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n13831), .ZN(n13641) );
  OAI22_X1 U17043 ( .A1(n19406), .A2(n13642), .B1(n19408), .B2(n13641), .ZN(
        n13643) );
  AOI211_X1 U17044 ( .C1(n16490), .C2(n14475), .A(n13644), .B(n13643), .ZN(
        n13653) );
  INV_X1 U17045 ( .A(n13645), .ZN(n13651) );
  INV_X1 U17046 ( .A(n13646), .ZN(n13649) );
  NAND2_X1 U17047 ( .A1(n13650), .A2(n13647), .ZN(n13648) );
  AOI22_X1 U17048 ( .A1(n13651), .A2(n13650), .B1(n13649), .B2(n13648), .ZN(
        n16492) );
  NAND2_X1 U17049 ( .A1(n16492), .A2(n19429), .ZN(n13652) );
  OAI211_X1 U17050 ( .C1(n16489), .C2(n19436), .A(n13653), .B(n13652), .ZN(
        P2_U3041) );
  INV_X1 U17051 ( .A(n13654), .ZN(n13657) );
  INV_X1 U17052 ( .A(n9885), .ZN(n13655) );
  OAI211_X1 U17053 ( .C1(n13657), .C2(n13656), .A(n13655), .B(n15346), .ZN(
        n13662) );
  AOI21_X1 U17054 ( .B1(n13660), .B2(n13659), .A(n13658), .ZN(n19193) );
  NAND2_X1 U17055 ( .A1(n15356), .A2(n19193), .ZN(n13661) );
  OAI211_X1 U17056 ( .C1(n15356), .C2(n13663), .A(n13662), .B(n13661), .ZN(
        P2_U2873) );
  NOR2_X1 U17057 ( .A1(n20042), .A2(n19496), .ZN(n13664) );
  NOR2_X1 U17058 ( .A1(n20042), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20036) );
  AOI21_X1 U17059 ( .B1(n19934), .B2(n13664), .A(n20036), .ZN(n13668) );
  NOR3_X2 U17060 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19501), .ZN(n19461) );
  INV_X1 U17061 ( .A(n19461), .ZN(n13665) );
  AND2_X1 U17062 ( .A1(n19889), .A2(n13665), .ZN(n13672) );
  INV_X1 U17063 ( .A(n13669), .ZN(n13666) );
  OAI21_X1 U17064 ( .B1(n13666), .B2(n19461), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13667) );
  OAI21_X1 U17065 ( .B1(n13668), .B2(n13672), .A(n13667), .ZN(n19467) );
  INV_X1 U17066 ( .A(n19467), .ZN(n13693) );
  INV_X1 U17067 ( .A(n13117), .ZN(n13708) );
  INV_X1 U17068 ( .A(n13668), .ZN(n13673) );
  AOI21_X1 U17069 ( .B1(n13669), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13670) );
  OAI21_X1 U17070 ( .B1(n13670), .B2(n19461), .A(n19737), .ZN(n13671) );
  INV_X1 U17071 ( .A(n19471), .ZN(n13690) );
  INV_X1 U17072 ( .A(n19894), .ZN(n19808) );
  AOI22_X1 U17073 ( .A1(n19805), .A2(n19496), .B1(n19885), .B2(n19461), .ZN(
        n13674) );
  OAI21_X1 U17074 ( .B1(n19808), .B2(n19934), .A(n13674), .ZN(n13675) );
  AOI21_X1 U17075 ( .B1(n13690), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n13675), .ZN(n13676) );
  OAI21_X1 U17076 ( .B1(n13693), .B2(n13708), .A(n13676), .ZN(P2_U3048) );
  INV_X1 U17077 ( .A(n13101), .ZN(n13680) );
  AOI22_X1 U17078 ( .A1(n19870), .A2(n19496), .B1(n19921), .B2(n19461), .ZN(
        n13677) );
  OAI21_X1 U17079 ( .B1(n19934), .B2(n19826), .A(n13677), .ZN(n13678) );
  AOI21_X1 U17080 ( .B1(n13690), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n13678), .ZN(n13679) );
  OAI21_X1 U17081 ( .B1(n13693), .B2(n13680), .A(n13679), .ZN(P2_U3054) );
  INV_X1 U17082 ( .A(n13681), .ZN(n13687) );
  AOI22_X1 U17083 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19466), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19465), .ZN(n19811) );
  AOI22_X1 U17084 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19466), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19465), .ZN(n19901) );
  AOI22_X1 U17085 ( .A1(n19853), .A2(n19496), .B1(n19461), .B2(n13683), .ZN(
        n13684) );
  OAI21_X1 U17086 ( .B1(n19811), .B2(n19934), .A(n13684), .ZN(n13685) );
  AOI21_X1 U17087 ( .B1(n13690), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n13685), .ZN(n13686) );
  OAI21_X1 U17088 ( .B1(n13693), .B2(n13687), .A(n13686), .ZN(P2_U3049) );
  INV_X1 U17089 ( .A(n13305), .ZN(n13692) );
  AOI22_X1 U17090 ( .A1(n19867), .A2(n19496), .B1(n19461), .B2(n13312), .ZN(
        n13688) );
  OAI21_X1 U17091 ( .B1(n19934), .B2(n19823), .A(n13688), .ZN(n13689) );
  AOI21_X1 U17092 ( .B1(n13690), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n13689), .ZN(n13691) );
  OAI21_X1 U17093 ( .B1(n13693), .B2(n13692), .A(n13691), .ZN(P2_U3053) );
  NOR2_X2 U17094 ( .A1(n19733), .A2(n20041), .ZN(n19930) );
  NOR3_X1 U17095 ( .A1(n19874), .A2(n19930), .A3(n20042), .ZN(n13694) );
  NOR2_X1 U17096 ( .A1(n13694), .A2(n20036), .ZN(n13698) );
  INV_X1 U17097 ( .A(n13695), .ZN(n19882) );
  NOR3_X2 U17098 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20048), .A3(
        n19882), .ZN(n19873) );
  NOR2_X1 U17099 ( .A1(n19873), .A2(n19846), .ZN(n13701) );
  INV_X1 U17100 ( .A(n13696), .ZN(n13699) );
  OAI21_X1 U17101 ( .B1(n13699), .B2(n19873), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13697) );
  OAI21_X1 U17102 ( .B1(n13698), .B2(n13701), .A(n13697), .ZN(n19876) );
  INV_X1 U17103 ( .A(n19876), .ZN(n13709) );
  INV_X1 U17104 ( .A(n13698), .ZN(n13702) );
  AOI211_X1 U17105 ( .C1(n13699), .C2(n13298), .A(n19873), .B(n20037), .ZN(
        n13700) );
  INV_X1 U17106 ( .A(n19880), .ZN(n13706) );
  INV_X1 U17107 ( .A(n19874), .ZN(n13704) );
  AOI22_X1 U17108 ( .A1(n19930), .A2(n19805), .B1(n19885), .B2(n19873), .ZN(
        n13703) );
  OAI21_X1 U17109 ( .B1(n13704), .B2(n19808), .A(n13703), .ZN(n13705) );
  AOI21_X1 U17110 ( .B1(n13706), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n13705), .ZN(n13707) );
  OAI21_X1 U17111 ( .B1(n13709), .B2(n13708), .A(n13707), .ZN(P2_U3160) );
  AOI22_X1 U17112 ( .A1(n14250), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n14439), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13723) );
  AOI22_X1 U17113 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13713) );
  AOI22_X1 U17114 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13712) );
  AOI22_X1 U17115 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13711) );
  AOI22_X1 U17116 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13710) );
  NAND4_X1 U17117 ( .A1(n13713), .A2(n13712), .A3(n13711), .A4(n13710), .ZN(
        n13719) );
  AOI22_X1 U17118 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14414), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13717) );
  AOI22_X1 U17119 ( .A1(n14352), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13716) );
  AOI22_X1 U17120 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U17121 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13714) );
  NAND4_X1 U17122 ( .A1(n13717), .A2(n13716), .A3(n13715), .A4(n13714), .ZN(
        n13718) );
  OR2_X1 U17123 ( .A1(n13719), .A2(n13718), .ZN(n13721) );
  XNOR2_X1 U17124 ( .A(n13720), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13792) );
  AOI22_X1 U17125 ( .A1(n14128), .A2(n13721), .B1(n14437), .B2(n13792), .ZN(
        n13722) );
  INV_X1 U17126 ( .A(n13822), .ZN(n13725) );
  AOI21_X1 U17127 ( .B1(n13726), .B2(n13724), .A(n13725), .ZN(n13794) );
  INV_X1 U17128 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n13944) );
  NOR2_X1 U17129 ( .A1(n13944), .A2(n20131), .ZN(n13730) );
  NAND3_X1 U17130 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_8__SCAN_IN), 
        .A3(n13728), .ZN(n13942) );
  NAND2_X1 U17131 ( .A1(n9798), .A2(n13942), .ZN(n20120) );
  INV_X1 U17132 ( .A(n20120), .ZN(n13729) );
  MUX2_X1 U17133 ( .A(n13730), .B(n13729), .S(P1_REIP_REG_8__SCAN_IN), .Z(
        n13743) );
  INV_X1 U17134 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21239) );
  INV_X1 U17135 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21034) );
  NAND2_X1 U17136 ( .A1(n14586), .A2(n21034), .ZN(n13733) );
  NAND2_X1 U17137 ( .A1(n14614), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13731) );
  OAI211_X1 U17138 ( .C1(n14593), .C2(P1_EBX_REG_7__SCAN_IN), .A(n14591), .B(
        n13731), .ZN(n13732) );
  MUX2_X1 U17139 ( .A(n9804), .B(n10135), .S(P1_EBX_REG_8__SCAN_IN), .Z(n13737) );
  AND2_X1 U17140 ( .A1(n14593), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13736) );
  NOR2_X1 U17141 ( .A1(n13737), .A2(n13736), .ZN(n13738) );
  AND2_X1 U17142 ( .A1(n16254), .A2(n13738), .ZN(n13739) );
  NOR2_X1 U17143 ( .A1(n16238), .A2(n13739), .ZN(n13802) );
  INV_X1 U17144 ( .A(n13802), .ZN(n13762) );
  OAI22_X1 U17145 ( .A1(n21239), .A2(n20156), .B1(n20162), .B2(n13762), .ZN(
        n13740) );
  AOI211_X1 U17146 ( .C1(n20153), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n13740), .B(n20138), .ZN(n13741) );
  OAI21_X1 U17147 ( .B1(n20140), .B2(n13792), .A(n13741), .ZN(n13742) );
  AOI211_X1 U17148 ( .C1(n13794), .C2(n20128), .A(n13743), .B(n13742), .ZN(
        n13744) );
  INV_X1 U17149 ( .A(n13744), .ZN(P1_U2832) );
  AOI21_X1 U17150 ( .B1(n13747), .B2(n13745), .A(n13746), .ZN(n13760) );
  NAND2_X1 U17151 ( .A1(n13760), .A2(n15346), .ZN(n13752) );
  NAND2_X1 U17152 ( .A1(n13749), .A2(n13748), .ZN(n13750) );
  NAND2_X1 U17153 ( .A1(n13766), .A2(n13750), .ZN(n15713) );
  INV_X1 U17154 ( .A(n15713), .ZN(n19182) );
  NAND2_X1 U17155 ( .A1(n19182), .A2(n15356), .ZN(n13751) );
  OAI211_X1 U17156 ( .C1(n15356), .C2(n10935), .A(n13752), .B(n13751), .ZN(
        P2_U2871) );
  OR2_X1 U17157 ( .A1(n13754), .A2(n13753), .ZN(n13755) );
  NAND2_X1 U17158 ( .A1(n13840), .A2(n13755), .ZN(n19186) );
  AOI22_X1 U17159 ( .A1(n19302), .A2(BUF2_REG_16__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n13758) );
  AOI22_X1 U17160 ( .A1(n16381), .A2(n13756), .B1(n19359), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n13757) );
  OAI211_X1 U17161 ( .C1(n19334), .C2(n19186), .A(n13758), .B(n13757), .ZN(
        n13759) );
  AOI21_X1 U17162 ( .B1(n13760), .B2(n19361), .A(n13759), .ZN(n13761) );
  INV_X1 U17163 ( .A(n13761), .ZN(P2_U2903) );
  INV_X1 U17164 ( .A(n13794), .ZN(n13763) );
  OAI222_X1 U17165 ( .A1(n13763), .A2(n14803), .B1(n20185), .B2(n21239), .C1(
        n13762), .C2(n20171), .ZN(P1_U2864) );
  OAI222_X1 U17166 ( .A1(n13763), .A2(n14881), .B1(n20199), .B2(n14879), .C1(
        n14878), .C2(n14832), .ZN(P1_U2896) );
  OAI21_X1 U17167 ( .B1(n13746), .B2(n13765), .A(n13764), .ZN(n13847) );
  NAND2_X1 U17168 ( .A1(n15352), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13769) );
  AOI21_X1 U17169 ( .B1(n13767), .B2(n13766), .A(n13851), .ZN(n19172) );
  NAND2_X1 U17170 ( .A1(n19172), .A2(n15356), .ZN(n13768) );
  OAI211_X1 U17171 ( .C1(n13847), .C2(n15359), .A(n13769), .B(n13768), .ZN(
        P2_U2870) );
  NAND2_X1 U17172 ( .A1(n13773), .A2(n13781), .ZN(n13778) );
  INV_X1 U17173 ( .A(n13774), .ZN(n13787) );
  NAND2_X1 U17174 ( .A1(n13787), .A2(n13785), .ZN(n13775) );
  XNOR2_X1 U17175 ( .A(n13775), .B(n13784), .ZN(n13776) );
  NAND2_X1 U17176 ( .A1(n13776), .A2(n13786), .ZN(n13777) );
  NAND2_X1 U17177 ( .A1(n13778), .A2(n13777), .ZN(n13779) );
  OR2_X1 U17178 ( .A1(n13779), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16101) );
  NAND2_X1 U17179 ( .A1(n16103), .A2(n16101), .ZN(n13780) );
  NAND2_X1 U17180 ( .A1(n13779), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16100) );
  AND2_X1 U17181 ( .A1(n13782), .A2(n13781), .ZN(n13783) );
  NAND4_X1 U17182 ( .A1(n13787), .A2(n13786), .A3(n13785), .A4(n13784), .ZN(
        n13788) );
  NAND2_X1 U17183 ( .A1(n16068), .A2(n13788), .ZN(n13904) );
  XOR2_X1 U17184 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n13904), .Z(
        n13789) );
  XNOR2_X1 U17185 ( .A(n13903), .B(n13789), .ZN(n13804) );
  INV_X1 U17186 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13790) );
  NOR2_X1 U17187 ( .A1(n12853), .A2(n13790), .ZN(n13801) );
  AOI21_X1 U17188 ( .B1(n16099), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n13801), .ZN(n13791) );
  OAI21_X1 U17189 ( .B1(n13792), .B2(n16110), .A(n13791), .ZN(n13793) );
  AOI21_X1 U17190 ( .B1(n13794), .B2(n16105), .A(n13793), .ZN(n13795) );
  OAI21_X1 U17191 ( .B1(n20095), .B2(n13804), .A(n13795), .ZN(P1_U2991) );
  INV_X1 U17192 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13798) );
  INV_X1 U17193 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16260) );
  NOR2_X1 U17194 ( .A1(n13798), .A2(n16260), .ZN(n16229) );
  INV_X1 U17195 ( .A(n16211), .ZN(n16181) );
  NOR2_X1 U17196 ( .A1(n13797), .A2(n16181), .ZN(n16256) );
  OAI21_X1 U17197 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16256), .ZN(n13799) );
  AOI21_X1 U17198 ( .B1(n13797), .B2(n16161), .A(n13796), .ZN(n16261) );
  OAI22_X1 U17199 ( .A1(n16229), .A2(n13799), .B1(n16261), .B2(n13798), .ZN(
        n13800) );
  AOI211_X1 U17200 ( .C1(n16263), .C2(n13802), .A(n13801), .B(n13800), .ZN(
        n13803) );
  OAI21_X1 U17201 ( .B1(n16215), .B2(n13804), .A(n13803), .ZN(P1_U3023) );
  XOR2_X1 U17202 ( .A(n20112), .B(n13805), .Z(n20115) );
  INV_X1 U17203 ( .A(n20115), .ZN(n13820) );
  AOI22_X1 U17204 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13809) );
  AOI22_X1 U17205 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13808) );
  AOI22_X1 U17206 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13807) );
  AOI22_X1 U17207 ( .A1(n14352), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13806) );
  NAND4_X1 U17208 ( .A1(n13809), .A2(n13808), .A3(n13807), .A4(n13806), .ZN(
        n13815) );
  AOI22_X1 U17209 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13813) );
  AOI22_X1 U17210 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13812) );
  AOI22_X1 U17211 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13811) );
  AOI22_X1 U17212 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13810) );
  NAND4_X1 U17213 ( .A1(n13813), .A2(n13812), .A3(n13811), .A4(n13810), .ZN(
        n13814) );
  OAI21_X1 U17214 ( .B1(n13815), .B2(n13814), .A(n14128), .ZN(n13818) );
  NAND2_X1 U17215 ( .A1(n14250), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13817) );
  NAND2_X1 U17216 ( .A1(n14439), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13816) );
  NAND3_X1 U17217 ( .A1(n13818), .A2(n13817), .A3(n13816), .ZN(n13819) );
  AOI21_X1 U17218 ( .B1(n13820), .B2(n14437), .A(n13819), .ZN(n13821) );
  AND2_X1 U17219 ( .A1(n13822), .A2(n13821), .ZN(n13823) );
  OR2_X1 U17220 ( .A1(n13823), .A2(n13879), .ZN(n20172) );
  INV_X1 U17221 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13824) );
  OAI222_X1 U17222 ( .A1(n20172), .A2(n14881), .B1(n13824), .B2(n14879), .C1(
        n14878), .C2(n14828), .ZN(P1_U2895) );
  OAI21_X1 U17223 ( .B1(n13826), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13825), .ZN(n16479) );
  OR2_X1 U17224 ( .A1(n13828), .A2(n13827), .ZN(n13829) );
  NAND2_X1 U17225 ( .A1(n13830), .A2(n13829), .ZN(n16481) );
  NOR2_X1 U17226 ( .A1(n16481), .A2(n19436), .ZN(n13837) );
  NOR2_X1 U17227 ( .A1(n13831), .A2(n19408), .ZN(n13833) );
  INV_X1 U17228 ( .A(n13832), .ZN(n16553) );
  MUX2_X1 U17229 ( .A(n13833), .B(n16553), .S(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n13836) );
  NOR2_X1 U17230 ( .A1(n19319), .A2(n16551), .ZN(n13835) );
  INV_X1 U17231 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19968) );
  OAI22_X1 U17232 ( .A1(n19411), .A2(n16485), .B1(n19968), .B2(n19254), .ZN(
        n13834) );
  NOR4_X1 U17233 ( .A1(n13837), .A2(n13836), .A3(n13835), .A4(n13834), .ZN(
        n13838) );
  OAI21_X1 U17234 ( .B1(n19419), .B2(n16479), .A(n13838), .ZN(P2_U3040) );
  AND2_X1 U17235 ( .A1(n13840), .A2(n13839), .ZN(n13841) );
  OR2_X1 U17236 ( .A1(n9897), .A2(n13841), .ZN(n19170) );
  AOI22_X1 U17237 ( .A1(n19302), .A2(BUF2_REG_17__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17238 ( .A1(n16381), .A2(n13842), .B1(n19359), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13843) );
  OAI211_X1 U17239 ( .C1(n19334), .C2(n19170), .A(n13844), .B(n13843), .ZN(
        n13845) );
  INV_X1 U17240 ( .A(n13845), .ZN(n13846) );
  OAI21_X1 U17241 ( .B1(n13847), .B2(n15425), .A(n13846), .ZN(P2_U2902) );
  AOI21_X1 U17242 ( .B1(n13848), .B2(n13764), .A(n9886), .ZN(n13862) );
  NAND2_X1 U17243 ( .A1(n13862), .A2(n15346), .ZN(n13854) );
  OR2_X1 U17244 ( .A1(n13851), .A2(n13850), .ZN(n13852) );
  NAND2_X1 U17245 ( .A1(n13849), .A2(n13852), .ZN(n15693) );
  INV_X1 U17246 ( .A(n15693), .ZN(n19157) );
  NAND2_X1 U17247 ( .A1(n19157), .A2(n15356), .ZN(n13853) );
  OAI211_X1 U17248 ( .C1(n15356), .C2(n11207), .A(n13854), .B(n13853), .ZN(
        P2_U2869) );
  OR2_X1 U17249 ( .A1(n9897), .A2(n13856), .ZN(n13857) );
  NAND2_X1 U17250 ( .A1(n13855), .A2(n13857), .ZN(n19161) );
  AOI22_X1 U17251 ( .A1(n19302), .A2(BUF2_REG_18__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n13860) );
  AOI22_X1 U17252 ( .A1(n16381), .A2(n13858), .B1(n19359), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n13859) );
  OAI211_X1 U17253 ( .C1(n19334), .C2(n19161), .A(n13860), .B(n13859), .ZN(
        n13861) );
  AOI21_X1 U17254 ( .B1(n13862), .B2(n19361), .A(n13861), .ZN(n13863) );
  INV_X1 U17255 ( .A(n13863), .ZN(P2_U2901) );
  AOI22_X1 U17256 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13867) );
  AOI22_X1 U17257 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13866) );
  AOI22_X1 U17258 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13865) );
  AOI22_X1 U17259 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13864) );
  NAND4_X1 U17260 ( .A1(n13867), .A2(n13866), .A3(n13865), .A4(n13864), .ZN(
        n13874) );
  AOI22_X1 U17261 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14368), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U17262 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13871) );
  AOI22_X1 U17263 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13870) );
  AOI22_X1 U17264 ( .A1(n14331), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13869) );
  NAND4_X1 U17265 ( .A1(n13872), .A2(n13871), .A3(n13870), .A4(n13869), .ZN(
        n13873) );
  NOR2_X1 U17266 ( .A1(n13874), .A2(n13873), .ZN(n13878) );
  XNOR2_X1 U17267 ( .A(n13875), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16033) );
  NAND2_X1 U17268 ( .A1(n16033), .A2(n14437), .ZN(n13877) );
  AOI22_X1 U17269 ( .A1(n14250), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n14439), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13876) );
  OAI211_X1 U17270 ( .C1(n13878), .C2(n10037), .A(n13877), .B(n13876), .ZN(
        n13917) );
  XOR2_X1 U17271 ( .A(n13917), .B(n13879), .Z(n16036) );
  INV_X1 U17272 ( .A(n16036), .ZN(n13901) );
  INV_X1 U17273 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13880) );
  NAND2_X1 U17274 ( .A1(n14591), .A2(n13880), .ZN(n13881) );
  OAI211_X1 U17275 ( .C1(n14593), .C2(P1_EBX_REG_10__SCAN_IN), .A(n14614), .B(
        n13881), .ZN(n13883) );
  INV_X1 U17276 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n21039) );
  NAND2_X1 U17277 ( .A1(n9804), .A2(n21039), .ZN(n13882) );
  INV_X1 U17278 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20175) );
  NAND2_X1 U17279 ( .A1(n14586), .A2(n20175), .ZN(n13886) );
  NAND2_X1 U17280 ( .A1(n14614), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13884) );
  OAI211_X1 U17281 ( .C1(n14593), .C2(P1_EBX_REG_9__SCAN_IN), .A(n14591), .B(
        n13884), .ZN(n13885) );
  AND2_X1 U17282 ( .A1(n13886), .A2(n13885), .ZN(n16237) );
  INV_X1 U17283 ( .A(n13939), .ZN(n13887) );
  AOI21_X1 U17284 ( .B1(n13888), .B2(n16240), .A(n13887), .ZN(n16032) );
  AOI22_X1 U17285 ( .A1(n16032), .A2(n20181), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14801), .ZN(n13889) );
  OAI21_X1 U17286 ( .B1(n13901), .B2(n14803), .A(n13889), .ZN(P1_U2862) );
  OAI21_X1 U17287 ( .B1(n9886), .B2(n13892), .A(n13891), .ZN(n15360) );
  NAND2_X1 U17288 ( .A1(n13855), .A2(n13893), .ZN(n13894) );
  NAND2_X1 U17289 ( .A1(n15428), .A2(n13894), .ZN(n19146) );
  AOI22_X1 U17290 ( .A1(n19302), .A2(BUF2_REG_19__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U17291 ( .A1(n16381), .A2(n13895), .B1(n19359), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n13896) );
  OAI211_X1 U17292 ( .C1(n19334), .C2(n19146), .A(n13897), .B(n13896), .ZN(
        n13898) );
  INV_X1 U17293 ( .A(n13898), .ZN(n13899) );
  OAI21_X1 U17294 ( .B1(n15360), .B2(n15425), .A(n13899), .ZN(P2_U2900) );
  INV_X1 U17295 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13900) );
  OAI222_X1 U17296 ( .A1(n14878), .A2(n14823), .B1(n14881), .B2(n13901), .C1(
        n13900), .C2(n14879), .ZN(P1_U2894) );
  NAND2_X1 U17297 ( .A1(n13904), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13905) );
  INV_X1 U17298 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14052) );
  MUX2_X1 U17299 ( .A(n14052), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .S(
        n16090), .Z(n13907) );
  XNOR2_X1 U17300 ( .A(n14051), .B(n13907), .ZN(n16235) );
  OAI22_X1 U17301 ( .A1(n16116), .A2(n20112), .B1(n12853), .B2(n20121), .ZN(
        n13909) );
  NOR2_X1 U17302 ( .A1(n20172), .A2(n16111), .ZN(n13908) );
  AOI211_X1 U17303 ( .C1(n16084), .C2(n20115), .A(n13909), .B(n13908), .ZN(
        n13910) );
  OAI21_X1 U17304 ( .B1(n20095), .B2(n16235), .A(n13910), .ZN(P1_U2990) );
  INV_X1 U17305 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13915) );
  OAI21_X1 U17306 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13912), .A(
        n13911), .ZN(n16098) );
  NAND2_X1 U17307 ( .A1(n16098), .A2(n14437), .ZN(n13913) );
  OAI21_X1 U17308 ( .B1(n13915), .B2(n13914), .A(n13913), .ZN(n13916) );
  AOI21_X1 U17309 ( .B1(n14250), .B2(P1_EAX_REG_11__SCAN_IN), .A(n13916), .ZN(
        n13920) );
  NAND2_X1 U17310 ( .A1(n13919), .A2(n13918), .ZN(n13922) );
  AOI22_X1 U17311 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13926) );
  AOI22_X1 U17312 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13925) );
  AOI22_X1 U17313 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13924) );
  AOI22_X1 U17314 ( .A1(n12252), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14368), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13923) );
  NAND4_X1 U17315 ( .A1(n13926), .A2(n13925), .A3(n13924), .A4(n13923), .ZN(
        n13932) );
  AOI22_X1 U17316 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13930) );
  AOI22_X1 U17317 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13929) );
  AOI22_X1 U17318 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13928) );
  INV_X1 U17319 ( .A(n13868), .ZN(n14295) );
  AOI22_X1 U17320 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13927) );
  NAND4_X1 U17321 ( .A1(n13930), .A2(n13929), .A3(n13928), .A4(n13927), .ZN(
        n13931) );
  OR2_X1 U17322 ( .A1(n13932), .A2(n13931), .ZN(n13933) );
  AND2_X1 U17323 ( .A1(n14128), .A2(n13933), .ZN(n13934) );
  NAND2_X1 U17324 ( .A1(n13935), .A2(n13934), .ZN(n14073) );
  OAI21_X1 U17325 ( .B1(n13935), .B2(n13934), .A(n14073), .ZN(n16094) );
  MUX2_X1 U17326 ( .A(n14586), .B(n9804), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13936) );
  INV_X1 U17327 ( .A(n13936), .ZN(n13938) );
  INV_X1 U17328 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16222) );
  NAND2_X1 U17329 ( .A1(n14567), .A2(n16222), .ZN(n13937) );
  NAND2_X1 U17330 ( .A1(n13938), .A2(n13937), .ZN(n13940) );
  AOI21_X1 U17331 ( .B1(n13940), .B2(n13939), .A(n14512), .ZN(n16217) );
  AOI22_X1 U17332 ( .A1(n16217), .A2(n20181), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14801), .ZN(n13941) );
  OAI21_X1 U17333 ( .B1(n16094), .B2(n14803), .A(n13941), .ZN(P1_U2861) );
  INV_X1 U17334 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21048) );
  NOR2_X1 U17335 ( .A1(n21048), .A2(n13942), .ZN(n13943) );
  AOI21_X1 U17336 ( .B1(n13943), .B2(P1_REIP_REG_9__SCAN_IN), .A(n15998), .ZN(
        n16035) );
  NAND2_X1 U17337 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20116), .ZN(n16039) );
  INV_X1 U17338 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21040) );
  AOI21_X1 U17339 ( .B1(n20153), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20138), .ZN(n13946) );
  AOI22_X1 U17340 ( .A1(n16217), .A2(n20144), .B1(n20110), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n13945) );
  OAI211_X1 U17341 ( .C1(n16098), .C2(n20140), .A(n13946), .B(n13945), .ZN(
        n13947) );
  AOI221_X1 U17342 ( .B1(n16035), .B2(P1_REIP_REG_11__SCAN_IN), .C1(n14516), 
        .C2(n21040), .A(n13947), .ZN(n13948) );
  OAI21_X1 U17343 ( .B1(n16094), .B2(n14774), .A(n13948), .ZN(P1_U2829) );
  INV_X1 U17344 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13949) );
  OAI222_X1 U17345 ( .A1(n16094), .A2(n14881), .B1(n13949), .B2(n14879), .C1(
        n14878), .C2(n14818), .ZN(P1_U2893) );
  INV_X1 U17346 ( .A(n19060), .ZN(n19095) );
  AOI21_X1 U17347 ( .B1(n18887), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15871) );
  INV_X1 U17348 ( .A(n15871), .ZN(n13950) );
  NAND2_X1 U17349 ( .A1(n18889), .A2(n13950), .ZN(n18876) );
  NOR2_X1 U17350 ( .A1(n19095), .A2(n18876), .ZN(n13961) );
  NAND2_X1 U17351 ( .A1(n18871), .A2(n19085), .ZN(n13959) );
  NAND2_X1 U17352 ( .A1(n19084), .A2(n9810), .ZN(n18923) );
  NAND2_X1 U17353 ( .A1(n13951), .A2(n18923), .ZN(n13952) );
  OAI211_X1 U17354 ( .C1(n13957), .C2(n13956), .A(n13955), .B(n13954), .ZN(
        n15887) );
  AOI211_X1 U17355 ( .C1(n13965), .C2(n18868), .A(n15989), .B(n15887), .ZN(
        n13958) );
  OAI21_X1 U17356 ( .B1(n13959), .B2(n17645), .A(n13958), .ZN(n18897) );
  INV_X1 U17357 ( .A(n18897), .ZN(n18908) );
  NAND2_X1 U17358 ( .A1(n13960), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18439) );
  INV_X1 U17359 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18432) );
  NAND3_X1 U17360 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19032)
         );
  OR2_X1 U17361 ( .A1(n18432), .A2(n19032), .ZN(n15872) );
  MUX2_X1 U17362 ( .A(n13961), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19065), .Z(P3_U3284) );
  AND2_X1 U17363 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17184) );
  NOR4_X1 U17364 ( .A1(n13962), .A2(n18478), .A3(n18452), .A4(n18467), .ZN(
        n13963) );
  NOR2_X1 U17365 ( .A1(n18478), .A2(n17488), .ZN(n17482) );
  INV_X1 U17366 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17291) );
  INV_X1 U17367 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17288) );
  INV_X1 U17368 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17111) );
  NAND2_X1 U17369 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17479) );
  NOR2_X1 U17370 ( .A1(n17111), .A2(n17479), .ZN(n17483) );
  NAND2_X1 U17371 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17483), .ZN(n17472) );
  AND3_X1 U17372 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n17456) );
  NAND4_X1 U17373 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .A3(P3_EBX_REG_8__SCAN_IN), .A4(n17456), .ZN(n15869) );
  NAND4_X1 U17374 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .A4(P3_EBX_REG_11__SCAN_IN), .ZN(n13966)
         );
  NOR3_X1 U17375 ( .A1(n16947), .A2(n15869), .A3(n13966), .ZN(n17289) );
  INV_X1 U17376 ( .A(n17289), .ZN(n13967) );
  NAND2_X1 U17377 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .ZN(n17290) );
  AND2_X1 U17378 ( .A1(n10430), .A2(n17272), .ZN(n17274) );
  NAND3_X1 U17379 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n17274), .ZN(n17206) );
  NAND3_X1 U17380 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .ZN(n17146) );
  NAND2_X1 U17381 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17211), .ZN(n17196) );
  NAND2_X1 U17382 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17200), .ZN(n17190) );
  NAND2_X1 U17383 ( .A1(n17468), .A2(n17190), .ZN(n17194) );
  OAI21_X1 U17384 ( .B1(n17184), .B2(n17491), .A(n17194), .ZN(n17185) );
  AOI22_X1 U17385 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13968) );
  OAI21_X1 U17386 ( .B1(n10412), .B2(n17233), .A(n13968), .ZN(n13977) );
  AOI22_X1 U17387 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13975) );
  OAI22_X1 U17388 ( .A1(n10416), .A2(n17229), .B1(n17453), .B2(n17469), .ZN(
        n13973) );
  AOI22_X1 U17389 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13971) );
  AOI22_X1 U17390 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13970) );
  AOI22_X1 U17391 ( .A1(n11665), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13969) );
  NAND3_X1 U17392 ( .A1(n13971), .A2(n13970), .A3(n13969), .ZN(n13972) );
  AOI211_X1 U17393 ( .C1(n17438), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n13973), .B(n13972), .ZN(n13974) );
  OAI211_X1 U17394 ( .C1(n17426), .C2(n17227), .A(n13975), .B(n13974), .ZN(
        n13976) );
  AOI211_X1 U17395 ( .C1(n11667), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n13977), .B(n13976), .ZN(n14046) );
  AOI22_X1 U17396 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13978) );
  OAI21_X1 U17397 ( .B1(n11496), .B2(n17260), .A(n13978), .ZN(n13988) );
  INV_X1 U17398 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17259) );
  AOI22_X1 U17399 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13986) );
  INV_X1 U17400 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13980) );
  AOI22_X1 U17401 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13979) );
  OAI21_X1 U17402 ( .B1(n17441), .B2(n13980), .A(n13979), .ZN(n13984) );
  INV_X1 U17403 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17379) );
  AOI22_X1 U17404 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13982) );
  AOI22_X1 U17405 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13981) );
  OAI211_X1 U17406 ( .C1(n17447), .C2(n17379), .A(n13982), .B(n13981), .ZN(
        n13983) );
  AOI211_X1 U17407 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n13984), .B(n13983), .ZN(n13985) );
  OAI211_X1 U17408 ( .C1(n10412), .C2(n17259), .A(n13986), .B(n13985), .ZN(
        n13987) );
  AOI211_X1 U17409 ( .C1(n17417), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n13988), .B(n13987), .ZN(n17192) );
  AOI22_X1 U17410 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17396), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17437), .ZN(n13989) );
  OAI21_X1 U17411 ( .B1(n9926), .B2(n17414), .A(n13989), .ZN(n13999) );
  AOI22_X1 U17412 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17410), .ZN(n13997) );
  OAI22_X1 U17413 ( .A1(n13990), .A2(n17426), .B1(n9847), .B2(n17412), .ZN(
        n13995) );
  AOI22_X1 U17414 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17442), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13993) );
  AOI22_X1 U17415 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11637), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13992) );
  AOI22_X1 U17416 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n9803), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n11665), .ZN(n13991) );
  NAND3_X1 U17417 ( .A1(n13993), .A2(n13992), .A3(n13991), .ZN(n13994) );
  AOI211_X1 U17418 ( .C1(n17438), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n13995), .B(n13994), .ZN(n13996) );
  OAI211_X1 U17419 ( .C1(n17484), .C2(n17453), .A(n13997), .B(n13996), .ZN(
        n13998) );
  AOI211_X1 U17420 ( .C1(n11667), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n13999), .B(n13998), .ZN(n17202) );
  AOI22_X1 U17421 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17442), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14010) );
  AOI22_X1 U17422 ( .A1(n14033), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14000) );
  OAI21_X1 U17423 ( .B1(n17453), .B2(n14001), .A(n14000), .ZN(n14008) );
  AOI22_X1 U17424 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U17425 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14003) );
  AOI22_X1 U17426 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14002) );
  OAI211_X1 U17427 ( .C1(n17441), .C2(n17320), .A(n14003), .B(n14002), .ZN(
        n14004) );
  AOI21_X1 U17428 ( .B1(n9803), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(n14004), .ZN(n14005) );
  OAI211_X1 U17429 ( .C1(n17426), .C2(n17435), .A(n14006), .B(n14005), .ZN(
        n14007) );
  AOI211_X1 U17430 ( .C1(n17396), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n14008), .B(n14007), .ZN(n14009) );
  OAI211_X1 U17431 ( .C1(n17415), .C2(n17446), .A(n14010), .B(n14009), .ZN(
        n17208) );
  AOI22_X1 U17432 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14020) );
  AOI22_X1 U17433 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14012) );
  AOI22_X1 U17434 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14011) );
  OAI211_X1 U17435 ( .C1(n17426), .C2(n17325), .A(n14012), .B(n14011), .ZN(
        n14018) );
  AOI22_X1 U17436 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14016) );
  AOI22_X1 U17437 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14015) );
  AOI22_X1 U17438 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14014) );
  NAND2_X1 U17439 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n14013) );
  NAND4_X1 U17440 ( .A1(n14016), .A2(n14015), .A3(n14014), .A4(n14013), .ZN(
        n14017) );
  AOI211_X1 U17441 ( .C1(n11665), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n14018), .B(n14017), .ZN(n14019) );
  OAI211_X1 U17442 ( .C1(n17415), .C2(n17459), .A(n14020), .B(n14019), .ZN(
        n17209) );
  NAND2_X1 U17443 ( .A1(n17208), .A2(n17209), .ZN(n17207) );
  NOR2_X1 U17444 ( .A1(n17202), .A2(n17207), .ZN(n17201) );
  AOI22_X1 U17445 ( .A1(n17396), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14032) );
  AOI22_X1 U17446 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14031) );
  OAI22_X1 U17447 ( .A1(n17441), .A2(n14021), .B1(n17453), .B2(n17278), .ZN(
        n14029) );
  AOI22_X1 U17448 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14027) );
  AOI22_X1 U17449 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14023) );
  AOI22_X1 U17450 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14022) );
  OAI211_X1 U17451 ( .C1(n17426), .C2(n14024), .A(n14023), .B(n14022), .ZN(
        n14025) );
  AOI21_X1 U17452 ( .B1(n9803), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(n14025), .ZN(n14026) );
  OAI211_X1 U17453 ( .C1(n17416), .C2(n17281), .A(n14027), .B(n14026), .ZN(
        n14028) );
  AOI211_X1 U17454 ( .C1(n17438), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n14029), .B(n14028), .ZN(n14030) );
  NAND3_X1 U17455 ( .A1(n14032), .A2(n14031), .A3(n14030), .ZN(n17198) );
  NAND2_X1 U17456 ( .A1(n17201), .A2(n17198), .ZN(n17197) );
  NOR2_X1 U17457 ( .A1(n17192), .A2(n17197), .ZN(n17191) );
  AOI22_X1 U17458 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14044) );
  AOI22_X1 U17459 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14035) );
  AOI22_X1 U17460 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14034) );
  OAI211_X1 U17461 ( .C1(n17426), .C2(n17361), .A(n14035), .B(n14034), .ZN(
        n14042) );
  AOI22_X1 U17462 ( .A1(n17396), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14040) );
  AOI22_X1 U17463 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14039) );
  AOI22_X1 U17464 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17442), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14038) );
  NAND2_X1 U17465 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n14037) );
  NAND4_X1 U17466 ( .A1(n14040), .A2(n14039), .A3(n14038), .A4(n14037), .ZN(
        n14041) );
  AOI211_X1 U17467 ( .C1(n9803), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n14042), .B(n14041), .ZN(n14043) );
  OAI211_X1 U17468 ( .C1(n17441), .C2(n14045), .A(n14044), .B(n14043), .ZN(
        n17188) );
  NAND2_X1 U17469 ( .A1(n17191), .A2(n17188), .ZN(n17187) );
  NOR2_X1 U17470 ( .A1(n14046), .A2(n17187), .ZN(n17182) );
  AOI21_X1 U17471 ( .B1(n14046), .B2(n17187), .A(n17182), .ZN(n17506) );
  AOI22_X1 U17472 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17185), .B1(n17506), 
        .B2(n17489), .ZN(n14050) );
  INV_X1 U17473 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14048) );
  INV_X1 U17474 ( .A(n17190), .ZN(n14047) );
  NAND3_X1 U17475 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14048), .A3(n14047), 
        .ZN(n14049) );
  NAND2_X1 U17476 ( .A1(n14050), .A2(n14049), .ZN(P3_U2675) );
  NAND2_X1 U17477 ( .A1(n16090), .A2(n14052), .ZN(n14053) );
  NOR2_X1 U17478 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14054) );
  INV_X1 U17479 ( .A(n14055), .ZN(n14066) );
  INV_X1 U17480 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16141) );
  INV_X1 U17481 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16183) );
  OR2_X1 U17482 ( .A1(n16090), .A2(n16183), .ZN(n14056) );
  INV_X1 U17483 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14060) );
  NAND2_X1 U17484 ( .A1(n16090), .A2(n16141), .ZN(n14058) );
  NAND2_X1 U17485 ( .A1(n16066), .A2(n14058), .ZN(n15012) );
  INV_X1 U17486 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16210) );
  AND2_X1 U17487 ( .A1(n16090), .A2(n16210), .ZN(n15011) );
  NOR2_X1 U17488 ( .A1(n15012), .A2(n15011), .ZN(n16064) );
  NAND2_X1 U17489 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14059) );
  NAND2_X1 U17490 ( .A1(n16068), .A2(n14059), .ZN(n16077) );
  OAI211_X1 U17491 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n10354), .A(
        n16064), .B(n16077), .ZN(n16042) );
  NOR2_X1 U17492 ( .A1(n16068), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15003) );
  AOI21_X1 U17493 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16068), .A(
        n15003), .ZN(n16049) );
  AOI211_X1 U17494 ( .C1(n14061), .C2(n16042), .A(n16048), .B(n16049), .ZN(
        n15000) );
  AND2_X1 U17495 ( .A1(n15000), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14064) );
  NOR2_X1 U17496 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14062) );
  AOI21_X1 U17497 ( .B1(n16046), .B2(n14064), .A(n14063), .ZN(n14065) );
  XOR2_X1 U17498 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n16090), .Z(
        n14994) );
  AND2_X1 U17499 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15132) );
  INV_X1 U17500 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15133) );
  NOR2_X1 U17501 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14963) );
  INV_X1 U17502 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14067) );
  NAND3_X1 U17503 ( .A1(n14963), .A2(n14067), .A3(n15134), .ZN(n14068) );
  AND2_X1 U17504 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15099) );
  NAND2_X1 U17505 ( .A1(n15099), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15041) );
  INV_X1 U17506 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15029) );
  NOR2_X1 U17507 ( .A1(n14070), .A2(n10354), .ZN(n14932) );
  AOI211_X2 U17508 ( .C1(n14948), .C2(n15041), .A(n15029), .B(n14932), .ZN(
        n14912) );
  NOR2_X1 U17509 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14899) );
  AND2_X1 U17510 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15035) );
  NAND2_X1 U17511 ( .A1(n15035), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15030) );
  INV_X1 U17512 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15062) );
  NAND2_X1 U17513 ( .A1(n10354), .A2(n15062), .ZN(n14889) );
  NOR2_X1 U17514 ( .A1(n14889), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14071) );
  NAND2_X1 U17515 ( .A1(n14073), .A2(n14072), .ZN(n14505) );
  XNOR2_X1 U17516 ( .A(n14074), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16026) );
  INV_X1 U17517 ( .A(n16026), .ZN(n15016) );
  AOI22_X1 U17518 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U17519 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14077) );
  AOI22_X1 U17520 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14076) );
  AOI22_X1 U17521 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14075) );
  NAND4_X1 U17522 ( .A1(n14078), .A2(n14077), .A3(n14076), .A4(n14075), .ZN(
        n14084) );
  AOI22_X1 U17523 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n12660), .B1(
        n9808), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17524 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n14198), .B1(
        n14367), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U17525 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14080) );
  AOI22_X1 U17526 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n14368), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14079) );
  NAND4_X1 U17527 ( .A1(n14082), .A2(n14081), .A3(n14080), .A4(n14079), .ZN(
        n14083) );
  OAI21_X1 U17528 ( .B1(n14084), .B2(n14083), .A(n14128), .ZN(n14087) );
  NAND2_X1 U17529 ( .A1(n14250), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n14086) );
  NAND2_X1 U17530 ( .A1(n14439), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14085) );
  NAND3_X1 U17531 ( .A1(n14087), .A2(n14086), .A3(n14085), .ZN(n14088) );
  AOI21_X1 U17532 ( .B1(n15016), .B2(n14437), .A(n14088), .ZN(n14794) );
  XOR2_X1 U17533 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n14089), .Z(
        n16083) );
  AOI22_X1 U17534 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14093) );
  AOI22_X1 U17535 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U17536 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14091) );
  AOI22_X1 U17537 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14090) );
  NAND4_X1 U17538 ( .A1(n14093), .A2(n14092), .A3(n14091), .A4(n14090), .ZN(
        n14099) );
  AOI22_X1 U17539 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14097) );
  AOI22_X1 U17540 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14096) );
  AOI22_X1 U17541 ( .A1(n14352), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14095) );
  AOI22_X1 U17542 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14241), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14094) );
  NAND4_X1 U17543 ( .A1(n14097), .A2(n14096), .A3(n14095), .A4(n14094), .ZN(
        n14098) );
  OR2_X1 U17544 ( .A1(n14099), .A2(n14098), .ZN(n14100) );
  AOI22_X1 U17545 ( .A1(n14128), .A2(n14100), .B1(n14439), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14102) );
  NAND2_X1 U17546 ( .A1(n14250), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n14101) );
  OAI211_X1 U17547 ( .C1(n16083), .C2(n14363), .A(n14102), .B(n14101), .ZN(
        n14506) );
  INV_X1 U17548 ( .A(n14506), .ZN(n14103) );
  NOR2_X1 U17549 ( .A1(n14794), .A2(n14103), .ZN(n14104) );
  XOR2_X1 U17550 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n14105), .Z(
        n16071) );
  AOI22_X1 U17551 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14109) );
  AOI22_X1 U17552 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14108) );
  AOI22_X1 U17553 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14107) );
  AOI22_X1 U17554 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14106) );
  NAND4_X1 U17555 ( .A1(n14109), .A2(n14108), .A3(n14107), .A4(n14106), .ZN(
        n14115) );
  AOI22_X1 U17556 ( .A1(n12255), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14113) );
  AOI22_X1 U17557 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14112) );
  AOI22_X1 U17558 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14111) );
  AOI22_X1 U17559 ( .A1(n14331), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14110) );
  NAND4_X1 U17560 ( .A1(n14113), .A2(n14112), .A3(n14111), .A4(n14110), .ZN(
        n14114) );
  OR2_X1 U17561 ( .A1(n14115), .A2(n14114), .ZN(n14116) );
  AOI22_X1 U17562 ( .A1(n14128), .A2(n14116), .B1(n14439), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14118) );
  NAND2_X1 U17563 ( .A1(n14250), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n14117) );
  OAI211_X1 U17564 ( .C1(n16071), .C2(n14363), .A(n14118), .B(n14117), .ZN(
        n14793) );
  NAND2_X1 U17565 ( .A1(n14790), .A2(n14793), .ZN(n14791) );
  XNOR2_X1 U17566 ( .A(n14119), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16059) );
  INV_X1 U17567 ( .A(n16059), .ZN(n14135) );
  AOI22_X1 U17568 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14123) );
  AOI22_X1 U17569 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U17570 ( .A1(n14352), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U17571 ( .A1(n14331), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14120) );
  NAND4_X1 U17572 ( .A1(n14123), .A2(n14122), .A3(n14121), .A4(n14120), .ZN(
        n14130) );
  AOI22_X1 U17573 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14127) );
  AOI22_X1 U17574 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14126) );
  AOI22_X1 U17575 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14125) );
  AOI22_X1 U17576 ( .A1(n12252), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14368), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14124) );
  NAND4_X1 U17577 ( .A1(n14127), .A2(n14126), .A3(n14125), .A4(n14124), .ZN(
        n14129) );
  OAI21_X1 U17578 ( .B1(n14130), .B2(n14129), .A(n14128), .ZN(n14133) );
  NAND2_X1 U17579 ( .A1(n14250), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n14132) );
  NAND2_X1 U17580 ( .A1(n14439), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14131) );
  NAND3_X1 U17581 ( .A1(n14133), .A2(n14132), .A3(n14131), .ZN(n14134) );
  AOI21_X1 U17582 ( .B1(n14135), .B2(n14437), .A(n14134), .ZN(n14869) );
  AOI22_X1 U17583 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14139) );
  AOI22_X1 U17584 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14138) );
  AOI22_X1 U17585 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14137) );
  AOI22_X1 U17586 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14136) );
  NAND4_X1 U17587 ( .A1(n14139), .A2(n14138), .A3(n14137), .A4(n14136), .ZN(
        n14145) );
  AOI22_X1 U17588 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14422), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14143) );
  AOI22_X1 U17589 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14142) );
  AOI22_X1 U17590 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14141) );
  AOI22_X1 U17591 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14140) );
  NAND4_X1 U17592 ( .A1(n14143), .A2(n14142), .A3(n14141), .A4(n14140), .ZN(
        n14144) );
  NOR2_X1 U17593 ( .A1(n14145), .A2(n14144), .ZN(n14149) );
  OAI21_X1 U17594 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20703), .A(
        n12749), .ZN(n14146) );
  INV_X1 U17595 ( .A(n14146), .ZN(n14147) );
  AOI21_X1 U17596 ( .B1(n14250), .B2(P1_EAX_REG_16__SCAN_IN), .A(n14147), .ZN(
        n14148) );
  OAI21_X1 U17597 ( .B1(n14434), .B2(n14149), .A(n14148), .ZN(n14153) );
  OAI21_X1 U17598 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n14151), .A(
        n14150), .ZN(n16054) );
  OR2_X1 U17599 ( .A1(n14363), .A2(n16054), .ZN(n14152) );
  NAND2_X1 U17600 ( .A1(n14153), .A2(n14152), .ZN(n14784) );
  INV_X1 U17601 ( .A(n14434), .ZN(n14402) );
  AOI22_X1 U17602 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14157) );
  AOI22_X1 U17603 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14156) );
  AOI22_X1 U17604 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14155) );
  AOI22_X1 U17605 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14368), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14154) );
  NAND4_X1 U17606 ( .A1(n14157), .A2(n14156), .A3(n14155), .A4(n14154), .ZN(
        n14163) );
  AOI22_X1 U17607 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14161) );
  AOI22_X1 U17608 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14331), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14160) );
  AOI22_X1 U17609 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14159) );
  AOI22_X1 U17610 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14158) );
  NAND4_X1 U17611 ( .A1(n14161), .A2(n14160), .A3(n14159), .A4(n14158), .ZN(
        n14162) );
  OR2_X1 U17612 ( .A1(n14163), .A2(n14162), .ZN(n14167) );
  XNOR2_X1 U17613 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n14164), .ZN(
        n15007) );
  AOI22_X1 U17614 ( .A1(n14437), .A2(n15007), .B1(n14439), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14165) );
  OAI21_X1 U17615 ( .B1(n9911), .B2(n13083), .A(n14165), .ZN(n14166) );
  AOI21_X1 U17616 ( .B1(n14402), .B2(n14167), .A(n14166), .ZN(n14765) );
  AOI22_X1 U17617 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14171) );
  AOI22_X1 U17618 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14170) );
  AOI22_X1 U17619 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14169) );
  AOI22_X1 U17620 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14168) );
  NAND4_X1 U17621 ( .A1(n14171), .A2(n14170), .A3(n14169), .A4(n14168), .ZN(
        n14177) );
  AOI22_X1 U17622 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14175) );
  AOI22_X1 U17623 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14174) );
  AOI22_X1 U17624 ( .A1(n14331), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14173) );
  AOI22_X1 U17625 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14172) );
  NAND4_X1 U17626 ( .A1(n14175), .A2(n14174), .A3(n14173), .A4(n14172), .ZN(
        n14176) );
  NOR2_X1 U17627 ( .A1(n14177), .A2(n14176), .ZN(n14179) );
  AOI22_X1 U17628 ( .A1(n14250), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12749), .ZN(n14178) );
  OAI21_X1 U17629 ( .B1(n14434), .B2(n14179), .A(n14178), .ZN(n14183) );
  INV_X1 U17630 ( .A(n14180), .ZN(n14181) );
  INV_X1 U17631 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14990) );
  NAND2_X1 U17632 ( .A1(n14181), .A2(n14990), .ZN(n14182) );
  NAND2_X1 U17633 ( .A1(n14196), .A2(n14182), .ZN(n14989) );
  MUX2_X1 U17634 ( .A(n14183), .B(n14989), .S(n14437), .Z(n14753) );
  AOI22_X1 U17635 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14187) );
  AOI22_X1 U17636 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14186) );
  AOI22_X1 U17637 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14185) );
  AOI22_X1 U17638 ( .A1(n12252), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14368), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14184) );
  NAND4_X1 U17639 ( .A1(n14187), .A2(n14186), .A3(n14185), .A4(n14184), .ZN(
        n14193) );
  AOI22_X1 U17640 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14191) );
  AOI22_X1 U17641 ( .A1(n12255), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14190) );
  AOI22_X1 U17642 ( .A1(n14352), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14189) );
  AOI22_X1 U17643 ( .A1(n14331), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14188) );
  NAND4_X1 U17644 ( .A1(n14191), .A2(n14190), .A3(n14189), .A4(n14188), .ZN(
        n14192) );
  NOR2_X1 U17645 ( .A1(n14193), .A2(n14192), .ZN(n14195) );
  AOI22_X1 U17646 ( .A1(n14250), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12749), .ZN(n14194) );
  OAI21_X1 U17647 ( .B1(n14434), .B2(n14195), .A(n14194), .ZN(n14197) );
  XNOR2_X1 U17648 ( .A(n14196), .B(n14743), .ZN(n14985) );
  MUX2_X1 U17649 ( .A(n14197), .B(n14985), .S(n14437), .Z(n14740) );
  AOI22_X1 U17650 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14203) );
  AOI22_X1 U17651 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14202) );
  AOI22_X1 U17652 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14201) );
  AOI22_X1 U17653 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14200) );
  NAND4_X1 U17654 ( .A1(n14203), .A2(n14202), .A3(n14201), .A4(n14200), .ZN(
        n14209) );
  AOI22_X1 U17655 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14207) );
  AOI22_X1 U17656 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14206) );
  AOI22_X1 U17657 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14205) );
  AOI22_X1 U17658 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14204) );
  NAND4_X1 U17659 ( .A1(n14207), .A2(n14206), .A3(n14205), .A4(n14204), .ZN(
        n14208) );
  NOR2_X1 U17660 ( .A1(n14209), .A2(n14208), .ZN(n14211) );
  AOI22_X1 U17661 ( .A1(n14250), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12749), .ZN(n14210) );
  OAI21_X1 U17662 ( .B1(n14434), .B2(n14211), .A(n14210), .ZN(n14212) );
  INV_X1 U17663 ( .A(n14212), .ZN(n14216) );
  INV_X1 U17664 ( .A(n14213), .ZN(n14214) );
  INV_X1 U17665 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14975) );
  NAND2_X1 U17666 ( .A1(n14214), .A2(n14975), .ZN(n14215) );
  AND2_X1 U17667 ( .A1(n14233), .A2(n14215), .ZN(n14979) );
  MUX2_X1 U17668 ( .A(n14216), .B(n14979), .S(n14437), .Z(n14730) );
  NAND2_X1 U17669 ( .A1(n14218), .A2(n14217), .ZN(n14717) );
  AOI22_X1 U17670 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n12660), .B1(
        n9808), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14222) );
  AOI22_X1 U17671 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n14198), .B1(
        n14367), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14221) );
  AOI22_X1 U17672 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14220) );
  AOI22_X1 U17673 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14219) );
  NAND4_X1 U17674 ( .A1(n14222), .A2(n14221), .A3(n14220), .A4(n14219), .ZN(
        n14229) );
  AOI22_X1 U17675 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n14368), .B1(
        n14331), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14227) );
  AOI22_X1 U17676 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14223), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14226) );
  AOI22_X1 U17677 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14225) );
  AOI22_X1 U17678 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14224) );
  NAND4_X1 U17679 ( .A1(n14227), .A2(n14226), .A3(n14225), .A4(n14224), .ZN(
        n14228) );
  NOR2_X1 U17680 ( .A1(n14229), .A2(n14228), .ZN(n14231) );
  AOI22_X1 U17681 ( .A1(n14250), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12749), .ZN(n14230) );
  OAI21_X1 U17682 ( .B1(n14434), .B2(n14231), .A(n14230), .ZN(n14232) );
  INV_X1 U17683 ( .A(n14232), .ZN(n14234) );
  XNOR2_X1 U17684 ( .A(n14233), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14969) );
  MUX2_X1 U17685 ( .A(n14234), .B(n14969), .S(n14437), .Z(n14719) );
  AOI22_X1 U17686 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14239) );
  AOI22_X1 U17687 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14238) );
  AOI22_X1 U17688 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14237) );
  AOI22_X1 U17689 ( .A1(n12252), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14368), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14236) );
  NAND4_X1 U17690 ( .A1(n14239), .A2(n14238), .A3(n14237), .A4(n14236), .ZN(
        n14247) );
  AOI22_X1 U17691 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14245) );
  AOI22_X1 U17692 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14244) );
  AOI22_X1 U17693 ( .A1(n14331), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14243) );
  AOI22_X1 U17694 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14242) );
  NAND4_X1 U17695 ( .A1(n14245), .A2(n14244), .A3(n14243), .A4(n14242), .ZN(
        n14246) );
  NOR2_X1 U17696 ( .A1(n14247), .A2(n14246), .ZN(n14252) );
  OAI21_X1 U17697 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20703), .A(
        n12749), .ZN(n14248) );
  INV_X1 U17698 ( .A(n14248), .ZN(n14249) );
  AOI21_X1 U17699 ( .B1(n14250), .B2(P1_EAX_REG_22__SCAN_IN), .A(n14249), .ZN(
        n14251) );
  OAI21_X1 U17700 ( .B1(n14434), .B2(n14252), .A(n14251), .ZN(n14258) );
  INV_X1 U17701 ( .A(n14253), .ZN(n14255) );
  INV_X1 U17702 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14254) );
  NAND2_X1 U17703 ( .A1(n14255), .A2(n14254), .ZN(n14256) );
  NAND2_X1 U17704 ( .A1(n14287), .A2(n14256), .ZN(n14959) );
  OR2_X1 U17705 ( .A1(n14959), .A2(n14363), .ZN(n14257) );
  INV_X1 U17706 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14268) );
  INV_X1 U17707 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14409) );
  INV_X1 U17708 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14259) );
  OAI22_X1 U17709 ( .A1(n14411), .A2(n14409), .B1(n12300), .B2(n14259), .ZN(
        n14265) );
  INV_X1 U17710 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14262) );
  INV_X1 U17711 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14260) );
  OAI22_X1 U17712 ( .A1(n14263), .A2(n14262), .B1(n14261), .B2(n14260), .ZN(
        n14264) );
  AOI211_X1 U17713 ( .C1(n13263), .C2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n14265), .B(n14264), .ZN(n14267) );
  AOI22_X1 U17714 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14266) );
  OAI211_X1 U17715 ( .C1(n12733), .C2(n14268), .A(n14267), .B(n14266), .ZN(
        n14274) );
  AOI22_X1 U17716 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14198), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14272) );
  AOI22_X1 U17717 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14271) );
  AOI22_X1 U17718 ( .A1(n14373), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14414), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14270) );
  AOI22_X1 U17719 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14331), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14269) );
  NAND4_X1 U17720 ( .A1(n14272), .A2(n14271), .A3(n14270), .A4(n14269), .ZN(
        n14273) );
  NOR2_X1 U17721 ( .A1(n14274), .A2(n14273), .ZN(n14290) );
  AOI22_X1 U17722 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14278) );
  AOI22_X1 U17723 ( .A1(n14418), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14277) );
  AOI22_X1 U17724 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14276) );
  AOI22_X1 U17725 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14275) );
  NAND4_X1 U17726 ( .A1(n14278), .A2(n14277), .A3(n14276), .A4(n14275), .ZN(
        n14284) );
  AOI22_X1 U17727 ( .A1(n14198), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14414), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14282) );
  AOI22_X1 U17728 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14281) );
  AOI22_X1 U17729 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14280) );
  AOI22_X1 U17730 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14279) );
  NAND4_X1 U17731 ( .A1(n14282), .A2(n14281), .A3(n14280), .A4(n14279), .ZN(
        n14283) );
  NOR2_X1 U17732 ( .A1(n14284), .A2(n14283), .ZN(n14289) );
  XOR2_X1 U17733 ( .A(n14290), .B(n14289), .Z(n14286) );
  INV_X1 U17734 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14950) );
  OAI22_X1 U17735 ( .A1(n9911), .A2(n12591), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14950), .ZN(n14285) );
  AOI21_X1 U17736 ( .B1(n14402), .B2(n14286), .A(n14285), .ZN(n14288) );
  XNOR2_X1 U17737 ( .A(n14287), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14952) );
  MUX2_X1 U17738 ( .A(n14288), .B(n14952), .S(n14437), .Z(n14696) );
  NOR2_X1 U17739 ( .A1(n14290), .A2(n14289), .ZN(n14310) );
  AOI22_X1 U17740 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14294) );
  AOI22_X1 U17741 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14293) );
  AOI22_X1 U17742 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14292) );
  AOI22_X1 U17743 ( .A1(n14394), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14291) );
  NAND4_X1 U17744 ( .A1(n14294), .A2(n14293), .A3(n14292), .A4(n14291), .ZN(
        n14301) );
  AOI22_X1 U17745 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14414), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14299) );
  AOI22_X1 U17746 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14298) );
  AOI22_X1 U17747 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14297) );
  AOI22_X1 U17748 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14296) );
  NAND4_X1 U17749 ( .A1(n14299), .A2(n14298), .A3(n14297), .A4(n14296), .ZN(
        n14300) );
  OR2_X1 U17750 ( .A1(n14301), .A2(n14300), .ZN(n14309) );
  XNOR2_X1 U17751 ( .A(n14310), .B(n14309), .ZN(n14303) );
  AOI22_X1 U17752 ( .A1(n14250), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12749), .ZN(n14302) );
  OAI21_X1 U17753 ( .B1(n14303), .B2(n14434), .A(n14302), .ZN(n14308) );
  INV_X1 U17754 ( .A(n14304), .ZN(n14306) );
  INV_X1 U17755 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14305) );
  NAND2_X1 U17756 ( .A1(n14306), .A2(n14305), .ZN(n14307) );
  NAND2_X1 U17757 ( .A1(n14323), .A2(n14307), .ZN(n14942) );
  MUX2_X1 U17758 ( .A(n14308), .B(n14942), .S(n14437), .Z(n14683) );
  NAND2_X1 U17759 ( .A1(n14310), .A2(n14309), .ZN(n14325) );
  AOI22_X1 U17760 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14314) );
  AOI22_X1 U17761 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14313) );
  AOI22_X1 U17762 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14368), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14312) );
  AOI22_X1 U17763 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14311) );
  NAND4_X1 U17764 ( .A1(n14314), .A2(n14313), .A3(n14312), .A4(n14311), .ZN(
        n14320) );
  AOI22_X1 U17765 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U17766 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14317) );
  AOI22_X1 U17767 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14316) );
  AOI22_X1 U17768 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14315) );
  NAND4_X1 U17769 ( .A1(n14318), .A2(n14317), .A3(n14316), .A4(n14315), .ZN(
        n14319) );
  NOR2_X1 U17770 ( .A1(n14320), .A2(n14319), .ZN(n14326) );
  XOR2_X1 U17771 ( .A(n14325), .B(n14326), .Z(n14322) );
  OAI22_X1 U17772 ( .A1(n9911), .A2(n21197), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14929), .ZN(n14321) );
  AOI21_X1 U17773 ( .B1(n14322), .B2(n14402), .A(n14321), .ZN(n14324) );
  XNOR2_X1 U17774 ( .A(n14323), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14931) );
  MUX2_X1 U17775 ( .A(n14324), .B(n14931), .S(n14437), .Z(n14673) );
  NOR2_X1 U17776 ( .A1(n14326), .A2(n14325), .ZN(n14347) );
  AOI22_X1 U17777 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12660), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14330) );
  AOI22_X1 U17778 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14329) );
  AOI22_X1 U17779 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14328) );
  AOI22_X1 U17780 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14327) );
  NAND4_X1 U17781 ( .A1(n14330), .A2(n14329), .A3(n14328), .A4(n14327), .ZN(
        n14337) );
  AOI22_X1 U17782 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14414), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14335) );
  AOI22_X1 U17783 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14334) );
  AOI22_X1 U17784 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14331), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14333) );
  AOI22_X1 U17785 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14240), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14332) );
  NAND4_X1 U17786 ( .A1(n14335), .A2(n14334), .A3(n14333), .A4(n14332), .ZN(
        n14336) );
  OR2_X1 U17787 ( .A1(n14337), .A2(n14336), .ZN(n14346) );
  XNOR2_X1 U17788 ( .A(n14347), .B(n14346), .ZN(n14339) );
  AOI22_X1 U17789 ( .A1(n14250), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n12749), .ZN(n14338) );
  OAI21_X1 U17790 ( .B1(n14339), .B2(n14434), .A(n14338), .ZN(n14343) );
  NAND2_X1 U17791 ( .A1(n14341), .A2(n14340), .ZN(n14342) );
  NAND2_X1 U17792 ( .A1(n14344), .A2(n14342), .ZN(n14924) );
  MUX2_X1 U17793 ( .A(n14343), .B(n14924), .S(n14437), .Z(n14660) );
  INV_X1 U17794 ( .A(n14344), .ZN(n14345) );
  XNOR2_X1 U17795 ( .A(n14345), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14915) );
  NAND2_X1 U17796 ( .A1(n14347), .A2(n14346), .ZN(n14364) );
  AOI22_X1 U17797 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14351) );
  AOI22_X1 U17798 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14350) );
  AOI22_X1 U17799 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14235), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14349) );
  AOI22_X1 U17800 ( .A1(n12252), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14348) );
  NAND4_X1 U17801 ( .A1(n14351), .A2(n14350), .A3(n14349), .A4(n14348), .ZN(
        n14358) );
  AOI22_X1 U17802 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14352), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14356) );
  AOI22_X1 U17803 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12236), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U17804 ( .A1(n12665), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14354) );
  AOI22_X1 U17805 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14353) );
  NAND4_X1 U17806 ( .A1(n14356), .A2(n14355), .A3(n14354), .A4(n14353), .ZN(
        n14357) );
  NOR2_X1 U17807 ( .A1(n14358), .A2(n14357), .ZN(n14365) );
  XOR2_X1 U17808 ( .A(n14364), .B(n14365), .Z(n14359) );
  NAND2_X1 U17809 ( .A1(n14359), .A2(n14402), .ZN(n14361) );
  OAI21_X1 U17810 ( .B1(n20703), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n12749), .ZN(n14360) );
  OAI211_X1 U17811 ( .C1(n9911), .C2(n21023), .A(n14361), .B(n14360), .ZN(
        n14362) );
  NOR2_X1 U17812 ( .A1(n14365), .A2(n14364), .ZN(n14388) );
  AOI22_X1 U17813 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n12660), .B1(
        n9808), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14372) );
  AOI22_X1 U17814 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n14367), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14371) );
  AOI22_X1 U17815 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14370) );
  AOI22_X1 U17816 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n14368), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14369) );
  NAND4_X1 U17817 ( .A1(n14372), .A2(n14371), .A3(n14370), .A4(n14369), .ZN(
        n14379) );
  AOI22_X1 U17818 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n14373), .B1(
        n12255), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U17819 ( .A1(n9800), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U17820 ( .A1(n14223), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14375) );
  AOI22_X1 U17821 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12236), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14374) );
  NAND4_X1 U17822 ( .A1(n14377), .A2(n14376), .A3(n14375), .A4(n14374), .ZN(
        n14378) );
  OR2_X1 U17823 ( .A1(n14379), .A2(n14378), .ZN(n14387) );
  XNOR2_X1 U17824 ( .A(n14388), .B(n14387), .ZN(n14381) );
  AOI22_X1 U17825 ( .A1(n14250), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n12749), .ZN(n14380) );
  OAI21_X1 U17826 ( .B1(n14381), .B2(n14434), .A(n14380), .ZN(n14386) );
  INV_X1 U17827 ( .A(n14382), .ZN(n14384) );
  INV_X1 U17828 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14383) );
  NAND2_X1 U17829 ( .A1(n14384), .A2(n14383), .ZN(n14385) );
  NAND2_X1 U17830 ( .A1(n14404), .A2(n14385), .ZN(n14907) );
  MUX2_X1 U17831 ( .A(n14386), .B(n14907), .S(n14437), .Z(n14636) );
  NAND2_X1 U17832 ( .A1(n14388), .A2(n14387), .ZN(n14429) );
  AOI22_X1 U17833 ( .A1(n9808), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13263), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14393) );
  AOI22_X1 U17834 ( .A1(n14367), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14422), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14392) );
  AOI22_X1 U17835 ( .A1(n12252), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14391) );
  AOI22_X1 U17836 ( .A1(n14240), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14295), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14390) );
  NAND4_X1 U17837 ( .A1(n14393), .A2(n14392), .A3(n14391), .A4(n14390), .ZN(
        n14400) );
  AOI22_X1 U17838 ( .A1(n14394), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14420), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14398) );
  AOI22_X1 U17839 ( .A1(n14198), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U17840 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12665), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14396) );
  AOI22_X1 U17841 ( .A1(n14235), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14199), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14395) );
  NAND4_X1 U17842 ( .A1(n14398), .A2(n14397), .A3(n14396), .A4(n14395), .ZN(
        n14399) );
  NOR2_X1 U17843 ( .A1(n14400), .A2(n14399), .ZN(n14430) );
  XOR2_X1 U17844 ( .A(n14429), .B(n14430), .Z(n14403) );
  INV_X1 U17845 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14895) );
  OAI22_X1 U17846 ( .A1(n9911), .A2(n21149), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14895), .ZN(n14401) );
  AOI21_X1 U17847 ( .B1(n14403), .B2(n14402), .A(n14401), .ZN(n14405) );
  XNOR2_X1 U17848 ( .A(n14404), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14893) );
  MUX2_X1 U17849 ( .A(n14405), .B(n14893), .S(n14437), .Z(n14624) );
  INV_X1 U17850 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14417) );
  INV_X1 U17851 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14407) );
  INV_X1 U17852 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14406) );
  OAI22_X1 U17853 ( .A1(n14408), .A2(n14407), .B1(n13868), .B2(n14406), .ZN(
        n14413) );
  INV_X1 U17854 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14410) );
  OAI22_X1 U17855 ( .A1(n14411), .A2(n14410), .B1(n12300), .B2(n14409), .ZN(
        n14412) );
  AOI211_X1 U17856 ( .C1(n13263), .C2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n14413), .B(n14412), .ZN(n14416) );
  AOI22_X1 U17857 ( .A1(n14414), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12665), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14415) );
  OAI211_X1 U17858 ( .C1(n12733), .C2(n14417), .A(n14416), .B(n14415), .ZN(
        n14428) );
  AOI22_X1 U17859 ( .A1(n14418), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14366), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14426) );
  AOI22_X1 U17860 ( .A1(n14368), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14425) );
  AOI22_X1 U17861 ( .A1(n14420), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12236), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14424) );
  AOI22_X1 U17862 ( .A1(n14422), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14421), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14423) );
  NAND4_X1 U17863 ( .A1(n14426), .A2(n14425), .A3(n14424), .A4(n14423), .ZN(
        n14427) );
  NOR2_X1 U17864 ( .A1(n14428), .A2(n14427), .ZN(n14432) );
  NOR2_X1 U17865 ( .A1(n14430), .A2(n14429), .ZN(n14431) );
  XOR2_X1 U17866 ( .A(n14432), .B(n14431), .Z(n14435) );
  AOI22_X1 U17867 ( .A1(n14250), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n12749), .ZN(n14433) );
  OAI21_X1 U17868 ( .B1(n14435), .B2(n14434), .A(n14433), .ZN(n14438) );
  XNOR2_X1 U17869 ( .A(n14436), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14885) );
  MUX2_X1 U17870 ( .A(n14438), .B(n14885), .S(n14437), .Z(n14612) );
  NAND2_X1 U17871 ( .A1(n14610), .A2(n14612), .ZN(n14611) );
  AOI22_X1 U17872 ( .A1(n14250), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n14439), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14440) );
  INV_X1 U17873 ( .A(n14440), .ZN(n14441) );
  XNOR2_X2 U17874 ( .A(n14611), .B(n14441), .ZN(n14536) );
  NAND2_X1 U17875 ( .A1(n14536), .A2(n16105), .ZN(n14445) );
  INV_X1 U17876 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21285) );
  NOR2_X1 U17877 ( .A1(n12853), .A2(n21285), .ZN(n15032) );
  NOR2_X1 U17878 ( .A1(n14442), .A2(n16110), .ZN(n14443) );
  AOI211_X1 U17879 ( .C1(n16099), .C2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15032), .B(n14443), .ZN(n14444) );
  OAI211_X1 U17880 ( .C1(n15048), .C2(n20095), .A(n14445), .B(n14444), .ZN(
        P1_U2968) );
  NOR2_X1 U17881 ( .A1(n14873), .A2(n14446), .ZN(n14448) );
  NAND2_X1 U17882 ( .A1(n14448), .A2(n20230), .ZN(n14827) );
  INV_X1 U17883 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20293) );
  AND2_X1 U17884 ( .A1(n14879), .A2(n20294), .ZN(n14447) );
  NAND2_X1 U17885 ( .A1(n14536), .A2(n14447), .ZN(n14450) );
  AOI22_X1 U17886 ( .A1(n14864), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14873), .ZN(n14449) );
  OAI211_X1 U17887 ( .C1(n14827), .C2(n20293), .A(n14450), .B(n14449), .ZN(
        P1_U2873) );
  NAND2_X1 U17888 ( .A1(n14459), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14454) );
  AOI21_X1 U17889 ( .B1(n16294), .B2(n14462), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15446) );
  INV_X1 U17890 ( .A(n16294), .ZN(n14456) );
  INV_X1 U17891 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14455) );
  INV_X1 U17892 ( .A(n14457), .ZN(n14461) );
  NOR2_X1 U17893 ( .A1(n14458), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14460) );
  MUX2_X1 U17894 ( .A(n14461), .B(n14460), .S(n14459), .Z(n16285) );
  NAND2_X1 U17895 ( .A1(n16285), .A2(n14462), .ZN(n14463) );
  XNOR2_X1 U17896 ( .A(n14463), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14464) );
  XNOR2_X1 U17897 ( .A(n14465), .B(n14464), .ZN(n15444) );
  AOI22_X1 U17898 ( .A1(n14468), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14470) );
  NAND2_X1 U17899 ( .A1(n11169), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14469) );
  OAI211_X1 U17900 ( .C1(n10615), .C2(n14471), .A(n14470), .B(n14469), .ZN(
        n14472) );
  INV_X1 U17901 ( .A(n14472), .ZN(n14473) );
  XNOR2_X1 U17902 ( .A(n14474), .B(n14473), .ZN(n16291) );
  INV_X1 U17903 ( .A(n14476), .ZN(n14478) );
  NAND2_X1 U17904 ( .A1(n14478), .A2(n14477), .ZN(n14481) );
  AOI222_X1 U17905 ( .A1(n11276), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11440), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n12080), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14479) );
  INV_X1 U17906 ( .A(n14479), .ZN(n14480) );
  NAND2_X1 U17907 ( .A1(n19404), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15438) );
  INV_X1 U17908 ( .A(n15438), .ZN(n14483) );
  NAND4_X1 U17909 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14484) );
  NOR3_X1 U17910 ( .A1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n14484), .A3(
        n15613), .ZN(n14482) );
  AOI211_X1 U17911 ( .C1(n19303), .C2(n19420), .A(n14483), .B(n14482), .ZN(
        n14488) );
  XNOR2_X1 U17912 ( .A(n15451), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15440) );
  INV_X1 U17913 ( .A(n14484), .ZN(n14486) );
  OAI21_X1 U17914 ( .B1(n15834), .B2(n14486), .A(n14485), .ZN(n15605) );
  NAND2_X1 U17915 ( .A1(n15605), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14487) );
  NAND3_X1 U17916 ( .A1(n14488), .A2(n10413), .A3(n14487), .ZN(n14489) );
  OAI21_X1 U17917 ( .B1(n15444), .B2(n19436), .A(n14490), .ZN(P2_U3015) );
  INV_X1 U17918 ( .A(n14492), .ZN(n14494) );
  NOR2_X1 U17919 ( .A1(n19277), .A2(n14493), .ZN(n15264) );
  OAI21_X1 U17920 ( .B1(n14495), .B2(n14494), .A(n15264), .ZN(n15279) );
  OAI21_X1 U17921 ( .B1(n9797), .B2(n19422), .A(n15279), .ZN(n14496) );
  INV_X1 U17922 ( .A(n14496), .ZN(n15855) );
  AOI22_X1 U17923 ( .A1(n19277), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19285), .B2(n14491), .ZN(n15849) );
  NOR2_X1 U17924 ( .A1(n15849), .A2(n14497), .ZN(n15854) );
  INV_X1 U17925 ( .A(n15854), .ZN(n14500) );
  INV_X1 U17926 ( .A(n20031), .ZN(n16563) );
  AOI22_X1 U17927 ( .A1(n20051), .A2(n16563), .B1(n20035), .B2(n14498), .ZN(
        n14499) );
  OAI21_X1 U17928 ( .B1(n15855), .B2(n14500), .A(n14499), .ZN(n14504) );
  OAI22_X1 U17929 ( .A1(n16562), .A2(n13298), .B1(n14502), .B2(n14501), .ZN(
        n14503) );
  AOI21_X1 U17930 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16561), .A(n14503), .ZN(
        n15880) );
  MUX2_X1 U17931 ( .A(n14504), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15880), .Z(P2_U3599) );
  NAND2_X1 U17932 ( .A1(n14505), .A2(n14506), .ZN(n14795) );
  INV_X1 U17933 ( .A(n14878), .ZN(n14875) );
  AOI22_X1 U17934 ( .A1(n14875), .A2(n14812), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14873), .ZN(n14507) );
  OAI21_X1 U17935 ( .B1(n16082), .B2(n14881), .A(n14507), .ZN(P1_U2892) );
  MUX2_X1 U17936 ( .A(n9804), .B(n10135), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n14508) );
  INV_X1 U17937 ( .A(n14508), .ZN(n14510) );
  NAND2_X1 U17938 ( .A1(n14593), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14509) );
  NAND2_X1 U17939 ( .A1(n14510), .A2(n14509), .ZN(n14511) );
  NAND2_X1 U17940 ( .A1(n14512), .A2(n14511), .ZN(n14799) );
  OAI21_X1 U17941 ( .B1(n14512), .B2(n14511), .A(n14799), .ZN(n16207) );
  INV_X1 U17942 ( .A(n16207), .ZN(n14519) );
  INV_X1 U17943 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14515) );
  AOI21_X1 U17944 ( .B1(n20110), .B2(P1_EBX_REG_12__SCAN_IN), .A(n20138), .ZN(
        n14514) );
  NAND2_X1 U17945 ( .A1(n20158), .A2(n16083), .ZN(n14513) );
  OAI211_X1 U17946 ( .C1(n20136), .C2(n14515), .A(n14514), .B(n14513), .ZN(
        n14518) );
  INV_X1 U17947 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21200) );
  NAND2_X1 U17948 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n14516), .ZN(n14602) );
  AOI21_X1 U17949 ( .B1(n21200), .B2(n14602), .A(n16031), .ZN(n14517) );
  AOI211_X1 U17950 ( .C1(n14519), .C2(n20144), .A(n14518), .B(n14517), .ZN(
        n14520) );
  OAI21_X1 U17951 ( .B1(n16082), .B2(n14774), .A(n14520), .ZN(P1_U2828) );
  XOR2_X1 U17952 ( .A(n14521), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n14527)
         );
  OR2_X1 U17953 ( .A1(n14523), .A2(n14522), .ZN(n14524) );
  NAND2_X1 U17954 ( .A1(n14525), .A2(n14524), .ZN(n19257) );
  MUX2_X1 U17955 ( .A(n19257), .B(n10885), .S(n15352), .Z(n14526) );
  OAI21_X1 U17956 ( .B1(n14527), .B2(n15359), .A(n14526), .ZN(P2_U2880) );
  INV_X1 U17957 ( .A(n14528), .ZN(n14530) );
  NOR2_X1 U17958 ( .A1(n14530), .A2(n14529), .ZN(n14531) );
  OAI211_X1 U17959 ( .C1(n14531), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15346), .B(n14521), .ZN(n14534) );
  NAND2_X1 U17960 ( .A1(n14532), .A2(n15356), .ZN(n14533) );
  OAI211_X1 U17961 ( .C1(n15356), .C2(n14535), .A(n14534), .B(n14533), .ZN(
        P2_U2881) );
  NAND2_X1 U17962 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14543) );
  INV_X1 U17963 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14905) );
  INV_X1 U17964 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21102) );
  NOR2_X1 U17965 ( .A1(n14905), .A2(n21102), .ZN(n14542) );
  NAND3_X1 U17966 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .A3(P1_REIP_REG_25__SCAN_IN), .ZN(n14607) );
  AND2_X1 U17967 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14603) );
  AND2_X1 U17968 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n15999) );
  NAND3_X1 U17969 ( .A1(n14603), .A2(P1_REIP_REG_15__SCAN_IN), .A3(n15999), 
        .ZN(n14537) );
  NAND2_X1 U17970 ( .A1(n9798), .A2(n14537), .ZN(n14538) );
  NAND3_X1 U17971 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .ZN(n14605) );
  NAND2_X1 U17972 ( .A1(n9798), .A2(n14605), .ZN(n14539) );
  NAND2_X1 U17973 ( .A1(n14766), .A2(n14539), .ZN(n14736) );
  INV_X1 U17974 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21148) );
  INV_X1 U17975 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21288) );
  INV_X1 U17976 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21209) );
  NOR3_X1 U17977 ( .A1(n21148), .A2(n21288), .A3(n21209), .ZN(n14606) );
  NOR2_X1 U17978 ( .A1(n14540), .A2(n14606), .ZN(n14541) );
  OAI21_X1 U17979 ( .B1(n15998), .B2(n14542), .A(n14649), .ZN(n14644) );
  AOI21_X1 U17980 ( .B1(n14543), .B2(n9798), .A(n14644), .ZN(n14618) );
  INV_X1 U17981 ( .A(n14618), .ZN(n14609) );
  INV_X1 U17982 ( .A(n14567), .ZN(n14599) );
  AOI22_X1 U17983 ( .A1(n14599), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14593), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14615) );
  MUX2_X1 U17984 ( .A(n14586), .B(n9804), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14544) );
  INV_X1 U17985 ( .A(n14544), .ZN(n14546) );
  NAND2_X1 U17986 ( .A1(n14567), .A2(n16141), .ZN(n14545) );
  NAND2_X1 U17987 ( .A1(n14546), .A2(n14545), .ZN(n14800) );
  MUX2_X1 U17988 ( .A(n9804), .B(n10135), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n14548) );
  AND2_X1 U17989 ( .A1(n14593), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14547) );
  NOR2_X1 U17990 ( .A1(n14548), .A2(n14547), .ZN(n14788) );
  MUX2_X1 U17991 ( .A(n14586), .B(n9804), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n14550) );
  NOR2_X1 U17992 ( .A1(n14599), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14549) );
  NOR2_X1 U17993 ( .A1(n14550), .A2(n14549), .ZN(n16003) );
  MUX2_X1 U17994 ( .A(n9804), .B(n10135), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n14551) );
  INV_X1 U17995 ( .A(n14551), .ZN(n14553) );
  NAND2_X1 U17996 ( .A1(n14593), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14552) );
  NAND2_X1 U17997 ( .A1(n14553), .A2(n14552), .ZN(n14785) );
  MUX2_X1 U17998 ( .A(n14586), .B(n9804), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14554) );
  INV_X1 U17999 ( .A(n14554), .ZN(n14556) );
  INV_X1 U18000 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15005) );
  NAND2_X1 U18001 ( .A1(n14567), .A2(n15005), .ZN(n14555) );
  INV_X1 U18002 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16145) );
  NAND2_X1 U18003 ( .A1(n14591), .A2(n16145), .ZN(n14557) );
  OAI211_X1 U18004 ( .C1(n14593), .C2(P1_EBX_REG_18__SCAN_IN), .A(n14614), .B(
        n14557), .ZN(n14559) );
  INV_X1 U18005 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21165) );
  NAND2_X1 U18006 ( .A1(n9804), .A2(n21165), .ZN(n14558) );
  AND2_X1 U18007 ( .A1(n14559), .A2(n14558), .ZN(n14754) );
  MUX2_X1 U18008 ( .A(n14586), .B(n9804), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n14560) );
  INV_X1 U18009 ( .A(n14560), .ZN(n14562) );
  INV_X1 U18010 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16123) );
  NAND2_X1 U18011 ( .A1(n14567), .A2(n16123), .ZN(n14561) );
  NAND2_X1 U18012 ( .A1(n14562), .A2(n14561), .ZN(n14742) );
  MUX2_X1 U18013 ( .A(n9804), .B(n10135), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n14563) );
  INV_X1 U18014 ( .A(n14563), .ZN(n14565) );
  NAND2_X1 U18015 ( .A1(n14593), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14564) );
  NAND2_X1 U18016 ( .A1(n14565), .A2(n14564), .ZN(n14731) );
  NAND2_X1 U18017 ( .A1(n14741), .A2(n14731), .ZN(n14733) );
  MUX2_X1 U18018 ( .A(n14586), .B(n9804), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n14566) );
  INV_X1 U18019 ( .A(n14566), .ZN(n14569) );
  INV_X1 U18020 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15134) );
  NAND2_X1 U18021 ( .A1(n14567), .A2(n15134), .ZN(n14568) );
  NAND2_X1 U18022 ( .A1(n14569), .A2(n14568), .ZN(n14720) );
  OR2_X2 U18023 ( .A1(n14733), .A2(n14720), .ZN(n14722) );
  NAND2_X1 U18024 ( .A1(n14591), .A2(n15133), .ZN(n14570) );
  OAI211_X1 U18025 ( .C1(n14593), .C2(P1_EBX_REG_22__SCAN_IN), .A(n14614), .B(
        n14570), .ZN(n14573) );
  INV_X1 U18026 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14571) );
  NAND2_X1 U18027 ( .A1(n9804), .A2(n14571), .ZN(n14572) );
  AND2_X1 U18028 ( .A1(n14573), .A2(n14572), .ZN(n14708) );
  INV_X1 U18029 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21224) );
  NAND2_X1 U18030 ( .A1(n14586), .A2(n21224), .ZN(n14576) );
  NAND2_X1 U18031 ( .A1(n14614), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14574) );
  OAI211_X1 U18032 ( .C1(n14593), .C2(P1_EBX_REG_23__SCAN_IN), .A(n14591), .B(
        n14574), .ZN(n14575) );
  AND2_X1 U18033 ( .A1(n14576), .A2(n14575), .ZN(n14697) );
  INV_X1 U18034 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15116) );
  NAND2_X1 U18035 ( .A1(n14591), .A2(n15116), .ZN(n14577) );
  OAI211_X1 U18036 ( .C1(n14593), .C2(P1_EBX_REG_24__SCAN_IN), .A(n14614), .B(
        n14577), .ZN(n14579) );
  INV_X1 U18037 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14778) );
  NAND2_X1 U18038 ( .A1(n9804), .A2(n14778), .ZN(n14578) );
  NAND2_X1 U18039 ( .A1(n14579), .A2(n14578), .ZN(n14685) );
  NAND2_X1 U18040 ( .A1(n14614), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14580) );
  OAI211_X1 U18041 ( .C1(n14593), .C2(P1_EBX_REG_25__SCAN_IN), .A(n14591), .B(
        n14580), .ZN(n14581) );
  OAI21_X1 U18042 ( .B1(n14582), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14581), .ZN(
        n14674) );
  NAND2_X1 U18043 ( .A1(n14591), .A2(n15029), .ZN(n14583) );
  OAI211_X1 U18044 ( .C1(n14593), .C2(P1_EBX_REG_26__SCAN_IN), .A(n14614), .B(
        n14583), .ZN(n14585) );
  INV_X1 U18045 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21072) );
  NAND2_X1 U18046 ( .A1(n9804), .A2(n21072), .ZN(n14584) );
  AND2_X1 U18047 ( .A1(n14585), .A2(n14584), .ZN(n14661) );
  NOR2_X2 U18048 ( .A1(n9816), .A2(n14661), .ZN(n14662) );
  INV_X1 U18049 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n21175) );
  NAND2_X1 U18050 ( .A1(n14586), .A2(n21175), .ZN(n14589) );
  NAND2_X1 U18051 ( .A1(n14614), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14587) );
  OAI211_X1 U18052 ( .C1(n14593), .C2(P1_EBX_REG_27__SCAN_IN), .A(n14591), .B(
        n14587), .ZN(n14588) );
  AND2_X1 U18053 ( .A1(n14589), .A2(n14588), .ZN(n14650) );
  AND2_X2 U18054 ( .A1(n14662), .A2(n14650), .ZN(n14652) );
  INV_X1 U18055 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14590) );
  NAND2_X1 U18056 ( .A1(n14591), .A2(n14590), .ZN(n14592) );
  OAI211_X1 U18057 ( .C1(n14593), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14614), .B(
        n14592), .ZN(n14595) );
  INV_X1 U18058 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n21009) );
  NAND2_X1 U18059 ( .A1(n9804), .A2(n21009), .ZN(n14594) );
  NAND2_X1 U18060 ( .A1(n14595), .A2(n14594), .ZN(n14637) );
  INV_X1 U18061 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U18062 ( .A1(n14597), .A2(n14596), .ZN(n14598) );
  OAI21_X1 U18063 ( .B1(n14599), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14598), .ZN(n14613) );
  MUX2_X1 U18064 ( .A(n14613), .B(n14598), .S(n9804), .Z(n14628) );
  MUX2_X1 U18065 ( .A(n14614), .B(n14615), .S(n14627), .Z(n14601) );
  AOI22_X1 U18066 ( .A1(n14599), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14593), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14600) );
  AOI22_X1 U18067 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n20110), .ZN(n14608) );
  NAND2_X1 U18068 ( .A1(n14603), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n14604) );
  OAI22_X1 U18069 ( .A1(n14627), .A2(n14614), .B1(n14613), .B2(n14639), .ZN(
        n14616) );
  XNOR2_X1 U18070 ( .A(n14616), .B(n14615), .ZN(n15053) );
  AOI22_X1 U18071 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n20110), .ZN(n14617) );
  OAI21_X1 U18072 ( .B1(n14885), .B2(n20140), .A(n14617), .ZN(n14621) );
  AOI21_X1 U18073 ( .B1(n14633), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14619) );
  NOR2_X1 U18074 ( .A1(n14619), .A2(n14618), .ZN(n14620) );
  AOI211_X1 U18075 ( .C1(n20144), .C2(n15053), .A(n14621), .B(n14620), .ZN(
        n14622) );
  OAI21_X1 U18076 ( .B1(n14888), .B2(n14774), .A(n14622), .ZN(P1_U2810) );
  INV_X1 U18077 ( .A(n14897), .ZN(n14811) );
  INV_X1 U18078 ( .A(n14893), .ZN(n14631) );
  AOI21_X1 U18079 ( .B1(n14628), .B2(n14639), .A(n14627), .ZN(n15061) );
  NAND2_X1 U18080 ( .A1(n15061), .A2(n20144), .ZN(n14630) );
  AOI22_X1 U18081 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n20110), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n14629) );
  OAI211_X1 U18082 ( .C1(n20140), .C2(n14631), .A(n14630), .B(n14629), .ZN(
        n14632) );
  AOI21_X1 U18083 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n14644), .A(n14632), 
        .ZN(n14635) );
  INV_X1 U18084 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20988) );
  NAND2_X1 U18085 ( .A1(n14633), .A2(n20988), .ZN(n14634) );
  OAI211_X1 U18086 ( .C1(n14811), .C2(n14774), .A(n14635), .B(n14634), .ZN(
        P1_U2811) );
  OAI21_X1 U18087 ( .B1(n14647), .B2(n14636), .A(n14623), .ZN(n14910) );
  OR2_X1 U18088 ( .A1(n14652), .A2(n14637), .ZN(n14638) );
  NAND2_X1 U18089 ( .A1(n15073), .A2(n20144), .ZN(n14641) );
  AOI22_X1 U18090 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n20110), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n14640) );
  OAI211_X1 U18091 ( .C1(n20140), .C2(n14907), .A(n14641), .B(n14640), .ZN(
        n14643) );
  NOR3_X1 U18092 ( .A1(n14658), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n21102), 
        .ZN(n14642) );
  AOI211_X1 U18093 ( .C1(P1_REIP_REG_28__SCAN_IN), .C2(n14644), .A(n14643), 
        .B(n14642), .ZN(n14645) );
  OAI21_X1 U18094 ( .B1(n14910), .B2(n14774), .A(n14645), .ZN(P1_U2812) );
  AOI21_X1 U18095 ( .B1(n14648), .B2(n14646), .A(n14647), .ZN(n14917) );
  NAND2_X1 U18096 ( .A1(n14917), .A2(n20128), .ZN(n14657) );
  INV_X1 U18097 ( .A(n14649), .ZN(n14669) );
  NOR2_X1 U18098 ( .A1(n14662), .A2(n14650), .ZN(n14651) );
  OR2_X1 U18099 ( .A1(n14652), .A2(n14651), .ZN(n15077) );
  NOR2_X1 U18100 ( .A1(n15077), .A2(n20162), .ZN(n14655) );
  AOI22_X1 U18101 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n20110), .B2(P1_EBX_REG_27__SCAN_IN), .ZN(n14653) );
  OAI21_X1 U18102 ( .B1(n14915), .B2(n20140), .A(n14653), .ZN(n14654) );
  AOI211_X1 U18103 ( .C1(n14669), .C2(P1_REIP_REG_27__SCAN_IN), .A(n14655), 
        .B(n14654), .ZN(n14656) );
  OAI211_X1 U18104 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14658), .A(n14657), 
        .B(n14656), .ZN(P1_U2813) );
  OAI21_X1 U18105 ( .B1(n14659), .B2(n14660), .A(n14646), .ZN(n14922) );
  AND2_X1 U18106 ( .A1(n9816), .A2(n14661), .ZN(n14663) );
  OR2_X1 U18107 ( .A1(n14663), .A2(n14662), .ZN(n15086) );
  AOI22_X1 U18108 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n20110), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n14666) );
  INV_X1 U18109 ( .A(n14924), .ZN(n14664) );
  NAND2_X1 U18110 ( .A1(n20158), .A2(n14664), .ZN(n14665) );
  OAI211_X1 U18111 ( .C1(n15086), .C2(n20162), .A(n14666), .B(n14665), .ZN(
        n14668) );
  INV_X1 U18112 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14928) );
  INV_X1 U18113 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21177) );
  NOR4_X1 U18114 ( .A1(n14694), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n14928), 
        .A4(n21177), .ZN(n14667) );
  AOI211_X1 U18115 ( .C1(P1_REIP_REG_26__SCAN_IN), .C2(n14669), .A(n14668), 
        .B(n14667), .ZN(n14670) );
  OAI21_X1 U18116 ( .B1(n14922), .B2(n14774), .A(n14670), .ZN(P1_U2814) );
  XNOR2_X1 U18118 ( .A(n14672), .B(n14673), .ZN(n14938) );
  INV_X1 U18119 ( .A(n14674), .ZN(n14675) );
  OAI21_X1 U18120 ( .B1(n10243), .B2(n14675), .A(n9816), .ZN(n15096) );
  AOI22_X1 U18121 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n20110), .B2(P1_EBX_REG_25__SCAN_IN), .ZN(n14677) );
  NAND2_X1 U18122 ( .A1(n20158), .A2(n14931), .ZN(n14676) );
  OAI211_X1 U18123 ( .C1(n15096), .C2(n20162), .A(n14677), .B(n14676), .ZN(
        n14680) );
  XNOR2_X1 U18124 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14678) );
  NOR2_X1 U18125 ( .A1(n14694), .A2(n14678), .ZN(n14679) );
  AOI211_X1 U18126 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14702), .A(n14680), 
        .B(n14679), .ZN(n14681) );
  OAI21_X1 U18127 ( .B1(n14938), .B2(n14774), .A(n14681), .ZN(P1_U2815) );
  OAI21_X1 U18128 ( .B1(n14682), .B2(n14683), .A(n14672), .ZN(n14946) );
  INV_X1 U18129 ( .A(n14946), .ZN(n14684) );
  NAND2_X1 U18130 ( .A1(n14684), .A2(n20128), .ZN(n14693) );
  OR2_X1 U18131 ( .A1(n14699), .A2(n14685), .ZN(n14686) );
  NAND2_X1 U18132 ( .A1(n14687), .A2(n14686), .ZN(n15109) );
  AOI22_X1 U18133 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n20110), .B2(P1_EBX_REG_24__SCAN_IN), .ZN(n14690) );
  INV_X1 U18134 ( .A(n14942), .ZN(n14688) );
  NAND2_X1 U18135 ( .A1(n20158), .A2(n14688), .ZN(n14689) );
  OAI211_X1 U18136 ( .C1(n15109), .C2(n20162), .A(n14690), .B(n14689), .ZN(
        n14691) );
  AOI21_X1 U18137 ( .B1(n14702), .B2(P1_REIP_REG_24__SCAN_IN), .A(n14691), 
        .ZN(n14692) );
  OAI211_X1 U18138 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(n14694), .A(n14693), 
        .B(n14692), .ZN(P1_U2816) );
  AOI21_X1 U18139 ( .B1(n14696), .B2(n14695), .A(n14682), .ZN(n14949) );
  INV_X1 U18140 ( .A(n14949), .ZN(n14839) );
  OAI22_X1 U18141 ( .A1(n20136), .A2(n14950), .B1(n20156), .B2(n21224), .ZN(
        n14701) );
  NOR2_X1 U18142 ( .A1(n14710), .A2(n14697), .ZN(n14698) );
  OR2_X1 U18143 ( .A1(n14699), .A2(n14698), .ZN(n15122) );
  NOR2_X1 U18144 ( .A1(n15122), .A2(n20162), .ZN(n14700) );
  AOI211_X1 U18145 ( .C1(n20158), .C2(n14952), .A(n14701), .B(n14700), .ZN(
        n14705) );
  NOR3_X1 U18146 ( .A1(n9848), .A2(n21288), .A3(n21209), .ZN(n14703) );
  OAI21_X1 U18147 ( .B1(n14703), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14702), 
        .ZN(n14704) );
  OAI211_X1 U18148 ( .C1(n14839), .C2(n14774), .A(n14705), .B(n14704), .ZN(
        P1_U2817) );
  OAI21_X1 U18149 ( .B1(n14706), .B2(n14707), .A(n14695), .ZN(n14957) );
  AND2_X1 U18150 ( .A1(n14722), .A2(n14708), .ZN(n14709) );
  NOR2_X1 U18151 ( .A1(n14710), .A2(n14709), .ZN(n15127) );
  NAND2_X1 U18152 ( .A1(n15127), .A2(n20144), .ZN(n14712) );
  AOI22_X1 U18153 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20110), .B2(P1_EBX_REG_22__SCAN_IN), .ZN(n14711) );
  OAI211_X1 U18154 ( .C1(n20140), .C2(n14959), .A(n14712), .B(n14711), .ZN(
        n14715) );
  XNOR2_X1 U18155 ( .A(P1_REIP_REG_21__SCAN_IN), .B(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14713) );
  NOR2_X1 U18156 ( .A1(n9848), .A2(n14713), .ZN(n14714) );
  AOI211_X1 U18157 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14736), .A(n14715), 
        .B(n14714), .ZN(n14716) );
  OAI21_X1 U18158 ( .B1(n14957), .B2(n14774), .A(n14716), .ZN(P1_U2818) );
  AOI21_X1 U18159 ( .B1(n14719), .B2(n14718), .A(n14706), .ZN(n14966) );
  NAND2_X1 U18160 ( .A1(n14966), .A2(n20128), .ZN(n14727) );
  NAND2_X1 U18161 ( .A1(n14733), .A2(n14720), .ZN(n14721) );
  NAND2_X1 U18162 ( .A1(n14722), .A2(n14721), .ZN(n15964) );
  AOI22_X1 U18163 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20110), .B2(P1_EBX_REG_21__SCAN_IN), .ZN(n14724) );
  NAND2_X1 U18164 ( .A1(n20158), .A2(n14969), .ZN(n14723) );
  OAI211_X1 U18165 ( .C1(n15964), .C2(n20162), .A(n14724), .B(n14723), .ZN(
        n14725) );
  AOI21_X1 U18166 ( .B1(n14736), .B2(P1_REIP_REG_21__SCAN_IN), .A(n14725), 
        .ZN(n14726) );
  OAI211_X1 U18167 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(n9848), .A(n14727), .B(
        n14726), .ZN(P1_U2819) );
  OAI21_X1 U18168 ( .B1(n14218), .B2(n14217), .A(n14718), .ZN(n14976) );
  INV_X1 U18169 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n21180) );
  OAI22_X1 U18170 ( .A1(n20136), .A2(n14975), .B1(n20156), .B2(n21180), .ZN(
        n14735) );
  OR2_X1 U18171 ( .A1(n14741), .A2(n14731), .ZN(n14732) );
  NAND2_X1 U18172 ( .A1(n14733), .A2(n14732), .ZN(n15147) );
  NOR2_X1 U18173 ( .A1(n15147), .A2(n20162), .ZN(n14734) );
  AOI211_X1 U18174 ( .C1(n20158), .C2(n14979), .A(n14735), .B(n14734), .ZN(
        n14739) );
  INV_X1 U18175 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21024) );
  INV_X1 U18176 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21237) );
  OR2_X1 U18177 ( .A1(n21024), .A2(n21237), .ZN(n14749) );
  NOR2_X1 U18178 ( .A1(n14748), .A2(n14749), .ZN(n14737) );
  OAI21_X1 U18179 ( .B1(n14737), .B2(P1_REIP_REG_20__SCAN_IN), .A(n14736), 
        .ZN(n14738) );
  OAI211_X1 U18180 ( .C1(n14976), .C2(n14774), .A(n14739), .B(n14738), .ZN(
        P1_U2820) );
  OAI21_X1 U18181 ( .B1(n9870), .B2(n14740), .A(n14729), .ZN(n14983) );
  AOI21_X1 U18182 ( .B1(n14742), .B2(n14756), .A(n14741), .ZN(n16118) );
  NOR2_X1 U18183 ( .A1(n20136), .A2(n14743), .ZN(n14744) );
  AOI211_X1 U18184 ( .C1(P1_EBX_REG_19__SCAN_IN), .C2(n20110), .A(n20138), .B(
        n14744), .ZN(n14745) );
  OAI21_X1 U18185 ( .B1(n14985), .B2(n20140), .A(n14745), .ZN(n14747) );
  NOR2_X1 U18186 ( .A1(n14766), .A2(n21024), .ZN(n14746) );
  AOI211_X1 U18187 ( .C1(n16118), .C2(n20144), .A(n14747), .B(n14746), .ZN(
        n14751) );
  INV_X1 U18188 ( .A(n14748), .ZN(n14762) );
  OAI211_X1 U18189 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(P1_REIP_REG_19__SCAN_IN), .A(n14762), .B(n14749), .ZN(n14750) );
  OAI211_X1 U18190 ( .C1(n14983), .C2(n14774), .A(n14751), .B(n14750), .ZN(
        P1_U2821) );
  INV_X1 U18191 ( .A(n9870), .ZN(n14752) );
  OAI21_X1 U18192 ( .B1(n9850), .B2(n14753), .A(n14752), .ZN(n14998) );
  NAND2_X1 U18193 ( .A1(n9817), .A2(n14754), .ZN(n14755) );
  NAND2_X1 U18194 ( .A1(n14756), .A2(n14755), .ZN(n16144) );
  OAI21_X1 U18195 ( .B1(n20156), .B2(n21165), .A(n20154), .ZN(n14758) );
  NOR2_X1 U18196 ( .A1(n20140), .A2(n14989), .ZN(n14757) );
  AOI211_X1 U18197 ( .C1(n20153), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n14758), .B(n14757), .ZN(n14759) );
  OAI21_X1 U18198 ( .B1(n16144), .B2(n20162), .A(n14759), .ZN(n14761) );
  NOR2_X1 U18199 ( .A1(n14766), .A2(n21237), .ZN(n14760) );
  AOI211_X1 U18200 ( .C1(n14762), .C2(n21237), .A(n14761), .B(n14760), .ZN(
        n14763) );
  OAI21_X1 U18201 ( .B1(n14998), .B2(n14774), .A(n14763), .ZN(P1_U2822) );
  AOI21_X1 U18202 ( .B1(n14765), .B2(n14764), .A(n9850), .ZN(n15009) );
  INV_X1 U18203 ( .A(n15009), .ZN(n14859) );
  NAND2_X1 U18204 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n15992) );
  INV_X1 U18205 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21210) );
  OAI21_X1 U18206 ( .B1(n16012), .B2(n15992), .A(n21210), .ZN(n14772) );
  INV_X1 U18207 ( .A(n14766), .ZN(n14771) );
  OAI21_X1 U18208 ( .B1(n10239), .B2(n9931), .A(n9817), .ZN(n16154) );
  INV_X1 U18209 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n21222) );
  OAI21_X1 U18210 ( .B1(n21222), .B2(n20156), .A(n20154), .ZN(n14768) );
  NOR2_X1 U18211 ( .A1(n20140), .A2(n15007), .ZN(n14767) );
  AOI211_X1 U18212 ( .C1(n20153), .C2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n14768), .B(n14767), .ZN(n14769) );
  OAI21_X1 U18213 ( .B1(n16154), .B2(n20162), .A(n14769), .ZN(n14770) );
  AOI21_X1 U18214 ( .B1(n14772), .B2(n14771), .A(n14770), .ZN(n14773) );
  OAI21_X1 U18215 ( .B1(n14859), .B2(n14774), .A(n14773), .ZN(P1_U2823) );
  INV_X1 U18216 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n21037) );
  OAI22_X1 U18217 ( .A1(n15024), .A2(n20171), .B1(n20185), .B2(n21037), .ZN(
        P1_U2841) );
  AOI22_X1 U18218 ( .A1(n15053), .A2(n20181), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n14801), .ZN(n14775) );
  OAI21_X1 U18219 ( .B1(n14888), .B2(n14803), .A(n14775), .ZN(P1_U2842) );
  AOI22_X1 U18220 ( .A1(n15061), .A2(n20181), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14801), .ZN(n14776) );
  OAI21_X1 U18221 ( .B1(n14811), .B2(n14803), .A(n14776), .ZN(P1_U2843) );
  INV_X1 U18222 ( .A(n15073), .ZN(n14777) );
  OAI222_X1 U18223 ( .A1(n14777), .A2(n20171), .B1(n21009), .B2(n20185), .C1(
        n14910), .C2(n14803), .ZN(P1_U2844) );
  INV_X1 U18224 ( .A(n14917), .ZN(n14822) );
  OAI222_X1 U18225 ( .A1(n14803), .A2(n14822), .B1(n21175), .B2(n20185), .C1(
        n15077), .C2(n20171), .ZN(P1_U2845) );
  OAI222_X1 U18226 ( .A1(n14922), .A2(n14803), .B1(n21072), .B2(n20185), .C1(
        n15086), .C2(n20171), .ZN(P1_U2846) );
  INV_X1 U18227 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21235) );
  OAI222_X1 U18228 ( .A1(n20171), .A2(n15096), .B1(n21235), .B2(n20185), .C1(
        n14803), .C2(n14938), .ZN(P1_U2847) );
  OAI222_X1 U18229 ( .A1(n14946), .A2(n14803), .B1(n14778), .B2(n20185), .C1(
        n15109), .C2(n20171), .ZN(P1_U2848) );
  OAI222_X1 U18230 ( .A1(n15122), .A2(n20171), .B1(n21224), .B2(n20185), .C1(
        n14839), .C2(n14803), .ZN(P1_U2849) );
  AOI22_X1 U18231 ( .A1(n15127), .A2(n20181), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14801), .ZN(n14779) );
  OAI21_X1 U18232 ( .B1(n14957), .B2(n14803), .A(n14779), .ZN(P1_U2850) );
  INV_X1 U18233 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14780) );
  INV_X1 U18234 ( .A(n14966), .ZN(n14846) );
  OAI222_X1 U18235 ( .A1(n15964), .A2(n20171), .B1(n14780), .B2(n20185), .C1(
        n14846), .C2(n14803), .ZN(P1_U2851) );
  OAI222_X1 U18236 ( .A1(n14976), .A2(n14803), .B1(n21180), .B2(n20185), .C1(
        n15147), .C2(n20171), .ZN(P1_U2852) );
  AOI22_X1 U18237 ( .A1(n16118), .A2(n20181), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14801), .ZN(n14781) );
  OAI21_X1 U18238 ( .B1(n14983), .B2(n14803), .A(n14781), .ZN(P1_U2853) );
  OAI222_X1 U18239 ( .A1(n16144), .A2(n20171), .B1(n21165), .B2(n20185), .C1(
        n14998), .C2(n14803), .ZN(P1_U2854) );
  OAI222_X1 U18240 ( .A1(n14859), .A2(n14803), .B1(n20185), .B2(n21222), .C1(
        n16154), .C2(n20171), .ZN(P1_U2855) );
  INV_X1 U18241 ( .A(n14764), .ZN(n14783) );
  AOI21_X1 U18242 ( .B1(n14784), .B2(n14782), .A(n14783), .ZN(n16051) );
  INV_X1 U18243 ( .A(n16051), .ZN(n14867) );
  INV_X1 U18244 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21164) );
  OR2_X1 U18245 ( .A1(n16006), .A2(n14785), .ZN(n14786) );
  NAND2_X1 U18246 ( .A1(n14787), .A2(n14786), .ZN(n16164) );
  OAI222_X1 U18247 ( .A1(n14867), .A2(n14803), .B1(n20185), .B2(n21164), .C1(
        n16164), .C2(n20171), .ZN(P1_U2856) );
  AND2_X1 U18248 ( .A1(n14797), .A2(n14788), .ZN(n14789) );
  NOR2_X1 U18249 ( .A1(n16004), .A2(n14789), .ZN(n16015) );
  INV_X1 U18250 ( .A(n16015), .ZN(n16178) );
  INV_X1 U18251 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n21127) );
  OAI21_X1 U18252 ( .B1(n14790), .B2(n14793), .A(n14792), .ZN(n16014) );
  OAI222_X1 U18253 ( .A1(n16178), .A2(n20171), .B1(n20185), .B2(n21127), .C1(
        n16014), .C2(n14803), .ZN(P1_U2858) );
  AND2_X1 U18254 ( .A1(n14795), .A2(n14794), .ZN(n14796) );
  OR2_X1 U18255 ( .A1(n14790), .A2(n14796), .ZN(n15014) );
  INV_X1 U18256 ( .A(n14797), .ZN(n14798) );
  AOI21_X1 U18257 ( .B1(n14800), .B2(n14799), .A(n14798), .ZN(n16189) );
  AOI22_X1 U18258 ( .A1(n16189), .A2(n20181), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14801), .ZN(n14802) );
  OAI21_X1 U18259 ( .B1(n15014), .B2(n14803), .A(n14802), .ZN(P1_U2859) );
  INV_X1 U18260 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n21125) );
  OAI222_X1 U18261 ( .A1(n16207), .A2(n20171), .B1(n20185), .B2(n21125), .C1(
        n16082), .C2(n14803), .ZN(P1_U2860) );
  INV_X1 U18262 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14805) );
  NOR3_X1 U18263 ( .A1(n14873), .A2(n20294), .A3(n20280), .ZN(n14813) );
  AOI22_X1 U18264 ( .A1(n14813), .A2(n14874), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n14873), .ZN(n14804) );
  OAI21_X1 U18265 ( .B1(n14805), .B2(n14827), .A(n14804), .ZN(n14806) );
  AOI21_X1 U18266 ( .B1(n14864), .B2(DATAI_30_), .A(n14806), .ZN(n14807) );
  OAI21_X1 U18267 ( .B1(n14888), .B2(n14881), .A(n14807), .ZN(P1_U2874) );
  OAI22_X1 U18268 ( .A1(n14861), .A2(n14877), .B1(n14879), .B2(n21149), .ZN(
        n14808) );
  AOI21_X1 U18269 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14863), .A(n14808), .ZN(
        n14810) );
  NAND2_X1 U18270 ( .A1(n14864), .A2(DATAI_29_), .ZN(n14809) );
  OAI211_X1 U18271 ( .C1(n14811), .C2(n14881), .A(n14810), .B(n14809), .ZN(
        P1_U2875) );
  INV_X1 U18272 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n14815) );
  AOI22_X1 U18273 ( .A1(n14813), .A2(n14812), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n14873), .ZN(n14814) );
  OAI21_X1 U18274 ( .B1(n14815), .B2(n14827), .A(n14814), .ZN(n14816) );
  AOI21_X1 U18275 ( .B1(n14864), .B2(DATAI_28_), .A(n14816), .ZN(n14817) );
  OAI21_X1 U18276 ( .B1(n14910), .B2(n14881), .A(n14817), .ZN(P1_U2876) );
  OAI22_X1 U18277 ( .A1(n14861), .A2(n14818), .B1(n14879), .B2(n21023), .ZN(
        n14819) );
  AOI21_X1 U18278 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14863), .A(n14819), .ZN(
        n14821) );
  NAND2_X1 U18279 ( .A1(n14864), .A2(DATAI_27_), .ZN(n14820) );
  OAI211_X1 U18280 ( .C1(n14822), .C2(n14881), .A(n14821), .B(n14820), .ZN(
        P1_U2877) );
  OAI22_X1 U18281 ( .A1(n14861), .A2(n14823), .B1(n14879), .B2(n21206), .ZN(
        n14824) );
  AOI21_X1 U18282 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14863), .A(n14824), .ZN(
        n14826) );
  NAND2_X1 U18283 ( .A1(n14864), .A2(DATAI_26_), .ZN(n14825) );
  OAI211_X1 U18284 ( .C1(n14922), .C2(n14881), .A(n14826), .B(n14825), .ZN(
        P1_U2878) );
  INV_X1 U18285 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20253) );
  NOR2_X1 U18286 ( .A1(n14827), .A2(n20253), .ZN(n14830) );
  OAI22_X1 U18287 ( .A1(n14861), .A2(n14828), .B1(n14879), .B2(n21197), .ZN(
        n14829) );
  AOI211_X1 U18288 ( .C1(DATAI_25_), .C2(n14864), .A(n14830), .B(n14829), .ZN(
        n14831) );
  OAI21_X1 U18289 ( .B1(n14938), .B2(n14881), .A(n14831), .ZN(P1_U2879) );
  OAI22_X1 U18290 ( .A1(n14861), .A2(n14832), .B1(n14879), .B2(n12607), .ZN(
        n14833) );
  AOI21_X1 U18291 ( .B1(n14863), .B2(BUF1_REG_24__SCAN_IN), .A(n14833), .ZN(
        n14835) );
  NAND2_X1 U18292 ( .A1(n14864), .A2(DATAI_24_), .ZN(n14834) );
  OAI211_X1 U18293 ( .C1(n14946), .C2(n14881), .A(n14835), .B(n14834), .ZN(
        P1_U2880) );
  OAI22_X1 U18294 ( .A1(n14861), .A2(n20297), .B1(n14879), .B2(n12591), .ZN(
        n14836) );
  AOI21_X1 U18295 ( .B1(n14863), .B2(BUF1_REG_23__SCAN_IN), .A(n14836), .ZN(
        n14838) );
  NAND2_X1 U18296 ( .A1(n14864), .A2(DATAI_23_), .ZN(n14837) );
  OAI211_X1 U18297 ( .C1(n14839), .C2(n14881), .A(n14838), .B(n14837), .ZN(
        P1_U2881) );
  OAI22_X1 U18298 ( .A1(n14861), .A2(n20287), .B1(n14879), .B2(n21191), .ZN(
        n14840) );
  AOI21_X1 U18299 ( .B1(n14863), .B2(BUF1_REG_22__SCAN_IN), .A(n14840), .ZN(
        n14842) );
  NAND2_X1 U18300 ( .A1(n14864), .A2(DATAI_22_), .ZN(n14841) );
  OAI211_X1 U18301 ( .C1(n14957), .C2(n14881), .A(n14842), .B(n14841), .ZN(
        P1_U2882) );
  OAI22_X1 U18302 ( .A1(n14861), .A2(n20281), .B1(n14879), .B2(n21132), .ZN(
        n14843) );
  AOI21_X1 U18303 ( .B1(n14863), .B2(BUF1_REG_21__SCAN_IN), .A(n14843), .ZN(
        n14845) );
  NAND2_X1 U18304 ( .A1(n14864), .A2(DATAI_21_), .ZN(n14844) );
  OAI211_X1 U18305 ( .C1(n14846), .C2(n14881), .A(n14845), .B(n14844), .ZN(
        P1_U2883) );
  OAI22_X1 U18306 ( .A1(n14861), .A2(n20274), .B1(n14879), .B2(n21155), .ZN(
        n14847) );
  AOI21_X1 U18307 ( .B1(n14863), .B2(BUF1_REG_20__SCAN_IN), .A(n14847), .ZN(
        n14849) );
  NAND2_X1 U18308 ( .A1(n14864), .A2(DATAI_20_), .ZN(n14848) );
  OAI211_X1 U18309 ( .C1(n14976), .C2(n14881), .A(n14849), .B(n14848), .ZN(
        P1_U2884) );
  OAI22_X1 U18310 ( .A1(n14861), .A2(n20269), .B1(n14879), .B2(n12588), .ZN(
        n14850) );
  AOI21_X1 U18311 ( .B1(n14863), .B2(BUF1_REG_19__SCAN_IN), .A(n14850), .ZN(
        n14852) );
  NAND2_X1 U18312 ( .A1(n14864), .A2(DATAI_19_), .ZN(n14851) );
  OAI211_X1 U18313 ( .C1(n14983), .C2(n14881), .A(n14852), .B(n14851), .ZN(
        P1_U2885) );
  OAI22_X1 U18314 ( .A1(n14861), .A2(n20262), .B1(n14879), .B2(n13088), .ZN(
        n14853) );
  AOI21_X1 U18315 ( .B1(n14863), .B2(BUF1_REG_18__SCAN_IN), .A(n14853), .ZN(
        n14855) );
  NAND2_X1 U18316 ( .A1(n14864), .A2(DATAI_18_), .ZN(n14854) );
  OAI211_X1 U18317 ( .C1(n14998), .C2(n14881), .A(n14855), .B(n14854), .ZN(
        P1_U2886) );
  OAI22_X1 U18318 ( .A1(n14861), .A2(n20255), .B1(n14879), .B2(n13083), .ZN(
        n14856) );
  AOI21_X1 U18319 ( .B1(n14863), .B2(BUF1_REG_17__SCAN_IN), .A(n14856), .ZN(
        n14858) );
  NAND2_X1 U18320 ( .A1(n14864), .A2(DATAI_17_), .ZN(n14857) );
  OAI211_X1 U18321 ( .C1(n14859), .C2(n14881), .A(n14858), .B(n14857), .ZN(
        P1_U2887) );
  OAI22_X1 U18322 ( .A1(n14861), .A2(n20244), .B1(n14879), .B2(n14860), .ZN(
        n14862) );
  AOI21_X1 U18323 ( .B1(n14863), .B2(BUF1_REG_16__SCAN_IN), .A(n14862), .ZN(
        n14866) );
  NAND2_X1 U18324 ( .A1(n14864), .A2(DATAI_16_), .ZN(n14865) );
  OAI211_X1 U18325 ( .C1(n14867), .C2(n14881), .A(n14866), .B(n14865), .ZN(
        P1_U2888) );
  INV_X1 U18326 ( .A(n14782), .ZN(n14868) );
  AOI21_X1 U18327 ( .B1(n14869), .B2(n14792), .A(n14868), .ZN(n16060) );
  INV_X1 U18328 ( .A(n16060), .ZN(n14872) );
  OAI222_X1 U18329 ( .A1(n14881), .A2(n14872), .B1(n14879), .B2(n14871), .C1(
        n14878), .C2(n14870), .ZN(P1_U2889) );
  AOI22_X1 U18330 ( .A1(n14875), .A2(n14874), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14873), .ZN(n14876) );
  OAI21_X1 U18331 ( .B1(n16014), .B2(n14881), .A(n14876), .ZN(P1_U2890) );
  INV_X1 U18332 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14880) );
  OAI222_X1 U18333 ( .A1(n15014), .A2(n14881), .B1(n14880), .B2(n14879), .C1(
        n14878), .C2(n14877), .ZN(P1_U2891) );
  XNOR2_X1 U18334 ( .A(n14883), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15049) );
  NAND2_X1 U18335 ( .A1(n16255), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15056) );
  NAND2_X1 U18336 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14884) );
  OAI211_X1 U18337 ( .C1(n16110), .C2(n14885), .A(n15056), .B(n14884), .ZN(
        n14886) );
  AOI21_X1 U18338 ( .B1(n15049), .B2(n16113), .A(n14886), .ZN(n14887) );
  INV_X1 U18339 ( .A(n14889), .ZN(n14890) );
  AOI21_X1 U18340 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16068), .A(
        n14890), .ZN(n14891) );
  XNOR2_X1 U18341 ( .A(n14892), .B(n14891), .ZN(n15066) );
  NAND2_X1 U18342 ( .A1(n16084), .A2(n14893), .ZN(n14894) );
  NAND2_X1 U18343 ( .A1(n16255), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15058) );
  OAI211_X1 U18344 ( .C1(n16116), .C2(n14895), .A(n14894), .B(n15058), .ZN(
        n14896) );
  AOI21_X1 U18345 ( .B1(n14897), .B2(n16105), .A(n14896), .ZN(n14898) );
  OAI21_X1 U18346 ( .B1(n15066), .B2(n20095), .A(n14898), .ZN(P1_U2970) );
  INV_X1 U18347 ( .A(n15041), .ZN(n15090) );
  OAI21_X1 U18348 ( .B1(n10354), .B2(n15090), .A(n14948), .ZN(n14903) );
  INV_X1 U18349 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15118) );
  NAND3_X1 U18350 ( .A1(n14899), .A2(n15029), .A3(n15118), .ZN(n14901) );
  MUX2_X1 U18351 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n15029), .S(
        n16090), .Z(n14900) );
  AOI21_X1 U18352 ( .B1(n14903), .B2(n14901), .A(n14900), .ZN(n14902) );
  OAI21_X1 U18353 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14903), .A(
        n14902), .ZN(n14904) );
  XNOR2_X1 U18354 ( .A(n14904), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15067) );
  NOR2_X1 U18355 ( .A1(n12853), .A2(n14905), .ZN(n15069) );
  AOI21_X1 U18356 ( .B1(n16099), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15069), .ZN(n14906) );
  OAI21_X1 U18357 ( .B1(n14907), .B2(n16110), .A(n14906), .ZN(n14908) );
  AOI21_X1 U18358 ( .B1(n15067), .B2(n16113), .A(n14908), .ZN(n14909) );
  OAI21_X1 U18359 ( .B1(n14910), .B2(n16111), .A(n14909), .ZN(P1_U2971) );
  MUX2_X1 U18360 ( .A(n14912), .B(n14911), .S(n10354), .Z(n14913) );
  XNOR2_X1 U18361 ( .A(n14913), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15085) );
  NOR2_X1 U18362 ( .A1(n12853), .A2(n21102), .ZN(n15080) );
  AOI21_X1 U18363 ( .B1(n16099), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15080), .ZN(n14914) );
  OAI21_X1 U18364 ( .B1(n14915), .B2(n16110), .A(n14914), .ZN(n14916) );
  AOI21_X1 U18365 ( .B1(n14917), .B2(n16105), .A(n14916), .ZN(n14918) );
  OAI21_X1 U18366 ( .B1(n20095), .B2(n15085), .A(n14918), .ZN(P1_U2972) );
  AOI21_X1 U18367 ( .B1(n14948), .B2(n15090), .A(n10354), .ZN(n14919) );
  NOR2_X1 U18368 ( .A1(n14920), .A2(n14919), .ZN(n14921) );
  XNOR2_X1 U18369 ( .A(n14921), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15094) );
  INV_X1 U18370 ( .A(n14922), .ZN(n14926) );
  INV_X1 U18371 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21139) );
  OR2_X1 U18372 ( .A1(n12853), .A2(n21139), .ZN(n15087) );
  NAND2_X1 U18373 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14923) );
  OAI211_X1 U18374 ( .C1(n16110), .C2(n14924), .A(n15087), .B(n14923), .ZN(
        n14925) );
  AOI21_X1 U18375 ( .B1(n14926), .B2(n16105), .A(n14925), .ZN(n14927) );
  OAI21_X1 U18376 ( .B1(n20095), .B2(n15094), .A(n14927), .ZN(P1_U2973) );
  NOR2_X1 U18377 ( .A1(n12853), .A2(n14928), .ZN(n15097) );
  NOR2_X1 U18378 ( .A1(n16116), .A2(n14929), .ZN(n14930) );
  AOI211_X1 U18379 ( .C1(n16084), .C2(n14931), .A(n15097), .B(n14930), .ZN(
        n14937) );
  NOR2_X1 U18380 ( .A1(n14932), .A2(n15118), .ZN(n14939) );
  MUX2_X1 U18381 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14933), .S(
        n10354), .Z(n14934) );
  OAI21_X1 U18382 ( .B1(n14939), .B2(n15116), .A(n14934), .ZN(n14935) );
  XNOR2_X1 U18383 ( .A(n14935), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15095) );
  NAND2_X1 U18384 ( .A1(n15095), .A2(n16113), .ZN(n14936) );
  OAI211_X1 U18385 ( .C1(n14938), .C2(n16111), .A(n14937), .B(n14936), .ZN(
        P1_U2974) );
  AOI21_X1 U18386 ( .B1(n9844), .B2(n14948), .A(n14939), .ZN(n14941) );
  XNOR2_X1 U18387 ( .A(n16068), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14940) );
  XNOR2_X1 U18388 ( .A(n14941), .B(n14940), .ZN(n15108) );
  NAND2_X1 U18389 ( .A1(n15108), .A2(n16113), .ZN(n14945) );
  NOR2_X1 U18390 ( .A1(n12853), .A2(n21177), .ZN(n15112) );
  NOR2_X1 U18391 ( .A1(n16110), .A2(n14942), .ZN(n14943) );
  AOI211_X1 U18392 ( .C1(n16099), .C2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15112), .B(n14943), .ZN(n14944) );
  OAI211_X1 U18393 ( .C1(n14946), .C2(n16111), .A(n14945), .B(n14944), .ZN(
        P1_U2975) );
  XNOR2_X1 U18394 ( .A(n16068), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14947) );
  XNOR2_X1 U18395 ( .A(n14948), .B(n14947), .ZN(n15126) );
  NAND2_X1 U18396 ( .A1(n14949), .A2(n16105), .ZN(n14954) );
  OR2_X1 U18397 ( .A1(n12853), .A2(n21148), .ZN(n15120) );
  OAI21_X1 U18398 ( .B1(n16116), .B2(n14950), .A(n15120), .ZN(n14951) );
  AOI21_X1 U18399 ( .B1(n16084), .B2(n14952), .A(n14951), .ZN(n14953) );
  OAI211_X1 U18400 ( .C1(n15126), .C2(n20095), .A(n14954), .B(n14953), .ZN(
        P1_U2976) );
  NOR2_X1 U18401 ( .A1(n14955), .A2(n14069), .ZN(n14956) );
  XNOR2_X1 U18402 ( .A(n14956), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15142) );
  INV_X1 U18403 ( .A(n14957), .ZN(n14961) );
  OR2_X1 U18404 ( .A1(n12853), .A2(n21209), .ZN(n15137) );
  NAND2_X1 U18405 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14958) );
  OAI211_X1 U18406 ( .C1(n16110), .C2(n14959), .A(n15137), .B(n14958), .ZN(
        n14960) );
  AOI21_X1 U18407 ( .B1(n14961), .B2(n16105), .A(n14960), .ZN(n14962) );
  OAI21_X1 U18408 ( .B1(n20095), .B2(n15142), .A(n14962), .ZN(P1_U2977) );
  NAND3_X1 U18409 ( .A1(n14995), .A2(n10354), .A3(n14963), .ZN(n14972) );
  NAND3_X1 U18410 ( .A1(n14993), .A2(n15132), .A3(n16090), .ZN(n14964) );
  OAI21_X1 U18411 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14972), .A(
        n14964), .ZN(n14965) );
  XNOR2_X1 U18412 ( .A(n14965), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15963) );
  NAND2_X1 U18413 ( .A1(n14966), .A2(n16105), .ZN(n14971) );
  INV_X1 U18414 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14967) );
  OAI22_X1 U18415 ( .A1(n16116), .A2(n14967), .B1(n12853), .B2(n21288), .ZN(
        n14968) );
  AOI21_X1 U18416 ( .B1(n16084), .B2(n14969), .A(n14968), .ZN(n14970) );
  OAI211_X1 U18417 ( .C1(n15963), .C2(n20095), .A(n14971), .B(n14970), .ZN(
        P1_U2978) );
  NAND3_X1 U18418 ( .A1(n14993), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16090), .ZN(n14973) );
  NAND2_X1 U18419 ( .A1(n14973), .A2(n14972), .ZN(n14974) );
  XNOR2_X1 U18420 ( .A(n14974), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15151) );
  NAND2_X1 U18421 ( .A1(n16255), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15145) );
  OAI21_X1 U18422 ( .B1(n16116), .B2(n14975), .A(n15145), .ZN(n14978) );
  NOR2_X1 U18423 ( .A1(n14976), .A2(n16111), .ZN(n14977) );
  AOI211_X1 U18424 ( .C1(n16084), .C2(n14979), .A(n14978), .B(n14977), .ZN(
        n14980) );
  OAI21_X1 U18425 ( .B1(n15151), .B2(n20095), .A(n14980), .ZN(P1_U2979) );
  NOR2_X1 U18426 ( .A1(n16068), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14981) );
  MUX2_X1 U18427 ( .A(n14981), .B(n16090), .S(n14993), .Z(n14982) );
  XNOR2_X1 U18428 ( .A(n14982), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16117) );
  INV_X1 U18429 ( .A(n14983), .ZN(n14987) );
  AOI22_X1 U18430 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n16255), .ZN(n14984) );
  OAI21_X1 U18431 ( .B1(n14985), .B2(n16110), .A(n14984), .ZN(n14986) );
  AOI21_X1 U18432 ( .B1(n14987), .B2(n16105), .A(n14986), .ZN(n14988) );
  OAI21_X1 U18433 ( .B1(n20095), .B2(n16117), .A(n14988), .ZN(P1_U2980) );
  INV_X1 U18434 ( .A(n14989), .ZN(n14992) );
  OAI22_X1 U18435 ( .A1(n16116), .A2(n14990), .B1(n21237), .B2(n12853), .ZN(
        n14991) );
  AOI21_X1 U18436 ( .B1(n16084), .B2(n14992), .A(n14991), .ZN(n14997) );
  INV_X1 U18437 ( .A(n14993), .ZN(n16128) );
  NAND2_X1 U18438 ( .A1(n14995), .A2(n14994), .ZN(n16127) );
  NAND3_X1 U18439 ( .A1(n16128), .A2(n16113), .A3(n16127), .ZN(n14996) );
  OAI211_X1 U18440 ( .C1(n14998), .C2(n16111), .A(n14997), .B(n14996), .ZN(
        P1_U2981) );
  NAND2_X1 U18441 ( .A1(n16089), .A2(n9849), .ZN(n16065) );
  OAI21_X1 U18442 ( .B1(n16065), .B2(n15001), .A(n15000), .ZN(n15002) );
  MUX2_X1 U18443 ( .A(n16090), .B(n15003), .S(n15002), .Z(n15004) );
  XOR2_X1 U18444 ( .A(n15005), .B(n15004), .Z(n16153) );
  AOI22_X1 U18445 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n16255), .ZN(n15006) );
  OAI21_X1 U18446 ( .B1(n15007), .B2(n16110), .A(n15006), .ZN(n15008) );
  AOI21_X1 U18447 ( .B1(n15009), .B2(n16105), .A(n15008), .ZN(n15010) );
  OAI21_X1 U18448 ( .B1(n16153), .B2(n20095), .A(n15010), .ZN(P1_U2982) );
  INV_X1 U18449 ( .A(n15011), .ZN(n16076) );
  NAND3_X1 U18450 ( .A1(n16065), .A2(n16076), .A3(n16077), .ZN(n15013) );
  XNOR2_X1 U18451 ( .A(n15013), .B(n15012), .ZN(n16192) );
  INV_X1 U18452 ( .A(n15014), .ZN(n16028) );
  AOI22_X1 U18453 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n16255), .ZN(n15015) );
  OAI21_X1 U18454 ( .B1(n15016), .B2(n16110), .A(n15015), .ZN(n15017) );
  AOI21_X1 U18455 ( .B1(n16028), .B2(n16105), .A(n15017), .ZN(n15018) );
  OAI21_X1 U18456 ( .B1(n20095), .B2(n16192), .A(n15018), .ZN(P1_U2986) );
  MUX2_X1 U18457 ( .A(n16088), .B(n16089), .S(n16090), .Z(n15019) );
  XOR2_X1 U18458 ( .A(n13880), .B(n15019), .Z(n16233) );
  INV_X1 U18459 ( .A(n16233), .ZN(n15023) );
  AOI22_X1 U18460 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n16255), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n15020) );
  OAI21_X1 U18461 ( .B1(n16033), .B2(n16110), .A(n15020), .ZN(n15021) );
  AOI21_X1 U18462 ( .B1(n16036), .B2(n16105), .A(n15021), .ZN(n15022) );
  OAI21_X1 U18463 ( .B1(n15023), .B2(n20095), .A(n15022), .ZN(P1_U2989) );
  INV_X1 U18464 ( .A(n15024), .ZN(n15034) );
  NAND4_X1 U18465 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n16229), .ZN(n16182) );
  NOR2_X1 U18466 ( .A1(n16222), .A2(n16182), .ZN(n16212) );
  NAND2_X1 U18467 ( .A1(n16226), .A2(n16212), .ZN(n16204) );
  NOR2_X1 U18468 ( .A1(n16210), .A2(n16204), .ZN(n16131) );
  NAND2_X1 U18469 ( .A1(n16205), .A2(n16131), .ZN(n15129) );
  NOR3_X1 U18470 ( .A1(n15026), .A2(n15025), .A3(n16182), .ZN(n16200) );
  NAND3_X1 U18471 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n16200), .ZN(n16198) );
  NOR2_X1 U18472 ( .A1(n16141), .A2(n16198), .ZN(n16132) );
  INV_X1 U18473 ( .A(n16132), .ZN(n15027) );
  OAI21_X1 U18474 ( .B1(n15129), .B2(n16141), .A(n15105), .ZN(n16162) );
  NAND4_X1 U18475 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16151) );
  NOR2_X1 U18476 ( .A1(n16145), .A2(n16151), .ZN(n15036) );
  AND4_X1 U18477 ( .A1(n15132), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n15036), .ZN(n15028) );
  NAND2_X1 U18478 ( .A1(n16162), .A2(n15028), .ZN(n15110) );
  OR2_X1 U18479 ( .A1(n15078), .A2(n15030), .ZN(n15050) );
  INV_X1 U18480 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15031) );
  NOR3_X1 U18481 ( .A1(n15050), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15031), .ZN(n15033) );
  AOI211_X1 U18482 ( .C1(n15034), .C2(n16263), .A(n15033), .B(n15032), .ZN(
        n15047) );
  INV_X1 U18483 ( .A(n15035), .ZN(n15068) );
  INV_X1 U18484 ( .A(n16198), .ZN(n15128) );
  AND2_X1 U18485 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15036), .ZN(
        n15130) );
  NAND2_X1 U18486 ( .A1(n15128), .A2(n15130), .ZN(n15131) );
  AOI21_X1 U18487 ( .B1(n15130), .B2(n16131), .A(n16130), .ZN(n15037) );
  AOI211_X1 U18488 ( .C1(n15038), .C2(n15131), .A(n15037), .B(n16202), .ZN(
        n16120) );
  NOR2_X1 U18489 ( .A1(n16161), .A2(n16202), .ZN(n16224) );
  AOI21_X1 U18490 ( .B1(n16120), .B2(n15132), .A(n16224), .ZN(n15962) );
  NAND2_X1 U18491 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15135) );
  AND2_X1 U18492 ( .A1(n16161), .A2(n15135), .ZN(n15039) );
  OR2_X1 U18493 ( .A1(n15962), .A2(n15039), .ZN(n15124) );
  NOR2_X1 U18494 ( .A1(n15124), .A2(n16161), .ZN(n15043) );
  INV_X1 U18495 ( .A(n15043), .ZN(n15045) );
  NOR2_X1 U18496 ( .A1(n16130), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15040) );
  OR2_X1 U18497 ( .A1(n15124), .A2(n15040), .ZN(n15106) );
  AND2_X1 U18498 ( .A1(n16161), .A2(n15041), .ZN(n15042) );
  NOR2_X1 U18499 ( .A1(n15106), .A2(n15042), .ZN(n15100) );
  AOI21_X1 U18500 ( .B1(n15100), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15043), .ZN(n15082) );
  AOI21_X1 U18501 ( .B1(n15068), .B2(n15045), .A(n15082), .ZN(n15063) );
  OAI211_X1 U18502 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15044), .A(
        n15063), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15051) );
  NAND3_X1 U18503 ( .A1(n15051), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15045), .ZN(n15046) );
  OAI211_X1 U18504 ( .C1(n15048), .C2(n16215), .A(n15047), .B(n15046), .ZN(
        P1_U3000) );
  NAND2_X1 U18505 ( .A1(n15049), .A2(n16268), .ZN(n15057) );
  INV_X1 U18506 ( .A(n15050), .ZN(n15052) );
  OAI21_X1 U18507 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15052), .A(
        n15051), .ZN(n15055) );
  NAND2_X1 U18508 ( .A1(n15053), .A2(n16263), .ZN(n15054) );
  NAND4_X1 U18509 ( .A1(n15057), .A2(n15056), .A3(n15055), .A4(n15054), .ZN(
        P1_U3001) );
  INV_X1 U18510 ( .A(n15058), .ZN(n15060) );
  NOR3_X1 U18511 ( .A1(n15078), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15068), .ZN(n15059) );
  AOI211_X1 U18512 ( .C1(n15061), .C2(n16263), .A(n15060), .B(n15059), .ZN(
        n15065) );
  OR2_X1 U18513 ( .A1(n15063), .A2(n15062), .ZN(n15064) );
  OAI211_X1 U18514 ( .C1(n15066), .C2(n16215), .A(n15065), .B(n15064), .ZN(
        P1_U3002) );
  INV_X1 U18515 ( .A(n15067), .ZN(n15076) );
  NAND2_X1 U18516 ( .A1(n9937), .A2(n15068), .ZN(n15071) );
  INV_X1 U18517 ( .A(n15069), .ZN(n15070) );
  OAI21_X1 U18518 ( .B1(n15078), .B2(n15071), .A(n15070), .ZN(n15072) );
  AOI21_X1 U18519 ( .B1(n15073), .B2(n16263), .A(n15072), .ZN(n15075) );
  NAND2_X1 U18520 ( .A1(n15082), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15074) );
  OAI211_X1 U18521 ( .C1(n15076), .C2(n16215), .A(n15075), .B(n15074), .ZN(
        P1_U3003) );
  INV_X1 U18522 ( .A(n15077), .ZN(n15081) );
  NOR2_X1 U18523 ( .A1(n15078), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15079) );
  AOI211_X1 U18524 ( .C1(n15081), .C2(n16263), .A(n15080), .B(n15079), .ZN(
        n15084) );
  NAND2_X1 U18525 ( .A1(n15082), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15083) );
  OAI211_X1 U18526 ( .C1(n15085), .C2(n16215), .A(n15084), .B(n15083), .ZN(
        P1_U3004) );
  INV_X1 U18527 ( .A(n15086), .ZN(n15089) );
  INV_X1 U18528 ( .A(n15087), .ZN(n15088) );
  AOI21_X1 U18529 ( .B1(n15089), .B2(n16263), .A(n15088), .ZN(n15093) );
  INV_X1 U18530 ( .A(n15110), .ZN(n15119) );
  NAND2_X1 U18531 ( .A1(n15119), .A2(n15090), .ZN(n15091) );
  MUX2_X1 U18532 ( .A(n15091), .B(n15100), .S(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n15092) );
  OAI211_X1 U18533 ( .C1(n15094), .C2(n16215), .A(n15093), .B(n15092), .ZN(
        P1_U3005) );
  INV_X1 U18534 ( .A(n15095), .ZN(n15104) );
  INV_X1 U18535 ( .A(n15096), .ZN(n15098) );
  AOI21_X1 U18536 ( .B1(n15098), .B2(n16263), .A(n15097), .ZN(n15103) );
  NAND2_X1 U18537 ( .A1(n15119), .A2(n15099), .ZN(n15101) );
  MUX2_X1 U18538 ( .A(n15101), .B(n15100), .S(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n15102) );
  OAI211_X1 U18539 ( .C1(n15104), .C2(n16215), .A(n15103), .B(n15102), .ZN(
        P1_U3006) );
  INV_X1 U18540 ( .A(n15105), .ZN(n15107) );
  AOI21_X1 U18541 ( .B1(n15107), .B2(n15118), .A(n15106), .ZN(n15117) );
  NAND2_X1 U18542 ( .A1(n15108), .A2(n16268), .ZN(n15115) );
  INV_X1 U18543 ( .A(n15109), .ZN(n15113) );
  NOR3_X1 U18544 ( .A1(n15110), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15118), .ZN(n15111) );
  AOI211_X1 U18545 ( .C1(n15113), .C2(n16263), .A(n15112), .B(n15111), .ZN(
        n15114) );
  OAI211_X1 U18546 ( .C1(n15117), .C2(n15116), .A(n15115), .B(n15114), .ZN(
        P1_U3007) );
  NAND2_X1 U18547 ( .A1(n15119), .A2(n15118), .ZN(n15121) );
  OAI211_X1 U18548 ( .C1(n15122), .C2(n16242), .A(n15121), .B(n15120), .ZN(
        n15123) );
  AOI21_X1 U18549 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15124), .A(
        n15123), .ZN(n15125) );
  OAI21_X1 U18550 ( .B1(n15126), .B2(n16215), .A(n15125), .ZN(P1_U3008) );
  INV_X1 U18551 ( .A(n15127), .ZN(n15139) );
  NAND2_X1 U18552 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15128), .ZN(
        n16134) );
  OAI21_X1 U18553 ( .B1(n16134), .B2(n16136), .A(n15129), .ZN(n16140) );
  NAND2_X1 U18554 ( .A1(n15130), .A2(n16140), .ZN(n15143) );
  OAI21_X1 U18555 ( .B1(n16133), .B2(n15131), .A(n15143), .ZN(n16124) );
  NAND2_X1 U18556 ( .A1(n15132), .A2(n16124), .ZN(n15969) );
  AOI21_X1 U18557 ( .B1(n15134), .B2(n15133), .A(n15969), .ZN(n15136) );
  NAND2_X1 U18558 ( .A1(n15136), .A2(n15135), .ZN(n15138) );
  OAI211_X1 U18559 ( .C1(n15139), .C2(n16242), .A(n15138), .B(n15137), .ZN(
        n15140) );
  AOI21_X1 U18560 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15962), .A(
        n15140), .ZN(n15141) );
  OAI21_X1 U18561 ( .B1(n15142), .B2(n16215), .A(n15141), .ZN(P1_U3009) );
  OAI221_X1 U18562 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16133), 
        .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15143), .A(n16120), .ZN(
        n15149) );
  NOR2_X1 U18563 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16123), .ZN(
        n15144) );
  NAND2_X1 U18564 ( .A1(n16124), .A2(n15144), .ZN(n15146) );
  OAI211_X1 U18565 ( .C1(n16242), .C2(n15147), .A(n15146), .B(n15145), .ZN(
        n15148) );
  AOI21_X1 U18566 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n15149), .A(
        n15148), .ZN(n15150) );
  OAI21_X1 U18567 ( .B1(n15151), .B2(n16215), .A(n15150), .ZN(P1_U3011) );
  NAND2_X1 U18568 ( .A1(n15152), .A2(n16268), .ZN(n15159) );
  AOI22_X1 U18569 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15154), .B1(
        n15153), .B2(n13259), .ZN(n15158) );
  NAND2_X1 U18570 ( .A1(n16263), .A2(n20180), .ZN(n15157) );
  INV_X1 U18571 ( .A(n15155), .ZN(n15156) );
  NAND4_X1 U18572 ( .A1(n15159), .A2(n15158), .A3(n15157), .A4(n15156), .ZN(
        P1_U3028) );
  OR2_X1 U18573 ( .A1(n20702), .A2(n15160), .ZN(n15168) );
  NAND2_X1 U18574 ( .A1(n15162), .A2(n15161), .ZN(n15163) );
  NOR2_X1 U18575 ( .A1(n15164), .A2(n15163), .ZN(n15165) );
  AOI21_X1 U18576 ( .B1(n15925), .B2(n15166), .A(n15165), .ZN(n15167) );
  NAND2_X1 U18577 ( .A1(n15168), .A2(n15167), .ZN(n15929) );
  INV_X1 U18578 ( .A(n15929), .ZN(n15176) );
  INV_X1 U18579 ( .A(n15169), .ZN(n20871) );
  NOR2_X1 U18580 ( .A1(n16272), .A2(n15170), .ZN(n20868) );
  INV_X1 U18581 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15171) );
  OAI22_X1 U18582 ( .A1(n15171), .A2(n12760), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20872) );
  NOR3_X1 U18583 ( .A1(n15173), .A2(n15172), .A3(n20875), .ZN(n15174) );
  AOI21_X1 U18584 ( .B1(n20868), .B2(n20872), .A(n15174), .ZN(n15175) );
  OAI21_X1 U18585 ( .B1(n15176), .B2(n20871), .A(n15175), .ZN(n15177) );
  MUX2_X1 U18586 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15177), .S(
        n20878), .Z(P1_U3473) );
  AOI21_X1 U18587 ( .B1(n15538), .B2(n15190), .A(n15514), .ZN(n15914) );
  AOI21_X1 U18588 ( .B1(n15188), .B2(n15563), .A(n15191), .ZN(n19142) );
  AOI21_X1 U18589 ( .B1(n11202), .B2(n15187), .A(n15189), .ZN(n19165) );
  AOI21_X1 U18590 ( .B1(n16415), .B2(n15185), .A(n9913), .ZN(n16406) );
  AOI21_X1 U18591 ( .B1(n19197), .B2(n15183), .A(n15186), .ZN(n19206) );
  AOI21_X1 U18592 ( .B1(n16448), .B2(n15182), .A(n15184), .ZN(n16433) );
  AOI21_X1 U18593 ( .B1(n16465), .B2(n15180), .A(n9888), .ZN(n16455) );
  AOI21_X1 U18594 ( .B1(n16473), .B2(n15178), .A(n15181), .ZN(n19251) );
  NAND2_X1 U18595 ( .A1(n15179), .A2(n16474), .ZN(n19250) );
  NOR2_X1 U18596 ( .A1(n19251), .A2(n19250), .ZN(n19239) );
  OAI21_X1 U18597 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n15181), .A(
        n15180), .ZN(n19240) );
  NAND2_X1 U18598 ( .A1(n19239), .A2(n19240), .ZN(n15234) );
  NOR2_X1 U18599 ( .A1(n16455), .A2(n15234), .ZN(n19229) );
  OAI21_X1 U18600 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n9888), .A(
        n15182), .ZN(n19230) );
  NAND2_X1 U18601 ( .A1(n19229), .A2(n19230), .ZN(n15219) );
  NOR2_X1 U18602 ( .A1(n16433), .A2(n15219), .ZN(n19217) );
  OAI21_X1 U18603 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n15184), .A(
        n15183), .ZN(n19218) );
  NAND2_X1 U18604 ( .A1(n19217), .A2(n19218), .ZN(n19207) );
  NOR2_X1 U18605 ( .A1(n19206), .A2(n19207), .ZN(n19191) );
  OAI21_X1 U18606 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n15186), .A(
        n15185), .ZN(n19192) );
  NAND2_X1 U18607 ( .A1(n19191), .A2(n19192), .ZN(n15214) );
  NOR2_X1 U18608 ( .A1(n16406), .A2(n15214), .ZN(n15213) );
  OAI21_X1 U18609 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n9913), .A(
        n15187), .ZN(n19180) );
  NAND2_X1 U18610 ( .A1(n15213), .A2(n19180), .ZN(n19164) );
  NOR2_X1 U18611 ( .A1(n19165), .A2(n19164), .ZN(n19163) );
  OAI21_X1 U18612 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n15189), .A(
        n15188), .ZN(n19155) );
  NAND2_X1 U18613 ( .A1(n19163), .A2(n19155), .ZN(n19140) );
  NOR2_X1 U18614 ( .A1(n19142), .A2(n19140), .ZN(n19129) );
  OAI21_X1 U18615 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n15191), .A(
        n15190), .ZN(n19133) );
  NAND2_X1 U18616 ( .A1(n19129), .A2(n19133), .ZN(n15913) );
  AOI21_X1 U18617 ( .B1(n9797), .B2(n15913), .A(n19301), .ZN(n15204) );
  NAND2_X1 U18618 ( .A1(n15349), .A2(n15192), .ZN(n15193) );
  NAND2_X1 U18619 ( .A1(n9887), .A2(n15193), .ZN(n15654) );
  NAND2_X1 U18620 ( .A1(n15194), .A2(n19288), .ZN(n15199) );
  AND2_X1 U18621 ( .A1(n15430), .A2(n15195), .ZN(n15196) );
  NOR2_X1 U18622 ( .A1(n15410), .A2(n15196), .ZN(n15659) );
  INV_X1 U18623 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19998) );
  OAI22_X1 U18624 ( .A1(n15538), .A2(n19264), .B1(n19998), .B2(n19256), .ZN(
        n15197) );
  AOI21_X1 U18625 ( .B1(n19203), .B2(n15659), .A(n15197), .ZN(n15198) );
  OAI211_X1 U18626 ( .C1(n19295), .C2(n15654), .A(n15199), .B(n15198), .ZN(
        n15203) );
  NAND2_X1 U18627 ( .A1(n19245), .A2(n9797), .ZN(n19162) );
  INV_X1 U18628 ( .A(n15913), .ZN(n15200) );
  NOR2_X1 U18629 ( .A1(n19162), .A2(n15200), .ZN(n19128) );
  INV_X1 U18630 ( .A(n19128), .ZN(n15201) );
  OAI22_X1 U18631 ( .A1(n15914), .A2(n15201), .B1(n19271), .B2(n9971), .ZN(
        n15202) );
  AOI211_X1 U18632 ( .C1(n15914), .C2(n15204), .A(n15203), .B(n15202), .ZN(
        n15205) );
  INV_X1 U18633 ( .A(n15205), .ZN(P2_U2834) );
  AOI22_X1 U18634 ( .A1(n16408), .A2(n19243), .B1(n19293), .B2(
        P2_EBX_REG_15__SCAN_IN), .ZN(n15212) );
  AOI21_X1 U18635 ( .B1(n15206), .B2(n15753), .A(n13753), .ZN(n19307) );
  INV_X1 U18636 ( .A(n19307), .ZN(n15208) );
  AOI22_X1 U18637 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n19286), .ZN(n15207) );
  OAI211_X1 U18638 ( .C1(n19290), .C2(n15208), .A(n15207), .B(n19254), .ZN(
        n15209) );
  INV_X1 U18639 ( .A(n15209), .ZN(n15211) );
  NAND2_X1 U18640 ( .A1(n16406), .A2(n19199), .ZN(n15210) );
  NAND3_X1 U18641 ( .A1(n15212), .A2(n15211), .A3(n15210), .ZN(n15216) );
  OR2_X1 U18642 ( .A1(n19277), .A2(n15213), .ZN(n19181) );
  AOI211_X1 U18643 ( .C1(n16406), .C2(n15214), .A(n19301), .B(n19181), .ZN(
        n15215) );
  AOI211_X1 U18644 ( .C1(n19288), .C2(n15217), .A(n15216), .B(n15215), .ZN(
        n15218) );
  INV_X1 U18645 ( .A(n15218), .ZN(P2_U2840) );
  NAND2_X1 U18646 ( .A1(n9797), .A2(n15219), .ZN(n15220) );
  XNOR2_X1 U18647 ( .A(n16433), .B(n15220), .ZN(n15221) );
  NAND2_X1 U18648 ( .A1(n15221), .A2(n19245), .ZN(n15232) );
  NAND2_X1 U18649 ( .A1(n15223), .A2(n15222), .ZN(n15226) );
  INV_X1 U18650 ( .A(n15224), .ZN(n15225) );
  NAND2_X1 U18651 ( .A1(n15226), .A2(n15225), .ZN(n16536) );
  OR2_X1 U18652 ( .A1(n19290), .A2(n16536), .ZN(n15229) );
  AOI22_X1 U18653 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n19293), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19298), .ZN(n15228) );
  NAND2_X1 U18654 ( .A1(n19286), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n15227) );
  NAND4_X1 U18655 ( .A1(n15229), .A2(n15228), .A3(n19254), .A4(n15227), .ZN(
        n15230) );
  AOI21_X1 U18656 ( .B1(n16539), .B2(n19243), .A(n15230), .ZN(n15231) );
  OAI211_X1 U18657 ( .C1(n19266), .C2(n15233), .A(n15232), .B(n15231), .ZN(
        P2_U2844) );
  NAND2_X1 U18658 ( .A1(n9797), .A2(n15234), .ZN(n15235) );
  XNOR2_X1 U18659 ( .A(n16455), .B(n15235), .ZN(n15242) );
  AOI22_X1 U18660 ( .A1(n15236), .A2(n19288), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19293), .ZN(n15237) );
  OAI21_X1 U18661 ( .B1(n16465), .B2(n19264), .A(n15237), .ZN(n15241) );
  AOI21_X1 U18662 ( .B1(n19286), .B2(P2_REIP_REG_9__SCAN_IN), .A(n19404), .ZN(
        n15239) );
  NAND2_X1 U18663 ( .A1(n19203), .A2(n15806), .ZN(n15238) );
  OAI211_X1 U18664 ( .C1(n15809), .C2(n19295), .A(n15239), .B(n15238), .ZN(
        n15240) );
  AOI211_X1 U18665 ( .C1(n15242), .C2(n19245), .A(n15241), .B(n15240), .ZN(
        n15243) );
  INV_X1 U18666 ( .A(n15243), .ZN(P2_U2846) );
  INV_X1 U18667 ( .A(n19297), .ZN(n19273) );
  NAND2_X1 U18668 ( .A1(n9797), .A2(n15244), .ZN(n15245) );
  XNOR2_X1 U18669 ( .A(n15246), .B(n15245), .ZN(n15247) );
  NAND2_X1 U18670 ( .A1(n15247), .A2(n19245), .ZN(n15255) );
  AOI22_X1 U18671 ( .A1(n20046), .A2(n19203), .B1(n19293), .B2(
        P2_EBX_REG_3__SCAN_IN), .ZN(n15248) );
  OAI21_X1 U18672 ( .B1(n15249), .B2(n19266), .A(n15248), .ZN(n15252) );
  INV_X1 U18673 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19963) );
  OAI22_X1 U18674 ( .A1(n15250), .A2(n19264), .B1(n19963), .B2(n19256), .ZN(
        n15251) );
  AOI211_X1 U18675 ( .C1(n19243), .C2(n15253), .A(n15252), .B(n15251), .ZN(
        n15254) );
  OAI211_X1 U18676 ( .C1(n19273), .C2(n20039), .A(n15255), .B(n15254), .ZN(
        P2_U2852) );
  AOI22_X1 U18677 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19286), .ZN(n15256) );
  OAI21_X1 U18678 ( .B1(n19266), .B2(n15257), .A(n15256), .ZN(n15259) );
  NOR2_X1 U18679 ( .A1(n19271), .A2(n10619), .ZN(n15258) );
  AOI211_X1 U18680 ( .C1(n19203), .C2(n20050), .A(n15259), .B(n15258), .ZN(
        n15260) );
  OAI21_X1 U18681 ( .B1(n15261), .B2(n19295), .A(n15260), .ZN(n15267) );
  INV_X1 U18682 ( .A(n15263), .ZN(n15265) );
  INV_X1 U18683 ( .A(n15264), .ZN(n15262) );
  AOI221_X1 U18684 ( .B1(n15265), .B2(n15264), .C1(n15263), .C2(n15262), .A(
        n19301), .ZN(n15266) );
  AOI211_X1 U18685 ( .C1(n20051), .C2(n19297), .A(n15267), .B(n15266), .ZN(
        n15268) );
  INV_X1 U18686 ( .A(n15268), .ZN(P2_U2853) );
  NAND2_X1 U18687 ( .A1(n19425), .A2(n19243), .ZN(n15277) );
  NAND2_X1 U18688 ( .A1(n15270), .A2(n15269), .ZN(n15271) );
  NAND2_X1 U18689 ( .A1(n15272), .A2(n15271), .ZN(n20062) );
  AOI22_X1 U18690 ( .A1(n19286), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19298), .ZN(n15273) );
  OAI21_X1 U18691 ( .B1(n19266), .B2(n15274), .A(n15273), .ZN(n15275) );
  AOI21_X1 U18692 ( .B1(n19203), .B2(n20062), .A(n15275), .ZN(n15276) );
  OAI211_X1 U18693 ( .C1(n19271), .C2(n15278), .A(n15277), .B(n15276), .ZN(
        n15281) );
  INV_X1 U18694 ( .A(n19199), .ZN(n19175) );
  OAI22_X1 U18695 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19175), .B1(
        n15279), .B2(n19301), .ZN(n15280) );
  AOI211_X1 U18696 ( .C1(n19297), .C2(n20060), .A(n15281), .B(n15280), .ZN(
        n15282) );
  INV_X1 U18697 ( .A(n15282), .ZN(P2_U2854) );
  MUX2_X1 U18698 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16291), .S(n15356), .Z(
        P2_U2856) );
  NAND2_X1 U18699 ( .A1(n15352), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15286) );
  NAND2_X1 U18700 ( .A1(n15288), .A2(n15287), .ZN(n15289) );
  XOR2_X1 U18701 ( .A(n15290), .B(n15289), .Z(n15367) );
  NAND2_X1 U18702 ( .A1(n15367), .A2(n15346), .ZN(n15292) );
  NAND2_X1 U18703 ( .A1(n15352), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15291) );
  OAI211_X1 U18704 ( .C1(n15323), .C2(n15468), .A(n15292), .B(n15291), .ZN(
        P2_U2859) );
  OAI21_X1 U18705 ( .B1(n15293), .B2(n15295), .A(n15294), .ZN(n15381) );
  NOR2_X1 U18706 ( .A1(n15306), .A2(n15296), .ZN(n15297) );
  NOR2_X1 U18707 ( .A1(n16329), .A2(n15352), .ZN(n15298) );
  AOI21_X1 U18708 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n15323), .A(n15298), .ZN(
        n15299) );
  OAI21_X1 U18709 ( .B1(n15381), .B2(n15359), .A(n15299), .ZN(P2_U2860) );
  OAI21_X1 U18710 ( .B1(n15301), .B2(n15303), .A(n15302), .ZN(n15390) );
  NAND2_X1 U18711 ( .A1(n15352), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15308) );
  AND2_X1 U18712 ( .A1(n9892), .A2(n15304), .ZN(n15305) );
  NOR2_X1 U18713 ( .A1(n15306), .A2(n15305), .ZN(n16506) );
  NAND2_X1 U18714 ( .A1(n16506), .A2(n15356), .ZN(n15307) );
  OAI211_X1 U18715 ( .C1(n15390), .C2(n15359), .A(n15308), .B(n15307), .ZN(
        P2_U2861) );
  OAI21_X1 U18716 ( .B1(n15309), .B2(n15311), .A(n15310), .ZN(n15398) );
  NAND2_X1 U18717 ( .A1(n9815), .A2(n15312), .ZN(n15313) );
  NAND2_X1 U18718 ( .A1(n9892), .A2(n15313), .ZN(n16348) );
  NOR2_X1 U18719 ( .A1(n16348), .A2(n15323), .ZN(n15314) );
  AOI21_X1 U18720 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n15323), .A(n15314), .ZN(
        n15315) );
  OAI21_X1 U18721 ( .B1(n15398), .B2(n15359), .A(n15315), .ZN(P2_U2862) );
  AOI21_X1 U18722 ( .B1(n15316), .B2(n15318), .A(n15317), .ZN(n15319) );
  XOR2_X1 U18723 ( .A(n15320), .B(n15319), .Z(n15408) );
  NAND2_X1 U18724 ( .A1(n9821), .A2(n15321), .ZN(n15322) );
  NAND2_X1 U18725 ( .A1(n9815), .A2(n15322), .ZN(n15629) );
  MUX2_X1 U18726 ( .A(n15629), .B(n16357), .S(n15323), .Z(n15324) );
  OAI21_X1 U18727 ( .B1(n15408), .B2(n15359), .A(n15324), .ZN(P2_U2863) );
  OR2_X1 U18728 ( .A1(n15325), .A2(n15336), .ZN(n15326) );
  NAND2_X1 U18729 ( .A1(n9821), .A2(n15326), .ZN(n16372) );
  AOI21_X1 U18730 ( .B1(n15327), .B2(n15329), .A(n15328), .ZN(n16382) );
  NAND2_X1 U18731 ( .A1(n16382), .A2(n15346), .ZN(n15331) );
  NAND2_X1 U18732 ( .A1(n15352), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15330) );
  OAI211_X1 U18733 ( .C1(n16372), .C2(n15352), .A(n15331), .B(n15330), .ZN(
        P2_U2864) );
  INV_X1 U18734 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15341) );
  AOI21_X1 U18735 ( .B1(n15334), .B2(n15333), .A(n11897), .ZN(n15417) );
  NAND2_X1 U18736 ( .A1(n15417), .A2(n15346), .ZN(n15340) );
  NAND2_X1 U18737 ( .A1(n9887), .A2(n15335), .ZN(n15338) );
  INV_X1 U18738 ( .A(n15336), .ZN(n15337) );
  NAND2_X1 U18739 ( .A1(n15338), .A2(n15337), .ZN(n15638) );
  INV_X1 U18740 ( .A(n15638), .ZN(n15920) );
  NAND2_X1 U18741 ( .A1(n15920), .A2(n15356), .ZN(n15339) );
  OAI211_X1 U18742 ( .C1(n15356), .C2(n15341), .A(n15340), .B(n15339), .ZN(
        P2_U2865) );
  OAI21_X1 U18743 ( .B1(n15342), .B2(n15343), .A(n15333), .ZN(n15426) );
  MUX2_X1 U18744 ( .A(n15654), .B(n9971), .S(n15352), .Z(n15344) );
  OAI21_X1 U18745 ( .B1(n15426), .B2(n15359), .A(n15344), .ZN(P2_U2866) );
  AOI21_X1 U18746 ( .B1(n15345), .B2(n13891), .A(n15342), .ZN(n15435) );
  NAND2_X1 U18747 ( .A1(n15435), .A2(n15346), .ZN(n15351) );
  NAND2_X1 U18748 ( .A1(n15355), .A2(n15347), .ZN(n15348) );
  NAND2_X1 U18749 ( .A1(n15349), .A2(n15348), .ZN(n15556) );
  NAND2_X1 U18750 ( .A1(n19136), .A2(n15356), .ZN(n15350) );
  OAI211_X1 U18751 ( .C1(n15356), .C2(n9973), .A(n15351), .B(n15350), .ZN(
        P2_U2867) );
  NAND2_X1 U18752 ( .A1(n15352), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15358) );
  NAND2_X1 U18753 ( .A1(n13849), .A2(n15353), .ZN(n15354) );
  AND2_X1 U18754 ( .A1(n15355), .A2(n15354), .ZN(n19148) );
  NAND2_X1 U18755 ( .A1(n19148), .A2(n15356), .ZN(n15357) );
  OAI211_X1 U18756 ( .C1(n15360), .C2(n15359), .A(n15358), .B(n15357), .ZN(
        P2_U2868) );
  NAND3_X1 U18757 ( .A1(n15283), .A2(n15361), .A3(n19361), .ZN(n15366) );
  AOI22_X1 U18758 ( .A1(n16307), .A2(n19360), .B1(n19359), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15365) );
  AOI22_X1 U18759 ( .A1(n19302), .A2(BUF2_REG_29__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15364) );
  NAND2_X1 U18760 ( .A1(n16381), .A2(n15362), .ZN(n15363) );
  NAND4_X1 U18761 ( .A1(n15366), .A2(n15365), .A3(n15364), .A4(n15363), .ZN(
        P2_U2890) );
  INV_X1 U18762 ( .A(n15367), .ZN(n15373) );
  OAI22_X1 U18763 ( .A1(n15404), .A2(n15369), .B1(n19333), .B2(n15368), .ZN(
        n15370) );
  AOI21_X1 U18764 ( .B1(n19360), .B2(n16319), .A(n15370), .ZN(n15372) );
  AOI22_X1 U18765 ( .A1(n19302), .A2(BUF2_REG_28__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15371) );
  OAI211_X1 U18766 ( .C1(n15373), .C2(n15425), .A(n15372), .B(n15371), .ZN(
        P2_U2891) );
  NOR2_X1 U18767 ( .A1(n15384), .A2(n15374), .ZN(n15375) );
  OAI22_X1 U18768 ( .A1(n15404), .A2(n19316), .B1(n19333), .B2(n15377), .ZN(
        n15378) );
  AOI21_X1 U18769 ( .B1(n19360), .B2(n10431), .A(n15378), .ZN(n15380) );
  AOI22_X1 U18770 ( .A1(n19302), .A2(BUF2_REG_27__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15379) );
  OAI211_X1 U18771 ( .C1(n15381), .C2(n15425), .A(n15380), .B(n15379), .ZN(
        P2_U2892) );
  NOR2_X1 U18772 ( .A1(n15392), .A2(n15382), .ZN(n15383) );
  OR2_X1 U18773 ( .A1(n15384), .A2(n15383), .ZN(n16501) );
  OAI22_X1 U18774 ( .A1(n19334), .A2(n16501), .B1(n19333), .B2(n15385), .ZN(
        n15386) );
  AOI21_X1 U18775 ( .B1(n16381), .B2(n15387), .A(n15386), .ZN(n15389) );
  AOI22_X1 U18776 ( .A1(n19302), .A2(BUF2_REG_26__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15388) );
  OAI211_X1 U18777 ( .C1(n15390), .C2(n15425), .A(n15389), .B(n15388), .ZN(
        P2_U2893) );
  AND2_X1 U18778 ( .A1(n15401), .A2(n15391), .ZN(n15393) );
  OR2_X1 U18779 ( .A1(n15393), .A2(n15392), .ZN(n16349) );
  OAI22_X1 U18780 ( .A1(n19334), .A2(n16349), .B1(n19333), .B2(n12821), .ZN(
        n15394) );
  AOI21_X1 U18781 ( .B1(n16381), .B2(n15395), .A(n15394), .ZN(n15397) );
  AOI22_X1 U18782 ( .A1(n19302), .A2(BUF2_REG_25__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15396) );
  OAI211_X1 U18783 ( .C1(n15398), .C2(n15425), .A(n15397), .B(n15396), .ZN(
        P2_U2894) );
  NAND2_X1 U18784 ( .A1(n16370), .A2(n15399), .ZN(n15400) );
  AND2_X1 U18785 ( .A1(n15401), .A2(n15400), .ZN(n16361) );
  OAI22_X1 U18786 ( .A1(n15404), .A2(n15403), .B1(n19333), .B2(n15402), .ZN(
        n15405) );
  AOI21_X1 U18787 ( .B1(n19360), .B2(n16361), .A(n15405), .ZN(n15407) );
  AOI22_X1 U18788 ( .A1(n19302), .A2(BUF2_REG_24__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15406) );
  OAI211_X1 U18789 ( .C1(n15408), .C2(n15425), .A(n15407), .B(n15406), .ZN(
        P2_U2895) );
  OR2_X1 U18790 ( .A1(n15410), .A2(n15409), .ZN(n15412) );
  NAND2_X1 U18791 ( .A1(n15412), .A2(n15411), .ZN(n15924) );
  AOI22_X1 U18792 ( .A1(n19302), .A2(BUF2_REG_22__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15415) );
  AOI22_X1 U18793 ( .A1(n16381), .A2(n15413), .B1(n19359), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n15414) );
  OAI211_X1 U18794 ( .C1(n19334), .C2(n15924), .A(n15415), .B(n15414), .ZN(
        n15416) );
  AOI21_X1 U18795 ( .B1(n15417), .B2(n19361), .A(n15416), .ZN(n15418) );
  INV_X1 U18796 ( .A(n15418), .ZN(P2_U2897) );
  INV_X1 U18797 ( .A(n15659), .ZN(n15422) );
  AOI22_X1 U18798 ( .A1(n19302), .A2(BUF2_REG_21__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n15421) );
  AOI22_X1 U18799 ( .A1(n16381), .A2(n15419), .B1(n19359), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15420) );
  OAI211_X1 U18800 ( .C1(n19334), .C2(n15422), .A(n15421), .B(n15420), .ZN(
        n15423) );
  INV_X1 U18801 ( .A(n15423), .ZN(n15424) );
  OAI21_X1 U18802 ( .B1(n15426), .B2(n15425), .A(n15424), .ZN(P2_U2898) );
  NAND2_X1 U18803 ( .A1(n15428), .A2(n15427), .ZN(n15429) );
  NAND2_X1 U18804 ( .A1(n15430), .A2(n15429), .ZN(n19139) );
  AOI22_X1 U18805 ( .A1(n19302), .A2(BUF2_REG_20__SCAN_IN), .B1(n19304), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n15433) );
  AOI22_X1 U18806 ( .A1(n16381), .A2(n15431), .B1(n19359), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n15432) );
  OAI211_X1 U18807 ( .C1(n19334), .C2(n19139), .A(n15433), .B(n15432), .ZN(
        n15434) );
  AOI21_X1 U18808 ( .B1(n15435), .B2(n19361), .A(n15434), .ZN(n15436) );
  INV_X1 U18809 ( .A(n15436), .ZN(P2_U2899) );
  NAND2_X1 U18810 ( .A1(n16477), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15437) );
  OAI211_X1 U18811 ( .C1(n16475), .C2(n15439), .A(n15438), .B(n15437), .ZN(
        n15442) );
  NOR2_X1 U18812 ( .A1(n15440), .A2(n16478), .ZN(n15441) );
  OAI21_X1 U18813 ( .B1(n15444), .B2(n16480), .A(n15443), .ZN(P2_U2983) );
  NOR2_X1 U18814 ( .A1(n15446), .A2(n9856), .ZN(n15447) );
  XNOR2_X1 U18815 ( .A(n15448), .B(n15447), .ZN(n15611) );
  INV_X1 U18816 ( .A(n15449), .ZN(n15450) );
  NOR2_X1 U18817 ( .A1(n15452), .A2(n15451), .ZN(n15610) );
  INV_X1 U18818 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20018) );
  NOR2_X1 U18819 ( .A1(n19254), .A2(n20018), .ZN(n15607) );
  XNOR2_X1 U18820 ( .A(n15453), .B(n15459), .ZN(n16301) );
  NOR2_X1 U18821 ( .A1(n16475), .A2(n16301), .ZN(n15454) );
  AOI211_X1 U18822 ( .C1(n16477), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15607), .B(n15454), .ZN(n15455) );
  OAI21_X1 U18823 ( .B1(n16295), .B2(n16486), .A(n15455), .ZN(n15456) );
  AOI21_X1 U18824 ( .B1(n15610), .B2(n16493), .A(n15456), .ZN(n15457) );
  OAI21_X1 U18825 ( .B1(n15611), .B2(n16480), .A(n15457), .ZN(P2_U2984) );
  AOI21_X1 U18826 ( .B1(n16477), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15458), .ZN(n15462) );
  INV_X1 U18827 ( .A(n15459), .ZN(n15460) );
  AOI21_X1 U18828 ( .B1(n15469), .B2(n10166), .A(n15460), .ZN(n16279) );
  NAND2_X1 U18829 ( .A1(n16488), .A2(n16279), .ZN(n15461) );
  OAI211_X1 U18830 ( .C1(n16309), .C2(n16486), .A(n15462), .B(n15461), .ZN(
        n15463) );
  AOI21_X1 U18831 ( .B1(n15464), .B2(n16493), .A(n15463), .ZN(n15465) );
  OAI21_X1 U18832 ( .B1(n15466), .B2(n16480), .A(n15465), .ZN(P2_U2985) );
  NAND2_X1 U18833 ( .A1(n15467), .A2(n16494), .ZN(n15474) );
  INV_X1 U18834 ( .A(n15468), .ZN(n16320) );
  OAI21_X1 U18835 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n15479), .A(
        n15469), .ZN(n16323) );
  NAND2_X1 U18836 ( .A1(n16477), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15470) );
  OAI211_X1 U18837 ( .C1(n16475), .C2(n16323), .A(n15471), .B(n15470), .ZN(
        n15472) );
  AOI21_X1 U18838 ( .B1(n16320), .B2(n16491), .A(n15472), .ZN(n15473) );
  OAI211_X1 U18839 ( .C1(n15475), .C2(n16478), .A(n15474), .B(n15473), .ZN(
        P2_U2986) );
  XNOR2_X1 U18840 ( .A(n15476), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15621) );
  OR2_X1 U18841 ( .A1(n15477), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15612) );
  NAND3_X1 U18842 ( .A1(n15612), .A2(n15478), .A3(n16494), .ZN(n15484) );
  AOI21_X1 U18843 ( .B1(n15493), .B2(n15480), .A(n15479), .ZN(n16280) );
  INV_X1 U18844 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20011) );
  NOR2_X1 U18845 ( .A1(n19254), .A2(n20011), .ZN(n15615) );
  AOI21_X1 U18846 ( .B1(n16477), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15615), .ZN(n15481) );
  OAI21_X1 U18847 ( .B1(n16329), .B2(n16486), .A(n15481), .ZN(n15482) );
  AOI21_X1 U18848 ( .B1(n16280), .B2(n16488), .A(n15482), .ZN(n15483) );
  OAI211_X1 U18849 ( .C1(n16478), .C2(n15621), .A(n15484), .B(n15483), .ZN(
        P2_U2987) );
  INV_X1 U18850 ( .A(n15485), .ZN(n16389) );
  NOR2_X1 U18851 ( .A1(n15486), .A2(n16389), .ZN(n15488) );
  MUX2_X1 U18852 ( .A(n15488), .B(n16389), .S(n15487), .Z(n15490) );
  NAND2_X1 U18853 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n16388), .ZN(
        n16387) );
  NAND2_X1 U18854 ( .A1(n16502), .A2(n16387), .ZN(n15491) );
  NAND2_X1 U18855 ( .A1(n15492), .A2(n15491), .ZN(n16508) );
  AOI22_X1 U18856 ( .A1(n16506), .A2(n16491), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n16477), .ZN(n15496) );
  INV_X1 U18857 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20008) );
  OAI21_X1 U18858 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n9914), .A(
        n15493), .ZN(n16342) );
  OAI22_X1 U18859 ( .A1(n20008), .A2(n19254), .B1(n16475), .B2(n16342), .ZN(
        n15494) );
  INV_X1 U18860 ( .A(n15494), .ZN(n15495) );
  OAI211_X1 U18861 ( .C1(n16508), .C2(n16478), .A(n15496), .B(n15495), .ZN(
        n15497) );
  INV_X1 U18862 ( .A(n15497), .ZN(n15498) );
  OAI21_X1 U18863 ( .B1(n16512), .B2(n16480), .A(n15498), .ZN(P2_U2988) );
  INV_X1 U18864 ( .A(n15499), .ZN(n15501) );
  NAND2_X1 U18865 ( .A1(n15501), .A2(n15500), .ZN(n15502) );
  XNOR2_X1 U18866 ( .A(n15503), .B(n15502), .ZN(n15622) );
  NOR2_X1 U18867 ( .A1(n16400), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15504) );
  OR2_X1 U18868 ( .A1(n16388), .A2(n15504), .ZN(n15634) );
  INV_X1 U18869 ( .A(n15629), .ZN(n16360) );
  AOI22_X1 U18870 ( .A1(n16360), .A2(n16491), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n16477), .ZN(n15507) );
  INV_X1 U18871 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20004) );
  OAI21_X1 U18872 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n16282), .A(
        n16281), .ZN(n16364) );
  OAI22_X1 U18873 ( .A1(n20004), .A2(n19254), .B1(n16475), .B2(n16364), .ZN(
        n15505) );
  INV_X1 U18874 ( .A(n15505), .ZN(n15506) );
  OAI211_X1 U18875 ( .C1(n15634), .C2(n16478), .A(n15507), .B(n15506), .ZN(
        n15508) );
  AOI21_X1 U18876 ( .B1(n15622), .B2(n16494), .A(n15508), .ZN(n15509) );
  INV_X1 U18877 ( .A(n15509), .ZN(P2_U2990) );
  NAND2_X1 U18878 ( .A1(n15511), .A2(n15510), .ZN(n15513) );
  XOR2_X1 U18879 ( .A(n15513), .B(n15512), .Z(n15646) );
  NOR2_X1 U18880 ( .A1(n15638), .A2(n16486), .ZN(n15516) );
  INV_X1 U18881 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20000) );
  OAI21_X1 U18882 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n15514), .A(
        n16283), .ZN(n15916) );
  OAI22_X1 U18883 ( .A1(n20000), .A2(n19254), .B1(n16475), .B2(n15916), .ZN(
        n15515) );
  AOI211_X1 U18884 ( .C1(n16477), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15516), .B(n15515), .ZN(n15519) );
  INV_X1 U18885 ( .A(n15521), .ZN(n15517) );
  NAND2_X1 U18886 ( .A1(n15517), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16401) );
  NAND2_X1 U18887 ( .A1(n15521), .A2(n15639), .ZN(n15643) );
  NAND3_X1 U18888 ( .A1(n16401), .A2(n16493), .A3(n15643), .ZN(n15518) );
  OAI211_X1 U18889 ( .C1(n15646), .C2(n16480), .A(n15519), .B(n15518), .ZN(
        P2_U2992) );
  AND2_X2 U18890 ( .A1(n15813), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16443) );
  INV_X1 U18891 ( .A(n15721), .ZN(n15740) );
  INV_X1 U18892 ( .A(n15520), .ZN(n15637) );
  NOR2_X1 U18893 ( .A1(n15740), .A2(n15637), .ZN(n15551) );
  OAI21_X1 U18894 ( .B1(n15551), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15521), .ZN(n15662) );
  INV_X1 U18895 ( .A(n15776), .ZN(n15522) );
  INV_X1 U18896 ( .A(n15523), .ZN(n15769) );
  AND3_X1 U18897 ( .A1(n15769), .A2(n15524), .A3(n15775), .ZN(n15526) );
  INV_X1 U18898 ( .A(n15768), .ZN(n15525) );
  AOI21_X1 U18899 ( .B1(n15527), .B2(n15526), .A(n15525), .ZN(n15745) );
  AND2_X1 U18900 ( .A1(n15745), .A2(n15743), .ZN(n15733) );
  OAI21_X1 U18901 ( .B1(n15733), .B2(n15528), .A(n15735), .ZN(n15590) );
  INV_X1 U18902 ( .A(n15589), .ZN(n15529) );
  NOR2_X1 U18903 ( .A1(n15590), .A2(n15529), .ZN(n15577) );
  OAI21_X1 U18904 ( .B1(n15577), .B2(n15530), .A(n15579), .ZN(n15569) );
  AND2_X1 U18905 ( .A1(n15569), .A2(n15531), .ZN(n15544) );
  INV_X1 U18906 ( .A(n15532), .ZN(n15533) );
  OAI21_X1 U18907 ( .B1(n15544), .B2(n15533), .A(n15545), .ZN(n15537) );
  NAND2_X1 U18908 ( .A1(n15535), .A2(n15534), .ZN(n15536) );
  XNOR2_X1 U18909 ( .A(n15537), .B(n15536), .ZN(n15647) );
  NAND2_X1 U18910 ( .A1(n15647), .A2(n16494), .ZN(n15542) );
  NAND2_X1 U18911 ( .A1(n19404), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15653) );
  OAI21_X1 U18912 ( .B1(n16498), .B2(n15538), .A(n15653), .ZN(n15540) );
  NOR2_X1 U18913 ( .A1(n15654), .A2(n16486), .ZN(n15539) );
  AOI211_X1 U18914 ( .C1(n16488), .C2(n15914), .A(n15540), .B(n15539), .ZN(
        n15541) );
  OAI211_X1 U18915 ( .C1(n16478), .C2(n15662), .A(n15542), .B(n15541), .ZN(
        P2_U2993) );
  NOR2_X1 U18916 ( .A1(n15544), .A2(n15543), .ZN(n15549) );
  INV_X1 U18917 ( .A(n15545), .ZN(n15547) );
  NOR2_X1 U18918 ( .A1(n15547), .A2(n15546), .ZN(n15548) );
  XNOR2_X1 U18919 ( .A(n15549), .B(n15548), .ZN(n15673) );
  NAND2_X1 U18920 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15550) );
  NAND2_X1 U18921 ( .A1(n15570), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15564) );
  AOI21_X1 U18922 ( .B1(n15564), .B2(n15669), .A(n15551), .ZN(n15671) );
  INV_X1 U18923 ( .A(n19133), .ZN(n15554) );
  INV_X1 U18924 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15552) );
  NAND2_X1 U18925 ( .A1(n19404), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15664) );
  OAI21_X1 U18926 ( .B1(n16498), .B2(n15552), .A(n15664), .ZN(n15553) );
  AOI21_X1 U18927 ( .B1(n16488), .B2(n15554), .A(n15553), .ZN(n15555) );
  OAI21_X1 U18928 ( .B1(n15556), .B2(n16486), .A(n15555), .ZN(n15557) );
  AOI21_X1 U18929 ( .B1(n15671), .B2(n16493), .A(n15557), .ZN(n15558) );
  OAI21_X1 U18930 ( .B1(n15673), .B2(n16480), .A(n15558), .ZN(P2_U2994) );
  INV_X1 U18931 ( .A(n15567), .ZN(n15561) );
  NAND2_X1 U18932 ( .A1(n19142), .A2(n16488), .ZN(n15562) );
  NAND2_X1 U18933 ( .A1(n19404), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15675) );
  OAI211_X1 U18934 ( .C1(n15563), .C2(n16498), .A(n15562), .B(n15675), .ZN(
        n15565) );
  NAND2_X1 U18935 ( .A1(n15567), .A2(n15566), .ZN(n15568) );
  XNOR2_X1 U18936 ( .A(n15569), .B(n15568), .ZN(n15699) );
  AOI21_X1 U18937 ( .B1(n15689), .B2(n15584), .A(n15570), .ZN(n15694) );
  INV_X1 U18938 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19992) );
  OAI22_X1 U18939 ( .A1(n19992), .A2(n19254), .B1(n16475), .B2(n19155), .ZN(
        n15573) );
  INV_X1 U18940 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15571) );
  OAI22_X1 U18941 ( .A1(n15693), .A2(n16486), .B1(n16498), .B2(n15571), .ZN(
        n15572) );
  AOI211_X1 U18942 ( .C1(n15694), .C2(n16493), .A(n15573), .B(n15572), .ZN(
        n15574) );
  OAI21_X1 U18943 ( .B1(n16480), .B2(n15699), .A(n15574), .ZN(P2_U2996) );
  INV_X1 U18944 ( .A(n15575), .ZN(n15576) );
  NOR2_X1 U18945 ( .A1(n15577), .A2(n15576), .ZN(n15581) );
  NAND2_X1 U18946 ( .A1(n15579), .A2(n15578), .ZN(n15580) );
  XNOR2_X1 U18947 ( .A(n15581), .B(n15580), .ZN(n15710) );
  INV_X1 U18948 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19990) );
  OAI22_X1 U18949 ( .A1(n16498), .A2(n11202), .B1(n19990), .B2(n19254), .ZN(
        n15583) );
  INV_X1 U18950 ( .A(n19165), .ZN(n19176) );
  NOR2_X1 U18951 ( .A1(n19176), .A2(n16475), .ZN(n15582) );
  AOI211_X1 U18952 ( .C1(n19172), .C2(n16491), .A(n15583), .B(n15582), .ZN(
        n15586) );
  NOR2_X1 U18953 ( .A1(n15723), .A2(n15719), .ZN(n15700) );
  OAI211_X1 U18954 ( .C1(n15700), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16493), .B(n15584), .ZN(n15585) );
  OAI211_X1 U18955 ( .C1(n15710), .C2(n16480), .A(n15586), .B(n15585), .ZN(
        P2_U2997) );
  XNOR2_X1 U18956 ( .A(n15723), .B(n15719), .ZN(n15593) );
  INV_X1 U18957 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19988) );
  NOR2_X1 U18958 ( .A1(n19988), .A2(n19254), .ZN(n15588) );
  OAI22_X1 U18959 ( .A1(n10179), .A2(n16498), .B1(n16475), .B2(n19180), .ZN(
        n15587) );
  AOI211_X1 U18960 ( .C1(n19182), .C2(n16491), .A(n15588), .B(n15587), .ZN(
        n15592) );
  XNOR2_X1 U18961 ( .A(n15590), .B(n15589), .ZN(n15717) );
  NAND2_X1 U18962 ( .A1(n15717), .A2(n16494), .ZN(n15591) );
  OAI211_X1 U18963 ( .C1(n15593), .C2(n16478), .A(n15592), .B(n15591), .ZN(
        P2_U2998) );
  NAND2_X1 U18964 ( .A1(n15594), .A2(n15818), .ZN(n15597) );
  XNOR2_X1 U18965 ( .A(n15787), .B(n15595), .ZN(n15596) );
  XNOR2_X1 U18966 ( .A(n15597), .B(n15596), .ZN(n16558) );
  OAI21_X1 U18967 ( .B1(n15600), .B2(n15599), .A(n15598), .ZN(n16554) );
  INV_X1 U18968 ( .A(n16554), .ZN(n15603) );
  INV_X1 U18969 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19972) );
  OAI22_X1 U18970 ( .A1(n19972), .A2(n19254), .B1(n16475), .B2(n19240), .ZN(
        n15602) );
  OAI22_X1 U18971 ( .A1(n16486), .A2(n19242), .B1(n16498), .B2(n10174), .ZN(
        n15601) );
  AOI211_X1 U18972 ( .C1(n15603), .C2(n16493), .A(n15602), .B(n15601), .ZN(
        n15604) );
  OAI21_X1 U18973 ( .B1(n16480), .B2(n16558), .A(n15604), .ZN(P2_U3006) );
  NAND2_X1 U18974 ( .A1(n15605), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15609) );
  NAND3_X1 U18975 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15606) );
  NOR3_X1 U18976 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15606), .A3(
        n15613), .ZN(n15608) );
  NAND3_X1 U18977 ( .A1(n15612), .A2(n15478), .A3(n19414), .ZN(n15620) );
  NOR2_X1 U18978 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15613), .ZN(
        n15614) );
  AOI211_X1 U18979 ( .C1(n19420), .C2(n10431), .A(n15615), .B(n15614), .ZN(
        n15616) );
  OAI21_X1 U18980 ( .B1(n16329), .B2(n19411), .A(n15616), .ZN(n15617) );
  AOI21_X1 U18981 ( .B1(n15618), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15617), .ZN(n15619) );
  OAI211_X1 U18982 ( .C1(n15621), .C2(n19419), .A(n15620), .B(n15619), .ZN(
        P2_U3019) );
  NAND2_X1 U18983 ( .A1(n15622), .A2(n19414), .ZN(n15633) );
  NAND2_X1 U18984 ( .A1(n19420), .A2(n16361), .ZN(n15628) );
  INV_X1 U18985 ( .A(n15623), .ZN(n15625) );
  NOR2_X1 U18986 ( .A1(n20004), .A2(n19254), .ZN(n15624) );
  AOI21_X1 U18987 ( .B1(n15626), .B2(n15625), .A(n15624), .ZN(n15627) );
  OAI211_X1 U18988 ( .C1(n15629), .C2(n19411), .A(n15628), .B(n15627), .ZN(
        n15630) );
  AOI21_X1 U18989 ( .B1(n15631), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15630), .ZN(n15632) );
  OAI211_X1 U18990 ( .C1(n15634), .C2(n19419), .A(n15633), .B(n15632), .ZN(
        P2_U3022) );
  NAND2_X1 U18991 ( .A1(n19427), .A2(n15635), .ZN(n15636) );
  AND2_X1 U18992 ( .A1(n15795), .A2(n15636), .ZN(n15686) );
  AOI21_X1 U18993 ( .B1(n15637), .B2(n19427), .A(n15731), .ZN(n15656) );
  OAI21_X1 U18994 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15834), .A(
        n15656), .ZN(n16526) );
  NOR2_X1 U18995 ( .A1(n15638), .A2(n19411), .ZN(n15642) );
  AOI22_X1 U18996 ( .A1(n19404), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n16531), 
        .B2(n15639), .ZN(n15640) );
  OAI21_X1 U18997 ( .B1(n16551), .B2(n15924), .A(n15640), .ZN(n15641) );
  AOI211_X1 U18998 ( .C1(n16526), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15642), .B(n15641), .ZN(n15645) );
  NAND3_X1 U18999 ( .A1(n16401), .A2(n19429), .A3(n15643), .ZN(n15644) );
  OAI211_X1 U19000 ( .C1(n15646), .C2(n19436), .A(n15645), .B(n15644), .ZN(
        P2_U3024) );
  NAND2_X1 U19001 ( .A1(n15647), .A2(n19414), .ZN(n15661) );
  NOR2_X1 U19002 ( .A1(n15814), .A2(n15794), .ZN(n16542) );
  NAND2_X1 U19003 ( .A1(n15648), .A2(n16542), .ZN(n15762) );
  NAND2_X1 U19004 ( .A1(n10314), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15649) );
  NOR2_X1 U19005 ( .A1(n15762), .A2(n15649), .ZN(n15726) );
  AND2_X1 U19006 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15687), .ZN(
        n15650) );
  NAND2_X1 U19007 ( .A1(n15726), .A2(n15650), .ZN(n15676) );
  OR3_X1 U19008 ( .A1(n15676), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15651), .ZN(n15652) );
  OAI211_X1 U19009 ( .C1(n15654), .C2(n19411), .A(n15653), .B(n15652), .ZN(
        n15658) );
  NOR2_X1 U19010 ( .A1(n15656), .A2(n15655), .ZN(n15657) );
  AOI211_X1 U19011 ( .C1(n19420), .C2(n15659), .A(n15658), .B(n15657), .ZN(
        n15660) );
  OAI211_X1 U19012 ( .C1(n15662), .C2(n19419), .A(n15661), .B(n15660), .ZN(
        P2_U3025) );
  AOI21_X1 U19013 ( .B1(n15663), .B2(n19427), .A(n15731), .ZN(n15681) );
  XNOR2_X1 U19014 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15665) );
  OAI21_X1 U19015 ( .B1(n15676), .B2(n15665), .A(n15664), .ZN(n15667) );
  NOR2_X1 U19016 ( .A1(n16551), .A2(n19139), .ZN(n15666) );
  AOI211_X1 U19017 ( .C1(n19136), .C2(n14475), .A(n15667), .B(n15666), .ZN(
        n15668) );
  OAI21_X1 U19018 ( .B1(n15681), .B2(n15669), .A(n15668), .ZN(n15670) );
  AOI21_X1 U19019 ( .B1(n15671), .B2(n19429), .A(n15670), .ZN(n15672) );
  OAI21_X1 U19020 ( .B1(n15673), .B2(n19436), .A(n15672), .ZN(P2_U3026) );
  INV_X1 U19021 ( .A(n15674), .ZN(n15683) );
  OAI21_X1 U19022 ( .B1(n15676), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15675), .ZN(n15678) );
  NOR2_X1 U19023 ( .A1(n16551), .A2(n19146), .ZN(n15677) );
  AOI211_X1 U19024 ( .C1(n19148), .C2(n14475), .A(n15678), .B(n15677), .ZN(
        n15679) );
  OAI21_X1 U19025 ( .B1(n15681), .B2(n15680), .A(n15679), .ZN(n15682) );
  AOI21_X1 U19026 ( .B1(n15683), .B2(n19429), .A(n15682), .ZN(n15684) );
  OAI21_X1 U19027 ( .B1(n15685), .B2(n19436), .A(n15684), .ZN(P2_U3027) );
  INV_X1 U19028 ( .A(n19161), .ZN(n15697) );
  OAI21_X1 U19029 ( .B1(n15687), .B2(n15834), .A(n15686), .ZN(n15690) );
  INV_X1 U19030 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15689) );
  AND2_X1 U19031 ( .A1(n15687), .A2(n15726), .ZN(n15688) );
  AOI22_X1 U19032 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15690), .B1(
        n15689), .B2(n15688), .ZN(n15692) );
  NAND2_X1 U19033 ( .A1(n19404), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15691) );
  OAI211_X1 U19034 ( .C1(n15693), .C2(n19411), .A(n15692), .B(n15691), .ZN(
        n15696) );
  AND2_X1 U19035 ( .A1(n15694), .A2(n19429), .ZN(n15695) );
  AOI211_X1 U19036 ( .C1(n19420), .C2(n15697), .A(n15696), .B(n15695), .ZN(
        n15698) );
  OAI21_X1 U19037 ( .B1(n19436), .B2(n15699), .A(n15698), .ZN(P2_U3028) );
  AOI21_X1 U19038 ( .B1(n19419), .B2(n15701), .A(n15700), .ZN(n15702) );
  OAI21_X1 U19039 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15834), .A(
        n15720), .ZN(n15708) );
  INV_X1 U19040 ( .A(n15723), .ZN(n15704) );
  AOI22_X1 U19041 ( .A1(n15704), .A2(n19429), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15726), .ZN(n15714) );
  NOR3_X1 U19042 ( .A1(n15714), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15719), .ZN(n15707) );
  AOI22_X1 U19043 ( .A1(n19172), .A2(n14475), .B1(n19404), .B2(
        P2_REIP_REG_17__SCAN_IN), .ZN(n15705) );
  OAI21_X1 U19044 ( .B1(n16551), .B2(n19170), .A(n15705), .ZN(n15706) );
  AOI211_X1 U19045 ( .C1(n15708), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15707), .B(n15706), .ZN(n15709) );
  OAI21_X1 U19046 ( .B1(n15710), .B2(n19436), .A(n15709), .ZN(P2_U3029) );
  INV_X1 U19047 ( .A(n19186), .ZN(n15711) );
  AOI22_X1 U19048 ( .A1(n19420), .A2(n15711), .B1(n19404), .B2(
        P2_REIP_REG_16__SCAN_IN), .ZN(n15712) );
  OAI21_X1 U19049 ( .B1(n19411), .B2(n15713), .A(n15712), .ZN(n15716) );
  NOR2_X1 U19050 ( .A1(n15714), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15715) );
  AOI211_X1 U19051 ( .C1(n15717), .C2(n19414), .A(n15716), .B(n15715), .ZN(
        n15718) );
  OAI21_X1 U19052 ( .B1(n15720), .B2(n15719), .A(n15718), .ZN(P2_U3030) );
  OR2_X1 U19053 ( .A1(n15721), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15722) );
  NAND2_X1 U19054 ( .A1(n15723), .A2(n15722), .ZN(n16411) );
  NAND2_X1 U19055 ( .A1(n19420), .A2(n19307), .ZN(n15728) );
  AND2_X1 U19056 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19404), .ZN(n15724) );
  AOI21_X1 U19057 ( .B1(n15726), .B2(n15725), .A(n15724), .ZN(n15727) );
  OAI211_X1 U19058 ( .C1(n15729), .C2(n19411), .A(n15728), .B(n15727), .ZN(
        n15730) );
  AOI21_X1 U19059 ( .B1(n15731), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15730), .ZN(n15739) );
  INV_X1 U19060 ( .A(n15742), .ZN(n15732) );
  OR2_X1 U19061 ( .A1(n15733), .A2(n15732), .ZN(n15737) );
  NAND2_X1 U19062 ( .A1(n15735), .A2(n15734), .ZN(n15736) );
  XNOR2_X1 U19063 ( .A(n15737), .B(n15736), .ZN(n16407) );
  NAND2_X1 U19064 ( .A1(n16407), .A2(n19414), .ZN(n15738) );
  OAI211_X1 U19065 ( .C1(n16411), .C2(n19419), .A(n15739), .B(n15738), .ZN(
        P2_U3031) );
  INV_X1 U19066 ( .A(n15760), .ZN(n15741) );
  OAI21_X1 U19067 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15741), .A(
        n15740), .ZN(n16417) );
  AND2_X1 U19068 ( .A1(n15743), .A2(n15742), .ZN(n15744) );
  XNOR2_X1 U19069 ( .A(n15745), .B(n15744), .ZN(n16416) );
  NOR2_X1 U19070 ( .A1(n15746), .A2(n15762), .ZN(n15751) );
  NOR2_X1 U19071 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15762), .ZN(
        n15780) );
  NOR2_X1 U19072 ( .A1(n15814), .A2(n16541), .ZN(n15747) );
  OAI21_X1 U19073 ( .B1(n15747), .B2(n15834), .A(n15795), .ZN(n15781) );
  NOR2_X1 U19074 ( .A1(n15780), .A2(n15781), .ZN(n15765) );
  OAI21_X1 U19075 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15762), .A(
        n15765), .ZN(n15749) );
  INV_X1 U19076 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19984) );
  NOR2_X1 U19077 ( .A1(n19984), .A2(n19254), .ZN(n15748) );
  AOI221_X1 U19078 ( .B1(n15751), .B2(n15750), .C1(n15749), .C2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n15748), .ZN(n15757) );
  OR2_X1 U19079 ( .A1(n15752), .A2(n13228), .ZN(n15754) );
  NAND2_X1 U19080 ( .A1(n15754), .A2(n15753), .ZN(n19313) );
  INV_X1 U19081 ( .A(n19313), .ZN(n15755) );
  AOI22_X1 U19082 ( .A1(n14475), .A2(n19193), .B1(n19420), .B2(n15755), .ZN(
        n15756) );
  OAI211_X1 U19083 ( .C1(n16416), .C2(n19436), .A(n15757), .B(n15756), .ZN(
        n15758) );
  INV_X1 U19084 ( .A(n15758), .ZN(n15759) );
  OAI21_X1 U19085 ( .B1(n16417), .B2(n19419), .A(n15759), .ZN(P2_U3032) );
  OAI21_X1 U19086 ( .B1(n16442), .B2(n15774), .A(n15764), .ZN(n15761) );
  NAND2_X1 U19087 ( .A1(n15761), .A2(n15760), .ZN(n16424) );
  INV_X1 U19088 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19982) );
  OAI22_X1 U19089 ( .A1(n16551), .A2(n19201), .B1(n19982), .B2(n19254), .ZN(
        n15767) );
  OR2_X1 U19090 ( .A1(n15762), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15763) );
  OAI22_X1 U19091 ( .A1(n15765), .A2(n15764), .B1(n15774), .B2(n15763), .ZN(
        n15766) );
  AOI211_X1 U19092 ( .C1(n19202), .C2(n14475), .A(n15767), .B(n15766), .ZN(
        n15773) );
  AND2_X1 U19093 ( .A1(n15769), .A2(n15768), .ZN(n15770) );
  XNOR2_X1 U19094 ( .A(n15771), .B(n15770), .ZN(n16421) );
  NAND2_X1 U19095 ( .A1(n16421), .A2(n19414), .ZN(n15772) );
  OAI211_X1 U19096 ( .C1(n16424), .C2(n19419), .A(n15773), .B(n15772), .ZN(
        P2_U3033) );
  XNOR2_X1 U19097 ( .A(n16442), .B(n15774), .ZN(n16429) );
  AND2_X1 U19098 ( .A1(n15776), .A2(n15775), .ZN(n15777) );
  XNOR2_X1 U19099 ( .A(n15778), .B(n15777), .ZN(n16428) );
  INV_X1 U19100 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19980) );
  NOR2_X1 U19101 ( .A1(n19980), .A2(n19254), .ZN(n15779) );
  AOI211_X1 U19102 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15781), .A(
        n15780), .B(n15779), .ZN(n15784) );
  INV_X1 U19103 ( .A(n19224), .ZN(n15782) );
  AOI22_X1 U19104 ( .A1(n14475), .A2(n19220), .B1(n19420), .B2(n15782), .ZN(
        n15783) );
  OAI211_X1 U19105 ( .C1(n16428), .C2(n19436), .A(n15784), .B(n15783), .ZN(
        n15785) );
  INV_X1 U19106 ( .A(n15785), .ZN(n15786) );
  OAI21_X1 U19107 ( .B1(n16429), .B2(n19419), .A(n15786), .ZN(P2_U3034) );
  XNOR2_X1 U19108 ( .A(n16443), .B(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16450) );
  NAND2_X1 U19109 ( .A1(n15594), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15788) );
  NAND2_X1 U19110 ( .A1(n15788), .A2(n15787), .ZN(n15789) );
  OAI211_X1 U19111 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n15594), .A(
        n15789), .B(n15818), .ZN(n15802) );
  INV_X1 U19112 ( .A(n15790), .ZN(n15803) );
  NOR2_X1 U19113 ( .A1(n16439), .A2(n16436), .ZN(n15793) );
  INV_X1 U19114 ( .A(n16438), .ZN(n15791) );
  NOR2_X1 U19115 ( .A1(n15791), .A2(n16437), .ZN(n15792) );
  XNOR2_X1 U19116 ( .A(n15793), .B(n15792), .ZN(n16449) );
  NOR2_X1 U19117 ( .A1(n15794), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15810) );
  INV_X1 U19118 ( .A(n15795), .ZN(n15812) );
  OR2_X1 U19119 ( .A1(n15810), .A2(n15812), .ZN(n16537) );
  INV_X1 U19120 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19976) );
  NOR2_X1 U19121 ( .A1(n19976), .A2(n19254), .ZN(n15796) );
  AOI221_X1 U19122 ( .B1(n16542), .B2(n15797), .C1(n16537), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15796), .ZN(n15799) );
  NAND2_X1 U19123 ( .A1(n9912), .A2(n14475), .ZN(n15798) );
  OAI211_X1 U19124 ( .C1(n16551), .C2(n19235), .A(n15799), .B(n15798), .ZN(
        n15800) );
  AOI21_X1 U19125 ( .B1(n16449), .B2(n19414), .A(n15800), .ZN(n15801) );
  OAI21_X1 U19126 ( .B1(n19419), .B2(n16450), .A(n15801), .ZN(P2_U3036) );
  OAI21_X1 U19127 ( .B1(n15803), .B2(n16436), .A(n15802), .ZN(n15804) );
  OAI21_X1 U19128 ( .B1(n15805), .B2(n16436), .A(n15804), .ZN(n16461) );
  NAND2_X1 U19129 ( .A1(n19420), .A2(n15806), .ZN(n15808) );
  NAND2_X1 U19130 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19404), .ZN(n15807) );
  OAI211_X1 U19131 ( .C1(n15809), .C2(n19411), .A(n15808), .B(n15807), .ZN(
        n15811) );
  AOI211_X1 U19132 ( .C1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15812), .A(
        n15811), .B(n15810), .ZN(n15817) );
  INV_X1 U19133 ( .A(n16443), .ZN(n16457) );
  INV_X1 U19134 ( .A(n15813), .ZN(n15815) );
  NAND2_X1 U19135 ( .A1(n15815), .A2(n15814), .ZN(n16456) );
  NAND3_X1 U19136 ( .A1(n16457), .A2(n19429), .A3(n16456), .ZN(n15816) );
  OAI211_X1 U19137 ( .C1(n16461), .C2(n19436), .A(n15817), .B(n15816), .ZN(
        P2_U3037) );
  INV_X1 U19138 ( .A(n15818), .ZN(n15820) );
  OR2_X1 U19139 ( .A1(n15820), .A2(n15819), .ZN(n15821) );
  XNOR2_X1 U19140 ( .A(n15822), .B(n15821), .ZN(n16466) );
  NAND2_X1 U19141 ( .A1(n16466), .A2(n19414), .ZN(n15833) );
  INV_X1 U19142 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19970) );
  NOR2_X1 U19143 ( .A1(n19970), .A2(n19254), .ZN(n15823) );
  AOI221_X1 U19144 ( .B1(n16548), .B2(n15826), .C1(n16553), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15823), .ZN(n15832) );
  INV_X1 U19145 ( .A(n19257), .ZN(n15824) );
  AOI22_X1 U19146 ( .A1(n15825), .A2(n19420), .B1(n14475), .B2(n15824), .ZN(
        n15831) );
  XNOR2_X1 U19147 ( .A(n15827), .B(n15826), .ZN(n15828) );
  XNOR2_X1 U19148 ( .A(n15829), .B(n15828), .ZN(n16467) );
  NAND2_X1 U19149 ( .A1(n16467), .A2(n19429), .ZN(n15830) );
  NAND4_X1 U19150 ( .A1(n15833), .A2(n15832), .A3(n15831), .A4(n15830), .ZN(
        P2_U3039) );
  MUX2_X1 U19151 ( .A(n15834), .B(n19423), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n15845) );
  OR2_X1 U19152 ( .A1(n15836), .A2(n15835), .ZN(n15837) );
  AND2_X1 U19153 ( .A1(n15838), .A2(n15837), .ZN(n19363) );
  AOI22_X1 U19154 ( .A1(n19429), .A2(n15839), .B1(n19420), .B2(n19363), .ZN(
        n15844) );
  OAI21_X1 U19155 ( .B1(n10384), .B2(n19411), .A(n15840), .ZN(n15841) );
  AOI21_X1 U19156 ( .B1(n19414), .B2(n15842), .A(n15841), .ZN(n15843) );
  NAND3_X1 U19157 ( .A1(n15845), .A2(n15844), .A3(n15843), .ZN(P2_U3046) );
  OAI22_X1 U19158 ( .A1(n15847), .A2(n20030), .B1(n15846), .B2(n20031), .ZN(
        n15848) );
  AOI21_X1 U19159 ( .B1(n15849), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n15848), 
        .ZN(n15851) );
  NAND2_X1 U19160 ( .A1(n15880), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15850) );
  OAI21_X1 U19161 ( .B1(n15851), .B2(n15880), .A(n15850), .ZN(P2_U3601) );
  OAI22_X1 U19162 ( .A1(n20038), .A2(n20031), .B1(n20030), .B2(n15852), .ZN(
        n15853) );
  AOI21_X1 U19163 ( .B1(n15855), .B2(n15854), .A(n15853), .ZN(n15857) );
  NAND2_X1 U19164 ( .A1(n15880), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15856) );
  OAI21_X1 U19165 ( .B1(n15857), .B2(n15880), .A(n15856), .ZN(P2_U3600) );
  AOI22_X1 U19166 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15858) );
  OAI21_X1 U19167 ( .B1(n11496), .B2(n17233), .A(n15858), .ZN(n15868) );
  AOI22_X1 U19168 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11665), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15866) );
  OAI22_X1 U19169 ( .A1(n17415), .A2(n15859), .B1(n17416), .B2(n17469), .ZN(
        n15864) );
  AOI22_X1 U19170 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15862) );
  AOI22_X1 U19171 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15861) );
  AOI22_X1 U19172 ( .A1(n11629), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15860) );
  NAND3_X1 U19173 ( .A1(n15862), .A2(n15861), .A3(n15860), .ZN(n15863) );
  AOI211_X1 U19174 ( .C1(n17396), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n15864), .B(n15863), .ZN(n15865) );
  OAI211_X1 U19175 ( .C1(n9926), .C2(n17227), .A(n15866), .B(n15865), .ZN(
        n15867) );
  AOI211_X1 U19176 ( .C1(n17442), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n15868), .B(n15867), .ZN(n17586) );
  NOR2_X1 U19177 ( .A1(n17462), .A2(n15869), .ZN(n17409) );
  NAND2_X1 U19178 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17409), .ZN(n17389) );
  INV_X1 U19179 ( .A(n17389), .ZN(n17359) );
  NAND2_X1 U19180 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17376), .ZN(n17339) );
  OAI21_X1 U19181 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17376), .A(n17339), .ZN(
        n15870) );
  AOI22_X1 U19182 ( .A1(n17489), .A2(n17586), .B1(n15870), .B2(n17468), .ZN(
        P3_U2690) );
  NAND2_X1 U19183 ( .A1(n18903), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18433) );
  NAND2_X1 U19184 ( .A1(n15871), .A2(n17415), .ZN(n18431) );
  INV_X1 U19185 ( .A(n18431), .ZN(n15873) );
  OAI211_X1 U19186 ( .C1(n19032), .C2(n15873), .A(n18488), .B(n15872), .ZN(
        n18438) );
  NAND2_X1 U19187 ( .A1(n18433), .A2(n18438), .ZN(n15876) );
  INV_X1 U19188 ( .A(n15876), .ZN(n15875) );
  OAI22_X1 U19189 ( .A1(n19078), .A2(n17935), .B1(n19034), .B2(n18903), .ZN(
        n15878) );
  NAND3_X1 U19190 ( .A1(n18905), .A2(n18438), .A3(n15878), .ZN(n15874) );
  OAI221_X1 U19191 ( .B1(n18905), .B2(n15875), .C1(n18905), .C2(n18599), .A(
        n15874), .ZN(P3_U2864) );
  NAND2_X1 U19192 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18621) );
  NOR2_X1 U19193 ( .A1(n19078), .A2(n17935), .ZN(n15877) );
  AOI221_X1 U19194 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18621), .C1(n15877), 
        .C2(n18621), .A(n15876), .ZN(n18437) );
  INV_X1 U19195 ( .A(n18599), .ZN(n18787) );
  OAI221_X1 U19196 ( .B1(n18787), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18787), .C2(n15878), .A(n18438), .ZN(n18435) );
  AOI22_X1 U19197 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18437), .B1(
        n18435), .B2(n18910), .ZN(P3_U2865) );
  INV_X1 U19198 ( .A(n15880), .ZN(n20032) );
  OR3_X1 U19199 ( .A1(n15880), .A2(n20030), .A3(n15879), .ZN(n15881) );
  OAI21_X1 U19200 ( .B1(n20032), .B2(n15882), .A(n15881), .ZN(P2_U3595) );
  INV_X1 U19201 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16619) );
  NAND3_X1 U19202 ( .A1(n16653), .A2(n16640), .A3(n17969), .ZN(n15971) );
  INV_X1 U19203 ( .A(n15883), .ZN(n15970) );
  XNOR2_X1 U19204 ( .A(n18448), .B(n18452), .ZN(n15885) );
  AOI21_X1 U19205 ( .B1(n19082), .B2(n15885), .A(n18932), .ZN(n16751) );
  AND3_X1 U19206 ( .A1(n15886), .A2(n18871), .A3(n16751), .ZN(n15888) );
  INV_X1 U19207 ( .A(n15890), .ZN(n15891) );
  OAI21_X1 U19208 ( .B1(n15891), .B2(n18462), .A(n18868), .ZN(n15892) );
  NOR2_X1 U19209 ( .A1(n17613), .A2(n18873), .ZN(n18296) );
  NOR2_X1 U19210 ( .A1(n18427), .A2(n18276), .ZN(n18340) );
  INV_X1 U19211 ( .A(n18340), .ZN(n15900) );
  NAND3_X1 U19212 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n18116), .ZN(n16646) );
  NAND2_X1 U19213 ( .A1(n18867), .A2(n18409), .ZN(n18385) );
  NAND3_X1 U19214 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18117), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16647) );
  NAND3_X1 U19215 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15895) );
  NAND2_X1 U19216 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18355) );
  NOR2_X1 U19217 ( .A1(n15894), .A2(n18355), .ZN(n18210) );
  NAND3_X1 U19218 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18210), .ZN(n18330) );
  NOR2_X1 U19219 ( .A1(n15895), .A2(n18330), .ZN(n18237) );
  INV_X1 U19220 ( .A(n18237), .ZN(n15896) );
  NOR2_X1 U19221 ( .A1(n18213), .A2(n15896), .ZN(n18214) );
  NAND2_X1 U19222 ( .A1(n18218), .A2(n18214), .ZN(n16633) );
  AOI21_X1 U19223 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18372) );
  INV_X1 U19224 ( .A(n18210), .ZN(n15897) );
  NOR2_X1 U19225 ( .A1(n18372), .A2(n15897), .ZN(n18332) );
  NAND4_X1 U19226 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n18332), .ZN(n15904) );
  NOR2_X1 U19227 ( .A1(n15904), .A2(n15898), .ZN(n18166) );
  NAND2_X1 U19228 ( .A1(n18890), .A2(n18166), .ZN(n16635) );
  OAI21_X1 U19229 ( .B1(n18900), .B2(n16633), .A(n16635), .ZN(n15899) );
  NAND2_X1 U19230 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18237), .ZN(
        n18299) );
  NOR2_X1 U19231 ( .A1(n18213), .A2(n18299), .ZN(n18235) );
  AND2_X1 U19232 ( .A1(n18218), .A2(n18171), .ZN(n18169) );
  NAND2_X1 U19233 ( .A1(n18235), .A2(n18169), .ZN(n18164) );
  NOR2_X1 U19234 ( .A1(n18173), .A2(n18164), .ZN(n15903) );
  AOI22_X1 U19235 ( .A1(n17801), .A2(n15899), .B1(n15903), .B2(n18304), .ZN(
        n18136) );
  OR3_X1 U19236 ( .A1(n18136), .A2(n16638), .A3(n16640), .ZN(n16625) );
  OAI222_X1 U19237 ( .A1(n15900), .A2(n16646), .B1(n18385), .B2(n16647), .C1(
        n18427), .C2(n16625), .ZN(n15973) );
  INV_X1 U19238 ( .A(n15973), .ZN(n15911) );
  NAND2_X1 U19239 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15901) );
  NOR2_X1 U19240 ( .A1(n15901), .A2(n16619), .ZN(n15974) );
  NAND2_X1 U19241 ( .A1(n18117), .A2(n15974), .ZN(n16594) );
  NAND2_X1 U19242 ( .A1(n18116), .A2(n15974), .ZN(n16595) );
  AOI22_X1 U19243 ( .A1(n16594), .A2(n18425), .B1(n16595), .B2(n18340), .ZN(
        n15902) );
  INV_X1 U19244 ( .A(n15902), .ZN(n15976) );
  NAND2_X1 U19245 ( .A1(n18409), .A2(n18334), .ZN(n18411) );
  INV_X1 U19246 ( .A(n18110), .ZN(n17752) );
  NOR2_X1 U19247 ( .A1(n16637), .A2(n16633), .ZN(n18111) );
  AOI21_X1 U19248 ( .B1(n17752), .B2(n18111), .A(n18900), .ZN(n15907) );
  AOI21_X1 U19249 ( .B1(n15903), .B2(n16603), .A(n18898), .ZN(n15906) );
  INV_X1 U19250 ( .A(n15904), .ZN(n18236) );
  AND2_X1 U19251 ( .A1(n18236), .A2(n15905), .ZN(n18149) );
  AOI21_X1 U19252 ( .B1(n18149), .B2(n17752), .A(n18393), .ZN(n18120) );
  NOR4_X1 U19253 ( .A1(n15907), .A2(n15906), .A3(n18120), .A4(n18427), .ZN(
        n15975) );
  OAI21_X1 U19254 ( .B1(n18317), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15975), .ZN(n16651) );
  INV_X1 U19255 ( .A(n16651), .ZN(n15908) );
  OAI22_X1 U19256 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18411), .B1(
        n18416), .B2(n15908), .ZN(n15909) );
  NOR2_X1 U19257 ( .A1(n15976), .A2(n15909), .ZN(n15910) );
  MUX2_X1 U19258 ( .A(n15911), .B(n15910), .S(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(n15912) );
  NAND2_X1 U19259 ( .A1(n18416), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16611) );
  OAI211_X1 U19260 ( .C1(n16616), .C2(n18344), .A(n15912), .B(n16611), .ZN(
        P3_U2833) );
  OAI21_X1 U19261 ( .B1(n15914), .B2(n15913), .A(n14491), .ZN(n15915) );
  NAND2_X1 U19262 ( .A1(n15916), .A2(n15915), .ZN(n16284) );
  OAI211_X1 U19263 ( .C1(n15916), .C2(n15915), .A(n19245), .B(n16284), .ZN(
        n15918) );
  AOI22_X1 U19264 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19293), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19286), .ZN(n15917) );
  NAND2_X1 U19265 ( .A1(n15918), .A2(n15917), .ZN(n15919) );
  AOI21_X1 U19266 ( .B1(n19298), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15919), .ZN(n15923) );
  AOI22_X1 U19267 ( .A1(n15921), .A2(n19288), .B1(n15920), .B2(n19243), .ZN(
        n15922) );
  OAI211_X1 U19268 ( .C1(n15924), .C2(n19290), .A(n15923), .B(n15922), .ZN(
        P2_U2833) );
  NAND2_X1 U19269 ( .A1(n15935), .A2(n12471), .ZN(n15933) );
  AOI21_X1 U19270 ( .B1(n15925), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20670), .ZN(n15926) );
  NAND2_X1 U19271 ( .A1(n15927), .A2(n15926), .ZN(n15930) );
  OAI211_X1 U19272 ( .C1(n15930), .C2(n20631), .A(n15929), .B(n15928), .ZN(
        n15932) );
  NAND2_X1 U19273 ( .A1(n15930), .A2(n20631), .ZN(n15931) );
  NAND3_X1 U19274 ( .A1(n15933), .A2(n15932), .A3(n15931), .ZN(n15934) );
  OAI21_X1 U19275 ( .B1(n12471), .B2(n15935), .A(n15934), .ZN(n15937) );
  INV_X1 U19276 ( .A(n15936), .ZN(n15938) );
  AND2_X1 U19277 ( .A1(n15937), .A2(n15938), .ZN(n15939) );
  OAI22_X1 U19278 ( .A1(n15939), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        n15938), .B2(n15937), .ZN(n15940) );
  AND2_X1 U19279 ( .A1(n15940), .A2(n20228), .ZN(n15948) );
  OAI21_X1 U19280 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15941), .ZN(n15944) );
  NAND4_X1 U19281 ( .A1(n15944), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n15943), 
        .A4(n15942), .ZN(n15945) );
  NOR3_X1 U19282 ( .A1(n12299), .A2(n20254), .A3(n15979), .ZN(n15951) );
  NAND3_X1 U19283 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20811), .A3(n20237), 
        .ZN(n15949) );
  AOI22_X1 U19284 ( .A1(n15951), .A2(n15950), .B1(n15952), .B2(n15949), .ZN(
        n15954) );
  INV_X1 U19285 ( .A(n15954), .ZN(n16275) );
  AOI21_X1 U19286 ( .B1(n16272), .B2(n15955), .A(n16275), .ZN(n15957) );
  NOR2_X1 U19287 ( .A1(n15957), .A2(n20237), .ZN(n16278) );
  NAND2_X1 U19288 ( .A1(n16278), .A2(n15952), .ZN(n20804) );
  AOI211_X1 U19289 ( .C1(n20804), .C2(n15955), .A(n15954), .B(n15953), .ZN(
        n15961) );
  AOI21_X1 U19290 ( .B1(n20811), .B2(n12749), .A(n15956), .ZN(n16273) );
  AOI21_X1 U19291 ( .B1(n20906), .B2(n15958), .A(n15957), .ZN(n15959) );
  INV_X1 U19292 ( .A(n15959), .ZN(n15960) );
  AOI22_X1 U19293 ( .A1(n15961), .A2(n16273), .B1(n20237), .B2(n15960), .ZN(
        P1_U3161) );
  AOI22_X1 U19294 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15962), .B1(
        n16255), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15968) );
  INV_X1 U19295 ( .A(n15963), .ZN(n15966) );
  INV_X1 U19296 ( .A(n15964), .ZN(n15965) );
  AOI22_X1 U19297 ( .A1(n15966), .A2(n16268), .B1(n16263), .B2(n15965), .ZN(
        n15967) );
  OAI211_X1 U19298 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15969), .A(
        n15968), .B(n15967), .ZN(P1_U3010) );
  NOR2_X1 U19299 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15971), .ZN(
        n16574) );
  NOR2_X1 U19300 ( .A1(n16575), .A2(n16574), .ZN(n15972) );
  XOR2_X1 U19301 ( .A(n15972), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16606) );
  NOR2_X1 U19302 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16619), .ZN(
        n16602) );
  AOI22_X1 U19303 ( .A1(n18308), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n16602), 
        .B2(n15973), .ZN(n15978) );
  INV_X1 U19304 ( .A(n18334), .ZN(n18241) );
  AOI221_X1 U19305 ( .B1(n18241), .B2(n15975), .C1(n15974), .C2(n15975), .A(
        n18308), .ZN(n16623) );
  OAI21_X1 U19306 ( .B1(n16623), .B2(n15976), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15977) );
  OAI211_X1 U19307 ( .C1(n16606), .C2(n18344), .A(n15978), .B(n15977), .ZN(
        P3_U2832) );
  INV_X1 U19308 ( .A(HOLD), .ZN(n20819) );
  INV_X1 U19309 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20820) );
  NAND2_X1 U19310 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20820), .ZN(n15981) );
  INV_X1 U19311 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20999) );
  AOI21_X1 U19312 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(HOLD), .A(n20999), .ZN(
        n20817) );
  AOI22_X1 U19313 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20811), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(n20817), .ZN(n15980) );
  OAI211_X1 U19314 ( .C1(n20819), .C2(n15981), .A(n15980), .B(n15979), .ZN(
        P1_U3195) );
  AND2_X1 U19315 ( .A1(n15982), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NAND2_X1 U19316 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATEBS16_REG_SCAN_IN), .ZN(n20057) );
  OAI21_X1 U19317 ( .B1(n16562), .B2(n20057), .A(n20067), .ZN(n15983) );
  AOI21_X1 U19318 ( .B1(n15984), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n15983), 
        .ZN(n15985) );
  NOR2_X1 U19319 ( .A1(n16561), .A2(n15985), .ZN(P2_U3178) );
  INV_X1 U19320 ( .A(n16560), .ZN(n20081) );
  AOI221_X1 U19321 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16561), .C1(n20081), .C2(
        n16561), .A(n19737), .ZN(n20072) );
  INV_X1 U19322 ( .A(n20072), .ZN(n20073) );
  NOR2_X1 U19323 ( .A1(n15986), .A2(n20073), .ZN(P2_U3047) );
  INV_X1 U19324 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17716) );
  OR2_X1 U19325 ( .A1(n18478), .A2(n17494), .ZN(n17536) );
  AOI22_X1 U19326 ( .A1(n17639), .A2(BUF2_REG_0__SCAN_IN), .B1(n17638), .B2(
        n18092), .ZN(n15991) );
  OAI221_X1 U19327 ( .B1(n17642), .B2(n17716), .C1(n17642), .C2(n17536), .A(
        n15991), .ZN(P3_U2735) );
  OAI21_X1 U19328 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), 
        .A(n15992), .ZN(n16002) );
  INV_X1 U19329 ( .A(n16164), .ZN(n15997) );
  NAND2_X1 U19330 ( .A1(n20110), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n15993) );
  AND2_X1 U19331 ( .A1(n20154), .A2(n15993), .ZN(n15995) );
  NAND2_X1 U19332 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15994) );
  OAI211_X1 U19333 ( .C1(n20140), .C2(n16054), .A(n15995), .B(n15994), .ZN(
        n15996) );
  AOI21_X1 U19334 ( .B1(n15997), .B2(n20144), .A(n15996), .ZN(n16001) );
  OAI21_X1 U19335 ( .B1(n15999), .B2(n15998), .A(n16031), .ZN(n16013) );
  AOI22_X1 U19336 ( .A1(n16051), .A2(n20128), .B1(P1_REIP_REG_16__SCAN_IN), 
        .B2(n16013), .ZN(n16000) );
  OAI211_X1 U19337 ( .C1(n16012), .C2(n16002), .A(n16001), .B(n16000), .ZN(
        P1_U2824) );
  NOR2_X1 U19338 ( .A1(n16004), .A2(n16003), .ZN(n16005) );
  OR2_X1 U19339 ( .A1(n16006), .A2(n16005), .ZN(n16173) );
  INV_X1 U19340 ( .A(n16173), .ZN(n16040) );
  AOI22_X1 U19341 ( .A1(n16040), .A2(n20144), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n20110), .ZN(n16007) );
  OAI211_X1 U19342 ( .C1(n20136), .C2(n16008), .A(n16007), .B(n20154), .ZN(
        n16009) );
  AOI21_X1 U19343 ( .B1(n16059), .B2(n20158), .A(n16009), .ZN(n16011) );
  AOI22_X1 U19344 ( .A1(n16060), .A2(n20128), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n16013), .ZN(n16010) );
  OAI211_X1 U19345 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n16012), .A(n16011), 
        .B(n16010), .ZN(P1_U2825) );
  INV_X1 U19346 ( .A(n16013), .ZN(n16022) );
  AOI21_X1 U19347 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n16027), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n16021) );
  AOI22_X1 U19348 ( .A1(n20158), .A2(n16071), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n20110), .ZN(n16020) );
  INV_X1 U19349 ( .A(n16014), .ZN(n16072) );
  INV_X1 U19350 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16017) );
  NAND2_X1 U19351 ( .A1(n16015), .A2(n20144), .ZN(n16016) );
  OAI211_X1 U19352 ( .C1(n16017), .C2(n20136), .A(n16016), .B(n20154), .ZN(
        n16018) );
  AOI21_X1 U19353 ( .B1(n16072), .B2(n20128), .A(n16018), .ZN(n16019) );
  OAI211_X1 U19354 ( .C1(n16022), .C2(n16021), .A(n16020), .B(n16019), .ZN(
        P1_U2826) );
  INV_X1 U19355 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n16190) );
  AOI22_X1 U19356 ( .A1(n16189), .A2(n20144), .B1(n20110), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n16023) );
  OAI211_X1 U19357 ( .C1(n20136), .C2(n16024), .A(n16023), .B(n20154), .ZN(
        n16025) );
  AOI21_X1 U19358 ( .B1(n16026), .B2(n20158), .A(n16025), .ZN(n16030) );
  AOI22_X1 U19359 ( .A1(n16028), .A2(n20128), .B1(n16027), .B2(n16190), .ZN(
        n16029) );
  OAI211_X1 U19360 ( .C1(n16031), .C2(n16190), .A(n16030), .B(n16029), .ZN(
        P1_U2827) );
  INV_X1 U19361 ( .A(n16032), .ZN(n16230) );
  OAI222_X1 U19362 ( .A1(n21039), .A2(n20156), .B1(n20140), .B2(n16033), .C1(
        n16230), .C2(n20162), .ZN(n16034) );
  AOI211_X1 U19363 ( .C1(n20153), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20138), .B(n16034), .ZN(n16038) );
  AOI22_X1 U19364 ( .A1(n16036), .A2(n20128), .B1(P1_REIP_REG_10__SCAN_IN), 
        .B2(n16035), .ZN(n16037) );
  OAI211_X1 U19365 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n16039), .A(n16038), 
        .B(n16037), .ZN(P1_U2830) );
  INV_X1 U19366 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n21161) );
  AOI22_X1 U19367 ( .A1(n16060), .A2(n20182), .B1(n20181), .B2(n16040), .ZN(
        n16041) );
  OAI21_X1 U19368 ( .B1(n20185), .B2(n21161), .A(n16041), .ZN(P1_U2857) );
  AOI22_X1 U19369 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16255), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16053) );
  INV_X1 U19370 ( .A(n16042), .ZN(n16045) );
  NAND2_X1 U19371 ( .A1(n9849), .A2(n16043), .ZN(n16044) );
  AOI21_X1 U19372 ( .B1(n16046), .B2(n16045), .A(n16044), .ZN(n16056) );
  NOR2_X1 U19373 ( .A1(n16068), .A2(n14060), .ZN(n16047) );
  NOR2_X1 U19374 ( .A1(n16048), .A2(n16047), .ZN(n16055) );
  AND2_X1 U19375 ( .A1(n16056), .A2(n16055), .ZN(n16058) );
  NOR2_X1 U19376 ( .A1(n16058), .A2(n16048), .ZN(n16050) );
  XNOR2_X1 U19377 ( .A(n16050), .B(n16049), .ZN(n16167) );
  AOI22_X1 U19378 ( .A1(n16051), .A2(n16105), .B1(n16113), .B2(n16167), .ZN(
        n16052) );
  OAI211_X1 U19379 ( .C1(n16110), .C2(n16054), .A(n16053), .B(n16052), .ZN(
        P1_U2983) );
  NOR2_X1 U19380 ( .A1(n16056), .A2(n16055), .ZN(n16057) );
  INV_X1 U19381 ( .A(n16175), .ZN(n16063) );
  AOI22_X1 U19382 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16255), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16062) );
  AOI22_X1 U19383 ( .A1(n16060), .A2(n16105), .B1(n16084), .B2(n16059), .ZN(
        n16061) );
  OAI211_X1 U19384 ( .C1(n16063), .C2(n20095), .A(n16062), .B(n16061), .ZN(
        P1_U2984) );
  NAND3_X1 U19385 ( .A1(n16065), .A2(n16064), .A3(n16077), .ZN(n16067) );
  NAND2_X1 U19386 ( .A1(n16067), .A2(n16066), .ZN(n16070) );
  XNOR2_X1 U19387 ( .A(n16068), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16069) );
  XNOR2_X1 U19388 ( .A(n16070), .B(n16069), .ZN(n16187) );
  AOI22_X1 U19389 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16255), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16074) );
  AOI22_X1 U19390 ( .A1(n16072), .A2(n16105), .B1(n16084), .B2(n16071), .ZN(
        n16073) );
  OAI211_X1 U19391 ( .C1(n16187), .C2(n20095), .A(n16074), .B(n16073), .ZN(
        P1_U2985) );
  NAND2_X1 U19392 ( .A1(n16076), .A2(n16075), .ZN(n16081) );
  INV_X1 U19393 ( .A(n16077), .ZN(n16079) );
  OAI21_X1 U19394 ( .B1(n16089), .B2(n16079), .A(n16078), .ZN(n16080) );
  XOR2_X1 U19395 ( .A(n16081), .B(n16080), .Z(n16216) );
  AOI22_X1 U19396 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16255), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16087) );
  INV_X1 U19397 ( .A(n16082), .ZN(n16085) );
  AOI22_X1 U19398 ( .A1(n16085), .A2(n16105), .B1(n16084), .B2(n16083), .ZN(
        n16086) );
  OAI211_X1 U19399 ( .C1(n16216), .C2(n20095), .A(n16087), .B(n16086), .ZN(
        P1_U2987) );
  AOI22_X1 U19400 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16255), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16097) );
  NOR2_X1 U19401 ( .A1(n16088), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16092) );
  NOR2_X1 U19402 ( .A1(n16089), .A2(n13880), .ZN(n16091) );
  MUX2_X1 U19403 ( .A(n16092), .B(n16091), .S(n16090), .Z(n16093) );
  XOR2_X1 U19404 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16093), .Z(
        n16219) );
  INV_X1 U19405 ( .A(n16094), .ZN(n16095) );
  AOI22_X1 U19406 ( .A1(n16219), .A2(n16113), .B1(n16105), .B2(n16095), .ZN(
        n16096) );
  OAI211_X1 U19407 ( .C1(n16110), .C2(n16098), .A(n16097), .B(n16096), .ZN(
        P1_U2988) );
  AOI22_X1 U19408 ( .A1(n16099), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16255), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16107) );
  NAND2_X1 U19409 ( .A1(n16101), .A2(n16100), .ZN(n16102) );
  XNOR2_X1 U19410 ( .A(n16103), .B(n16102), .ZN(n16257) );
  INV_X1 U19411 ( .A(n16104), .ZN(n20177) );
  AOI22_X1 U19412 ( .A1(n16257), .A2(n16113), .B1(n16105), .B2(n20177), .ZN(
        n16106) );
  OAI211_X1 U19413 ( .C1(n16110), .C2(n20125), .A(n16107), .B(n16106), .ZN(
        P1_U2992) );
  INV_X1 U19414 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20135) );
  XOR2_X1 U19415 ( .A(n16109), .B(n16108), .Z(n16269) );
  OAI22_X1 U19416 ( .A1(n20134), .A2(n16111), .B1(n20141), .B2(n16110), .ZN(
        n16112) );
  AOI21_X1 U19417 ( .B1(n16269), .B2(n16113), .A(n16112), .ZN(n16115) );
  NOR2_X1 U19418 ( .A1(n12853), .A2(n21162), .ZN(n16262) );
  INV_X1 U19419 ( .A(n16262), .ZN(n16114) );
  OAI211_X1 U19420 ( .C1(n20135), .C2(n16116), .A(n16115), .B(n16114), .ZN(
        P1_U2994) );
  INV_X1 U19421 ( .A(n16117), .ZN(n16119) );
  AOI22_X1 U19422 ( .A1(n16119), .A2(n16268), .B1(n16263), .B2(n16118), .ZN(
        n16126) );
  INV_X1 U19423 ( .A(n16120), .ZN(n16122) );
  NOR2_X1 U19424 ( .A1(n12853), .A2(n21024), .ZN(n16121) );
  AOI221_X1 U19425 ( .B1(n16124), .B2(n16123), .C1(n16122), .C2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n16121), .ZN(n16125) );
  NAND2_X1 U19426 ( .A1(n16126), .A2(n16125), .ZN(P1_U3012) );
  NAND2_X1 U19427 ( .A1(n16145), .A2(n16162), .ZN(n16150) );
  AND3_X1 U19428 ( .A1(n16128), .A2(n16268), .A3(n16127), .ZN(n16147) );
  OAI21_X1 U19429 ( .B1(n16131), .B2(n16130), .A(n16129), .ZN(n16139) );
  NOR2_X1 U19430 ( .A1(n16133), .A2(n16132), .ZN(n16188) );
  INV_X1 U19431 ( .A(n16134), .ZN(n16135) );
  NOR2_X1 U19432 ( .A1(n16136), .A2(n16135), .ZN(n16137) );
  OR2_X1 U19433 ( .A1(n16188), .A2(n16137), .ZN(n16138) );
  OR2_X1 U19434 ( .A1(n16139), .A2(n16138), .ZN(n16195) );
  INV_X1 U19435 ( .A(n16195), .ZN(n16142) );
  NAND2_X1 U19436 ( .A1(n16141), .A2(n16140), .ZN(n16196) );
  NAND2_X1 U19437 ( .A1(n16142), .A2(n16196), .ZN(n16180) );
  AND2_X1 U19438 ( .A1(n16161), .A2(n16151), .ZN(n16143) );
  NOR2_X1 U19439 ( .A1(n16180), .A2(n16143), .ZN(n16160) );
  OAI22_X1 U19440 ( .A1(n16160), .A2(n16145), .B1(n16242), .B2(n16144), .ZN(
        n16146) );
  NOR2_X1 U19441 ( .A1(n16147), .A2(n16146), .ZN(n16149) );
  NAND2_X1 U19442 ( .A1(n16255), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16148) );
  OAI211_X1 U19443 ( .C1(n16151), .C2(n16150), .A(n16149), .B(n16148), .ZN(
        P1_U3013) );
  INV_X1 U19444 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16169) );
  NOR3_X1 U19445 ( .A1(n16183), .A2(n14060), .A3(n16169), .ZN(n16152) );
  AOI21_X1 U19446 ( .B1(n16152), .B2(n16162), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16159) );
  INV_X1 U19447 ( .A(n16153), .ZN(n16156) );
  INV_X1 U19448 ( .A(n16154), .ZN(n16155) );
  AOI22_X1 U19449 ( .A1(n16156), .A2(n16268), .B1(n16263), .B2(n16155), .ZN(
        n16158) );
  NAND2_X1 U19450 ( .A1(n16255), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16157) );
  OAI211_X1 U19451 ( .C1(n16160), .C2(n16159), .A(n16158), .B(n16157), .ZN(
        P1_U3014) );
  AOI21_X1 U19452 ( .B1(n16183), .B2(n16161), .A(n16180), .ZN(n16177) );
  NAND2_X1 U19453 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16162), .ZN(
        n16170) );
  AOI221_X1 U19454 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n14060), .C2(n16169), .A(
        n16170), .ZN(n16166) );
  INV_X1 U19455 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n16163) );
  OAI22_X1 U19456 ( .A1(n16164), .A2(n16242), .B1(n16163), .B2(n12853), .ZN(
        n16165) );
  AOI211_X1 U19457 ( .C1(n16167), .C2(n16268), .A(n16166), .B(n16165), .ZN(
        n16168) );
  OAI21_X1 U19458 ( .B1(n16177), .B2(n16169), .A(n16168), .ZN(P1_U3015) );
  INV_X1 U19459 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21058) );
  OAI22_X1 U19460 ( .A1(n12853), .A2(n21058), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16170), .ZN(n16171) );
  INV_X1 U19461 ( .A(n16171), .ZN(n16172) );
  OAI21_X1 U19462 ( .B1(n16173), .B2(n16242), .A(n16172), .ZN(n16174) );
  AOI21_X1 U19463 ( .B1(n16175), .B2(n16268), .A(n16174), .ZN(n16176) );
  OAI21_X1 U19464 ( .B1(n16177), .B2(n14060), .A(n16176), .ZN(P1_U3016) );
  INV_X1 U19465 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20963) );
  OAI22_X1 U19466 ( .A1(n16178), .A2(n16242), .B1(n20963), .B2(n12853), .ZN(
        n16179) );
  AOI21_X1 U19467 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16180), .A(
        n16179), .ZN(n16186) );
  NOR2_X1 U19468 ( .A1(n16222), .A2(n16210), .ZN(n16184) );
  NOR2_X1 U19469 ( .A1(n16182), .A2(n16181), .ZN(n16218) );
  NAND4_X1 U19470 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16184), .A3(
        n16218), .A4(n16183), .ZN(n16185) );
  OAI211_X1 U19471 ( .C1(n16187), .C2(n16215), .A(n16186), .B(n16185), .ZN(
        P1_U3017) );
  INV_X1 U19472 ( .A(n16188), .ZN(n16199) );
  INV_X1 U19473 ( .A(n16189), .ZN(n16191) );
  OAI22_X1 U19474 ( .A1(n16191), .A2(n16242), .B1(n16190), .B2(n12853), .ZN(
        n16194) );
  NOR2_X1 U19475 ( .A1(n16192), .A2(n16215), .ZN(n16193) );
  AOI211_X1 U19476 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16195), .A(
        n16194), .B(n16193), .ZN(n16197) );
  OAI211_X1 U19477 ( .C1(n16199), .C2(n16198), .A(n16197), .B(n16196), .ZN(
        P1_U3018) );
  NOR2_X1 U19478 ( .A1(n16201), .A2(n16200), .ZN(n16203) );
  AOI211_X1 U19479 ( .C1(n16205), .C2(n16204), .A(n16203), .B(n16202), .ZN(
        n16223) );
  OAI21_X1 U19480 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16206), .A(
        n16223), .ZN(n16209) );
  OAI22_X1 U19481 ( .A1(n16207), .A2(n16242), .B1(n21200), .B2(n12853), .ZN(
        n16208) );
  AOI21_X1 U19482 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16209), .A(
        n16208), .ZN(n16214) );
  NAND3_X1 U19483 ( .A1(n16212), .A2(n16211), .A3(n16210), .ZN(n16213) );
  OAI211_X1 U19484 ( .C1(n16216), .C2(n16215), .A(n16214), .B(n16213), .ZN(
        P1_U3019) );
  AOI22_X1 U19485 ( .A1(n16217), .A2(n16263), .B1(n16255), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16221) );
  AOI22_X1 U19486 ( .A1(n16219), .A2(n16268), .B1(n16218), .B2(n16222), .ZN(
        n16220) );
  OAI211_X1 U19487 ( .C1(n16223), .C2(n16222), .A(n16221), .B(n16220), .ZN(
        P1_U3020) );
  INV_X1 U19488 ( .A(n16224), .ZN(n16228) );
  NAND4_X1 U19489 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16229), .A3(
        n16226), .A4(n16225), .ZN(n16227) );
  NAND2_X1 U19490 ( .A1(n16228), .A2(n16227), .ZN(n16247) );
  NAND2_X1 U19491 ( .A1(n16229), .A2(n16256), .ZN(n16236) );
  AOI221_X1 U19492 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n13880), .C2(n14052), .A(
        n16236), .ZN(n16232) );
  OAI22_X1 U19493 ( .A1(n16230), .A2(n16242), .B1(n21048), .B2(n12853), .ZN(
        n16231) );
  AOI211_X1 U19494 ( .C1(n16233), .C2(n16268), .A(n16232), .B(n16231), .ZN(
        n16234) );
  OAI21_X1 U19495 ( .B1(n13880), .B2(n16247), .A(n16234), .ZN(P1_U3021) );
  INV_X1 U19496 ( .A(n16235), .ZN(n16245) );
  NOR2_X1 U19497 ( .A1(n16236), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16244) );
  OR2_X1 U19498 ( .A1(n16238), .A2(n16237), .ZN(n16239) );
  NAND2_X1 U19499 ( .A1(n16240), .A2(n16239), .ZN(n20170) );
  INV_X1 U19500 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20121) );
  OAI22_X1 U19501 ( .A1(n20170), .A2(n16242), .B1(n20121), .B2(n12853), .ZN(
        n16243) );
  AOI211_X1 U19502 ( .C1(n16245), .C2(n16268), .A(n16244), .B(n16243), .ZN(
        n16246) );
  OAI21_X1 U19503 ( .B1(n14052), .B2(n16247), .A(n16246), .ZN(P1_U3022) );
  INV_X1 U19504 ( .A(n16248), .ZN(n16251) );
  INV_X1 U19505 ( .A(n16249), .ZN(n16250) );
  OAI21_X1 U19506 ( .B1(n16252), .B2(n16251), .A(n16250), .ZN(n16253) );
  AND2_X1 U19507 ( .A1(n16254), .A2(n16253), .ZN(n20176) );
  AOI22_X1 U19508 ( .A1(n20176), .A2(n16263), .B1(n16255), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16259) );
  AOI22_X1 U19509 ( .A1(n16257), .A2(n16268), .B1(n16256), .B2(n16260), .ZN(
        n16258) );
  OAI211_X1 U19510 ( .C1(n16261), .C2(n16260), .A(n16259), .B(n16258), .ZN(
        P1_U3024) );
  AOI21_X1 U19511 ( .B1(n20143), .B2(n16263), .A(n16262), .ZN(n16264) );
  OAI21_X1 U19512 ( .B1(n16266), .B2(n16265), .A(n16264), .ZN(n16267) );
  AOI21_X1 U19513 ( .B1(n16269), .B2(n16268), .A(n16267), .ZN(n16270) );
  OAI21_X1 U19514 ( .B1(n16271), .B2(n13614), .A(n16270), .ZN(P1_U3026) );
  AOI221_X1 U19515 ( .B1(n20811), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20703), 
        .C2(n20237), .A(n16272), .ZN(n20803) );
  AOI21_X1 U19516 ( .B1(n16273), .B2(n16278), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n16274) );
  AOI221_X1 U19517 ( .B1(n16276), .B2(n16275), .C1(n20803), .C2(n16275), .A(
        n16274), .ZN(P1_U3162) );
  OAI21_X1 U19518 ( .B1(n16278), .B2(n20637), .A(n16277), .ZN(P1_U3466) );
  INV_X1 U19519 ( .A(n16279), .ZN(n16313) );
  INV_X1 U19520 ( .A(n16280), .ZN(n16333) );
  AOI21_X1 U19521 ( .B1(n11229), .B2(n16281), .A(n9914), .ZN(n16386) );
  INV_X1 U19522 ( .A(n16386), .ZN(n16352) );
  AOI21_X1 U19523 ( .B1(n16405), .B2(n16283), .A(n16282), .ZN(n16395) );
  INV_X1 U19524 ( .A(n16395), .ZN(n16375) );
  NAND2_X1 U19525 ( .A1(n14491), .A2(n16284), .ZN(n16374) );
  NAND2_X1 U19526 ( .A1(n16375), .A2(n16374), .ZN(n16373) );
  NAND2_X1 U19527 ( .A1(n14491), .A2(n16373), .ZN(n16363) );
  NAND2_X1 U19528 ( .A1(n16364), .A2(n16363), .ZN(n16362) );
  NAND2_X1 U19529 ( .A1(n14491), .A2(n16362), .ZN(n16351) );
  NAND2_X1 U19530 ( .A1(n16352), .A2(n16351), .ZN(n16350) );
  NAND2_X1 U19531 ( .A1(n14491), .A2(n16350), .ZN(n16341) );
  NAND2_X1 U19532 ( .A1(n16342), .A2(n16341), .ZN(n16340) );
  NAND2_X1 U19533 ( .A1(n14491), .A2(n16340), .ZN(n16332) );
  NAND2_X1 U19534 ( .A1(n16333), .A2(n16332), .ZN(n16331) );
  NAND2_X1 U19535 ( .A1(n14491), .A2(n16331), .ZN(n16322) );
  NAND2_X1 U19536 ( .A1(n16323), .A2(n16322), .ZN(n16321) );
  NAND2_X1 U19537 ( .A1(n9797), .A2(n16321), .ZN(n16312) );
  NAND2_X1 U19538 ( .A1(n16313), .A2(n16312), .ZN(n16311) );
  NAND2_X1 U19539 ( .A1(n9797), .A2(n16311), .ZN(n16300) );
  NAND2_X1 U19540 ( .A1(n16301), .A2(n16300), .ZN(n16299) );
  INV_X1 U19541 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20020) );
  NAND2_X1 U19542 ( .A1(n16285), .A2(n19288), .ZN(n16289) );
  NAND3_X1 U19543 ( .A1(n16287), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n16286), 
        .ZN(n16288) );
  OAI211_X1 U19544 ( .C1(n19256), .C2(n20020), .A(n16289), .B(n16288), .ZN(
        n16290) );
  AOI21_X1 U19545 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19298), .A(
        n16290), .ZN(n16293) );
  AOI22_X1 U19546 ( .A1(n16291), .A2(n19243), .B1(n19203), .B2(n19303), .ZN(
        n16292) );
  OAI211_X1 U19547 ( .C1(n19162), .C2(n16299), .A(n16293), .B(n16292), .ZN(
        P2_U2824) );
  AOI22_X1 U19548 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19286), .ZN(n16305) );
  AOI22_X1 U19549 ( .A1(n16294), .A2(n19288), .B1(P2_EBX_REG_30__SCAN_IN), 
        .B2(n19293), .ZN(n16304) );
  OR2_X1 U19550 ( .A1(n16295), .A2(n19295), .ZN(n16298) );
  NAND2_X1 U19551 ( .A1(n16296), .A2(n19203), .ZN(n16297) );
  AND2_X1 U19552 ( .A1(n16298), .A2(n16297), .ZN(n16303) );
  OAI211_X1 U19553 ( .C1(n16301), .C2(n16300), .A(n19245), .B(n16299), .ZN(
        n16302) );
  AOI22_X1 U19554 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19286), .ZN(n16317) );
  AOI22_X1 U19555 ( .A1(n16306), .A2(n19288), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n19293), .ZN(n16316) );
  INV_X1 U19556 ( .A(n16307), .ZN(n16308) );
  OAI22_X1 U19557 ( .A1(n16309), .A2(n19295), .B1(n16308), .B2(n19290), .ZN(
        n16310) );
  INV_X1 U19558 ( .A(n16310), .ZN(n16315) );
  OAI211_X1 U19559 ( .C1(n16313), .C2(n16312), .A(n19245), .B(n16311), .ZN(
        n16314) );
  NAND4_X1 U19560 ( .A1(n16317), .A2(n16316), .A3(n16315), .A4(n16314), .ZN(
        P2_U2826) );
  AOI22_X1 U19561 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19286), .ZN(n16327) );
  AOI22_X1 U19562 ( .A1(n16318), .A2(n19288), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n19293), .ZN(n16326) );
  AOI22_X1 U19563 ( .A1(n16320), .A2(n19243), .B1(n16319), .B2(n19203), .ZN(
        n16325) );
  OAI211_X1 U19564 ( .C1(n16323), .C2(n16322), .A(n19245), .B(n16321), .ZN(
        n16324) );
  NAND4_X1 U19565 ( .A1(n16327), .A2(n16326), .A3(n16325), .A4(n16324), .ZN(
        P2_U2827) );
  AOI22_X1 U19566 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19286), .ZN(n16337) );
  AOI22_X1 U19567 ( .A1(n16328), .A2(n19288), .B1(P2_EBX_REG_27__SCAN_IN), 
        .B2(n19293), .ZN(n16336) );
  INV_X1 U19568 ( .A(n16329), .ZN(n16330) );
  AOI22_X1 U19569 ( .A1(n16330), .A2(n19243), .B1(n10431), .B2(n19203), .ZN(
        n16335) );
  OAI211_X1 U19570 ( .C1(n16333), .C2(n16332), .A(n19245), .B(n16331), .ZN(
        n16334) );
  NAND4_X1 U19571 ( .A1(n16337), .A2(n16336), .A3(n16335), .A4(n16334), .ZN(
        P2_U2828) );
  AOI22_X1 U19572 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19286), .ZN(n16346) );
  AOI22_X1 U19573 ( .A1(n16338), .A2(n19288), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n19293), .ZN(n16345) );
  INV_X1 U19574 ( .A(n16501), .ZN(n16339) );
  AOI22_X1 U19575 ( .A1(n16506), .A2(n19243), .B1(n16339), .B2(n19203), .ZN(
        n16344) );
  OAI211_X1 U19576 ( .C1(n16342), .C2(n16341), .A(n19245), .B(n16340), .ZN(
        n16343) );
  NAND4_X1 U19577 ( .A1(n16346), .A2(n16345), .A3(n16344), .A4(n16343), .ZN(
        P2_U2829) );
  AOI22_X1 U19578 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19286), .ZN(n16356) );
  AOI22_X1 U19579 ( .A1(n16347), .A2(n19288), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n19293), .ZN(n16355) );
  INV_X1 U19580 ( .A(n16348), .ZN(n16520) );
  INV_X1 U19581 ( .A(n16349), .ZN(n16519) );
  AOI22_X1 U19582 ( .A1(n16520), .A2(n19243), .B1(n19203), .B2(n16519), .ZN(
        n16354) );
  OAI211_X1 U19583 ( .C1(n16352), .C2(n16351), .A(n19245), .B(n16350), .ZN(
        n16353) );
  NAND4_X1 U19584 ( .A1(n16356), .A2(n16355), .A3(n16354), .A4(n16353), .ZN(
        P2_U2830) );
  AOI22_X1 U19585 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19286), .ZN(n16368) );
  OAI22_X1 U19586 ( .A1(n16358), .A2(n19266), .B1(n19271), .B2(n16357), .ZN(
        n16359) );
  INV_X1 U19587 ( .A(n16359), .ZN(n16367) );
  AOI22_X1 U19588 ( .A1(n16361), .A2(n19203), .B1(n19243), .B2(n16360), .ZN(
        n16366) );
  OAI211_X1 U19589 ( .C1(n16364), .C2(n16363), .A(n19245), .B(n16362), .ZN(
        n16365) );
  NAND4_X1 U19590 ( .A1(n16368), .A2(n16367), .A3(n16366), .A4(n16365), .ZN(
        P2_U2831) );
  AOI22_X1 U19591 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19286), .ZN(n16379) );
  AOI22_X1 U19592 ( .A1(n16369), .A2(n19288), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n19293), .ZN(n16378) );
  INV_X1 U19593 ( .A(n16370), .ZN(n16371) );
  AOI21_X1 U19594 ( .B1(n9929), .B2(n15411), .A(n16371), .ZN(n16525) );
  INV_X1 U19595 ( .A(n16372), .ZN(n16527) );
  AOI22_X1 U19596 ( .A1(n16525), .A2(n19203), .B1(n19243), .B2(n16527), .ZN(
        n16377) );
  OAI211_X1 U19597 ( .C1(n16375), .C2(n16374), .A(n19245), .B(n16373), .ZN(
        n16376) );
  NAND4_X1 U19598 ( .A1(n16379), .A2(n16378), .A3(n16377), .A4(n16376), .ZN(
        P2_U2832) );
  AOI22_X1 U19599 ( .A1(n16381), .A2(n16380), .B1(n19359), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16385) );
  AOI22_X1 U19600 ( .A1(n19304), .A2(BUF1_REG_23__SCAN_IN), .B1(n19302), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n16384) );
  AOI22_X1 U19601 ( .A1(n16382), .A2(n19361), .B1(n19360), .B2(n16525), .ZN(
        n16383) );
  NAND3_X1 U19602 ( .A1(n16385), .A2(n16384), .A3(n16383), .ZN(P2_U2896) );
  AOI22_X1 U19603 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19404), .B1(n16488), 
        .B2(n16386), .ZN(n16394) );
  OAI21_X1 U19604 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16388), .A(
        n16387), .ZN(n16524) );
  INV_X1 U19605 ( .A(n16524), .ZN(n16392) );
  NOR2_X1 U19606 ( .A1(n16390), .A2(n16389), .ZN(n16391) );
  OAI211_X1 U19607 ( .C1(n11229), .C2(n16498), .A(n16394), .B(n16393), .ZN(
        P2_U2989) );
  AOI22_X1 U19608 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19404), .B1(n16488), 
        .B2(n16395), .ZN(n16404) );
  OAI21_X1 U19609 ( .B1(n16398), .B2(n16397), .A(n16396), .ZN(n16399) );
  INV_X1 U19610 ( .A(n16399), .ZN(n16529) );
  INV_X1 U19611 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16402) );
  AOI21_X1 U19612 ( .B1(n16402), .B2(n16401), .A(n16400), .ZN(n16528) );
  AOI222_X1 U19613 ( .A1(n16529), .A2(n16494), .B1(n16493), .B2(n16528), .C1(
        n16491), .C2(n16527), .ZN(n16403) );
  OAI211_X1 U19614 ( .C1(n16405), .C2(n16498), .A(n16404), .B(n16403), .ZN(
        P2_U2991) );
  AOI22_X1 U19615 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19404), .B1(n16488), 
        .B2(n16406), .ZN(n16414) );
  NAND2_X1 U19616 ( .A1(n16407), .A2(n16494), .ZN(n16410) );
  NAND2_X1 U19617 ( .A1(n16491), .A2(n16408), .ZN(n16409) );
  OAI211_X1 U19618 ( .C1(n16411), .C2(n16478), .A(n16410), .B(n16409), .ZN(
        n16412) );
  INV_X1 U19619 ( .A(n16412), .ZN(n16413) );
  OAI211_X1 U19620 ( .C1(n16415), .C2(n16498), .A(n16414), .B(n16413), .ZN(
        P2_U2999) );
  AOI22_X1 U19621 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16477), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19404), .ZN(n16420) );
  OAI22_X1 U19622 ( .A1(n16417), .A2(n16478), .B1(n16480), .B2(n16416), .ZN(
        n16418) );
  AOI21_X1 U19623 ( .B1(n16491), .B2(n19193), .A(n16418), .ZN(n16419) );
  OAI211_X1 U19624 ( .C1(n16475), .C2(n19192), .A(n16420), .B(n16419), .ZN(
        P2_U3000) );
  AOI22_X1 U19625 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19404), .B1(n16488), 
        .B2(n19206), .ZN(n16427) );
  NAND2_X1 U19626 ( .A1(n16421), .A2(n16494), .ZN(n16423) );
  NAND2_X1 U19627 ( .A1(n16491), .A2(n19202), .ZN(n16422) );
  OAI211_X1 U19628 ( .C1(n16424), .C2(n16478), .A(n16423), .B(n16422), .ZN(
        n16425) );
  INV_X1 U19629 ( .A(n16425), .ZN(n16426) );
  OAI211_X1 U19630 ( .C1(n19197), .C2(n16498), .A(n16427), .B(n16426), .ZN(
        P2_U3001) );
  AOI22_X1 U19631 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16477), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19404), .ZN(n16432) );
  OAI22_X1 U19632 ( .A1(n16429), .A2(n16478), .B1(n16428), .B2(n16480), .ZN(
        n16430) );
  AOI21_X1 U19633 ( .B1(n16491), .B2(n19220), .A(n16430), .ZN(n16431) );
  OAI211_X1 U19634 ( .C1(n16475), .C2(n19218), .A(n16432), .B(n16431), .ZN(
        P2_U3002) );
  AOI22_X1 U19635 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19404), .B1(n16488), 
        .B2(n16433), .ZN(n16447) );
  NAND2_X1 U19636 ( .A1(n16435), .A2(n16434), .ZN(n16441) );
  AOI211_X1 U19637 ( .C1(n16439), .C2(n16438), .A(n16437), .B(n16436), .ZN(
        n16440) );
  XOR2_X1 U19638 ( .A(n16441), .B(n16440), .Z(n16540) );
  INV_X1 U19639 ( .A(n16442), .ZN(n16445) );
  AOI21_X1 U19640 ( .B1(n16443), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16444) );
  NOR2_X1 U19641 ( .A1(n16445), .A2(n16444), .ZN(n16538) );
  AOI222_X1 U19642 ( .A1(n16540), .A2(n16494), .B1(n16491), .B2(n16539), .C1(
        n16493), .C2(n16538), .ZN(n16446) );
  OAI211_X1 U19643 ( .C1(n16448), .C2(n16498), .A(n16447), .B(n16446), .ZN(
        P2_U3003) );
  AOI22_X1 U19644 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16477), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19404), .ZN(n16454) );
  INV_X1 U19645 ( .A(n16449), .ZN(n16451) );
  OAI22_X1 U19646 ( .A1(n16451), .A2(n16480), .B1(n16478), .B2(n16450), .ZN(
        n16452) );
  AOI21_X1 U19647 ( .B1(n16491), .B2(n9912), .A(n16452), .ZN(n16453) );
  OAI211_X1 U19648 ( .C1(n16475), .C2(n19230), .A(n16454), .B(n16453), .ZN(
        P2_U3004) );
  AOI22_X1 U19649 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19404), .B1(n16488), 
        .B2(n16455), .ZN(n16464) );
  NAND3_X1 U19650 ( .A1(n16457), .A2(n16493), .A3(n16456), .ZN(n16460) );
  NAND2_X1 U19651 ( .A1(n16458), .A2(n16491), .ZN(n16459) );
  OAI211_X1 U19652 ( .C1(n16461), .C2(n16480), .A(n16460), .B(n16459), .ZN(
        n16462) );
  INV_X1 U19653 ( .A(n16462), .ZN(n16463) );
  OAI211_X1 U19654 ( .C1(n16465), .C2(n16498), .A(n16464), .B(n16463), .ZN(
        P2_U3005) );
  AOI22_X1 U19655 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19404), .B1(n16488), 
        .B2(n19251), .ZN(n16472) );
  NAND2_X1 U19656 ( .A1(n16466), .A2(n16494), .ZN(n16469) );
  NAND2_X1 U19657 ( .A1(n16467), .A2(n16493), .ZN(n16468) );
  OAI211_X1 U19658 ( .C1(n16486), .C2(n19257), .A(n16469), .B(n16468), .ZN(
        n16470) );
  INV_X1 U19659 ( .A(n16470), .ZN(n16471) );
  OAI211_X1 U19660 ( .C1(n16473), .C2(n16498), .A(n16472), .B(n16471), .ZN(
        P2_U3007) );
  OAI22_X1 U19661 ( .A1(n19968), .A2(n19254), .B1(n16475), .B2(n16474), .ZN(
        n16476) );
  AOI21_X1 U19662 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16477), .A(
        n16476), .ZN(n16484) );
  OAI22_X1 U19663 ( .A1(n16481), .A2(n16480), .B1(n16479), .B2(n16478), .ZN(
        n16482) );
  INV_X1 U19664 ( .A(n16482), .ZN(n16483) );
  OAI211_X1 U19665 ( .C1(n16486), .C2(n16485), .A(n16484), .B(n16483), .ZN(
        P2_U3008) );
  AOI22_X1 U19666 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19404), .B1(n16488), 
        .B2(n16487), .ZN(n16497) );
  INV_X1 U19667 ( .A(n16489), .ZN(n16495) );
  AOI222_X1 U19668 ( .A1(n16495), .A2(n16494), .B1(n16493), .B2(n16492), .C1(
        n16491), .C2(n16490), .ZN(n16496) );
  OAI211_X1 U19669 ( .C1(n16499), .C2(n16498), .A(n16497), .B(n16496), .ZN(
        P2_U3009) );
  AOI21_X1 U19670 ( .B1(n16516), .B2(n16502), .A(n16500), .ZN(n16505) );
  NOR2_X1 U19671 ( .A1(n20008), .A2(n19254), .ZN(n16504) );
  OAI22_X1 U19672 ( .A1(n16515), .A2(n16502), .B1(n16551), .B2(n16501), .ZN(
        n16503) );
  AOI211_X1 U19673 ( .C1(n16513), .C2(n16505), .A(n16504), .B(n16503), .ZN(
        n16511) );
  INV_X1 U19674 ( .A(n16506), .ZN(n16507) );
  OAI22_X1 U19675 ( .A1(n16508), .A2(n19419), .B1(n19411), .B2(n16507), .ZN(
        n16509) );
  INV_X1 U19676 ( .A(n16509), .ZN(n16510) );
  OAI211_X1 U19677 ( .C1(n16512), .C2(n19436), .A(n16511), .B(n16510), .ZN(
        P2_U3020) );
  INV_X1 U19678 ( .A(n16513), .ZN(n16517) );
  NAND2_X1 U19679 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19404), .ZN(n16514) );
  OAI221_X1 U19680 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16517), 
        .C1(n16516), .C2(n16515), .A(n16514), .ZN(n16518) );
  AOI21_X1 U19681 ( .B1(n16519), .B2(n19420), .A(n16518), .ZN(n16523) );
  AOI22_X1 U19682 ( .A1(n16521), .A2(n19414), .B1(n14475), .B2(n16520), .ZN(
        n16522) );
  OAI211_X1 U19683 ( .C1(n19419), .C2(n16524), .A(n16523), .B(n16522), .ZN(
        P2_U3021) );
  AOI22_X1 U19684 ( .A1(n16526), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n19420), .B2(n16525), .ZN(n16535) );
  AOI222_X1 U19685 ( .A1(n16529), .A2(n19414), .B1(n19429), .B2(n16528), .C1(
        n14475), .C2(n16527), .ZN(n16534) );
  NAND2_X1 U19686 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19404), .ZN(n16533) );
  OAI211_X1 U19687 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n16531), .B(n16530), .ZN(
        n16532) );
  NAND4_X1 U19688 ( .A1(n16535), .A2(n16534), .A3(n16533), .A4(n16532), .ZN(
        P2_U3023) );
  INV_X1 U19689 ( .A(n16536), .ZN(n19314) );
  AOI22_X1 U19690 ( .A1(n16537), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19420), .B2(n19314), .ZN(n16546) );
  AOI222_X1 U19691 ( .A1(n16540), .A2(n19414), .B1(n14475), .B2(n16539), .C1(
        n19429), .C2(n16538), .ZN(n16545) );
  NAND2_X1 U19692 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19404), .ZN(n16544) );
  OAI211_X1 U19693 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16542), .B(n16541), .ZN(
        n16543) );
  NAND4_X1 U19694 ( .A1(n16546), .A2(n16545), .A3(n16544), .A4(n16543), .ZN(
        P2_U3035) );
  OAI211_X1 U19695 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16548), .B(n16547), .ZN(n16550) );
  NAND2_X1 U19696 ( .A1(n19404), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16549) );
  OAI211_X1 U19697 ( .C1(n16551), .C2(n19249), .A(n16550), .B(n16549), .ZN(
        n16552) );
  AOI21_X1 U19698 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16553), .A(
        n16552), .ZN(n16557) );
  OAI22_X1 U19699 ( .A1(n16554), .A2(n19419), .B1(n19411), .B2(n19242), .ZN(
        n16555) );
  INV_X1 U19700 ( .A(n16555), .ZN(n16556) );
  OAI211_X1 U19701 ( .C1(n19436), .C2(n16558), .A(n16557), .B(n16556), .ZN(
        P2_U3038) );
  INV_X1 U19702 ( .A(n19103), .ZN(n16573) );
  AOI21_X1 U19703 ( .B1(n16561), .B2(n16560), .A(n16559), .ZN(n16572) );
  NOR2_X1 U19704 ( .A1(n16563), .A2(n16562), .ZN(n16564) );
  OAI22_X1 U19705 ( .A1(n16567), .A2(n19937), .B1(n16565), .B2(n16564), .ZN(
        n16566) );
  OAI21_X1 U19706 ( .B1(n16567), .B2(n11751), .A(n16566), .ZN(n16568) );
  AOI21_X1 U19707 ( .B1(n16570), .B2(n16569), .A(n16568), .ZN(n16571) );
  OAI211_X1 U19708 ( .C1(n19937), .C2(n16573), .A(n16572), .B(n16571), .ZN(
        P2_U3176) );
  NOR2_X1 U19709 ( .A1(n18002), .A2(n16574), .ZN(n16583) );
  INV_X1 U19710 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16596) );
  INV_X1 U19711 ( .A(n16575), .ZN(n16577) );
  OAI21_X1 U19712 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18002), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16576) );
  OAI221_X1 U19713 ( .B1(n16596), .B2(n16577), .C1(n18002), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n16576), .ZN(n16582) );
  OAI21_X1 U19714 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16596), .A(
        n16577), .ZN(n16580) );
  NAND2_X1 U19715 ( .A1(n18002), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16578) );
  OAI22_X1 U19716 ( .A1(n18002), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n16578), .B2(n16596), .ZN(n16579) );
  OAI21_X1 U19717 ( .B1(n16583), .B2(n16580), .A(n16579), .ZN(n16581) );
  OAI21_X1 U19718 ( .B1(n16583), .B2(n16582), .A(n16581), .ZN(n16632) );
  INV_X1 U19719 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19021) );
  NOR2_X1 U19720 ( .A1(n18426), .A2(n19021), .ZN(n16621) );
  NAND2_X1 U19721 ( .A1(n16584), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16586) );
  OR2_X1 U19722 ( .A1(n16586), .A2(n17891), .ZN(n16599) );
  XNOR2_X1 U19723 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16588) );
  NOR2_X1 U19724 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16585), .ZN(
        n16609) );
  NAND2_X1 U19725 ( .A1(n18815), .A2(n16586), .ZN(n16613) );
  OAI211_X1 U19726 ( .C1(n16587), .C2(n18104), .A(n18103), .B(n16613), .ZN(
        n16618) );
  NOR2_X1 U19727 ( .A1(n16609), .A2(n16618), .ZN(n16598) );
  OAI22_X1 U19728 ( .A1(n16599), .A2(n16588), .B1(n16598), .B2(n16779), .ZN(
        n16589) );
  AOI211_X1 U19729 ( .C1(n17952), .C2(n9807), .A(n16621), .B(n16589), .ZN(
        n16593) );
  INV_X1 U19730 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19043) );
  NAND3_X1 U19731 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n19043), .ZN(n16626) );
  OAI21_X1 U19732 ( .B1(n16596), .B2(n16595), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16590) );
  OAI21_X1 U19733 ( .B1(n16626), .B2(n16646), .A(n16590), .ZN(n16624) );
  OAI21_X1 U19734 ( .B1(n16596), .B2(n16594), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16591) );
  OAI21_X1 U19735 ( .B1(n16626), .B2(n16647), .A(n16591), .ZN(n16628) );
  AOI22_X1 U19736 ( .A1(n18012), .A2(n16624), .B1(n18040), .B2(n16628), .ZN(
        n16592) );
  OAI211_X1 U19737 ( .C1(n18015), .C2(n16632), .A(n16593), .B(n16592), .ZN(
        P3_U2799) );
  INV_X1 U19738 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16783) );
  XNOR2_X1 U19739 ( .A(n16783), .B(n16607), .ZN(n16782) );
  NAND2_X1 U19740 ( .A1(n18040), .A2(n16594), .ZN(n16620) );
  NAND2_X1 U19741 ( .A1(n18012), .A2(n16595), .ZN(n16614) );
  AOI21_X1 U19742 ( .B1(n16620), .B2(n16614), .A(n16596), .ZN(n16601) );
  NAND2_X1 U19743 ( .A1(n18416), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16597) );
  OAI221_X1 U19744 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16599), .C1(
        n16783), .C2(n16598), .A(n16597), .ZN(n16600) );
  AOI211_X1 U19745 ( .C1(n17952), .C2(n16782), .A(n16601), .B(n16600), .ZN(
        n16605) );
  INV_X1 U19746 ( .A(n17770), .ZN(n17812) );
  NAND4_X1 U19747 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16603), .A3(
        n17812), .A4(n16602), .ZN(n16604) );
  OAI211_X1 U19748 ( .C1(n16606), .C2(n18015), .A(n16605), .B(n16604), .ZN(
        P3_U2800) );
  AOI21_X1 U19749 ( .B1(n16794), .B2(n16608), .A(n16607), .ZN(n16793) );
  OAI21_X1 U19750 ( .B1(n16609), .B2(n17952), .A(n16793), .ZN(n16610) );
  OAI211_X1 U19751 ( .C1(n16613), .C2(n16612), .A(n16611), .B(n16610), .ZN(
        n16617) );
  AND2_X1 U19752 ( .A1(n16646), .A2(n16619), .ZN(n16615) );
  NOR2_X1 U19753 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18411), .ZN(
        n16622) );
  AOI221_X1 U19754 ( .B1(n16623), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), 
        .C1(n16622), .C2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n16621), .ZN(
        n16631) );
  INV_X1 U19755 ( .A(n16624), .ZN(n16627) );
  OAI22_X1 U19756 ( .A1(n16627), .A2(n18276), .B1(n16626), .B2(n16625), .ZN(
        n16629) );
  AOI22_X1 U19757 ( .A1(n18409), .A2(n16629), .B1(n18425), .B2(n16628), .ZN(
        n16630) );
  OAI211_X1 U19758 ( .C1(n18344), .C2(n16632), .A(n16631), .B(n16630), .ZN(
        P3_U2831) );
  INV_X1 U19759 ( .A(n18867), .ZN(n18401) );
  OAI22_X1 U19760 ( .A1(n18297), .A2(n18401), .B1(n18276), .B2(n18295), .ZN(
        n18212) );
  INV_X1 U19761 ( .A(n16633), .ZN(n16634) );
  NOR2_X1 U19762 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18878), .ZN(
        n18412) );
  NAND2_X1 U19763 ( .A1(n18900), .A2(n18898), .ZN(n18374) );
  NOR2_X1 U19764 ( .A1(n18412), .A2(n18394), .ZN(n18209) );
  AOI22_X1 U19765 ( .A1(n17797), .A2(n18212), .B1(n16634), .B2(n18209), .ZN(
        n16636) );
  NAND2_X1 U19766 ( .A1(n16636), .A2(n16635), .ZN(n18170) );
  NAND2_X1 U19767 ( .A1(n18409), .A2(n18170), .ZN(n18180) );
  OAI33_X1 U19768 ( .A1(n16638), .A2(n16637), .A3(n18180), .B1(n17969), .B2(
        n18420), .B3(n16642), .ZN(n16641) );
  AOI21_X1 U19769 ( .B1(n16641), .B2(n16640), .A(n16639), .ZN(n16656) );
  INV_X1 U19770 ( .A(n16642), .ZN(n16643) );
  OAI211_X1 U19771 ( .C1(n16645), .C2(n16644), .A(n17613), .B(n16643), .ZN(
        n16649) );
  AOI22_X1 U19772 ( .A1(n18867), .A2(n16647), .B1(n18296), .B2(n16646), .ZN(
        n16648) );
  OAI21_X1 U19773 ( .B1(n18873), .B2(n16649), .A(n16648), .ZN(n16650) );
  OAI211_X1 U19774 ( .C1(n16651), .C2(n16650), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18426), .ZN(n16655) );
  NAND3_X1 U19775 ( .A1(n16653), .A2(n18325), .A3(n16652), .ZN(n16654) );
  NAND3_X1 U19776 ( .A1(n16656), .A2(n16655), .A3(n16654), .ZN(P3_U2834) );
  NOR3_X1 U19777 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16658) );
  NOR4_X1 U19778 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16657) );
  INV_X2 U19779 ( .A(n16739), .ZN(U215) );
  NAND4_X1 U19780 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16658), .A3(n16657), .A4(
        U215), .ZN(U213) );
  INV_X1 U19781 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16741) );
  INV_X2 U19782 ( .A(U214), .ZN(n16702) );
  INV_X1 U19783 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16742) );
  OAI222_X1 U19784 ( .A1(U212), .A2(n16741), .B1(n16704), .B2(n20293), .C1(
        U214), .C2(n16742), .ZN(U216) );
  AOI22_X1 U19785 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16692), .ZN(n16660) );
  OAI21_X1 U19786 ( .B1(n14805), .B2(n16704), .A(n16660), .ZN(U217) );
  INV_X1 U19787 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20279) );
  AOI22_X1 U19788 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16692), .ZN(n16661) );
  OAI21_X1 U19789 ( .B1(n20279), .B2(n16704), .A(n16661), .ZN(U218) );
  AOI22_X1 U19790 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16692), .ZN(n16662) );
  OAI21_X1 U19791 ( .B1(n14815), .B2(n16704), .A(n16662), .ZN(U219) );
  INV_X1 U19792 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20266) );
  AOI22_X1 U19793 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16692), .ZN(n16663) );
  OAI21_X1 U19794 ( .B1(n20266), .B2(n16704), .A(n16663), .ZN(U220) );
  INV_X1 U19795 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20259) );
  AOI22_X1 U19796 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16692), .ZN(n16664) );
  OAI21_X1 U19797 ( .B1(n20259), .B2(n16704), .A(n16664), .ZN(U221) );
  AOI22_X1 U19798 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16692), .ZN(n16665) );
  OAI21_X1 U19799 ( .B1(n20253), .B2(n16704), .A(n16665), .ZN(U222) );
  AOI22_X1 U19800 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16692), .ZN(n16666) );
  OAI21_X1 U19801 ( .B1(n20235), .B2(n16704), .A(n16666), .ZN(U223) );
  INV_X1 U19802 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20290) );
  AOI22_X1 U19803 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16692), .ZN(n16667) );
  OAI21_X1 U19804 ( .B1(n20290), .B2(n16704), .A(n16667), .ZN(U224) );
  INV_X1 U19805 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20284) );
  AOI22_X1 U19806 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16692), .ZN(n16668) );
  OAI21_X1 U19807 ( .B1(n20284), .B2(n16704), .A(n16668), .ZN(U225) );
  AOI22_X1 U19808 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16692), .ZN(n16669) );
  OAI21_X1 U19809 ( .B1(n20277), .B2(n16704), .A(n16669), .ZN(U226) );
  INV_X1 U19810 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20273) );
  AOI22_X1 U19811 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16692), .ZN(n16670) );
  OAI21_X1 U19812 ( .B1(n20273), .B2(n16704), .A(n16670), .ZN(U227) );
  INV_X1 U19813 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20265) );
  AOI22_X1 U19814 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16692), .ZN(n16671) );
  OAI21_X1 U19815 ( .B1(n20265), .B2(n16704), .A(n16671), .ZN(U228) );
  INV_X1 U19816 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20258) );
  AOI22_X1 U19817 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16692), .ZN(n16672) );
  OAI21_X1 U19818 ( .B1(n20258), .B2(n16704), .A(n16672), .ZN(U229) );
  INV_X1 U19819 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20252) );
  AOI22_X1 U19820 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16692), .ZN(n16673) );
  OAI21_X1 U19821 ( .B1(n20252), .B2(n16704), .A(n16673), .ZN(U230) );
  INV_X1 U19822 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20231) );
  AOI22_X1 U19823 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16692), .ZN(n16674) );
  OAI21_X1 U19824 ( .B1(n20231), .B2(n16704), .A(n16674), .ZN(U231) );
  AOI22_X1 U19825 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16692), .ZN(n16675) );
  OAI21_X1 U19826 ( .B1(n12621), .B2(n16704), .A(n16675), .ZN(U232) );
  AOI22_X1 U19827 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16692), .ZN(n16676) );
  OAI21_X1 U19828 ( .B1(n16677), .B2(n16704), .A(n16676), .ZN(U233) );
  AOI22_X1 U19829 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16692), .ZN(n16678) );
  OAI21_X1 U19830 ( .B1(n16679), .B2(n16704), .A(n16678), .ZN(U234) );
  INV_X1 U19831 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16681) );
  AOI22_X1 U19832 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16692), .ZN(n16680) );
  OAI21_X1 U19833 ( .B1(n16681), .B2(n16704), .A(n16680), .ZN(U235) );
  AOI22_X1 U19834 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16692), .ZN(n16682) );
  OAI21_X1 U19835 ( .B1(n16683), .B2(n16704), .A(n16682), .ZN(U236) );
  AOI22_X1 U19836 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16692), .ZN(n16684) );
  OAI21_X1 U19837 ( .B1(n16685), .B2(n16704), .A(n16684), .ZN(U237) );
  AOI22_X1 U19838 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16692), .ZN(n16686) );
  OAI21_X1 U19839 ( .B1(n16687), .B2(n16704), .A(n16686), .ZN(U238) );
  AOI22_X1 U19840 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16692), .ZN(n16688) );
  OAI21_X1 U19841 ( .B1(n16689), .B2(n16704), .A(n16688), .ZN(U239) );
  INV_X1 U19842 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16691) );
  AOI22_X1 U19843 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16692), .ZN(n16690) );
  OAI21_X1 U19844 ( .B1(n16691), .B2(n16704), .A(n16690), .ZN(U240) );
  AOI22_X1 U19845 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16692), .ZN(n16693) );
  OAI21_X1 U19846 ( .B1(n12522), .B2(n16704), .A(n16693), .ZN(U241) );
  AOI22_X1 U19847 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16692), .ZN(n16694) );
  OAI21_X1 U19848 ( .B1(n12537), .B2(n16704), .A(n16694), .ZN(U242) );
  INV_X1 U19849 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16696) );
  AOI22_X1 U19850 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16692), .ZN(n16695) );
  OAI21_X1 U19851 ( .B1(n16696), .B2(n16704), .A(n16695), .ZN(U243) );
  AOI22_X1 U19852 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16692), .ZN(n16697) );
  OAI21_X1 U19853 ( .B1(n12516), .B2(n16704), .A(n16697), .ZN(U244) );
  INV_X1 U19854 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16699) );
  AOI22_X1 U19855 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16692), .ZN(n16698) );
  OAI21_X1 U19856 ( .B1(n16699), .B2(n16704), .A(n16698), .ZN(U245) );
  INV_X1 U19857 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16701) );
  AOI22_X1 U19858 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16692), .ZN(n16700) );
  OAI21_X1 U19859 ( .B1(n16701), .B2(n16704), .A(n16700), .ZN(U246) );
  INV_X1 U19860 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16705) );
  AOI22_X1 U19861 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16702), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16692), .ZN(n16703) );
  OAI21_X1 U19862 ( .B1(n16705), .B2(n16704), .A(n16703), .ZN(U247) );
  OAI22_X1 U19863 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16739), .ZN(n16706) );
  INV_X1 U19864 ( .A(n16706), .ZN(U251) );
  OAI22_X1 U19865 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16739), .ZN(n16707) );
  INV_X1 U19866 ( .A(n16707), .ZN(U252) );
  OAI22_X1 U19867 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16739), .ZN(n16708) );
  INV_X1 U19868 ( .A(n16708), .ZN(U253) );
  OAI22_X1 U19869 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16739), .ZN(n16709) );
  INV_X1 U19870 ( .A(n16709), .ZN(U254) );
  OAI22_X1 U19871 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16739), .ZN(n16710) );
  INV_X1 U19872 ( .A(n16710), .ZN(U255) );
  OAI22_X1 U19873 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16739), .ZN(n16711) );
  INV_X1 U19874 ( .A(n16711), .ZN(U256) );
  OAI22_X1 U19875 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16739), .ZN(n16712) );
  INV_X1 U19876 ( .A(n16712), .ZN(U257) );
  OAI22_X1 U19877 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16739), .ZN(n16713) );
  INV_X1 U19878 ( .A(n16713), .ZN(U258) );
  OAI22_X1 U19879 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16739), .ZN(n16714) );
  INV_X1 U19880 ( .A(n16714), .ZN(U259) );
  OAI22_X1 U19881 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16733), .ZN(n16715) );
  INV_X1 U19882 ( .A(n16715), .ZN(U260) );
  OAI22_X1 U19883 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16733), .ZN(n16716) );
  INV_X1 U19884 ( .A(n16716), .ZN(U261) );
  OAI22_X1 U19885 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16739), .ZN(n16717) );
  INV_X1 U19886 ( .A(n16717), .ZN(U262) );
  OAI22_X1 U19887 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16739), .ZN(n16718) );
  INV_X1 U19888 ( .A(n16718), .ZN(U263) );
  OAI22_X1 U19889 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16739), .ZN(n16719) );
  INV_X1 U19890 ( .A(n16719), .ZN(U264) );
  OAI22_X1 U19891 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16739), .ZN(n16720) );
  INV_X1 U19892 ( .A(n16720), .ZN(U265) );
  OAI22_X1 U19893 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16733), .ZN(n16721) );
  INV_X1 U19894 ( .A(n16721), .ZN(U266) );
  OAI22_X1 U19895 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16733), .ZN(n16722) );
  INV_X1 U19896 ( .A(n16722), .ZN(U267) );
  OAI22_X1 U19897 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16733), .ZN(n16723) );
  INV_X1 U19898 ( .A(n16723), .ZN(U268) );
  OAI22_X1 U19899 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16733), .ZN(n16724) );
  INV_X1 U19900 ( .A(n16724), .ZN(U269) );
  OAI22_X1 U19901 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16733), .ZN(n16725) );
  INV_X1 U19902 ( .A(n16725), .ZN(U270) );
  OAI22_X1 U19903 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16733), .ZN(n16726) );
  INV_X1 U19904 ( .A(n16726), .ZN(U271) );
  OAI22_X1 U19905 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16739), .ZN(n16727) );
  INV_X1 U19906 ( .A(n16727), .ZN(U272) );
  OAI22_X1 U19907 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16739), .ZN(n16728) );
  INV_X1 U19908 ( .A(n16728), .ZN(U273) );
  OAI22_X1 U19909 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16733), .ZN(n16729) );
  INV_X1 U19910 ( .A(n16729), .ZN(U274) );
  OAI22_X1 U19911 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16739), .ZN(n16730) );
  INV_X1 U19912 ( .A(n16730), .ZN(U275) );
  OAI22_X1 U19913 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16739), .ZN(n16731) );
  INV_X1 U19914 ( .A(n16731), .ZN(U276) );
  OAI22_X1 U19915 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16739), .ZN(n16732) );
  INV_X1 U19916 ( .A(n16732), .ZN(U277) );
  OAI22_X1 U19917 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16733), .ZN(n16734) );
  INV_X1 U19918 ( .A(n16734), .ZN(U278) );
  OAI22_X1 U19919 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16739), .ZN(n16735) );
  INV_X1 U19920 ( .A(n16735), .ZN(U279) );
  OAI22_X1 U19921 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16739), .ZN(n16736) );
  INV_X1 U19922 ( .A(n16736), .ZN(U280) );
  OAI22_X1 U19923 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16739), .ZN(n16738) );
  INV_X1 U19924 ( .A(n16738), .ZN(U281) );
  INV_X1 U19925 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19457) );
  AOI22_X1 U19926 ( .A1(n16739), .A2(n16741), .B1(n19457), .B2(U215), .ZN(U282) );
  INV_X1 U19927 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16740) );
  AOI222_X1 U19928 ( .A1(n16742), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16741), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16740), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16743) );
  INV_X2 U19929 ( .A(n16745), .ZN(n16744) );
  INV_X1 U19930 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18979) );
  INV_X1 U19931 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19977) );
  AOI22_X1 U19932 ( .A1(n16744), .A2(n18979), .B1(n19977), .B2(n16745), .ZN(
        U347) );
  INV_X1 U19933 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18977) );
  INV_X1 U19934 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19975) );
  AOI22_X1 U19935 ( .A1(n16744), .A2(n18977), .B1(n19975), .B2(n16745), .ZN(
        U348) );
  INV_X1 U19936 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18974) );
  INV_X1 U19937 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19973) );
  AOI22_X1 U19938 ( .A1(n16744), .A2(n18974), .B1(n19973), .B2(n16745), .ZN(
        U349) );
  INV_X1 U19939 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18973) );
  INV_X1 U19940 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19971) );
  AOI22_X1 U19941 ( .A1(n16744), .A2(n18973), .B1(n19971), .B2(n16745), .ZN(
        U350) );
  INV_X1 U19942 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18971) );
  INV_X1 U19943 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19969) );
  AOI22_X1 U19944 ( .A1(n16744), .A2(n18971), .B1(n19969), .B2(n16745), .ZN(
        U351) );
  INV_X1 U19945 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18969) );
  INV_X1 U19946 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19967) );
  AOI22_X1 U19947 ( .A1(n16744), .A2(n18969), .B1(n19967), .B2(n16745), .ZN(
        U352) );
  INV_X1 U19948 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18967) );
  INV_X1 U19949 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19965) );
  AOI22_X1 U19950 ( .A1(n16744), .A2(n18967), .B1(n19965), .B2(n16745), .ZN(
        U353) );
  INV_X1 U19951 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18965) );
  AOI22_X1 U19952 ( .A1(n16744), .A2(n18965), .B1(n19962), .B2(n16745), .ZN(
        U354) );
  INV_X1 U19953 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19017) );
  INV_X1 U19954 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20016) );
  AOI22_X1 U19955 ( .A1(n16744), .A2(n19017), .B1(n20016), .B2(n16745), .ZN(
        U356) );
  INV_X1 U19956 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19015) );
  INV_X1 U19957 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20013) );
  AOI22_X1 U19958 ( .A1(n16744), .A2(n19015), .B1(n20013), .B2(n16745), .ZN(
        U357) );
  INV_X1 U19959 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19012) );
  INV_X1 U19960 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20010) );
  AOI22_X1 U19961 ( .A1(n16744), .A2(n19012), .B1(n20010), .B2(n16745), .ZN(
        U358) );
  INV_X1 U19962 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19011) );
  INV_X1 U19963 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20009) );
  AOI22_X1 U19964 ( .A1(n16744), .A2(n19011), .B1(n20009), .B2(n16745), .ZN(
        U359) );
  INV_X1 U19965 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19009) );
  INV_X1 U19966 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20007) );
  AOI22_X1 U19967 ( .A1(n16744), .A2(n19009), .B1(n20007), .B2(n16745), .ZN(
        U360) );
  INV_X1 U19968 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19007) );
  INV_X1 U19969 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20005) );
  AOI22_X1 U19970 ( .A1(n16744), .A2(n19007), .B1(n20005), .B2(n16745), .ZN(
        U361) );
  INV_X1 U19971 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19005) );
  INV_X1 U19972 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20003) );
  AOI22_X1 U19973 ( .A1(n16744), .A2(n19005), .B1(n20003), .B2(n16745), .ZN(
        U362) );
  INV_X1 U19974 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19003) );
  INV_X1 U19975 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20001) );
  AOI22_X1 U19976 ( .A1(n16744), .A2(n19003), .B1(n20001), .B2(n16745), .ZN(
        U363) );
  INV_X1 U19977 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19001) );
  INV_X1 U19978 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19999) );
  AOI22_X1 U19979 ( .A1(n16744), .A2(n19001), .B1(n19999), .B2(n16745), .ZN(
        U364) );
  INV_X1 U19980 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18962) );
  INV_X1 U19981 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19960) );
  AOI22_X1 U19982 ( .A1(n16744), .A2(n18962), .B1(n19960), .B2(n16745), .ZN(
        U365) );
  INV_X1 U19983 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18998) );
  INV_X1 U19984 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19997) );
  AOI22_X1 U19985 ( .A1(n16744), .A2(n18998), .B1(n19997), .B2(n16745), .ZN(
        U366) );
  INV_X1 U19986 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18997) );
  INV_X1 U19987 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19995) );
  AOI22_X1 U19988 ( .A1(n16744), .A2(n18997), .B1(n19995), .B2(n16745), .ZN(
        U367) );
  INV_X1 U19989 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18995) );
  INV_X1 U19990 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19993) );
  AOI22_X1 U19991 ( .A1(n16744), .A2(n18995), .B1(n19993), .B2(n16745), .ZN(
        U368) );
  INV_X1 U19992 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18993) );
  INV_X1 U19993 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19991) );
  AOI22_X1 U19994 ( .A1(n16744), .A2(n18993), .B1(n19991), .B2(n16745), .ZN(
        U369) );
  INV_X1 U19995 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18991) );
  INV_X1 U19996 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19989) );
  AOI22_X1 U19997 ( .A1(n16744), .A2(n18991), .B1(n19989), .B2(n16745), .ZN(
        U370) );
  INV_X1 U19998 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18989) );
  INV_X1 U19999 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19987) );
  AOI22_X1 U20000 ( .A1(n16744), .A2(n18989), .B1(n19987), .B2(n16745), .ZN(
        U371) );
  INV_X1 U20001 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18986) );
  INV_X1 U20002 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19985) );
  AOI22_X1 U20003 ( .A1(n16744), .A2(n18986), .B1(n19985), .B2(n16745), .ZN(
        U372) );
  INV_X1 U20004 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18985) );
  INV_X1 U20005 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19983) );
  AOI22_X1 U20006 ( .A1(n16744), .A2(n18985), .B1(n19983), .B2(n16745), .ZN(
        U373) );
  INV_X1 U20007 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18983) );
  INV_X1 U20008 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U20009 ( .A1(n16744), .A2(n18983), .B1(n19981), .B2(n16745), .ZN(
        U374) );
  INV_X1 U20010 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18981) );
  INV_X1 U20011 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19979) );
  AOI22_X1 U20012 ( .A1(n16744), .A2(n18981), .B1(n19979), .B2(n16745), .ZN(
        U375) );
  INV_X1 U20013 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18960) );
  INV_X1 U20014 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19959) );
  AOI22_X1 U20015 ( .A1(n16744), .A2(n18960), .B1(n19959), .B2(n16745), .ZN(
        U376) );
  INV_X1 U20016 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18957) );
  NOR2_X1 U20017 ( .A1(n18944), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18949) );
  OAI22_X1 U20018 ( .A1(n18957), .A2(n18949), .B1(n18944), .B2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18942) );
  INV_X1 U20019 ( .A(n18942), .ZN(n19031) );
  AOI21_X1 U20020 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19031), .ZN(n16746) );
  INV_X1 U20021 ( .A(n16746), .ZN(P3_U2633) );
  NAND2_X1 U20022 ( .A1(n19034), .A2(n18931), .ZN(n16748) );
  OAI21_X1 U20023 ( .B1(n16752), .B2(n17683), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16747) );
  OAI21_X1 U20024 ( .B1(n16748), .B2(n18935), .A(n16747), .ZN(P3_U2634) );
  INV_X1 U20025 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18959) );
  AOI21_X1 U20026 ( .B1(n18957), .B2(n18959), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16749) );
  AOI22_X1 U20027 ( .A1(n19026), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16749), 
        .B2(n19093), .ZN(P3_U2635) );
  OAI21_X1 U20028 ( .B1(n18945), .B2(BS16), .A(n19031), .ZN(n19029) );
  OAI21_X1 U20029 ( .B1(n19031), .B2(n19083), .A(n19029), .ZN(P3_U2636) );
  NOR3_X1 U20030 ( .A1(n16752), .A2(n16751), .A3(n16750), .ZN(n18874) );
  NOR2_X1 U20031 ( .A1(n18874), .A2(n18929), .ZN(n19076) );
  OAI21_X1 U20032 ( .B1(n19076), .B2(n18432), .A(n16753), .ZN(P3_U2637) );
  NOR4_X1 U20033 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16757) );
  NOR4_X1 U20034 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16756) );
  NOR4_X1 U20035 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16755) );
  NOR4_X1 U20036 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16754) );
  NAND4_X1 U20037 ( .A1(n16757), .A2(n16756), .A3(n16755), .A4(n16754), .ZN(
        n16763) );
  NOR4_X1 U20038 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16761) );
  AOI211_X1 U20039 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16760) );
  NOR4_X1 U20040 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16759) );
  NOR4_X1 U20041 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16758) );
  NAND4_X1 U20042 ( .A1(n16761), .A2(n16760), .A3(n16759), .A4(n16758), .ZN(
        n16762) );
  NOR2_X1 U20043 ( .A1(n16763), .A2(n16762), .ZN(n19070) );
  INV_X1 U20044 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16765) );
  NOR3_X1 U20045 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16766) );
  OAI21_X1 U20046 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16766), .A(n19070), .ZN(
        n16764) );
  OAI21_X1 U20047 ( .B1(n19070), .B2(n16765), .A(n16764), .ZN(P3_U2638) );
  INV_X1 U20048 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19030) );
  AOI21_X1 U20049 ( .B1(n19066), .B2(n19030), .A(n16766), .ZN(n16768) );
  INV_X1 U20050 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16767) );
  INV_X1 U20051 ( .A(n19070), .ZN(n19073) );
  AOI22_X1 U20052 ( .A1(n19070), .A2(n16768), .B1(n16767), .B2(n19073), .ZN(
        P3_U2639) );
  INV_X1 U20053 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19018) );
  NOR2_X1 U20054 ( .A1(n19010), .A2(n16769), .ZN(n16813) );
  NAND4_X1 U20055 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16813), .ZN(n16775) );
  NOR3_X1 U20056 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19018), .A3(n16775), 
        .ZN(n16770) );
  AOI21_X1 U20057 ( .B1(n17136), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16770), .ZN(
        n16778) );
  INV_X1 U20058 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16821) );
  NAND2_X1 U20059 ( .A1(n16822), .A2(n16821), .ZN(n16820) );
  NOR2_X1 U20060 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16820), .ZN(n16803) );
  INV_X1 U20061 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17147) );
  NAND2_X1 U20062 ( .A1(n16803), .A2(n17147), .ZN(n16780) );
  NOR2_X1 U20063 ( .A1(n17139), .A2(n16780), .ZN(n16787) );
  INV_X1 U20064 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17152) );
  OAI21_X1 U20065 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16772), .A(
        n16771), .ZN(n17762) );
  INV_X1 U20066 ( .A(n17762), .ZN(n16816) );
  NOR2_X1 U20067 ( .A1(n16773), .A2(n17116), .ZN(n16815) );
  NOR2_X1 U20068 ( .A1(n16816), .A2(n16815), .ZN(n16814) );
  NOR2_X1 U20069 ( .A1(n16814), .A2(n17116), .ZN(n16805) );
  NOR2_X1 U20070 ( .A1(n16806), .A2(n16805), .ZN(n16804) );
  NOR2_X1 U20071 ( .A1(n16804), .A2(n17116), .ZN(n16792) );
  NAND2_X1 U20072 ( .A1(n9807), .A2(n17084), .ZN(n17049) );
  NAND2_X1 U20073 ( .A1(n17143), .A2(n17132), .ZN(n17141) );
  NAND3_X1 U20074 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16774) );
  AOI21_X1 U20075 ( .B1(n17141), .B2(n16774), .A(n16819), .ZN(n16802) );
  NOR2_X1 U20076 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16775), .ZN(n16785) );
  INV_X1 U20077 ( .A(n16785), .ZN(n16776) );
  AOI21_X1 U20078 ( .B1(n16802), .B2(n16776), .A(n19021), .ZN(n16777) );
  NAND2_X1 U20079 ( .A1(n17110), .A2(n16780), .ZN(n16798) );
  XOR2_X1 U20080 ( .A(n16782), .B(n16781), .Z(n16786) );
  OAI22_X1 U20081 ( .A1(n16802), .A2(n19018), .B1(n16783), .B2(n17127), .ZN(
        n16784) );
  AOI211_X1 U20082 ( .C1(n16786), .C2(n17084), .A(n16785), .B(n16784), .ZN(
        n16789) );
  OAI21_X1 U20083 ( .B1(n17136), .B2(n16787), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16788) );
  OAI211_X1 U20084 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16798), .A(n16789), .B(
        n16788), .ZN(P3_U2641) );
  INV_X1 U20085 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19016) );
  INV_X1 U20086 ( .A(n16790), .ZN(n16791) );
  AOI211_X1 U20087 ( .C1(n16793), .C2(n16792), .A(n16791), .B(n18938), .ZN(
        n16797) );
  NAND3_X1 U20088 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16813), .ZN(n16795) );
  OAI22_X1 U20089 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16795), .B1(n16794), 
        .B2(n17127), .ZN(n16796) );
  AOI211_X1 U20090 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17136), .A(n16797), .B(
        n16796), .ZN(n16801) );
  INV_X1 U20091 ( .A(n16798), .ZN(n16799) );
  OAI21_X1 U20092 ( .B1(n16803), .B2(n17147), .A(n16799), .ZN(n16800) );
  OAI211_X1 U20093 ( .C1(n16802), .C2(n19016), .A(n16801), .B(n16800), .ZN(
        P3_U2642) );
  AOI22_X1 U20094 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16819), .B1(n17136), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16811) );
  INV_X1 U20095 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19013) );
  INV_X1 U20096 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19014) );
  AOI22_X1 U20097 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .B1(n19013), .B2(n19014), .ZN(n16809) );
  AOI211_X1 U20098 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16820), .A(n16803), .B(
        n17139), .ZN(n16808) );
  AOI211_X1 U20099 ( .C1(n16806), .C2(n16805), .A(n16804), .B(n18938), .ZN(
        n16807) );
  AOI211_X1 U20100 ( .C1(n16813), .C2(n16809), .A(n16808), .B(n16807), .ZN(
        n16810) );
  OAI211_X1 U20101 ( .C1(n16812), .C2(n17127), .A(n16811), .B(n16810), .ZN(
        P3_U2643) );
  INV_X1 U20102 ( .A(n16813), .ZN(n16825) );
  AOI211_X1 U20103 ( .C1(n16816), .C2(n16815), .A(n16814), .B(n18938), .ZN(
        n16818) );
  OAI22_X1 U20104 ( .A1(n17758), .A2(n17127), .B1(n17140), .B2(n16821), .ZN(
        n16817) );
  AOI211_X1 U20105 ( .C1(n16819), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16818), 
        .B(n16817), .ZN(n16824) );
  OAI211_X1 U20106 ( .C1(n16822), .C2(n16821), .A(n17110), .B(n16820), .ZN(
        n16823) );
  OAI211_X1 U20107 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16825), .A(n16824), 
        .B(n16823), .ZN(P3_U2644) );
  INV_X1 U20108 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17782) );
  OAI21_X1 U20109 ( .B1(n17132), .B2(n16845), .A(n17143), .ZN(n16826) );
  INV_X1 U20110 ( .A(n16826), .ZN(n16859) );
  OAI21_X1 U20111 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n17132), .A(n16859), 
        .ZN(n16834) );
  AOI211_X1 U20112 ( .C1(n16829), .C2(n16828), .A(n16827), .B(n18938), .ZN(
        n16833) );
  NAND2_X1 U20113 ( .A1(n17121), .A2(n19008), .ZN(n16830) );
  OAI22_X1 U20114 ( .A1(n17140), .A2(n16836), .B1(n16831), .B2(n16830), .ZN(
        n16832) );
  AOI211_X1 U20115 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16834), .A(n16833), 
        .B(n16832), .ZN(n16838) );
  OAI211_X1 U20116 ( .C1(n16842), .C2(n16836), .A(n17110), .B(n16835), .ZN(
        n16837) );
  OAI211_X1 U20117 ( .C1(n17127), .C2(n17782), .A(n16838), .B(n16837), .ZN(
        P3_U2646) );
  INV_X1 U20118 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19006) );
  AOI22_X1 U20119 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17092), .B1(
        n17136), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16848) );
  NOR2_X1 U20120 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17132), .ZN(n16846) );
  INV_X1 U20121 ( .A(n16839), .ZN(n16840) );
  AOI211_X1 U20122 ( .C1(n17793), .C2(n16841), .A(n16840), .B(n18938), .ZN(
        n16844) );
  AOI211_X1 U20123 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16850), .A(n16842), .B(
        n17139), .ZN(n16843) );
  AOI211_X1 U20124 ( .C1(n16846), .C2(n16845), .A(n16844), .B(n16843), .ZN(
        n16847) );
  OAI211_X1 U20125 ( .C1(n19006), .C2(n16859), .A(n16848), .B(n16847), .ZN(
        P3_U2647) );
  AOI21_X1 U20126 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n16849), .A(n17139), .ZN(
        n16851) );
  AOI22_X1 U20127 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17092), .B1(
        n16851), .B2(n16850), .ZN(n16858) );
  AOI211_X1 U20128 ( .C1(n17804), .C2(n16853), .A(n16852), .B(n18938), .ZN(
        n16856) );
  NOR4_X1 U20129 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17132), .A3(n16866), 
        .A4(n16854), .ZN(n16855) );
  AOI211_X1 U20130 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n17136), .A(n16856), .B(
        n16855), .ZN(n16857) );
  OAI211_X1 U20131 ( .C1(n19004), .C2(n16859), .A(n16858), .B(n16857), .ZN(
        P3_U2648) );
  NOR3_X1 U20132 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16866), .A3(n17132), 
        .ZN(n16860) );
  AOI22_X1 U20133 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17092), .B1(
        P3_REIP_REG_21__SCAN_IN), .B2(n16860), .ZN(n16869) );
  AOI211_X1 U20134 ( .C1(n17823), .C2(n16862), .A(n16861), .B(n18938), .ZN(
        n16865) );
  AOI211_X1 U20135 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16871), .A(n16863), .B(
        n17139), .ZN(n16864) );
  AOI211_X1 U20136 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17136), .A(n16865), .B(
        n16864), .ZN(n16868) );
  AOI21_X1 U20137 ( .B1(n16866), .B2(n17121), .A(n17073), .ZN(n16880) );
  INV_X1 U20138 ( .A(n16880), .ZN(n16885) );
  NOR3_X1 U20139 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16866), .A3(n17132), 
        .ZN(n16877) );
  OAI21_X1 U20140 ( .B1(n16885), .B2(n16877), .A(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n16867) );
  NAND3_X1 U20141 ( .A1(n16869), .A2(n16868), .A3(n16867), .ZN(P3_U2649) );
  INV_X1 U20142 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19000) );
  OAI21_X1 U20143 ( .B1(n17241), .B2(n16881), .A(n17110), .ZN(n16870) );
  INV_X1 U20144 ( .A(n16870), .ZN(n16872) );
  AOI22_X1 U20145 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17092), .B1(
        n16872), .B2(n16871), .ZN(n16879) );
  INV_X1 U20146 ( .A(n16873), .ZN(n16874) );
  AOI211_X1 U20147 ( .C1(n17837), .C2(n16875), .A(n16874), .B(n18938), .ZN(
        n16876) );
  AOI211_X1 U20148 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n17136), .A(n16877), .B(
        n16876), .ZN(n16878) );
  OAI211_X1 U20149 ( .C1(n19000), .C2(n16880), .A(n16879), .B(n16878), .ZN(
        P3_U2650) );
  AOI211_X1 U20150 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16902), .A(n16881), .B(
        n17139), .ZN(n16884) );
  AOI211_X1 U20151 ( .C1(n17846), .C2(n16895), .A(n16882), .B(n18938), .ZN(
        n16883) );
  AOI211_X1 U20152 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17136), .A(n16884), .B(
        n16883), .ZN(n16888) );
  NAND2_X1 U20153 ( .A1(n17121), .A2(n16889), .ZN(n16952) );
  INV_X1 U20154 ( .A(n16952), .ZN(n16938) );
  OAI221_X1 U20155 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n16886), .C1(
        P3_REIP_REG_20__SCAN_IN), .C2(n16938), .A(n16885), .ZN(n16887) );
  OAI211_X1 U20156 ( .C1(n17127), .C2(n17841), .A(n16888), .B(n16887), .ZN(
        P3_U2651) );
  INV_X1 U20157 ( .A(n16891), .ZN(n16890) );
  NAND2_X1 U20158 ( .A1(n16889), .A2(n17143), .ZN(n16955) );
  OAI21_X1 U20159 ( .B1(n16890), .B2(n16955), .A(n17141), .ZN(n16918) );
  INV_X1 U20160 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18994) );
  NAND3_X1 U20161 ( .A1(n16891), .A2(n16938), .A3(n18994), .ZN(n16912) );
  AOI21_X1 U20162 ( .B1(n16918), .B2(n16912), .A(n18996), .ZN(n16901) );
  NOR3_X1 U20163 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16892), .A3(n16952), 
        .ZN(n16900) );
  NOR3_X1 U20164 ( .A1(n18097), .A2(n17879), .A3(n16927), .ZN(n17856) );
  NAND2_X1 U20165 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17856), .ZN(
        n16906) );
  INV_X1 U20166 ( .A(n16906), .ZN(n16894) );
  OAI21_X1 U20167 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16894), .A(
        n16893), .ZN(n17860) );
  AOI211_X1 U20168 ( .C1(n16894), .C2(n16914), .A(n17116), .B(n17860), .ZN(
        n16898) );
  INV_X1 U20169 ( .A(n17860), .ZN(n16896) );
  OAI21_X1 U20170 ( .B1(n16896), .B2(n16895), .A(n17084), .ZN(n16897) );
  INV_X1 U20171 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17858) );
  OAI22_X1 U20172 ( .A1(n16898), .A2(n16897), .B1(n17858), .B2(n17127), .ZN(
        n16899) );
  NOR4_X1 U20173 ( .A1(n18416), .A2(n16901), .A3(n16900), .A4(n16899), .ZN(
        n16904) );
  OAI211_X1 U20174 ( .C1(n16905), .C2(n17273), .A(n17110), .B(n16902), .ZN(
        n16903) );
  OAI211_X1 U20175 ( .C1(n17273), .C2(n17140), .A(n16904), .B(n16903), .ZN(
        P3_U2652) );
  AOI211_X1 U20176 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16923), .A(n16905), .B(
        n17139), .ZN(n16911) );
  OAI21_X1 U20177 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17856), .A(
        n16906), .ZN(n17870) );
  INV_X1 U20178 ( .A(n16914), .ZN(n16945) );
  INV_X1 U20179 ( .A(n17856), .ZN(n16915) );
  OAI21_X1 U20180 ( .B1(n16945), .B2(n16915), .A(n9807), .ZN(n16908) );
  AOI21_X1 U20181 ( .B1(n17870), .B2(n16908), .A(n18938), .ZN(n16907) );
  OAI21_X1 U20182 ( .B1(n17870), .B2(n16908), .A(n16907), .ZN(n16909) );
  OAI211_X1 U20183 ( .C1(n17140), .C2(n17291), .A(n18426), .B(n16909), .ZN(
        n16910) );
  AOI211_X1 U20184 ( .C1(n17092), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16911), .B(n16910), .ZN(n16913) );
  OAI211_X1 U20185 ( .C1(n16918), .C2(n18994), .A(n16913), .B(n16912), .ZN(
        P3_U2653) );
  AOI21_X1 U20186 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16914), .A(
        n17116), .ZN(n16916) );
  NOR2_X1 U20187 ( .A1(n18097), .A2(n17879), .ZN(n16929) );
  OAI21_X1 U20188 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16929), .A(
        n16915), .ZN(n17883) );
  XOR2_X1 U20189 ( .A(n16916), .B(n17883), .Z(n16917) );
  OAI21_X1 U20190 ( .B1(n18938), .B2(n16917), .A(n18426), .ZN(n16922) );
  NOR2_X1 U20191 ( .A1(n16937), .A2(n16952), .ZN(n16920) );
  INV_X1 U20192 ( .A(n16918), .ZN(n16919) );
  MUX2_X1 U20193 ( .A(n16920), .B(n16919), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n16921) );
  AOI211_X1 U20194 ( .C1(n17136), .C2(P3_EBX_REG_17__SCAN_IN), .A(n16922), .B(
        n16921), .ZN(n16926) );
  OAI211_X1 U20195 ( .C1(n16928), .C2(n16924), .A(n17110), .B(n16923), .ZN(
        n16925) );
  OAI211_X1 U20196 ( .C1(n17127), .C2(n16927), .A(n16926), .B(n16925), .ZN(
        P3_U2654) );
  NAND2_X1 U20197 ( .A1(n17141), .A2(n16955), .ZN(n16963) );
  INV_X1 U20198 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18990) );
  AOI211_X1 U20199 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16943), .A(n16928), .B(
        n17139), .ZN(n16936) );
  NAND2_X1 U20200 ( .A1(n16945), .A2(n9807), .ZN(n16930) );
  INV_X1 U20201 ( .A(n16930), .ZN(n16932) );
  INV_X1 U20202 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16933) );
  AOI21_X1 U20203 ( .B1(n16933), .B2(n16941), .A(n16929), .ZN(n16931) );
  INV_X1 U20204 ( .A(n16931), .ZN(n17895) );
  AOI221_X1 U20205 ( .B1(n16932), .B2(n16931), .C1(n16930), .C2(n17895), .A(
        n18938), .ZN(n16935) );
  INV_X1 U20206 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17294) );
  OAI22_X1 U20207 ( .A1(n16933), .A2(n17127), .B1(n17140), .B2(n17294), .ZN(
        n16934) );
  NOR4_X1 U20208 ( .A1(n18416), .A2(n16936), .A3(n16935), .A4(n16934), .ZN(
        n16940) );
  OAI211_X1 U20209 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16938), .B(n16937), .ZN(n16939) );
  OAI211_X1 U20210 ( .C1(n16963), .C2(n18990), .A(n16940), .B(n16939), .ZN(
        P3_U2655) );
  INV_X1 U20211 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18988) );
  OAI21_X1 U20212 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17890), .A(
        n16941), .ZN(n17915) );
  NAND2_X1 U20213 ( .A1(n9807), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17128) );
  NAND2_X1 U20214 ( .A1(n17084), .A2(n17128), .ZN(n17129) );
  AOI211_X1 U20215 ( .C1(n9807), .C2(n16942), .A(n17915), .B(n17129), .ZN(
        n16950) );
  INV_X1 U20216 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17905) );
  OAI211_X1 U20217 ( .C1(n16958), .C2(n16947), .A(n17110), .B(n16943), .ZN(
        n16944) );
  OAI21_X1 U20218 ( .B1(n17127), .B2(n17905), .A(n16944), .ZN(n16949) );
  NAND2_X1 U20219 ( .A1(n16945), .A2(n17915), .ZN(n16946) );
  OAI22_X1 U20220 ( .A1(n17140), .A2(n16947), .B1(n17049), .B2(n16946), .ZN(
        n16948) );
  NOR4_X1 U20221 ( .A1(n18416), .A2(n16950), .A3(n16949), .A4(n16948), .ZN(
        n16951) );
  OAI221_X1 U20222 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16952), .C1(n18988), 
        .C2(n16963), .A(n16951), .ZN(P3_U2656) );
  OR2_X1 U20223 ( .A1(n18097), .A2(n17921), .ZN(n16964) );
  AOI21_X1 U20224 ( .B1(n17920), .B2(n16964), .A(n17890), .ZN(n17923) );
  NAND3_X1 U20225 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17961), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16992) );
  NOR2_X1 U20226 ( .A1(n17934), .A2(n16992), .ZN(n17937) );
  INV_X1 U20227 ( .A(n17937), .ZN(n16980) );
  OAI21_X1 U20228 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16980), .A(
        n9807), .ZN(n16982) );
  OAI21_X1 U20229 ( .B1(n10426), .B2(n17116), .A(n16982), .ZN(n16974) );
  OAI21_X1 U20230 ( .B1(n17923), .B2(n16974), .A(n17084), .ZN(n16953) );
  AOI21_X1 U20231 ( .B1(n17923), .B2(n16974), .A(n16953), .ZN(n16954) );
  AOI211_X1 U20232 ( .C1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n17092), .A(
        n18308), .B(n16954), .ZN(n16962) );
  INV_X1 U20233 ( .A(n16955), .ZN(n16957) );
  NOR3_X1 U20234 ( .A1(n16957), .A2(n16956), .A3(n17132), .ZN(n16960) );
  AOI211_X1 U20235 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16972), .A(n16958), .B(
        n17139), .ZN(n16959) );
  AOI211_X1 U20236 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17136), .A(n16960), .B(
        n16959), .ZN(n16961) );
  OAI211_X1 U20237 ( .C1(n18987), .C2(n16963), .A(n16962), .B(n16961), .ZN(
        P3_U2657) );
  NOR2_X1 U20238 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17132), .ZN(n16967) );
  NAND2_X1 U20239 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17937), .ZN(
        n16965) );
  INV_X1 U20240 ( .A(n16965), .ZN(n16979) );
  OAI21_X1 U20241 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16979), .A(
        n16964), .ZN(n17939) );
  AOI211_X1 U20242 ( .C1(n9807), .C2(n16965), .A(n17939), .B(n17129), .ZN(
        n16966) );
  AOI211_X1 U20243 ( .C1(n16968), .C2(n16967), .A(n18308), .B(n16966), .ZN(
        n16978) );
  NOR2_X1 U20244 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17132), .ZN(n16986) );
  INV_X1 U20245 ( .A(n16969), .ZN(n16987) );
  OAI21_X1 U20246 ( .B1(n16987), .B2(n17132), .A(n17143), .ZN(n16998) );
  INV_X1 U20247 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16970) );
  OAI22_X1 U20248 ( .A1(n16970), .A2(n17127), .B1(n17140), .B2(n16973), .ZN(
        n16971) );
  AOI221_X1 U20249 ( .B1(n16986), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n16998), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n16971), .ZN(n16977) );
  OAI211_X1 U20250 ( .C1(n16983), .C2(n16973), .A(n17110), .B(n16972), .ZN(
        n16976) );
  NAND3_X1 U20251 ( .A1(n17084), .A2(n17939), .A3(n16974), .ZN(n16975) );
  NAND4_X1 U20252 ( .A1(n16978), .A2(n16977), .A3(n16976), .A4(n16975), .ZN(
        P3_U2658) );
  INV_X1 U20253 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16981) );
  AOI21_X1 U20254 ( .B1(n16981), .B2(n16980), .A(n16979), .ZN(n17951) );
  XNOR2_X1 U20255 ( .A(n17951), .B(n16982), .ZN(n16985) );
  AOI211_X1 U20256 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16999), .A(n16983), .B(
        n17139), .ZN(n16984) );
  AOI211_X1 U20257 ( .C1(n17084), .C2(n16985), .A(n18308), .B(n16984), .ZN(
        n16990) );
  AOI22_X1 U20258 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17092), .B1(
        n17136), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20259 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16998), .B1(n16987), 
        .B2(n16986), .ZN(n16988) );
  NAND3_X1 U20260 ( .A1(n16990), .A2(n16989), .A3(n16988), .ZN(P3_U2659) );
  INV_X1 U20261 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17964) );
  NAND2_X1 U20262 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16991) );
  NAND2_X1 U20263 ( .A1(n17121), .A2(n17010), .ZN(n17011) );
  INV_X1 U20264 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18980) );
  OAI21_X1 U20265 ( .B1(n16991), .B2(n17011), .A(n18980), .ZN(n16997) );
  INV_X1 U20266 ( .A(n16992), .ZN(n17048) );
  NAND2_X1 U20267 ( .A1(n17962), .A2(n17048), .ZN(n16993) );
  AOI21_X1 U20268 ( .B1(n17964), .B2(n16993), .A(n17937), .ZN(n17966) );
  INV_X1 U20269 ( .A(n16993), .ZN(n17003) );
  OAI21_X1 U20270 ( .B1(n17003), .B2(n17116), .A(n17128), .ZN(n16994) );
  XNOR2_X1 U20271 ( .A(n17966), .B(n16994), .ZN(n16995) );
  OAI22_X1 U20272 ( .A1(n17140), .A2(n17000), .B1(n18938), .B2(n16995), .ZN(
        n16996) );
  AOI211_X1 U20273 ( .C1(n16998), .C2(n16997), .A(n18308), .B(n16996), .ZN(
        n17002) );
  OAI211_X1 U20274 ( .C1(n17006), .C2(n17000), .A(n17110), .B(n16999), .ZN(
        n17001) );
  OAI211_X1 U20275 ( .C1(n17127), .C2(n17964), .A(n17002), .B(n17001), .ZN(
        P3_U2660) );
  NOR2_X1 U20276 ( .A1(n17933), .A2(n18023), .ZN(n18006) );
  NAND2_X1 U20277 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18006), .ZN(
        n17036) );
  NOR2_X1 U20278 ( .A1(n18009), .A2(n17036), .ZN(n17027) );
  NAND2_X1 U20279 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17027), .ZN(
        n17020) );
  AOI21_X1 U20280 ( .B1(n17004), .B2(n17020), .A(n17003), .ZN(n17981) );
  OAI21_X1 U20281 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17020), .A(
        n9807), .ZN(n17022) );
  XNOR2_X1 U20282 ( .A(n17981), .B(n17022), .ZN(n17005) );
  AOI22_X1 U20283 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17092), .B1(
        n17084), .B2(n17005), .ZN(n17014) );
  INV_X1 U20284 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18976) );
  NOR3_X1 U20285 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18976), .A3(n17011), 
        .ZN(n17009) );
  AOI211_X1 U20286 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17007), .A(n17006), .B(
        n17139), .ZN(n17008) );
  AOI211_X1 U20287 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17136), .A(n17009), .B(
        n17008), .ZN(n17013) );
  OAI21_X1 U20288 ( .B1(n17010), .B2(n17132), .A(n17143), .ZN(n17032) );
  NOR2_X1 U20289 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17011), .ZN(n17019) );
  OAI21_X1 U20290 ( .B1(n17032), .B2(n17019), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n17012) );
  NAND4_X1 U20291 ( .A1(n17014), .A2(n17013), .A3(n18426), .A4(n17012), .ZN(
        P3_U2661) );
  NOR2_X1 U20292 ( .A1(n17015), .A2(n17139), .ZN(n17030) );
  AOI21_X1 U20293 ( .B1(n17110), .B2(n17015), .A(n17136), .ZN(n17017) );
  INV_X1 U20294 ( .A(n17032), .ZN(n17016) );
  OAI22_X1 U20295 ( .A1(n17430), .A2(n17017), .B1(n18976), .B2(n17016), .ZN(
        n17018) );
  AOI211_X1 U20296 ( .C1(n17030), .C2(n17430), .A(n17019), .B(n17018), .ZN(
        n17026) );
  OAI21_X1 U20297 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17027), .A(
        n17020), .ZN(n17992) );
  INV_X1 U20298 ( .A(n17992), .ZN(n17023) );
  NOR2_X1 U20299 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18097), .ZN(
        n17078) );
  NAND4_X1 U20300 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18006), .A3(
        n17078), .A4(n17974), .ZN(n17021) );
  OAI221_X1 U20301 ( .B1(n17023), .B2(n17022), .C1(n17992), .C2(n9807), .A(
        n17021), .ZN(n17024) );
  AOI21_X1 U20302 ( .B1(n17084), .B2(n17024), .A(n18308), .ZN(n17025) );
  OAI211_X1 U20303 ( .C1(n17127), .C2(n17974), .A(n17026), .B(n17025), .ZN(
        P3_U2662) );
  AOI21_X1 U20304 ( .B1(n18009), .B2(n17036), .A(n17027), .ZN(n18011) );
  AOI21_X1 U20305 ( .B1(n18006), .B2(n17078), .A(n17116), .ZN(n17038) );
  XOR2_X1 U20306 ( .A(n18011), .B(n17038), .Z(n17028) );
  AOI22_X1 U20307 ( .A1(n17136), .A2(P3_EBX_REG_8__SCAN_IN), .B1(n17084), .B2(
        n17028), .ZN(n17035) );
  NAND2_X1 U20308 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17044), .ZN(n17029) );
  AOI22_X1 U20309 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17092), .B1(
        n17030), .B2(n17029), .ZN(n17034) );
  NOR2_X1 U20310 ( .A1(n17132), .A2(n17031), .ZN(n17043) );
  OAI221_X1 U20311 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(P3_REIP_REG_7__SCAN_IN), 
        .C1(P3_REIP_REG_8__SCAN_IN), .C2(n17043), .A(n17032), .ZN(n17033) );
  NAND4_X1 U20312 ( .A1(n17035), .A2(n17034), .A3(n18426), .A4(n17033), .ZN(
        P3_U2663) );
  OAI221_X1 U20313 ( .B1(n17132), .B2(P3_REIP_REG_6__SCAN_IN), .C1(n17132), 
        .C2(n17055), .A(n17143), .ZN(n17042) );
  OAI21_X1 U20314 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17048), .A(
        n17036), .ZN(n18025) );
  INV_X1 U20315 ( .A(n18025), .ZN(n17039) );
  INV_X1 U20316 ( .A(n17078), .ZN(n17114) );
  OAI21_X1 U20317 ( .B1(n17933), .B2(n17114), .A(n9807), .ZN(n17037) );
  OAI221_X1 U20318 ( .B1(n17039), .B2(n17038), .C1(n18025), .C2(n17037), .A(
        n17084), .ZN(n17040) );
  OAI211_X1 U20319 ( .C1(n18023), .C2(n17127), .A(n18426), .B(n17040), .ZN(
        n17041) );
  AOI221_X1 U20320 ( .B1(n17043), .B2(n18972), .C1(n17042), .C2(
        P3_REIP_REG_7__SCAN_IN), .A(n17041), .ZN(n17046) );
  OAI211_X1 U20321 ( .C1(n17053), .C2(n17047), .A(n17110), .B(n17044), .ZN(
        n17045) );
  OAI211_X1 U20322 ( .C1(n17047), .C2(n17140), .A(n17046), .B(n17045), .ZN(
        P3_U2664) );
  AOI22_X1 U20323 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17092), .B1(
        n17136), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n17059) );
  INV_X1 U20324 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18043) );
  NAND2_X1 U20325 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17961), .ZN(
        n17061) );
  AOI21_X1 U20326 ( .B1(n18043), .B2(n17061), .A(n17048), .ZN(n18039) );
  AOI21_X1 U20327 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9807), .A(
        n17129), .ZN(n17052) );
  INV_X1 U20328 ( .A(n17933), .ZN(n17050) );
  AOI211_X1 U20329 ( .C1(n17050), .C2(n17078), .A(n18039), .B(n17049), .ZN(
        n17051) );
  AOI211_X1 U20330 ( .C1(n18039), .C2(n17052), .A(n18308), .B(n17051), .ZN(
        n17058) );
  OAI21_X1 U20331 ( .B1(n17055), .B2(n17132), .A(n17143), .ZN(n17069) );
  AOI211_X1 U20332 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17070), .A(n17053), .B(
        n17139), .ZN(n17054) );
  AOI21_X1 U20333 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n17069), .A(n17054), .ZN(
        n17057) );
  INV_X1 U20334 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18970) );
  NAND3_X1 U20335 ( .A1(n17121), .A2(n17055), .A3(n18970), .ZN(n17056) );
  NAND4_X1 U20336 ( .A1(n17059), .A2(n17058), .A3(n17057), .A4(n17056), .ZN(
        P3_U2665) );
  OAI21_X1 U20337 ( .B1(n17132), .B2(n17060), .A(n18968), .ZN(n17068) );
  NOR2_X1 U20338 ( .A1(n18097), .A2(n18048), .ZN(n17062) );
  OAI21_X1 U20339 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17062), .A(
        n17061), .ZN(n17063) );
  INV_X1 U20340 ( .A(n17063), .ZN(n18054) );
  INV_X1 U20341 ( .A(n17062), .ZN(n17074) );
  OAI21_X1 U20342 ( .B1(n17074), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n9807), .ZN(n17064) );
  INV_X1 U20343 ( .A(n17064), .ZN(n17077) );
  AOI221_X1 U20344 ( .B1(n18054), .B2(n17064), .C1(n17063), .C2(n17077), .A(
        n18416), .ZN(n17065) );
  OAI22_X1 U20345 ( .A1(n17066), .A2(n17065), .B1(n18049), .B2(n17127), .ZN(
        n17067) );
  AOI21_X1 U20346 ( .B1(n17069), .B2(n17068), .A(n17067), .ZN(n17072) );
  OAI211_X1 U20347 ( .C1(n17085), .C2(n17463), .A(n17110), .B(n17070), .ZN(
        n17071) );
  OAI211_X1 U20348 ( .C1(n17463), .C2(n17140), .A(n17072), .B(n17071), .ZN(
        P3_U2666) );
  NOR2_X1 U20349 ( .A1(n17086), .A2(n17132), .ZN(n17106) );
  NOR2_X1 U20350 ( .A1(n17073), .A2(n17106), .ZN(n17109) );
  INV_X1 U20351 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18966) );
  NAND2_X1 U20352 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18061), .ZN(
        n17095) );
  INV_X1 U20353 ( .A(n17095), .ZN(n17075) );
  OAI21_X1 U20354 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17075), .A(
        n17074), .ZN(n18065) );
  NOR2_X1 U20355 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17076), .ZN(
        n18059) );
  AOI22_X1 U20356 ( .A1(n17078), .A2(n18059), .B1(n17077), .B2(n18065), .ZN(
        n17079) );
  OAI21_X1 U20357 ( .B1(n9807), .B2(n18065), .A(n17079), .ZN(n17083) );
  INV_X1 U20358 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18877) );
  NAND2_X1 U20359 ( .A1(n17081), .A2(n17080), .ZN(n19099) );
  AOI21_X1 U20360 ( .B1(n11517), .B2(n18877), .A(n19099), .ZN(n17082) );
  AOI211_X1 U20361 ( .C1(n17084), .C2(n17083), .A(n18308), .B(n17082), .ZN(
        n17091) );
  AOI211_X1 U20362 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17099), .A(n17085), .B(
        n17139), .ZN(n17089) );
  NAND2_X1 U20363 ( .A1(n17121), .A2(n17086), .ZN(n17087) );
  OAI22_X1 U20364 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17087), .B1(n17140), 
        .B2(n17288), .ZN(n17088) );
  AOI211_X1 U20365 ( .C1(n17092), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n17089), .B(n17088), .ZN(n17090) );
  OAI211_X1 U20366 ( .C1(n17109), .C2(n18966), .A(n17091), .B(n17090), .ZN(
        P3_U2667) );
  AOI22_X1 U20367 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17092), .B1(
        n17136), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n17093) );
  INV_X1 U20368 ( .A(n17093), .ZN(n17105) );
  NAND2_X1 U20369 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18887), .ZN(
        n18882) );
  AOI21_X1 U20370 ( .B1(n17094), .B2(n18882), .A(n9803), .ZN(n19037) );
  INV_X1 U20371 ( .A(n19037), .ZN(n17103) );
  NAND2_X1 U20372 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17097) );
  INV_X1 U20373 ( .A(n17097), .ZN(n17112) );
  OAI21_X1 U20374 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17112), .A(
        n17095), .ZN(n18074) );
  OAI21_X1 U20375 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17097), .A(
        n9807), .ZN(n17113) );
  AOI21_X1 U20376 ( .B1(n18074), .B2(n17113), .A(n18938), .ZN(n17098) );
  OAI21_X1 U20377 ( .B1(n18074), .B2(n17113), .A(n17098), .ZN(n17102) );
  OAI211_X1 U20378 ( .C1(n17125), .C2(n17100), .A(n17110), .B(n17099), .ZN(
        n17101) );
  OAI211_X1 U20379 ( .C1(n17103), .C2(n19099), .A(n17102), .B(n17101), .ZN(
        n17104) );
  AOI211_X1 U20380 ( .C1(n17107), .C2(n17106), .A(n17105), .B(n17104), .ZN(
        n17108) );
  OAI21_X1 U20381 ( .B1(n17109), .B2(n18964), .A(n17108), .ZN(P3_U2668) );
  NOR2_X1 U20382 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17130) );
  OAI21_X1 U20383 ( .B1(n17130), .B2(n17111), .A(n17110), .ZN(n17124) );
  INV_X1 U20384 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18090) );
  AOI21_X1 U20385 ( .B1(n18097), .B2(n18090), .A(n17112), .ZN(n18082) );
  AOI21_X1 U20386 ( .B1(n17114), .B2(n18082), .A(n17113), .ZN(n17115) );
  AOI21_X1 U20387 ( .B1(n18082), .B2(n17116), .A(n17115), .ZN(n17117) );
  NAND2_X1 U20388 ( .A1(n19050), .A2(n18886), .ZN(n18880) );
  NAND2_X1 U20389 ( .A1(n18882), .A2(n18880), .ZN(n19045) );
  OAI22_X1 U20390 ( .A1(n17117), .A2(n18938), .B1(n19045), .B2(n19099), .ZN(
        n17119) );
  OAI22_X1 U20391 ( .A1(n18090), .A2(n17127), .B1(n17143), .B2(n18961), .ZN(
        n17118) );
  AOI211_X1 U20392 ( .C1(n17136), .C2(P3_EBX_REG_2__SCAN_IN), .A(n17119), .B(
        n17118), .ZN(n17123) );
  OAI211_X1 U20393 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17121), .B(n17120), .ZN(n17122) );
  OAI211_X1 U20394 ( .C1(n17125), .C2(n17124), .A(n17123), .B(n17122), .ZN(
        P3_U2669) );
  NAND2_X1 U20395 ( .A1(n17126), .A2(n18886), .ZN(n19051) );
  OAI21_X1 U20396 ( .B1(n18938), .B2(n17128), .A(n17127), .ZN(n17135) );
  OAI22_X1 U20397 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17129), .B1(
        n19066), .B2(n17143), .ZN(n17134) );
  INV_X1 U20398 ( .A(n17130), .ZN(n17131) );
  NAND2_X1 U20399 ( .A1(n17131), .A2(n17479), .ZN(n17487) );
  OAI22_X1 U20400 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17132), .B1(n17139), 
        .B2(n17487), .ZN(n17133) );
  AOI211_X1 U20401 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n17135), .A(
        n17134), .B(n17133), .ZN(n17138) );
  NAND2_X1 U20402 ( .A1(n17136), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(n17137) );
  OAI211_X1 U20403 ( .C1(n19099), .C2(n19051), .A(n17138), .B(n17137), .ZN(
        P3_U2670) );
  NAND2_X1 U20404 ( .A1(n17140), .A2(n17139), .ZN(n17142) );
  AOI22_X1 U20405 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17142), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17141), .ZN(n17145) );
  NAND3_X1 U20406 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19095), .A3(
        n17143), .ZN(n17144) );
  OAI211_X1 U20407 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n19099), .A(
        n17145), .B(n17144), .ZN(P3_U2671) );
  NAND3_X1 U20408 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n17272), .ZN(n17240) );
  NOR4_X1 U20409 ( .A1(n17147), .A2(n17195), .A3(n17146), .A4(n17240), .ZN(
        n17148) );
  NAND4_X1 U20410 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n17184), .A4(n17148), .ZN(n17151) );
  NOR2_X1 U20411 ( .A1(n17152), .A2(n17151), .ZN(n17179) );
  NAND2_X1 U20412 ( .A1(n17468), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17150) );
  NAND2_X1 U20413 ( .A1(n17179), .A2(n10430), .ZN(n17149) );
  OAI22_X1 U20414 ( .A1(n17179), .A2(n17150), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17149), .ZN(P3_U2672) );
  NAND2_X1 U20415 ( .A1(n17152), .A2(n17151), .ZN(n17153) );
  NAND2_X1 U20416 ( .A1(n17153), .A2(n17468), .ZN(n17178) );
  AOI22_X1 U20417 ( .A1(n11629), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17163) );
  INV_X1 U20418 ( .A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U20419 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20420 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17154) );
  OAI211_X1 U20421 ( .C1(n11517), .C2(n17346), .A(n17155), .B(n17154), .ZN(
        n17161) );
  AOI22_X1 U20422 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17159) );
  AOI22_X1 U20423 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U20424 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17157) );
  NAND2_X1 U20425 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n17156) );
  NAND4_X1 U20426 ( .A1(n17159), .A2(n17158), .A3(n17157), .A4(n17156), .ZN(
        n17160) );
  AOI211_X1 U20427 ( .C1(n11665), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17161), .B(n17160), .ZN(n17162) );
  OAI211_X1 U20428 ( .C1(n17415), .C2(n17164), .A(n17163), .B(n17162), .ZN(
        n17181) );
  NAND2_X1 U20429 ( .A1(n17182), .A2(n17181), .ZN(n17180) );
  AOI22_X1 U20430 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11626), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17176) );
  INV_X1 U20431 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17168) );
  AOI22_X1 U20432 ( .A1(n14033), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14036), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17167) );
  AOI22_X1 U20433 ( .A1(n17396), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17166) );
  OAI211_X1 U20434 ( .C1(n11517), .C2(n17168), .A(n17167), .B(n17166), .ZN(
        n17174) );
  AOI22_X1 U20435 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17172) );
  AOI22_X1 U20436 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17171) );
  AOI22_X1 U20437 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17170) );
  NAND2_X1 U20438 ( .A1(n11665), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n17169) );
  NAND4_X1 U20439 ( .A1(n17172), .A2(n17171), .A3(n17170), .A4(n17169), .ZN(
        n17173) );
  AOI211_X1 U20440 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n17174), .B(n17173), .ZN(n17175) );
  OAI211_X1 U20441 ( .C1(n17230), .C2(n17327), .A(n17176), .B(n17175), .ZN(
        n17177) );
  XOR2_X1 U20442 ( .A(n17180), .B(n17177), .Z(n17501) );
  OAI22_X1 U20443 ( .A1(n17179), .A2(n17178), .B1(n17501), .B2(n17468), .ZN(
        P3_U2673) );
  OAI21_X1 U20444 ( .B1(n17182), .B2(n17181), .A(n17180), .ZN(n17505) );
  NOR2_X1 U20445 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17190), .ZN(n17183) );
  AOI22_X1 U20446 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17185), .B1(n17184), 
        .B2(n17183), .ZN(n17186) );
  OAI21_X1 U20447 ( .B1(n17505), .B2(n17468), .A(n17186), .ZN(P3_U2674) );
  OAI21_X1 U20448 ( .B1(n17191), .B2(n17188), .A(n17187), .ZN(n17514) );
  NAND3_X1 U20449 ( .A1(n17190), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17468), 
        .ZN(n17189) );
  OAI221_X1 U20450 ( .B1(n17190), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17468), 
        .C2(n17514), .A(n17189), .ZN(P3_U2676) );
  AOI21_X1 U20451 ( .B1(n17192), .B2(n17197), .A(n17191), .ZN(n17515) );
  AOI22_X1 U20452 ( .A1(n17489), .A2(n17515), .B1(n17200), .B2(n17195), .ZN(
        n17193) );
  OAI21_X1 U20453 ( .B1(n17195), .B2(n17194), .A(n17193), .ZN(P3_U2677) );
  INV_X1 U20454 ( .A(n17196), .ZN(n17205) );
  AOI21_X1 U20455 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17468), .A(n17205), .ZN(
        n17199) );
  OAI21_X1 U20456 ( .B1(n17201), .B2(n17198), .A(n17197), .ZN(n17523) );
  OAI22_X1 U20457 ( .A1(n17200), .A2(n17199), .B1(n17523), .B2(n17468), .ZN(
        P3_U2678) );
  AOI21_X1 U20458 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17468), .A(n17211), .ZN(
        n17204) );
  AOI21_X1 U20459 ( .B1(n17202), .B2(n17207), .A(n17201), .ZN(n17524) );
  INV_X1 U20460 ( .A(n17524), .ZN(n17203) );
  OAI22_X1 U20461 ( .A1(n17205), .A2(n17204), .B1(n17203), .B2(n17468), .ZN(
        P3_U2679) );
  INV_X1 U20462 ( .A(n17206), .ZN(n17242) );
  AND3_X1 U20463 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17242), .ZN(n17225) );
  AOI21_X1 U20464 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17468), .A(n17225), .ZN(
        n17210) );
  OAI21_X1 U20465 ( .B1(n17209), .B2(n17208), .A(n17207), .ZN(n17533) );
  OAI22_X1 U20466 ( .A1(n17211), .A2(n17210), .B1(n17533), .B2(n17468), .ZN(
        P3_U2680) );
  AOI22_X1 U20467 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17468), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n17242), .ZN(n17224) );
  AOI22_X1 U20468 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20469 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17213) );
  AOI22_X1 U20470 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17212) );
  OAI211_X1 U20471 ( .C1(n17426), .C2(n17214), .A(n17213), .B(n17212), .ZN(
        n17220) );
  AOI22_X1 U20472 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17218) );
  AOI22_X1 U20473 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20474 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17216) );
  NAND2_X1 U20475 ( .A1(n11665), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n17215) );
  NAND4_X1 U20476 ( .A1(n17218), .A2(n17217), .A3(n17216), .A4(n17215), .ZN(
        n17219) );
  AOI211_X1 U20477 ( .C1(n9803), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n17220), .B(n17219), .ZN(n17221) );
  OAI211_X1 U20478 ( .C1(n17415), .C2(n17464), .A(n17222), .B(n17221), .ZN(
        n17534) );
  INV_X1 U20479 ( .A(n17534), .ZN(n17223) );
  OAI22_X1 U20480 ( .A1(n17225), .A2(n17224), .B1(n17223), .B2(n17468), .ZN(
        P3_U2681) );
  AOI22_X1 U20481 ( .A1(n11637), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17226) );
  OAI21_X1 U20482 ( .B1(n11496), .B2(n17227), .A(n17226), .ZN(n17239) );
  AOI22_X1 U20483 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U20484 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17228) );
  OAI21_X1 U20485 ( .B1(n17230), .B2(n17229), .A(n17228), .ZN(n17235) );
  AOI22_X1 U20486 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17232) );
  AOI22_X1 U20487 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17231) );
  OAI211_X1 U20488 ( .C1(n17426), .C2(n17233), .A(n17232), .B(n17231), .ZN(
        n17234) );
  AOI211_X1 U20489 ( .C1(n11665), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n17235), .B(n17234), .ZN(n17236) );
  OAI211_X1 U20490 ( .C1(n17415), .C2(n17469), .A(n17237), .B(n17236), .ZN(
        n17238) );
  AOI211_X1 U20491 ( .C1(n17437), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n17239), .B(n17238), .ZN(n17542) );
  AND2_X1 U20492 ( .A1(n17468), .A2(n17240), .ZN(n17255) );
  AOI22_X1 U20493 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17255), .B1(n17242), 
        .B2(n17241), .ZN(n17243) );
  OAI21_X1 U20494 ( .B1(n17542), .B2(n17468), .A(n17243), .ZN(P3_U2682) );
  AOI22_X1 U20495 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17254) );
  AOI22_X1 U20496 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17245) );
  AOI22_X1 U20497 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11684), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17244) );
  OAI211_X1 U20498 ( .C1(n11517), .C2(n17246), .A(n17245), .B(n17244), .ZN(
        n17252) );
  AOI22_X1 U20499 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17250) );
  AOI22_X1 U20500 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11637), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17249) );
  AOI22_X1 U20501 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17248) );
  NAND2_X1 U20502 ( .A1(n11629), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n17247) );
  NAND4_X1 U20503 ( .A1(n17250), .A2(n17249), .A3(n17248), .A4(n17247), .ZN(
        n17251) );
  AOI211_X1 U20504 ( .C1(n11665), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n17252), .B(n17251), .ZN(n17253) );
  OAI211_X1 U20505 ( .C1(n17415), .C2(n17473), .A(n17254), .B(n17253), .ZN(
        n17546) );
  INV_X1 U20506 ( .A(n17546), .ZN(n17257) );
  OAI221_X1 U20507 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(P3_EBX_REG_19__SCAN_IN), 
        .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17274), .A(n17255), .ZN(n17256) );
  OAI21_X1 U20508 ( .B1(n17257), .B2(n17468), .A(n17256), .ZN(P3_U2683) );
  OAI22_X1 U20509 ( .A1(n17258), .A2(n17379), .B1(n17415), .B2(n17476), .ZN(
        n17271) );
  AOI22_X1 U20510 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U20511 ( .A1(n17396), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17268) );
  OAI22_X1 U20512 ( .A1(n9926), .A2(n17260), .B1(n17426), .B2(n17259), .ZN(
        n17266) );
  AOI22_X1 U20513 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17261), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17264) );
  AOI22_X1 U20514 ( .A1(n14033), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17263) );
  AOI22_X1 U20515 ( .A1(n11665), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17262) );
  NAND3_X1 U20516 ( .A1(n17264), .A2(n17263), .A3(n17262), .ZN(n17265) );
  AOI211_X1 U20517 ( .C1(n17413), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n17266), .B(n17265), .ZN(n17267) );
  NAND3_X1 U20518 ( .A1(n17269), .A2(n17268), .A3(n17267), .ZN(n17270) );
  AOI211_X1 U20519 ( .C1(n17442), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n17271), .B(n17270), .ZN(n17554) );
  NOR2_X1 U20520 ( .A1(n17489), .A2(n17272), .ZN(n17292) );
  AOI22_X1 U20521 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17292), .B1(n17274), 
        .B2(n17273), .ZN(n17275) );
  OAI21_X1 U20522 ( .B1(n17554), .B2(n17468), .A(n17275), .ZN(P3_U2684) );
  AOI22_X1 U20523 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17276) );
  OAI21_X1 U20524 ( .B1(n17453), .B2(n17405), .A(n17276), .ZN(n17287) );
  AOI22_X1 U20525 ( .A1(n11626), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17285) );
  AOI22_X1 U20526 ( .A1(n11665), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17277) );
  OAI21_X1 U20527 ( .B1(n17415), .B2(n17278), .A(n17277), .ZN(n17283) );
  AOI22_X1 U20528 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11637), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17280) );
  AOI22_X1 U20529 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17442), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17279) );
  OAI211_X1 U20530 ( .C1(n11517), .C2(n17281), .A(n17280), .B(n17279), .ZN(
        n17282) );
  AOI211_X1 U20531 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n17283), .B(n17282), .ZN(n17284) );
  OAI211_X1 U20532 ( .C1(n9926), .C2(n17393), .A(n17285), .B(n17284), .ZN(
        n17286) );
  AOI211_X1 U20533 ( .C1(n17433), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n17287), .B(n17286), .ZN(n17560) );
  NOR3_X1 U20534 ( .A1(n17288), .A2(n17472), .A3(n17491), .ZN(n17475) );
  NAND2_X1 U20535 ( .A1(n17289), .A2(n17475), .ZN(n17340) );
  NOR2_X1 U20536 ( .A1(n17290), .A2(n17340), .ZN(n17307) );
  AOI22_X1 U20537 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17292), .B1(n17307), 
        .B2(n17291), .ZN(n17293) );
  OAI21_X1 U20538 ( .B1(n17560), .B2(n17468), .A(n17293), .ZN(P3_U2685) );
  NOR2_X1 U20539 ( .A1(n17294), .A2(n17340), .ZN(n17324) );
  AOI21_X1 U20540 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17468), .A(n17324), .ZN(
        n17306) );
  AOI22_X1 U20541 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17304) );
  AOI22_X1 U20542 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17410), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17394), .ZN(n17303) );
  AOI22_X1 U20543 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n9803), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n11665), .ZN(n17302) );
  OAI22_X1 U20544 ( .A1(n17484), .A2(n17415), .B1(n17372), .B2(n17412), .ZN(
        n17300) );
  AOI22_X1 U20545 ( .A1(n11626), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17396), .ZN(n17298) );
  AOI22_X1 U20546 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n14033), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17165), .ZN(n17297) );
  AOI22_X1 U20547 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17296) );
  NAND2_X1 U20548 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17413), .ZN(
        n17295) );
  NAND4_X1 U20549 ( .A1(n17298), .A2(n17297), .A3(n17296), .A4(n17295), .ZN(
        n17299) );
  AOI211_X1 U20550 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n17300), .B(n17299), .ZN(n17301) );
  NAND4_X1 U20551 ( .A1(n17304), .A2(n17303), .A3(n17302), .A4(n17301), .ZN(
        n17561) );
  INV_X1 U20552 ( .A(n17561), .ZN(n17305) );
  OAI22_X1 U20553 ( .A1(n17307), .A2(n17306), .B1(n17305), .B2(n17468), .ZN(
        P3_U2686) );
  INV_X1 U20554 ( .A(n17340), .ZN(n17308) );
  AOI21_X1 U20555 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17468), .A(n17308), .ZN(
        n17323) );
  AOI22_X1 U20556 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11629), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17319) );
  AOI22_X1 U20557 ( .A1(n17396), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U20558 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17309) );
  OAI211_X1 U20559 ( .C1(n11517), .C2(n17311), .A(n17310), .B(n17309), .ZN(
        n17317) );
  AOI22_X1 U20560 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17315) );
  AOI22_X1 U20561 ( .A1(n11626), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U20562 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17313) );
  NAND2_X1 U20563 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n17312) );
  NAND4_X1 U20564 ( .A1(n17315), .A2(n17314), .A3(n17313), .A4(n17312), .ZN(
        n17316) );
  AOI211_X1 U20565 ( .C1(n11665), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17317), .B(n17316), .ZN(n17318) );
  OAI211_X1 U20566 ( .C1(n17321), .C2(n17320), .A(n17319), .B(n17318), .ZN(
        n17566) );
  INV_X1 U20567 ( .A(n17566), .ZN(n17322) );
  OAI22_X1 U20568 ( .A1(n17324), .A2(n17323), .B1(n17322), .B2(n17468), .ZN(
        P3_U2687) );
  AOI22_X1 U20569 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20570 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17417), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17337) );
  OAI22_X1 U20571 ( .A1(n9847), .A2(n17326), .B1(n11496), .B2(n17325), .ZN(
        n17335) );
  OAI22_X1 U20572 ( .A1(n17415), .A2(n17328), .B1(n17372), .B2(n17327), .ZN(
        n17329) );
  AOI21_X1 U20573 ( .B1(n11665), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n17329), .ZN(n17333) );
  AOI22_X1 U20574 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17332) );
  AOI22_X1 U20575 ( .A1(n17396), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17331) );
  AOI22_X1 U20576 ( .A1(n11629), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17330) );
  NAND4_X1 U20577 ( .A1(n17333), .A2(n17332), .A3(n17331), .A4(n17330), .ZN(
        n17334) );
  AOI211_X1 U20578 ( .C1(n17413), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n17335), .B(n17334), .ZN(n17336) );
  NAND3_X1 U20579 ( .A1(n17338), .A2(n17337), .A3(n17336), .ZN(n17576) );
  INV_X1 U20580 ( .A(n17576), .ZN(n17342) );
  INV_X1 U20581 ( .A(n17339), .ZN(n17343) );
  AND2_X1 U20582 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17343), .ZN(n17358) );
  OAI21_X1 U20583 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17358), .A(n17340), .ZN(
        n17341) );
  AOI22_X1 U20584 ( .A1(n17489), .A2(n17342), .B1(n17341), .B2(n17468), .ZN(
        P3_U2688) );
  OAI21_X1 U20585 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17343), .A(n17468), .ZN(
        n17357) );
  AOI22_X1 U20586 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17354) );
  AOI22_X1 U20587 ( .A1(n14033), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17345) );
  AOI22_X1 U20588 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17433), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17344) );
  OAI211_X1 U20589 ( .C1(n17441), .C2(n17346), .A(n17345), .B(n17344), .ZN(
        n17352) );
  AOI22_X1 U20590 ( .A1(n17437), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17350) );
  AOI22_X1 U20591 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17349) );
  AOI22_X1 U20592 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17348) );
  NAND2_X1 U20593 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n17347) );
  NAND4_X1 U20594 ( .A1(n17350), .A2(n17349), .A3(n17348), .A4(n17347), .ZN(
        n17351) );
  AOI211_X1 U20595 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n17352), .B(n17351), .ZN(n17353) );
  OAI211_X1 U20596 ( .C1(n17415), .C2(n17355), .A(n17354), .B(n17353), .ZN(
        n17581) );
  INV_X1 U20597 ( .A(n17581), .ZN(n17356) );
  OAI22_X1 U20598 ( .A1(n17358), .A2(n17357), .B1(n17356), .B2(n17468), .ZN(
        P3_U2689) );
  OAI21_X1 U20599 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17359), .A(n17468), .ZN(
        n17375) );
  AOI22_X1 U20600 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17360) );
  OAI21_X1 U20601 ( .B1(n9926), .B2(n17361), .A(n17360), .ZN(n17374) );
  AOI22_X1 U20602 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17370) );
  AOI22_X1 U20603 ( .A1(n11665), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17362) );
  OAI21_X1 U20604 ( .B1(n17415), .B2(n17363), .A(n17362), .ZN(n17368) );
  INV_X1 U20605 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17366) );
  AOI22_X1 U20606 ( .A1(n17396), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20607 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17364) );
  OAI211_X1 U20608 ( .C1(n11517), .C2(n17366), .A(n17365), .B(n17364), .ZN(
        n17367) );
  AOI211_X1 U20609 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17368), .B(n17367), .ZN(n17369) );
  OAI211_X1 U20610 ( .C1(n17372), .C2(n17371), .A(n17370), .B(n17369), .ZN(
        n17373) );
  AOI211_X1 U20611 ( .C1(n11626), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n17374), .B(n17373), .ZN(n17591) );
  OAI22_X1 U20612 ( .A1(n17376), .A2(n17375), .B1(n17591), .B2(n17468), .ZN(
        P3_U2691) );
  AOI22_X1 U20613 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17438), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U20614 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17378) );
  AOI22_X1 U20615 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17377) );
  OAI211_X1 U20616 ( .C1(n17441), .C2(n17379), .A(n17378), .B(n17377), .ZN(
        n17385) );
  AOI22_X1 U20617 ( .A1(n17410), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17383) );
  AOI22_X1 U20618 ( .A1(n17396), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17394), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U20619 ( .A1(n11667), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17413), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17381) );
  NAND2_X1 U20620 ( .A1(n11629), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n17380) );
  NAND4_X1 U20621 ( .A1(n17383), .A2(n17382), .A3(n17381), .A4(n17380), .ZN(
        n17384) );
  AOI211_X1 U20622 ( .C1(n9803), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n17385), .B(n17384), .ZN(n17386) );
  OAI211_X1 U20623 ( .C1(n10412), .C2(n17388), .A(n17387), .B(n17386), .ZN(
        n17595) );
  INV_X1 U20624 ( .A(n17595), .ZN(n17391) );
  OAI21_X1 U20625 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17409), .A(n17389), .ZN(
        n17390) );
  AOI22_X1 U20626 ( .A1(n17489), .A2(n17391), .B1(n17390), .B2(n17468), .ZN(
        P3_U2692) );
  AOI22_X1 U20627 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17392) );
  OAI21_X1 U20628 ( .B1(n17453), .B2(n17393), .A(n17392), .ZN(n17407) );
  AOI22_X1 U20629 ( .A1(n17394), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17404) );
  AOI22_X1 U20630 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11665), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17395) );
  INV_X1 U20631 ( .A(n17395), .ZN(n17402) );
  AOI22_X1 U20632 ( .A1(n17397), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17400) );
  AOI22_X1 U20633 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20634 ( .A1(n11629), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9803), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17398) );
  NAND3_X1 U20635 ( .A1(n17400), .A2(n17399), .A3(n17398), .ZN(n17401) );
  AOI211_X1 U20636 ( .C1(n17442), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n17402), .B(n17401), .ZN(n17403) );
  OAI211_X1 U20637 ( .C1(n17415), .C2(n17405), .A(n17404), .B(n17403), .ZN(
        n17406) );
  AOI211_X1 U20638 ( .C1(n11667), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17407), .B(n17406), .ZN(n17598) );
  NAND3_X1 U20639 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17467), .A3(n17456), .ZN(
        n17457) );
  OAI21_X1 U20640 ( .B1(n17430), .B2(n17457), .A(n17468), .ZN(n17431) );
  NOR2_X1 U20641 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17431), .ZN(n17408) );
  AOI221_X1 U20642 ( .B1(n17598), .B2(n17489), .C1(n17409), .C2(n17468), .A(
        n17408), .ZN(P3_U2693) );
  AOI22_X1 U20643 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17394), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17411) );
  OAI21_X1 U20644 ( .B1(n10412), .B2(n17412), .A(n17411), .ZN(n17429) );
  INV_X1 U20645 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17427) );
  AOI22_X1 U20646 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17413), .ZN(n17425) );
  OAI22_X1 U20647 ( .A1(n17484), .A2(n17416), .B1(n17415), .B2(n17414), .ZN(
        n17422) );
  AOI22_X1 U20648 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17417), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U20649 ( .A1(n17396), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17165), .ZN(n17419) );
  AOI22_X1 U20650 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11665), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n9803), .ZN(n17418) );
  NAND3_X1 U20651 ( .A1(n17420), .A2(n17419), .A3(n17418), .ZN(n17421) );
  AOI211_X1 U20652 ( .C1(n11667), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n17422), .B(n17421), .ZN(n17424) );
  OAI211_X1 U20653 ( .C1(n17427), .C2(n17426), .A(n17425), .B(n17424), .ZN(
        n17428) );
  AOI211_X1 U20654 ( .C1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(n11626), .A(
        n17429), .B(n17428), .ZN(n17604) );
  AND2_X1 U20655 ( .A1(n17430), .A2(n17457), .ZN(n17432) );
  OAI22_X1 U20656 ( .A1(n17604), .A2(n17468), .B1(n17432), .B2(n17431), .ZN(
        P3_U2694) );
  AOI22_X1 U20657 ( .A1(n17433), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14033), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17434) );
  OAI21_X1 U20658 ( .B1(n9926), .B2(n17435), .A(n17434), .ZN(n17455) );
  AOI22_X1 U20659 ( .A1(n17413), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17436), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17451) );
  INV_X1 U20660 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U20661 ( .A1(n17438), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17437), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17439) );
  OAI21_X1 U20662 ( .B1(n17441), .B2(n17440), .A(n17439), .ZN(n17449) );
  AOI22_X1 U20663 ( .A1(n17442), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17396), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17445) );
  AOI22_X1 U20664 ( .A1(n17443), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17410), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17444) );
  OAI211_X1 U20665 ( .C1(n17447), .C2(n17446), .A(n17445), .B(n17444), .ZN(
        n17448) );
  AOI211_X1 U20666 ( .C1(n11629), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17449), .B(n17448), .ZN(n17450) );
  OAI211_X1 U20667 ( .C1(n17453), .C2(n17452), .A(n17451), .B(n17450), .ZN(
        n17454) );
  AOI211_X1 U20668 ( .C1(n11667), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17455), .B(n17454), .ZN(n17612) );
  AND2_X1 U20669 ( .A1(n17467), .A2(n17456), .ZN(n17461) );
  OAI21_X1 U20670 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17461), .A(n17457), .ZN(
        n17458) );
  AOI22_X1 U20671 ( .A1(n17489), .A2(n17612), .B1(n17458), .B2(n17468), .ZN(
        P3_U2695) );
  AND3_X1 U20672 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17475), .ZN(n17466) );
  AOI21_X1 U20673 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17468), .A(n17466), .ZN(
        n17460) );
  OAI22_X1 U20674 ( .A1(n17461), .A2(n17460), .B1(n17459), .B2(n17468), .ZN(
        P3_U2696) );
  NOR2_X1 U20675 ( .A1(n17463), .A2(n17462), .ZN(n17471) );
  OAI21_X1 U20676 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17471), .A(n17468), .ZN(
        n17465) );
  OAI22_X1 U20677 ( .A1(n17466), .A2(n17465), .B1(n17464), .B2(n17468), .ZN(
        P3_U2697) );
  OAI21_X1 U20678 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17467), .A(n17468), .ZN(
        n17470) );
  OAI22_X1 U20679 ( .A1(n17471), .A2(n17470), .B1(n17469), .B2(n17468), .ZN(
        P3_U2698) );
  NOR2_X1 U20680 ( .A1(n17472), .A2(n17491), .ZN(n17478) );
  AOI21_X1 U20681 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17468), .A(n17478), .ZN(
        n17474) );
  OAI22_X1 U20682 ( .A1(n17475), .A2(n17474), .B1(n17473), .B2(n17468), .ZN(
        P3_U2699) );
  AOI22_X1 U20683 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17468), .B1(n17483), .B2(
        n17482), .ZN(n17477) );
  OAI22_X1 U20684 ( .A1(n17478), .A2(n17477), .B1(n17476), .B2(n17468), .ZN(
        P3_U2700) );
  AOI21_X1 U20685 ( .B1(n10430), .B2(n17479), .A(n17488), .ZN(n17480) );
  OAI22_X1 U20686 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17480), .B1(
        P3_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n17468), .ZN(n17481) );
  AOI21_X1 U20687 ( .B1(n17483), .B2(n17482), .A(n17481), .ZN(P3_U2701) );
  INV_X1 U20688 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17486) );
  OAI222_X1 U20689 ( .A1(n17491), .A2(n17487), .B1(n17486), .B2(n17485), .C1(
        n17484), .C2(n17468), .ZN(P3_U2702) );
  AOI22_X1 U20690 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17489), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17488), .ZN(n17490) );
  OAI21_X1 U20691 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17491), .A(n17490), .ZN(
        P3_U2703) );
  INV_X1 U20692 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17710) );
  INV_X1 U20693 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17706) );
  INV_X1 U20694 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17699) );
  INV_X1 U20695 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17689) );
  INV_X1 U20696 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17750) );
  INV_X1 U20697 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17730) );
  INV_X1 U20698 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17728) );
  INV_X1 U20699 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17726) );
  INV_X1 U20700 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17724) );
  NOR4_X1 U20701 ( .A1(n17730), .A2(n17728), .A3(n17726), .A4(n17724), .ZN(
        n17492) );
  NAND3_X1 U20702 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(n17492), .ZN(n17573) );
  INV_X1 U20703 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17732) );
  NAND2_X1 U20704 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .ZN(n17579) );
  NAND4_X1 U20705 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .A4(P3_EAX_REG_11__SCAN_IN), .ZN(n17493)
         );
  NOR3_X1 U20706 ( .A1(n17732), .A2(n17579), .A3(n17493), .ZN(n17574) );
  NAND2_X1 U20707 ( .A1(n17608), .A2(n17574), .ZN(n17575) );
  NAND4_X1 U20708 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_18__SCAN_IN), .ZN(n17541)
         );
  NAND2_X1 U20709 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17525), .ZN(n17526) );
  NAND2_X1 U20710 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17507), .ZN(n17502) );
  NAND2_X1 U20711 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17498), .ZN(n17497) );
  NAND2_X1 U20712 ( .A1(n17497), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n17496) );
  NAND2_X1 U20713 ( .A1(n18473), .A2(n17609), .ZN(n17572) );
  NAND2_X1 U20714 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17555), .ZN(n17495) );
  OAI221_X1 U20715 ( .B1(n17497), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n17496), 
        .C2(n17609), .A(n17495), .ZN(P3_U2704) );
  AOI22_X1 U20716 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17555), .ZN(n17500) );
  OAI211_X1 U20717 ( .C1(n17498), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17641), .B(
        n17497), .ZN(n17499) );
  OAI211_X1 U20718 ( .C1(n17501), .C2(n17633), .A(n17500), .B(n17499), .ZN(
        P3_U2705) );
  AOI22_X1 U20719 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17555), .ZN(n17504) );
  OAI211_X1 U20720 ( .C1(n17507), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17641), .B(
        n17502), .ZN(n17503) );
  OAI211_X1 U20721 ( .C1(n17505), .C2(n17633), .A(n17504), .B(n17503), .ZN(
        P3_U2706) );
  INV_X1 U20722 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19450) );
  AOI22_X1 U20723 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17567), .B1(n17638), .B2(
        n17506), .ZN(n17510) );
  AOI211_X1 U20724 ( .C1(n17710), .C2(n17511), .A(n17507), .B(n17609), .ZN(
        n17508) );
  INV_X1 U20725 ( .A(n17508), .ZN(n17509) );
  OAI211_X1 U20726 ( .C1(n17572), .C2(n19450), .A(n17510), .B(n17509), .ZN(
        P3_U2707) );
  AOI22_X1 U20727 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17555), .ZN(n17513) );
  OAI211_X1 U20728 ( .C1(n9852), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17641), .B(
        n17511), .ZN(n17512) );
  OAI211_X1 U20729 ( .C1(n17514), .C2(n17633), .A(n17513), .B(n17512), .ZN(
        P3_U2708) );
  INV_X1 U20730 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19438) );
  AOI22_X1 U20731 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17567), .B1(n17638), .B2(
        n17515), .ZN(n17518) );
  AOI211_X1 U20732 ( .C1(n17706), .C2(n17519), .A(n9852), .B(n17609), .ZN(
        n17516) );
  INV_X1 U20733 ( .A(n17516), .ZN(n17517) );
  OAI211_X1 U20734 ( .C1(n17572), .C2(n19438), .A(n17518), .B(n17517), .ZN(
        P3_U2709) );
  AOI22_X1 U20735 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17555), .ZN(n17522) );
  OAI211_X1 U20736 ( .C1(n17520), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17641), .B(
        n17519), .ZN(n17521) );
  OAI211_X1 U20737 ( .C1(n17523), .C2(n17633), .A(n17522), .B(n17521), .ZN(
        P3_U2710) );
  AOI22_X1 U20738 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17567), .B1(n17638), .B2(
        n17524), .ZN(n17528) );
  OAI211_X1 U20739 ( .C1(n17525), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17641), .B(
        n17526), .ZN(n17527) );
  OAI211_X1 U20740 ( .C1(n17572), .C2(n18442), .A(n17528), .B(n17527), .ZN(
        P3_U2711) );
  AOI22_X1 U20741 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17555), .ZN(n17532) );
  OAI211_X1 U20742 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17530), .A(n17641), .B(
        n17529), .ZN(n17531) );
  OAI211_X1 U20743 ( .C1(n17533), .C2(n17633), .A(n17532), .B(n17531), .ZN(
        P3_U2712) );
  NAND2_X1 U20744 ( .A1(n17557), .A2(n17699), .ZN(n17540) );
  AOI22_X1 U20745 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17555), .B1(n17638), .B2(
        n17534), .ZN(n17539) );
  NAND2_X1 U20746 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n17535) );
  INV_X1 U20747 ( .A(n17557), .ZN(n17562) );
  NAND2_X1 U20748 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17551), .ZN(n17547) );
  NAND2_X1 U20749 ( .A1(n17641), .A2(n17547), .ZN(n17545) );
  OAI21_X1 U20750 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17536), .A(n17545), .ZN(
        n17537) );
  AOI22_X1 U20751 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17567), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17537), .ZN(n17538) );
  OAI211_X1 U20752 ( .C1(n17541), .C2(n17540), .A(n17539), .B(n17538), .ZN(
        P3_U2713) );
  INV_X1 U20753 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17697) );
  OAI22_X1 U20754 ( .A1(n17542), .A2(n17633), .B1(n18470), .B2(n17572), .ZN(
        n17543) );
  AOI21_X1 U20755 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17567), .A(n17543), .ZN(
        n17544) );
  OAI221_X1 U20756 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17547), .C1(n17697), 
        .C2(n17545), .A(n17544), .ZN(P3_U2714) );
  INV_X1 U20757 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18464) );
  AOI22_X1 U20758 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17567), .B1(n17638), .B2(
        n17546), .ZN(n17549) );
  OAI211_X1 U20759 ( .C1(n17551), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17641), .B(
        n17547), .ZN(n17548) );
  OAI211_X1 U20760 ( .C1(n17572), .C2(n18464), .A(n17549), .B(n17548), .ZN(
        P3_U2715) );
  AOI22_X1 U20761 ( .A1(n17557), .A2(P3_EAX_REG_18__SCAN_IN), .B1(
        P3_EAX_REG_19__SCAN_IN), .B2(n17641), .ZN(n17550) );
  INV_X1 U20762 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18459) );
  OAI22_X1 U20763 ( .A1(n17551), .A2(n17550), .B1(n18459), .B2(n17572), .ZN(
        n17552) );
  AOI21_X1 U20764 ( .B1(BUF2_REG_3__SCAN_IN), .B2(n17567), .A(n17552), .ZN(
        n17553) );
  OAI21_X1 U20765 ( .B1(n17554), .B2(n17633), .A(n17553), .ZN(P3_U2716) );
  AOI22_X1 U20766 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17567), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17555), .ZN(n17559) );
  NAND2_X1 U20767 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17557), .ZN(n17556) );
  OAI211_X1 U20768 ( .C1(n17557), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17641), .B(
        n17556), .ZN(n17558) );
  OAI211_X1 U20769 ( .C1(n17560), .C2(n17633), .A(n17559), .B(n17558), .ZN(
        P3_U2717) );
  INV_X1 U20770 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18449) );
  AOI22_X1 U20771 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17567), .B1(n17638), .B2(
        n17561), .ZN(n17565) );
  INV_X1 U20772 ( .A(n17568), .ZN(n17563) );
  OAI211_X1 U20773 ( .C1(n17563), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17641), .B(
        n17562), .ZN(n17564) );
  OAI211_X1 U20774 ( .C1(n17572), .C2(n18449), .A(n17565), .B(n17564), .ZN(
        P3_U2718) );
  INV_X1 U20775 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18443) );
  AOI22_X1 U20776 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17567), .B1(n17638), .B2(
        n17566), .ZN(n17571) );
  OAI211_X1 U20777 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17569), .A(n17641), .B(
        n17568), .ZN(n17570) );
  OAI211_X1 U20778 ( .C1(n17572), .C2(n18443), .A(n17571), .B(n17570), .ZN(
        P3_U2719) );
  NAND2_X1 U20779 ( .A1(n17574), .A2(n17616), .ZN(n17578) );
  NAND2_X1 U20780 ( .A1(n17641), .A2(n17575), .ZN(n17583) );
  AOI22_X1 U20781 ( .A1(n17638), .A2(n17576), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n17639), .ZN(n17577) );
  OAI221_X1 U20782 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17578), .C1(n17750), 
        .C2(n17583), .A(n17577), .ZN(P3_U2720) );
  NAND2_X1 U20783 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .ZN(n17580) );
  INV_X1 U20784 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17738) );
  NAND2_X1 U20785 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17616), .ZN(n17602) );
  INV_X1 U20786 ( .A(n17590), .ZN(n17585) );
  NOR2_X1 U20787 ( .A1(n17580), .A2(n17585), .ZN(n17588) );
  INV_X1 U20788 ( .A(n17588), .ZN(n17584) );
  INV_X1 U20789 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17746) );
  AOI22_X1 U20790 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17639), .B1(n17638), .B2(
        n17581), .ZN(n17582) );
  OAI221_X1 U20791 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17584), .C1(n17746), 
        .C2(n17583), .A(n17582), .ZN(P3_U2721) );
  INV_X1 U20792 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17589) );
  INV_X1 U20793 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17741) );
  NOR2_X1 U20794 ( .A1(n17741), .A2(n17585), .ZN(n17593) );
  AOI21_X1 U20795 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17641), .A(n17593), .ZN(
        n17587) );
  OAI222_X1 U20796 ( .A1(n17636), .A2(n17589), .B1(n17588), .B2(n17587), .C1(
        n17633), .C2(n17586), .ZN(P3_U2722) );
  INV_X1 U20797 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17594) );
  AOI21_X1 U20798 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17641), .A(n17590), .ZN(
        n17592) );
  OAI222_X1 U20799 ( .A1(n17636), .A2(n17594), .B1(n17593), .B2(n17592), .C1(
        n17633), .C2(n17591), .ZN(P3_U2723) );
  NAND2_X1 U20800 ( .A1(n17641), .A2(n17597), .ZN(n17600) );
  AOI22_X1 U20801 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17639), .B1(n17638), .B2(
        n17595), .ZN(n17596) );
  OAI221_X1 U20802 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17597), .C1(n17738), 
        .C2(n17600), .A(n17596), .ZN(P3_U2724) );
  INV_X1 U20803 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17601) );
  INV_X1 U20804 ( .A(n17602), .ZN(n17603) );
  AOI21_X1 U20805 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17603), .A(
        P3_EAX_REG_10__SCAN_IN), .ZN(n17599) );
  OAI222_X1 U20806 ( .A1(n17636), .A2(n17601), .B1(n17600), .B2(n17599), .C1(
        n17633), .C2(n17598), .ZN(P3_U2725) );
  INV_X1 U20807 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17607) );
  INV_X1 U20808 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17734) );
  NOR2_X1 U20809 ( .A1(n17734), .A2(n17602), .ZN(n17606) );
  AOI21_X1 U20810 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17641), .A(n17603), .ZN(
        n17605) );
  OAI222_X1 U20811 ( .A1(n17636), .A2(n17607), .B1(n17606), .B2(n17605), .C1(
        n17633), .C2(n17604), .ZN(P3_U2726) );
  AOI22_X1 U20812 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17639), .B1(n17616), .B2(
        n17732), .ZN(n17611) );
  OR3_X1 U20813 ( .A1(n17609), .A2(n17608), .A3(n17732), .ZN(n17610) );
  OAI211_X1 U20814 ( .C1(n17612), .C2(n17633), .A(n17611), .B(n17610), .ZN(
        P3_U2727) );
  INV_X1 U20815 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17720) );
  NOR3_X1 U20816 ( .A1(n18478), .A2(n17640), .A3(n17720), .ZN(n17635) );
  NAND2_X1 U20817 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17635), .ZN(n17624) );
  NOR2_X1 U20818 ( .A1(n17724), .A2(n17624), .ZN(n17626) );
  NAND2_X1 U20819 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17626), .ZN(n17617) );
  NOR2_X1 U20820 ( .A1(n17728), .A2(n17617), .ZN(n17619) );
  OAI21_X1 U20821 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17619), .A(n17641), .ZN(
        n17615) );
  AOI22_X1 U20822 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17639), .B1(n17638), .B2(
        n17613), .ZN(n17614) );
  OAI21_X1 U20823 ( .B1(n17616), .B2(n17615), .A(n17614), .ZN(P3_U2728) );
  INV_X1 U20824 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18474) );
  INV_X1 U20825 ( .A(n17617), .ZN(n17622) );
  AOI21_X1 U20826 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17641), .A(n17622), .ZN(
        n17620) );
  OAI222_X1 U20827 ( .A1(n17636), .A2(n18474), .B1(n17620), .B2(n17619), .C1(
        n17633), .C2(n17618), .ZN(P3_U2729) );
  INV_X1 U20828 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18469) );
  AOI21_X1 U20829 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17641), .A(n17626), .ZN(
        n17623) );
  OAI222_X1 U20830 ( .A1(n17636), .A2(n18469), .B1(n17623), .B2(n17622), .C1(
        n17633), .C2(n17621), .ZN(P3_U2730) );
  INV_X1 U20831 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18463) );
  INV_X1 U20832 ( .A(n17624), .ZN(n17629) );
  AOI21_X1 U20833 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17641), .A(n17629), .ZN(
        n17627) );
  OAI222_X1 U20834 ( .A1(n17636), .A2(n18463), .B1(n17627), .B2(n17626), .C1(
        n17633), .C2(n17625), .ZN(P3_U2731) );
  INV_X1 U20835 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18458) );
  AOI21_X1 U20836 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17641), .A(n17635), .ZN(
        n17630) );
  OAI222_X1 U20837 ( .A1(n17636), .A2(n18458), .B1(n17630), .B2(n17629), .C1(
        n17633), .C2(n17628), .ZN(P3_U2732) );
  INV_X1 U20838 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18454) );
  NOR2_X1 U20839 ( .A1(n18478), .A2(n17640), .ZN(n17631) );
  AOI21_X1 U20840 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17641), .A(n17631), .ZN(
        n17634) );
  OAI222_X1 U20841 ( .A1(n18454), .A2(n17636), .B1(n17635), .B2(n17634), .C1(
        n17633), .C2(n17632), .ZN(P3_U2733) );
  AOI22_X1 U20842 ( .A1(n17639), .A2(BUF2_REG_1__SCAN_IN), .B1(n17638), .B2(
        n17637), .ZN(n17644) );
  OAI211_X1 U20843 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17642), .A(n17641), .B(
        n17640), .ZN(n17643) );
  NAND2_X1 U20844 ( .A1(n17644), .A2(n17643), .ZN(P3_U2734) );
  AND2_X1 U20845 ( .A1(n17660), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20846 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17714) );
  NAND2_X1 U20847 ( .A1(n17663), .A2(n18441), .ZN(n17662) );
  AOI22_X1 U20848 ( .A1(n19081), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17679), .ZN(n17646) );
  OAI21_X1 U20849 ( .B1(n17714), .B2(n17662), .A(n17646), .ZN(P3_U2737) );
  INV_X1 U20850 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17712) );
  AOI22_X1 U20851 ( .A1(n19081), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17647) );
  OAI21_X1 U20852 ( .B1(n17712), .B2(n17662), .A(n17647), .ZN(P3_U2738) );
  AOI22_X1 U20853 ( .A1(n19081), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17648) );
  OAI21_X1 U20854 ( .B1(n17710), .B2(n17662), .A(n17648), .ZN(P3_U2739) );
  INV_X1 U20855 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17708) );
  AOI22_X1 U20856 ( .A1(n19081), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17660), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17649) );
  OAI21_X1 U20857 ( .B1(n17708), .B2(n17662), .A(n17649), .ZN(P3_U2740) );
  AOI22_X1 U20858 ( .A1(n19081), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17650) );
  OAI21_X1 U20859 ( .B1(n17706), .B2(n17662), .A(n17650), .ZN(P3_U2741) );
  AOI22_X1 U20860 ( .A1(n19081), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17660), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17651) );
  OAI21_X1 U20861 ( .B1(n10080), .B2(n17662), .A(n17651), .ZN(P3_U2742) );
  INV_X1 U20862 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17703) );
  AOI22_X1 U20863 ( .A1(n19081), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17660), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17652) );
  OAI21_X1 U20864 ( .B1(n17703), .B2(n17662), .A(n17652), .ZN(P3_U2743) );
  INV_X1 U20865 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17701) );
  CLKBUF_X1 U20866 ( .A(n19081), .Z(n17680) );
  AOI22_X1 U20867 ( .A1(n17680), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17653) );
  OAI21_X1 U20868 ( .B1(n17701), .B2(n17662), .A(n17653), .ZN(P3_U2744) );
  AOI22_X1 U20869 ( .A1(n17680), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17660), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17654) );
  OAI21_X1 U20870 ( .B1(n17699), .B2(n17662), .A(n17654), .ZN(P3_U2745) );
  AOI22_X1 U20871 ( .A1(n17680), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17660), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17655) );
  OAI21_X1 U20872 ( .B1(n17697), .B2(n17662), .A(n17655), .ZN(P3_U2746) );
  INV_X1 U20873 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17695) );
  AOI22_X1 U20874 ( .A1(n17680), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17660), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17656) );
  OAI21_X1 U20875 ( .B1(n17695), .B2(n17662), .A(n17656), .ZN(P3_U2747) );
  INV_X1 U20876 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17693) );
  AOI22_X1 U20877 ( .A1(n17680), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17660), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17657) );
  OAI21_X1 U20878 ( .B1(n17693), .B2(n17662), .A(n17657), .ZN(P3_U2748) );
  INV_X1 U20879 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17691) );
  AOI22_X1 U20880 ( .A1(n17680), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17660), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17658) );
  OAI21_X1 U20881 ( .B1(n17691), .B2(n17662), .A(n17658), .ZN(P3_U2749) );
  AOI22_X1 U20882 ( .A1(n17680), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17660), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17659) );
  OAI21_X1 U20883 ( .B1(n17689), .B2(n17662), .A(n17659), .ZN(P3_U2750) );
  INV_X1 U20884 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17687) );
  AOI22_X1 U20885 ( .A1(n17680), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17660), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17661) );
  OAI21_X1 U20886 ( .B1(n17687), .B2(n17662), .A(n17661), .ZN(P3_U2751) );
  AOI22_X1 U20887 ( .A1(n17680), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17664) );
  OAI21_X1 U20888 ( .B1(n17750), .B2(n17682), .A(n17664), .ZN(P3_U2752) );
  AOI22_X1 U20889 ( .A1(n17680), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17665) );
  OAI21_X1 U20890 ( .B1(n17746), .B2(n17682), .A(n17665), .ZN(P3_U2753) );
  INV_X1 U20891 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17743) );
  AOI22_X1 U20892 ( .A1(n17680), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17666) );
  OAI21_X1 U20893 ( .B1(n17743), .B2(n17682), .A(n17666), .ZN(P3_U2754) );
  AOI22_X1 U20894 ( .A1(n17680), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17667) );
  OAI21_X1 U20895 ( .B1(n17741), .B2(n17682), .A(n17667), .ZN(P3_U2755) );
  AOI22_X1 U20896 ( .A1(n17680), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17668) );
  OAI21_X1 U20897 ( .B1(n17738), .B2(n17682), .A(n17668), .ZN(P3_U2756) );
  INV_X1 U20898 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17736) );
  AOI22_X1 U20899 ( .A1(n17680), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17669) );
  OAI21_X1 U20900 ( .B1(n17736), .B2(n17682), .A(n17669), .ZN(P3_U2757) );
  AOI22_X1 U20901 ( .A1(n17680), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17670) );
  OAI21_X1 U20902 ( .B1(n17734), .B2(n17682), .A(n17670), .ZN(P3_U2758) );
  AOI22_X1 U20903 ( .A1(n17680), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17671) );
  OAI21_X1 U20904 ( .B1(n17732), .B2(n17682), .A(n17671), .ZN(P3_U2759) );
  AOI22_X1 U20905 ( .A1(n17680), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17672) );
  OAI21_X1 U20906 ( .B1(n17730), .B2(n17682), .A(n17672), .ZN(P3_U2760) );
  AOI22_X1 U20907 ( .A1(n17680), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17673) );
  OAI21_X1 U20908 ( .B1(n17728), .B2(n17682), .A(n17673), .ZN(P3_U2761) );
  AOI22_X1 U20909 ( .A1(n17680), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17674) );
  OAI21_X1 U20910 ( .B1(n17726), .B2(n17682), .A(n17674), .ZN(P3_U2762) );
  AOI22_X1 U20911 ( .A1(n17680), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17675) );
  OAI21_X1 U20912 ( .B1(n17724), .B2(n17682), .A(n17675), .ZN(P3_U2763) );
  INV_X1 U20913 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17722) );
  AOI22_X1 U20914 ( .A1(n17680), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17676) );
  OAI21_X1 U20915 ( .B1(n17722), .B2(n17682), .A(n17676), .ZN(P3_U2764) );
  AOI22_X1 U20916 ( .A1(n17680), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17677) );
  OAI21_X1 U20917 ( .B1(n17720), .B2(n17682), .A(n17677), .ZN(P3_U2765) );
  INV_X1 U20918 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17718) );
  AOI22_X1 U20919 ( .A1(n17680), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17678) );
  OAI21_X1 U20920 ( .B1(n17718), .B2(n17682), .A(n17678), .ZN(P3_U2766) );
  AOI22_X1 U20921 ( .A1(n17680), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17679), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17681) );
  OAI21_X1 U20922 ( .B1(n17716), .B2(n17682), .A(n17681), .ZN(P3_U2767) );
  AOI22_X1 U20923 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17739), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17747), .ZN(n17686) );
  OAI21_X1 U20924 ( .B1(n17687), .B2(n17749), .A(n17686), .ZN(P3_U2768) );
  AOI22_X1 U20925 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17739), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17747), .ZN(n17688) );
  OAI21_X1 U20926 ( .B1(n17689), .B2(n17749), .A(n17688), .ZN(P3_U2769) );
  AOI22_X1 U20927 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17739), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17747), .ZN(n17690) );
  OAI21_X1 U20928 ( .B1(n17691), .B2(n17749), .A(n17690), .ZN(P3_U2770) );
  AOI22_X1 U20929 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n9812), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17747), .ZN(n17692) );
  OAI21_X1 U20930 ( .B1(n17693), .B2(n17749), .A(n17692), .ZN(P3_U2771) );
  AOI22_X1 U20931 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n9812), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17747), .ZN(n17694) );
  OAI21_X1 U20932 ( .B1(n17695), .B2(n17749), .A(n17694), .ZN(P3_U2772) );
  AOI22_X1 U20933 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n9812), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17747), .ZN(n17696) );
  OAI21_X1 U20934 ( .B1(n17697), .B2(n17749), .A(n17696), .ZN(P3_U2773) );
  AOI22_X1 U20935 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n9812), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17747), .ZN(n17698) );
  OAI21_X1 U20936 ( .B1(n17699), .B2(n17749), .A(n17698), .ZN(P3_U2774) );
  AOI22_X1 U20937 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n9812), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17747), .ZN(n17700) );
  OAI21_X1 U20938 ( .B1(n17701), .B2(n17749), .A(n17700), .ZN(P3_U2775) );
  AOI22_X1 U20939 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n9812), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17747), .ZN(n17702) );
  OAI21_X1 U20940 ( .B1(n17703), .B2(n17749), .A(n17702), .ZN(P3_U2776) );
  AOI22_X1 U20941 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n9812), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17747), .ZN(n17704) );
  OAI21_X1 U20942 ( .B1(n10080), .B2(n17749), .A(n17704), .ZN(P3_U2777) );
  AOI22_X1 U20943 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9812), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17747), .ZN(n17705) );
  OAI21_X1 U20944 ( .B1(n17706), .B2(n17749), .A(n17705), .ZN(P3_U2778) );
  AOI22_X1 U20945 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n9812), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17747), .ZN(n17707) );
  OAI21_X1 U20946 ( .B1(n17708), .B2(n17749), .A(n17707), .ZN(P3_U2779) );
  AOI22_X1 U20947 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17739), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17747), .ZN(n17709) );
  OAI21_X1 U20948 ( .B1(n17710), .B2(n17749), .A(n17709), .ZN(P3_U2780) );
  AOI22_X1 U20949 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17739), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17747), .ZN(n17711) );
  OAI21_X1 U20950 ( .B1(n17712), .B2(n17749), .A(n17711), .ZN(P3_U2781) );
  AOI22_X1 U20951 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17739), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17747), .ZN(n17713) );
  OAI21_X1 U20952 ( .B1(n17714), .B2(n17749), .A(n17713), .ZN(P3_U2782) );
  AOI22_X1 U20953 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17747), .ZN(n17715) );
  OAI21_X1 U20954 ( .B1(n17716), .B2(n17749), .A(n17715), .ZN(P3_U2783) );
  AOI22_X1 U20955 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17747), .ZN(n17717) );
  OAI21_X1 U20956 ( .B1(n17718), .B2(n17749), .A(n17717), .ZN(P3_U2784) );
  AOI22_X1 U20957 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17747), .ZN(n17719) );
  OAI21_X1 U20958 ( .B1(n17720), .B2(n17749), .A(n17719), .ZN(P3_U2785) );
  AOI22_X1 U20959 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17744), .ZN(n17721) );
  OAI21_X1 U20960 ( .B1(n17722), .B2(n17749), .A(n17721), .ZN(P3_U2786) );
  AOI22_X1 U20961 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17744), .ZN(n17723) );
  OAI21_X1 U20962 ( .B1(n17724), .B2(n17749), .A(n17723), .ZN(P3_U2787) );
  AOI22_X1 U20963 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17744), .ZN(n17725) );
  OAI21_X1 U20964 ( .B1(n17726), .B2(n17749), .A(n17725), .ZN(P3_U2788) );
  AOI22_X1 U20965 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17744), .ZN(n17727) );
  OAI21_X1 U20966 ( .B1(n17728), .B2(n17749), .A(n17727), .ZN(P3_U2789) );
  AOI22_X1 U20967 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17744), .ZN(n17729) );
  OAI21_X1 U20968 ( .B1(n17730), .B2(n17749), .A(n17729), .ZN(P3_U2790) );
  AOI22_X1 U20969 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17744), .ZN(n17731) );
  OAI21_X1 U20970 ( .B1(n17732), .B2(n17749), .A(n17731), .ZN(P3_U2791) );
  AOI22_X1 U20971 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17744), .ZN(n17733) );
  OAI21_X1 U20972 ( .B1(n17734), .B2(n17749), .A(n17733), .ZN(P3_U2792) );
  AOI22_X1 U20973 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9812), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17747), .ZN(n17735) );
  OAI21_X1 U20974 ( .B1(n17736), .B2(n17749), .A(n17735), .ZN(P3_U2793) );
  AOI22_X1 U20975 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17744), .ZN(n17737) );
  OAI21_X1 U20976 ( .B1(n17738), .B2(n17749), .A(n17737), .ZN(P3_U2794) );
  AOI22_X1 U20977 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n9812), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17747), .ZN(n17740) );
  OAI21_X1 U20978 ( .B1(n17741), .B2(n17749), .A(n17740), .ZN(P3_U2795) );
  AOI22_X1 U20979 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17744), .ZN(n17742) );
  OAI21_X1 U20980 ( .B1(n17743), .B2(n17749), .A(n17742), .ZN(P3_U2796) );
  AOI22_X1 U20981 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17744), .ZN(n17745) );
  OAI21_X1 U20982 ( .B1(n17746), .B2(n17749), .A(n17745), .ZN(P3_U2797) );
  AOI22_X1 U20983 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17739), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17747), .ZN(n17748) );
  OAI21_X1 U20984 ( .B1(n17750), .B2(n17749), .A(n17748), .ZN(P3_U2798) );
  AOI22_X1 U20985 ( .A1(n18308), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17751), .ZN(n17761) );
  AOI21_X1 U20986 ( .B1(n17752), .B2(n17812), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17755) );
  AOI21_X1 U20987 ( .B1(n17969), .B2(n17754), .A(n17753), .ZN(n18125) );
  OAI22_X1 U20988 ( .A1(n17756), .A2(n17755), .B1(n18125), .B2(n18015), .ZN(
        n17757) );
  AOI21_X1 U20989 ( .B1(n17759), .B2(n17758), .A(n17757), .ZN(n17760) );
  OAI211_X1 U20990 ( .C1(n17938), .C2(n17762), .A(n17761), .B(n17760), .ZN(
        P3_U2803) );
  INV_X1 U20991 ( .A(n17763), .ZN(n17764) );
  AOI21_X1 U20992 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17765), .A(
        n17764), .ZN(n18129) );
  NOR2_X2 U20993 ( .A1(n17819), .A2(n17952), .ZN(n18087) );
  INV_X1 U20994 ( .A(n18087), .ZN(n17845) );
  NAND3_X1 U20995 ( .A1(n18815), .A2(n9927), .A3(n17778), .ZN(n17767) );
  AOI21_X1 U20996 ( .B1(n10273), .B2(n17767), .A(n17766), .ZN(n17768) );
  AOI211_X1 U20997 ( .C1(n17769), .C2(n17845), .A(n9934), .B(n17768), .ZN(
        n17774) );
  INV_X1 U20998 ( .A(n18130), .ZN(n18126) );
  OAI21_X1 U20999 ( .B1(n18126), .B2(n17770), .A(n10200), .ZN(n17772) );
  NAND2_X1 U21000 ( .A1(n17772), .A2(n17771), .ZN(n17773) );
  OAI211_X1 U21001 ( .C1(n18129), .C2(n18015), .A(n17774), .B(n17773), .ZN(
        P3_U2804) );
  OAI21_X1 U21002 ( .B1(n17969), .B2(n17776), .A(n17775), .ZN(n17777) );
  XOR2_X1 U21003 ( .A(n17777), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18143) );
  AOI211_X1 U21004 ( .C1(n17790), .C2(n17782), .A(n17778), .B(n17791), .ZN(
        n17784) );
  OR2_X1 U21005 ( .A1(n18482), .A2(n9927), .ZN(n17808) );
  OAI211_X1 U21006 ( .C1(n17779), .C2(n18104), .A(n18103), .B(n17808), .ZN(
        n17805) );
  AOI21_X1 U21007 ( .B1(n17819), .B2(n17780), .A(n17805), .ZN(n17789) );
  OAI22_X1 U21008 ( .A1(n17789), .A2(n17782), .B1(n17938), .B2(n17781), .ZN(
        n17783) );
  AOI211_X1 U21009 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n18308), .A(n17784), 
        .B(n17783), .ZN(n17788) );
  XOR2_X1 U21010 ( .A(n18135), .B(n17785), .Z(n18139) );
  XOR2_X1 U21011 ( .A(n18135), .B(n17786), .Z(n18140) );
  AOI22_X1 U21012 ( .A1(n18012), .A2(n18139), .B1(n18040), .B2(n18140), .ZN(
        n17787) );
  OAI211_X1 U21013 ( .C1(n18015), .C2(n18143), .A(n17788), .B(n17787), .ZN(
        P3_U2805) );
  NAND2_X1 U21014 ( .A1(n18308), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18155) );
  OAI221_X1 U21015 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17791), .C1(
        n17790), .C2(n17789), .A(n18155), .ZN(n17792) );
  AOI21_X1 U21016 ( .B1(n17952), .B2(n17793), .A(n17792), .ZN(n17800) );
  OAI22_X1 U21017 ( .A1(n17794), .A2(n17943), .B1(n18146), .B2(n18108), .ZN(
        n17810) );
  OAI21_X1 U21018 ( .B1(n17796), .B2(n18151), .A(n17795), .ZN(n18154) );
  AOI22_X1 U21019 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17810), .B1(
        n17997), .B2(n18154), .ZN(n17799) );
  NAND4_X1 U21020 ( .A1(n18144), .A2(n17797), .A3(n18151), .A4(n17984), .ZN(
        n17798) );
  NAND3_X1 U21021 ( .A1(n17800), .A2(n17799), .A3(n17798), .ZN(P3_U2806) );
  AOI21_X1 U21022 ( .B1(n17801), .B2(n17868), .A(n17815), .ZN(n17802) );
  AOI211_X1 U21023 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17969), .A(
        n17848), .B(n17802), .ZN(n17803) );
  XOR2_X1 U21024 ( .A(n17811), .B(n17803), .Z(n18163) );
  AOI22_X1 U21025 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17805), .B1(
        n17804), .B2(n17845), .ZN(n17806) );
  NAND2_X1 U21026 ( .A1(n18416), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18162) );
  OAI211_X1 U21027 ( .C1(n17808), .C2(n17807), .A(n17806), .B(n18162), .ZN(
        n17809) );
  AOI221_X1 U21028 ( .B1(n17812), .B2(n17811), .C1(n17810), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17809), .ZN(n17813) );
  OAI21_X1 U21029 ( .B1(n18015), .B2(n18163), .A(n17813), .ZN(P3_U2807) );
  OAI221_X1 U21030 ( .B1(n17815), .B2(n17897), .C1(n17815), .C2(n18169), .A(
        n17814), .ZN(n17816) );
  XOR2_X1 U21031 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17816), .Z(
        n18179) );
  AOI22_X1 U21032 ( .A1(n18012), .A2(n18249), .B1(n18040), .B2(n18246), .ZN(
        n17903) );
  OAI21_X1 U21033 ( .B1(n18169), .B2(n17847), .A(n17903), .ZN(n17838) );
  OR2_X1 U21034 ( .A1(n18104), .A2(n17817), .ZN(n17818) );
  OAI211_X1 U21035 ( .C1(n17820), .C2(n18060), .A(n18103), .B(n17818), .ZN(
        n17844) );
  AOI21_X1 U21036 ( .B1(n17819), .B2(n17841), .A(n17844), .ZN(n17833) );
  NAND2_X1 U21037 ( .A1(n17820), .A2(n17949), .ZN(n17835) );
  AOI21_X1 U21038 ( .B1(n17834), .B2(n17825), .A(n17835), .ZN(n17822) );
  AOI22_X1 U21039 ( .A1(n17823), .A2(n17952), .B1(n17822), .B2(n17821), .ZN(
        n17824) );
  NAND2_X1 U21040 ( .A1(n18416), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18177) );
  OAI211_X1 U21041 ( .C1(n17833), .C2(n17825), .A(n17824), .B(n18177), .ZN(
        n17826) );
  AOI21_X1 U21042 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17838), .A(
        n17826), .ZN(n17828) );
  NAND3_X1 U21043 ( .A1(n18169), .A2(n17885), .A3(n18173), .ZN(n17827) );
  OAI211_X1 U21044 ( .C1(n18179), .C2(n18015), .A(n17828), .B(n17827), .ZN(
        P3_U2808) );
  INV_X1 U21045 ( .A(n17829), .ZN(n17830) );
  NAND3_X1 U21046 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18002), .A3(
        n17830), .ZN(n17853) );
  OAI22_X1 U21047 ( .A1(n18184), .A2(n17853), .B1(n17831), .B2(n17868), .ZN(
        n17832) );
  XOR2_X1 U21048 ( .A(n18185), .B(n17832), .Z(n18191) );
  NAND2_X1 U21049 ( .A1(n18416), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18189) );
  OAI221_X1 U21050 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17835), .C1(
        n17834), .C2(n17833), .A(n18189), .ZN(n17836) );
  AOI21_X1 U21051 ( .B1(n17952), .B2(n17837), .A(n17836), .ZN(n17840) );
  NOR2_X1 U21052 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18184), .ZN(
        n18188) );
  AOI22_X1 U21053 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17838), .B1(
        n18188), .B2(n17863), .ZN(n17839) );
  OAI211_X1 U21054 ( .C1(n18191), .C2(n18015), .A(n17840), .B(n17839), .ZN(
        P3_U2809) );
  OAI21_X1 U21055 ( .B1(n17842), .B2(n18482), .A(n17841), .ZN(n17843) );
  AOI22_X1 U21056 ( .A1(n17846), .A2(n17845), .B1(n17844), .B2(n17843), .ZN(
        n17852) );
  NAND3_X1 U21057 ( .A1(n18218), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18193) );
  INV_X1 U21058 ( .A(n18193), .ZN(n18165) );
  OAI21_X1 U21059 ( .B1(n17847), .B2(n18165), .A(n17903), .ZN(n17864) );
  INV_X1 U21060 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18204) );
  AOI221_X1 U21061 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17853), 
        .C1(n18204), .C2(n17867), .A(n17848), .ZN(n17849) );
  XOR2_X1 U21062 ( .A(n17849), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n18198) );
  AOI22_X1 U21063 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17864), .B1(
        n17997), .B2(n18198), .ZN(n17851) );
  NAND2_X1 U21064 ( .A1(n18308), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18199) );
  NOR2_X1 U21065 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18204), .ZN(
        n18197) );
  NAND2_X1 U21066 ( .A1(n17863), .A2(n18197), .ZN(n17850) );
  NAND4_X1 U21067 ( .A1(n17852), .A2(n17851), .A3(n18199), .A4(n17850), .ZN(
        P3_U2810) );
  OAI21_X1 U21068 ( .B1(n17868), .B2(n17867), .A(n17853), .ZN(n17854) );
  XOR2_X1 U21069 ( .A(n17854), .B(n18204), .Z(n18208) );
  OAI21_X1 U21070 ( .B1(n18060), .B2(n17857), .A(n18103), .ZN(n17880) );
  INV_X1 U21071 ( .A(n17880), .ZN(n17855) );
  OAI21_X1 U21072 ( .B1(n17856), .B2(n18104), .A(n17855), .ZN(n17874) );
  INV_X1 U21073 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17859) );
  NAND2_X1 U21074 ( .A1(n17857), .A2(n17949), .ZN(n17871) );
  AOI221_X1 U21075 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(n17859), .C2(n17858), .A(
        n17871), .ZN(n17862) );
  OAI22_X1 U21076 ( .A1(n18426), .A2(n18996), .B1(n17938), .B2(n17860), .ZN(
        n17861) );
  AOI211_X1 U21077 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17874), .A(
        n17862), .B(n17861), .ZN(n17866) );
  AOI22_X1 U21078 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17864), .B1(
        n17863), .B2(n18204), .ZN(n17865) );
  OAI211_X1 U21079 ( .C1(n18208), .C2(n18015), .A(n17866), .B(n17865), .ZN(
        P3_U2811) );
  OAI21_X1 U21080 ( .B1(n17969), .B2(n18221), .A(n17867), .ZN(n17869) );
  XNOR2_X1 U21081 ( .A(n17869), .B(n17868), .ZN(n18226) );
  NAND2_X1 U21082 ( .A1(n18416), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18224) );
  INV_X1 U21083 ( .A(n18224), .ZN(n17873) );
  OAI22_X1 U21084 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17871), .B1(
        n17870), .B2(n17938), .ZN(n17872) );
  AOI211_X1 U21085 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17874), .A(
        n17873), .B(n17872), .ZN(n17876) );
  OAI21_X1 U21086 ( .B1(n18218), .B2(n17899), .A(n17903), .ZN(n17886) );
  NOR2_X1 U21087 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18181), .ZN(
        n18223) );
  AOI22_X1 U21088 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17886), .B1(
        n17885), .B2(n18223), .ZN(n17875) );
  OAI211_X1 U21089 ( .C1(n18015), .C2(n18226), .A(n17876), .B(n17875), .ZN(
        P3_U2812) );
  AOI21_X1 U21090 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17878), .A(
        n17877), .ZN(n18232) );
  NAND2_X1 U21091 ( .A1(n18416), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18230) );
  INV_X1 U21092 ( .A(n17879), .ZN(n17881) );
  OAI221_X1 U21093 ( .B1(n18815), .B2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C1(
        n17881), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(n17880), .ZN(
        n17882) );
  OAI211_X1 U21094 ( .C1(n17883), .C2(n18087), .A(n18230), .B(n17882), .ZN(
        n17884) );
  INV_X1 U21095 ( .A(n17884), .ZN(n17888) );
  NOR2_X1 U21096 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18233), .ZN(
        n18228) );
  AOI22_X1 U21097 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17886), .B1(
        n17885), .B2(n18228), .ZN(n17887) );
  OAI211_X1 U21098 ( .C1(n18232), .C2(n18015), .A(n17888), .B(n17887), .ZN(
        P3_U2813) );
  AOI21_X1 U21099 ( .B1(n17935), .B2(n10271), .A(n18089), .ZN(n17919) );
  OAI21_X1 U21100 ( .B1(n17890), .B2(n18104), .A(n17919), .ZN(n17904) );
  NAND2_X1 U21101 ( .A1(n18416), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17894) );
  NOR2_X1 U21102 ( .A1(n17891), .A2(n10271), .ZN(n17906) );
  OAI211_X1 U21103 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17906), .B(n17892), .ZN(n17893) );
  OAI211_X1 U21104 ( .C1(n17938), .C2(n17895), .A(n17894), .B(n17893), .ZN(
        n17901) );
  OAI21_X1 U21105 ( .B1(n17969), .B2(n17897), .A(n17896), .ZN(n17898) );
  XOR2_X1 U21106 ( .A(n17898), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(
        n18245) );
  OAI22_X1 U21107 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17899), .B1(
        n18245), .B2(n18015), .ZN(n17900) );
  AOI211_X1 U21108 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n17904), .A(
        n17901), .B(n17900), .ZN(n17902) );
  OAI21_X1 U21109 ( .B1(n17903), .B2(n18233), .A(n17902), .ZN(P3_U2814) );
  NOR2_X1 U21110 ( .A1(n18426), .A2(n18988), .ZN(n18247) );
  AOI221_X1 U21111 ( .B1(n17906), .B2(n17905), .C1(n17904), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18247), .ZN(n17914) );
  INV_X1 U21112 ( .A(n18295), .ZN(n18001) );
  NAND2_X1 U21113 ( .A1(n17907), .A2(n18001), .ZN(n17925) );
  NAND2_X1 U21114 ( .A1(n18002), .A2(n18277), .ZN(n17917) );
  NAND2_X1 U21115 ( .A1(n17908), .A2(n17969), .ZN(n17916) );
  NOR2_X1 U21116 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18294), .ZN(
        n18275) );
  AOI221_X1 U21117 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17917), 
        .C1(n18268), .C2(n17916), .A(n18275), .ZN(n17909) );
  XOR2_X1 U21118 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17909), .Z(
        n18254) );
  NOR2_X1 U21119 ( .A1(n17927), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18259) );
  NAND2_X1 U21120 ( .A1(n18040), .A2(n18246), .ZN(n17911) );
  NOR2_X1 U21121 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17924), .ZN(
        n18251) );
  NAND2_X1 U21122 ( .A1(n18012), .A2(n18249), .ZN(n17910) );
  OAI22_X1 U21123 ( .A1(n18259), .A2(n17911), .B1(n18251), .B2(n17910), .ZN(
        n17912) );
  AOI21_X1 U21124 ( .B1(n17997), .B2(n18254), .A(n17912), .ZN(n17913) );
  OAI211_X1 U21125 ( .C1(n17938), .C2(n17915), .A(n17914), .B(n17913), .ZN(
        P3_U2815) );
  AOI21_X1 U21126 ( .B1(n17917), .B2(n17916), .A(n18275), .ZN(n17918) );
  XOR2_X1 U21127 ( .A(n18268), .B(n17918), .Z(n18274) );
  AOI221_X1 U21128 ( .B1(n17921), .B2(n17920), .C1(n18482), .C2(n17920), .A(
        n17919), .ZN(n17922) );
  NOR2_X1 U21129 ( .A1(n18426), .A2(n18987), .ZN(n18260) );
  AOI211_X1 U21130 ( .C1(n17923), .C2(n17845), .A(n17922), .B(n18260), .ZN(
        n17930) );
  INV_X1 U21131 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17926) );
  AOI221_X1 U21132 ( .B1(n17926), .B2(n18268), .C1(n17925), .C2(n18268), .A(
        n17924), .ZN(n18270) );
  AOI21_X1 U21133 ( .B1(n18268), .B2(n17928), .A(n17927), .ZN(n18266) );
  AOI22_X1 U21134 ( .A1(n18012), .A2(n18270), .B1(n18040), .B2(n18266), .ZN(
        n17929) );
  OAI211_X1 U21135 ( .C1(n18015), .C2(n18274), .A(n17930), .B(n17929), .ZN(
        P3_U2816) );
  NAND2_X1 U21136 ( .A1(n17969), .A2(n17931), .ZN(n17946) );
  OAI221_X1 U21137 ( .B1(n18277), .B2(n18294), .C1(n18277), .C2(n17969), .A(
        n17946), .ZN(n17932) );
  XOR2_X1 U21138 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17932), .Z(
        n18284) );
  AOI21_X1 U21139 ( .B1(n17935), .B2(n17933), .A(n18089), .ZN(n18024) );
  NAND2_X1 U21140 ( .A1(n17935), .A2(n17934), .ZN(n17936) );
  OAI211_X1 U21141 ( .C1(n17937), .C2(n18104), .A(n18024), .B(n17936), .ZN(
        n17953) );
  INV_X1 U21142 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18984) );
  NOR2_X1 U21143 ( .A1(n18426), .A2(n18984), .ZN(n17942) );
  OAI211_X1 U21144 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17950), .B(n17949), .ZN(n17940) );
  OAI22_X1 U21145 ( .A1(n10426), .A2(n17940), .B1(n17939), .B2(n17938), .ZN(
        n17941) );
  AOI211_X1 U21146 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17953), .A(
        n17942), .B(n17941), .ZN(n17945) );
  OAI22_X1 U21147 ( .A1(n18278), .A2(n18108), .B1(n18277), .B2(n17943), .ZN(
        n17958) );
  INV_X1 U21148 ( .A(n17947), .ZN(n18305) );
  NOR2_X1 U21149 ( .A1(n18000), .A2(n18305), .ZN(n17959) );
  AOI22_X1 U21150 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17958), .B1(
        n18275), .B2(n17959), .ZN(n17944) );
  OAI211_X1 U21151 ( .C1(n18015), .C2(n18284), .A(n17945), .B(n17944), .ZN(
        P3_U2817) );
  OAI221_X1 U21152 ( .B1(n17969), .B2(n17947), .C1(n17969), .C2(n18001), .A(
        n17946), .ZN(n17948) );
  XNOR2_X1 U21153 ( .A(n18294), .B(n17948), .ZN(n18285) );
  NAND2_X1 U21154 ( .A1(n17950), .A2(n17949), .ZN(n17956) );
  AOI22_X1 U21155 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17953), .B1(
        n17952), .B2(n17951), .ZN(n17955) );
  NAND2_X1 U21156 ( .A1(n18416), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17954) );
  OAI211_X1 U21157 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17956), .A(
        n17955), .B(n17954), .ZN(n17957) );
  AOI221_X1 U21158 ( .B1(n17959), .B2(n18294), .C1(n17958), .C2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17957), .ZN(n17960) );
  OAI21_X1 U21159 ( .B1(n18015), .B2(n18285), .A(n17960), .ZN(P3_U2818) );
  INV_X1 U21160 ( .A(n18303), .ZN(n17979) );
  NAND2_X1 U21161 ( .A1(n17979), .A2(n18307), .ZN(n18314) );
  NAND2_X1 U21162 ( .A1(n18815), .A2(n17961), .ZN(n18032) );
  NOR2_X1 U21163 ( .A1(n18043), .A2(n18032), .ZN(n17990) );
  NAND2_X1 U21164 ( .A1(n17962), .A2(n17990), .ZN(n17975) );
  NAND2_X1 U21165 ( .A1(n18098), .A2(n17975), .ZN(n17963) );
  NAND2_X1 U21166 ( .A1(n18308), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18312) );
  OAI221_X1 U21167 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17975), .C1(
        n17964), .C2(n17963), .A(n18312), .ZN(n17965) );
  AOI21_X1 U21168 ( .B1(n17966), .B2(n17845), .A(n17965), .ZN(n17973) );
  AOI22_X1 U21169 ( .A1(n18297), .A2(n18040), .B1(n18012), .B2(n18295), .ZN(
        n17999) );
  OAI21_X1 U21170 ( .B1(n17979), .B2(n18000), .A(n17999), .ZN(n17983) );
  NAND2_X1 U21171 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18211) );
  NOR3_X1 U21172 ( .A1(n17967), .A2(n18211), .A3(n17969), .ZN(n17980) );
  AND2_X1 U21173 ( .A1(n17968), .A2(n17969), .ZN(n17976) );
  AOI22_X1 U21174 ( .A1(n17979), .A2(n17980), .B1(n17970), .B2(n17976), .ZN(
        n17971) );
  XOR2_X1 U21175 ( .A(n18307), .B(n17971), .Z(n18311) );
  AOI22_X1 U21176 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17983), .B1(
        n17997), .B2(n18311), .ZN(n17972) );
  OAI211_X1 U21177 ( .C1(n18000), .C2(n18314), .A(n17973), .B(n17972), .ZN(
        P3_U2819) );
  INV_X1 U21178 ( .A(n17990), .ZN(n18022) );
  NOR3_X1 U21179 ( .A1(n18005), .A2(n17974), .A3(n18022), .ZN(n17994) );
  OAI211_X1 U21180 ( .C1(n17994), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18098), .B(n17975), .ZN(n17987) );
  OR2_X1 U21181 ( .A1(n17980), .A2(n17976), .ZN(n17989) );
  NAND2_X1 U21182 ( .A1(n18328), .A2(n17989), .ZN(n17988) );
  NOR3_X1 U21183 ( .A1(n18315), .A2(n11729), .A3(n17988), .ZN(n17978) );
  AOI221_X1 U21184 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17980), .C1(
        n18328), .C2(n17976), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17977) );
  AOI211_X1 U21185 ( .C1(n17980), .C2(n17979), .A(n17978), .B(n17977), .ZN(
        n18319) );
  AOI22_X1 U21186 ( .A1(n17997), .A2(n18319), .B1(n17981), .B2(n17845), .ZN(
        n17986) );
  NAND2_X1 U21187 ( .A1(n18416), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18320) );
  OAI211_X1 U21188 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17984), .A(
        n17983), .B(n17982), .ZN(n17985) );
  NAND4_X1 U21189 ( .A1(n17987), .A2(n17986), .A3(n18320), .A4(n17985), .ZN(
        P3_U2820) );
  OAI21_X1 U21190 ( .B1(n17989), .B2(n18328), .A(n17988), .ZN(n18324) );
  NOR2_X1 U21191 ( .A1(n18426), .A2(n18976), .ZN(n17996) );
  AOI22_X1 U21192 ( .A1(n17991), .A2(n17990), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18098), .ZN(n17993) );
  OAI22_X1 U21193 ( .A1(n17994), .A2(n17993), .B1(n18087), .B2(n17992), .ZN(
        n17995) );
  AOI211_X1 U21194 ( .C1(n17997), .C2(n18324), .A(n17996), .B(n17995), .ZN(
        n17998) );
  OAI221_X1 U21195 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18000), .C1(
        n18328), .C2(n17999), .A(n17998), .ZN(P3_U2821) );
  NOR2_X1 U21196 ( .A1(n18001), .A2(n17968), .ZN(n18339) );
  XOR2_X1 U21197 ( .A(n18339), .B(n18002), .Z(n18345) );
  AOI21_X1 U21198 ( .B1(n18004), .B2(n18337), .A(n18003), .ZN(n18341) );
  AOI22_X1 U21199 ( .A1(n18308), .A2(P3_REIP_REG_8__SCAN_IN), .B1(n18040), 
        .B2(n18341), .ZN(n18008) );
  OAI211_X1 U21200 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18006), .A(
        n18815), .B(n18005), .ZN(n18007) );
  OAI211_X1 U21201 ( .C1(n18024), .C2(n18009), .A(n18008), .B(n18007), .ZN(
        n18010) );
  AOI21_X1 U21202 ( .B1(n18011), .B2(n17845), .A(n18010), .ZN(n18014) );
  NAND2_X1 U21203 ( .A1(n18345), .A2(n18012), .ZN(n18013) );
  OAI211_X1 U21204 ( .C1(n18345), .C2(n18015), .A(n18014), .B(n18013), .ZN(
        P3_U2822) );
  OAI21_X1 U21205 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18017), .A(
        n18016), .ZN(n18349) );
  OAI21_X1 U21206 ( .B1(n18020), .B2(n18019), .A(n18018), .ZN(n18021) );
  XOR2_X1 U21207 ( .A(n18021), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18348) );
  OAI22_X1 U21208 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18022), .B1(
        n18108), .B2(n18348), .ZN(n18027) );
  OAI22_X1 U21209 ( .A1(n18087), .A2(n18025), .B1(n18024), .B2(n18023), .ZN(
        n18026) );
  AOI211_X1 U21210 ( .C1(n18308), .C2(P3_REIP_REG_7__SCAN_IN), .A(n18027), .B(
        n18026), .ZN(n18028) );
  OAI21_X1 U21211 ( .B1(n18107), .B2(n18349), .A(n18028), .ZN(P3_U2823) );
  NAND2_X1 U21212 ( .A1(n18098), .A2(n18032), .ZN(n18047) );
  OAI21_X1 U21213 ( .B1(n18031), .B2(n18030), .A(n18029), .ZN(n18363) );
  OAI22_X1 U21214 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18032), .B1(
        n18107), .B2(n18363), .ZN(n18033) );
  AOI21_X1 U21215 ( .B1(n18416), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18033), .ZN(
        n18042) );
  AOI22_X1 U21216 ( .A1(n18036), .A2(n18044), .B1(n18035), .B2(n18034), .ZN(
        n18037) );
  XNOR2_X1 U21217 ( .A(n18038), .B(n18037), .ZN(n18361) );
  AOI22_X1 U21218 ( .A1(n18040), .A2(n18361), .B1(n18039), .B2(n17845), .ZN(
        n18041) );
  OAI211_X1 U21219 ( .C1(n18043), .C2(n18047), .A(n18042), .B(n18041), .ZN(
        P3_U2824) );
  OAI21_X1 U21220 ( .B1(n18046), .B2(n18045), .A(n18044), .ZN(n18371) );
  AOI221_X1 U21221 ( .B1(n18089), .B2(n18049), .C1(n18048), .C2(n18049), .A(
        n18047), .ZN(n18053) );
  OAI21_X1 U21222 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18051), .A(
        n18050), .ZN(n18364) );
  OAI22_X1 U21223 ( .A1(n18426), .A2(n18968), .B1(n18107), .B2(n18364), .ZN(
        n18052) );
  AOI211_X1 U21224 ( .C1(n18054), .C2(n17845), .A(n18053), .B(n18052), .ZN(
        n18055) );
  OAI21_X1 U21225 ( .B1(n18108), .B2(n18371), .A(n18055), .ZN(P3_U2825) );
  OAI21_X1 U21226 ( .B1(n18058), .B2(n18057), .A(n18056), .ZN(n18382) );
  AOI22_X1 U21227 ( .A1(n18308), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18815), 
        .B2(n18059), .ZN(n18068) );
  OAI21_X1 U21228 ( .B1(n18061), .B2(n18060), .A(n18103), .ZN(n18077) );
  OAI21_X1 U21229 ( .B1(n18064), .B2(n18063), .A(n18062), .ZN(n18376) );
  OAI22_X1 U21230 ( .A1(n18087), .A2(n18065), .B1(n18108), .B2(n18376), .ZN(
        n18066) );
  AOI21_X1 U21231 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18077), .A(
        n18066), .ZN(n18067) );
  OAI211_X1 U21232 ( .C1(n18107), .C2(n18382), .A(n18068), .B(n18067), .ZN(
        P3_U2826) );
  OAI21_X1 U21233 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18070), .A(
        n18069), .ZN(n18391) );
  NOR2_X1 U21234 ( .A1(n18089), .A2(n18090), .ZN(n18076) );
  OAI21_X1 U21235 ( .B1(n18073), .B2(n18072), .A(n18071), .ZN(n18384) );
  OAI22_X1 U21236 ( .A1(n18087), .A2(n18074), .B1(n18108), .B2(n18384), .ZN(
        n18075) );
  AOI221_X1 U21237 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18077), .C1(
        n18076), .C2(n18077), .A(n18075), .ZN(n18078) );
  NAND2_X1 U21238 ( .A1(n18416), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18389) );
  OAI211_X1 U21239 ( .C1(n18107), .C2(n18391), .A(n18078), .B(n18389), .ZN(
        P3_U2827) );
  OAI21_X1 U21240 ( .B1(n18081), .B2(n18080), .A(n18079), .ZN(n18407) );
  INV_X1 U21241 ( .A(n18082), .ZN(n18086) );
  OAI21_X1 U21242 ( .B1(n18085), .B2(n18084), .A(n18083), .ZN(n18402) );
  OAI22_X1 U21243 ( .A1(n18087), .A2(n18086), .B1(n18108), .B2(n18402), .ZN(
        n18088) );
  AOI221_X1 U21244 ( .B1(n18815), .B2(n18090), .C1(n18089), .C2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n18088), .ZN(n18091) );
  NAND2_X1 U21245 ( .A1(n18416), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18405) );
  OAI211_X1 U21246 ( .C1(n18107), .C2(n18407), .A(n18091), .B(n18405), .ZN(
        P3_U2828) );
  NOR2_X1 U21247 ( .A1(n18092), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18093) );
  XOR2_X1 U21248 ( .A(n18093), .B(n18095), .Z(n18415) );
  INV_X1 U21249 ( .A(n18415), .ZN(n18100) );
  OAI21_X1 U21250 ( .B1(n18095), .B2(n18101), .A(n18094), .ZN(n18419) );
  OAI22_X1 U21251 ( .A1(n18426), .A2(n19066), .B1(n18107), .B2(n18419), .ZN(
        n18096) );
  AOI221_X1 U21252 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18098), .C1(
        n18097), .C2(n17845), .A(n18096), .ZN(n18099) );
  OAI21_X1 U21253 ( .B1(n18100), .B2(n18108), .A(n18099), .ZN(P3_U2829) );
  AOI21_X1 U21254 ( .B1(n18102), .B2(n19061), .A(n18101), .ZN(n18422) );
  INV_X1 U21255 ( .A(n18422), .ZN(n18424) );
  NAND3_X1 U21256 ( .A1(n19042), .A2(n18104), .A3(n18103), .ZN(n18105) );
  AOI22_X1 U21257 ( .A1(n18308), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18105), .ZN(n18106) );
  OAI221_X1 U21258 ( .B1(n18422), .B2(n18108), .C1(n18424), .C2(n18107), .A(
        n18106), .ZN(P3_U2830) );
  NAND3_X1 U21259 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18171), .A3(
        n18170), .ZN(n18158) );
  AOI221_X1 U21260 ( .B1(n18110), .B2(n18109), .C1(n18158), .C2(n18109), .A(
        n18427), .ZN(n18122) );
  NAND2_X1 U21261 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18134) );
  INV_X1 U21262 ( .A(n18134), .ZN(n18113) );
  INV_X1 U21263 ( .A(n18111), .ZN(n18112) );
  OAI221_X1 U21264 ( .B1(n18112), .B2(n18304), .C1(n18112), .C2(n18164), .A(
        n18374), .ZN(n18145) );
  OAI21_X1 U21265 ( .B1(n18113), .B2(n18394), .A(n18145), .ZN(n18131) );
  INV_X1 U21266 ( .A(n18114), .ZN(n18115) );
  OAI22_X1 U21267 ( .A1(n18900), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18898), .B2(n18115), .ZN(n18119) );
  OAI22_X1 U21268 ( .A1(n18117), .A2(n18401), .B1(n18116), .B2(n18276), .ZN(
        n18118) );
  NOR4_X1 U21269 ( .A1(n18120), .A2(n18131), .A3(n18119), .A4(n18118), .ZN(
        n18127) );
  OAI211_X1 U21270 ( .C1(n18900), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n18127), .ZN(n18121) );
  AOI22_X1 U21271 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18404), .B1(
        n18122), .B2(n18121), .ZN(n18124) );
  NAND2_X1 U21272 ( .A1(n18416), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18123) );
  OAI211_X1 U21273 ( .C1(n18125), .C2(n18344), .A(n18124), .B(n18123), .ZN(
        P3_U2835) );
  NOR2_X1 U21274 ( .A1(n18126), .A2(n18158), .ZN(n18128) );
  NOR2_X1 U21275 ( .A1(n18426), .A2(n19008), .ZN(n18138) );
  AOI22_X1 U21276 ( .A1(n18130), .A2(n18149), .B1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18393), .ZN(n18132) );
  OAI21_X1 U21277 ( .B1(n18132), .B2(n18131), .A(n18409), .ZN(n18133) );
  AOI221_X1 U21278 ( .B1(n18136), .B2(n18135), .C1(n18134), .C2(n18135), .A(
        n18133), .ZN(n18137) );
  AOI211_X1 U21279 ( .C1(n18404), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18138), .B(n18137), .ZN(n18142) );
  AOI22_X1 U21280 ( .A1(n18425), .A2(n18140), .B1(n18340), .B2(n18139), .ZN(
        n18141) );
  OAI211_X1 U21281 ( .C1(n18344), .C2(n18143), .A(n18142), .B(n18141), .ZN(
        P3_U2837) );
  NAND2_X1 U21282 ( .A1(n18144), .A2(n18151), .ZN(n18157) );
  OAI21_X1 U21283 ( .B1(n18146), .B2(n18401), .A(n18145), .ZN(n18147) );
  AOI211_X1 U21284 ( .C1(n18296), .C2(n18148), .A(n18404), .B(n18147), .ZN(
        n18152) );
  OAI211_X1 U21285 ( .C1(n18149), .C2(n18393), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n18152), .ZN(n18150) );
  AND2_X1 U21286 ( .A1(n18426), .A2(n18150), .ZN(n18159) );
  AOI21_X1 U21287 ( .B1(n18241), .B2(n18152), .A(n18151), .ZN(n18153) );
  AOI22_X1 U21288 ( .A1(n18325), .A2(n18154), .B1(n18159), .B2(n18153), .ZN(
        n18156) );
  OAI211_X1 U21289 ( .C1(n18157), .C2(n18180), .A(n18156), .B(n18155), .ZN(
        P3_U2838) );
  INV_X1 U21290 ( .A(n18158), .ZN(n18160) );
  OAI221_X1 U21291 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18160), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18410), .A(n18159), .ZN(
        n18161) );
  OAI211_X1 U21292 ( .C1(n18163), .C2(n18344), .A(n18162), .B(n18161), .ZN(
        P3_U2839) );
  INV_X1 U21293 ( .A(n18317), .ZN(n18306) );
  AOI22_X1 U21294 ( .A1(n18306), .A2(n18185), .B1(n18304), .B2(n18164), .ZN(
        n18175) );
  NAND2_X1 U21295 ( .A1(n18401), .A2(n18276), .ZN(n18302) );
  INV_X1 U21296 ( .A(n18302), .ZN(n18217) );
  AOI21_X1 U21297 ( .B1(n18214), .B2(n18165), .A(n18900), .ZN(n18167) );
  AOI22_X1 U21298 ( .A1(n18867), .A2(n18246), .B1(n18296), .B2(n18249), .ZN(
        n18240) );
  OAI21_X1 U21299 ( .B1(n18166), .B2(n18393), .A(n18240), .ZN(n18220) );
  AOI211_X1 U21300 ( .C1(n18890), .C2(n18221), .A(n18167), .B(n18220), .ZN(
        n18195) );
  NAND2_X1 U21301 ( .A1(n18878), .A2(n18201), .ZN(n18168) );
  OAI211_X1 U21302 ( .C1(n18169), .C2(n18217), .A(n18195), .B(n18168), .ZN(
        n18183) );
  AOI211_X1 U21303 ( .C1(n18890), .C2(n18184), .A(n18173), .B(n18183), .ZN(
        n18174) );
  NAND2_X1 U21304 ( .A1(n18171), .A2(n18170), .ZN(n18172) );
  AOI22_X1 U21305 ( .A1(n18175), .A2(n18174), .B1(n18173), .B2(n18172), .ZN(
        n18176) );
  AOI22_X1 U21306 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18404), .B1(
        n18409), .B2(n18176), .ZN(n18178) );
  OAI211_X1 U21307 ( .C1(n18179), .C2(n18344), .A(n18178), .B(n18177), .ZN(
        P3_U2840) );
  NOR2_X1 U21308 ( .A1(n18221), .A2(n18180), .ZN(n18205) );
  NOR2_X1 U21309 ( .A1(n18304), .A2(n18890), .ZN(n18261) );
  INV_X1 U21310 ( .A(n18261), .ZN(n18408) );
  NOR2_X1 U21311 ( .A1(n18181), .A2(n18221), .ZN(n18182) );
  OAI221_X1 U21312 ( .B1(n18898), .B2(n18235), .C1(n18898), .C2(n18182), .A(
        n18409), .ZN(n18192) );
  AOI211_X1 U21313 ( .C1(n18184), .C2(n18408), .A(n18192), .B(n18183), .ZN(
        n18186) );
  NOR3_X1 U21314 ( .A1(n18308), .A2(n18186), .A3(n18185), .ZN(n18187) );
  AOI21_X1 U21315 ( .B1(n18205), .B2(n18188), .A(n18187), .ZN(n18190) );
  OAI211_X1 U21316 ( .C1(n18191), .C2(n18344), .A(n18190), .B(n18189), .ZN(
        P3_U2841) );
  NOR2_X1 U21317 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18931), .ZN(
        n18196) );
  AOI21_X1 U21318 ( .B1(n18193), .B2(n18302), .A(n18192), .ZN(n18194) );
  AOI21_X1 U21319 ( .B1(n18195), .B2(n18194), .A(n18308), .ZN(n18206) );
  AOI21_X1 U21320 ( .B1(n18196), .B2(n18408), .A(n18206), .ZN(n18202) );
  AOI22_X1 U21321 ( .A1(n18325), .A2(n18198), .B1(n18205), .B2(n18197), .ZN(
        n18200) );
  OAI211_X1 U21322 ( .C1(n18202), .C2(n18201), .A(n18200), .B(n18199), .ZN(
        P3_U2842) );
  NOR2_X1 U21323 ( .A1(n18426), .A2(n18996), .ZN(n18203) );
  AOI221_X1 U21324 ( .B1(n18206), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), 
        .C1(n18205), .C2(n18204), .A(n18203), .ZN(n18207) );
  OAI21_X1 U21325 ( .B1(n18208), .B2(n18344), .A(n18207), .ZN(P3_U2843) );
  NAND2_X1 U21326 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18375) );
  INV_X1 U21327 ( .A(n18209), .ZN(n18395) );
  OAI22_X1 U21328 ( .A1(n18372), .A2(n18393), .B1(n18375), .B2(n18395), .ZN(
        n18383) );
  NAND3_X1 U21329 ( .A1(n18210), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18383), .ZN(n18347) );
  NOR2_X1 U21330 ( .A1(n18213), .A2(n18329), .ZN(n18234) );
  NOR2_X1 U21331 ( .A1(n18898), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18398) );
  INV_X1 U21332 ( .A(n18214), .ZN(n18215) );
  NOR3_X1 U21333 ( .A1(n18398), .A2(n18215), .A3(n18233), .ZN(n18216) );
  OAI22_X1 U21334 ( .A1(n18218), .A2(n18217), .B1(n18394), .B2(n18216), .ZN(
        n18219) );
  NOR3_X1 U21335 ( .A1(n18427), .A2(n18220), .A3(n18219), .ZN(n18227) );
  AOI221_X1 U21336 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18227), 
        .C1(n18394), .C2(n18227), .A(n18221), .ZN(n18222) );
  AOI22_X1 U21337 ( .A1(n18234), .A2(n18223), .B1(n18222), .B2(n18426), .ZN(
        n18225) );
  OAI211_X1 U21338 ( .C1(n18226), .C2(n18344), .A(n18225), .B(n18224), .ZN(
        P3_U2844) );
  NOR2_X1 U21339 ( .A1(n18416), .A2(n18227), .ZN(n18229) );
  AOI22_X1 U21340 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18229), .B1(
        n18234), .B2(n18228), .ZN(n18231) );
  OAI211_X1 U21341 ( .C1(n18232), .C2(n18344), .A(n18231), .B(n18230), .ZN(
        P3_U2845) );
  AOI22_X1 U21342 ( .A1(n18308), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18234), 
        .B2(n18233), .ZN(n18244) );
  AOI21_X1 U21343 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18898), .A(
        n18235), .ZN(n18238) );
  OAI22_X1 U21344 ( .A1(n18900), .A2(n18237), .B1(n18236), .B2(n18393), .ZN(
        n18298) );
  AOI211_X1 U21345 ( .C1(n18306), .C2(n18239), .A(n18238), .B(n18298), .ZN(
        n18253) );
  OAI211_X1 U21346 ( .C1(n18241), .C2(n18253), .A(n18409), .B(n18240), .ZN(
        n18242) );
  NAND3_X1 U21347 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18426), .A3(
        n18242), .ZN(n18243) );
  OAI211_X1 U21348 ( .C1(n18245), .C2(n18344), .A(n18244), .B(n18243), .ZN(
        P3_U2846) );
  NAND2_X1 U21349 ( .A1(n18425), .A2(n18246), .ZN(n18258) );
  AOI21_X1 U21350 ( .B1(n18404), .B2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n18247), .ZN(n18257) );
  AOI21_X1 U21351 ( .B1(n18248), .B2(n18265), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18252) );
  NAND2_X1 U21352 ( .A1(n18296), .A2(n18249), .ZN(n18250) );
  OAI22_X1 U21353 ( .A1(n18253), .A2(n18252), .B1(n18251), .B2(n18250), .ZN(
        n18255) );
  AOI22_X1 U21354 ( .A1(n18409), .A2(n18255), .B1(n18325), .B2(n18254), .ZN(
        n18256) );
  OAI211_X1 U21355 ( .C1(n18259), .C2(n18258), .A(n18257), .B(n18256), .ZN(
        P3_U2847) );
  AOI21_X1 U21356 ( .B1(n18404), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n18260), .ZN(n18273) );
  OAI21_X1 U21357 ( .B1(n18287), .B2(n18299), .A(n18304), .ZN(n18280) );
  OAI21_X1 U21358 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18261), .A(
        n18280), .ZN(n18262) );
  AOI211_X1 U21359 ( .C1(n18306), .C2(n18263), .A(n18298), .B(n18262), .ZN(
        n18269) );
  NOR2_X1 U21360 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18263), .ZN(
        n18264) );
  AOI22_X1 U21361 ( .A1(n18867), .A2(n18266), .B1(n18265), .B2(n18264), .ZN(
        n18267) );
  OAI21_X1 U21362 ( .B1(n18269), .B2(n18268), .A(n18267), .ZN(n18271) );
  AOI22_X1 U21363 ( .A1(n18409), .A2(n18271), .B1(n18340), .B2(n18270), .ZN(
        n18272) );
  OAI211_X1 U21364 ( .C1(n18344), .C2(n18274), .A(n18273), .B(n18272), .ZN(
        P3_U2848) );
  NOR2_X1 U21365 ( .A1(n18305), .A2(n18329), .ZN(n18291) );
  AOI22_X1 U21366 ( .A1(n18308), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18275), 
        .B2(n18291), .ZN(n18283) );
  OAI22_X1 U21367 ( .A1(n18278), .A2(n18401), .B1(n18277), .B2(n18276), .ZN(
        n18279) );
  AOI211_X1 U21368 ( .C1(n18306), .C2(n18305), .A(n18298), .B(n18279), .ZN(
        n18288) );
  OAI211_X1 U21369 ( .C1(n18317), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18288), .B(n18280), .ZN(n18281) );
  OAI211_X1 U21370 ( .C1(n18427), .C2(n18281), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18426), .ZN(n18282) );
  OAI211_X1 U21371 ( .C1(n18284), .C2(n18344), .A(n18283), .B(n18282), .ZN(
        P3_U2849) );
  INV_X1 U21372 ( .A(n18285), .ZN(n18286) );
  AOI22_X1 U21373 ( .A1(n18308), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n18325), 
        .B2(n18286), .ZN(n18293) );
  NOR2_X1 U21374 ( .A1(n18287), .A2(n18299), .ZN(n18289) );
  OAI211_X1 U21375 ( .C1(n18289), .C2(n18898), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18288), .ZN(n18290) );
  OAI211_X1 U21376 ( .C1(n18291), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18409), .B(n18290), .ZN(n18292) );
  OAI211_X1 U21377 ( .C1(n18410), .C2(n18294), .A(n18293), .B(n18292), .ZN(
        P3_U2850) );
  AOI22_X1 U21378 ( .A1(n18867), .A2(n18297), .B1(n18296), .B2(n18295), .ZN(
        n18301) );
  AOI211_X1 U21379 ( .C1(n18304), .C2(n18299), .A(n18427), .B(n18298), .ZN(
        n18300) );
  NAND2_X1 U21380 ( .A1(n18301), .A2(n18300), .ZN(n18323) );
  AOI221_X1 U21381 ( .B1(n18304), .B2(n18303), .C1(n18302), .C2(n18303), .A(
        n18323), .ZN(n18316) );
  NAND2_X1 U21382 ( .A1(n18306), .A2(n18305), .ZN(n18309) );
  AOI211_X1 U21383 ( .C1(n18316), .C2(n18309), .A(n18308), .B(n18307), .ZN(
        n18310) );
  AOI21_X1 U21384 ( .B1(n18325), .B2(n18311), .A(n18310), .ZN(n18313) );
  OAI211_X1 U21385 ( .C1(n18314), .C2(n18329), .A(n18313), .B(n18312), .ZN(
        P3_U2851) );
  NAND2_X1 U21386 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18315), .ZN(
        n18322) );
  AOI221_X1 U21387 ( .B1(n18317), .B2(n18316), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18316), .A(n18315), .ZN(
        n18318) );
  AOI22_X1 U21388 ( .A1(n18319), .A2(n18325), .B1(n18318), .B2(n18426), .ZN(
        n18321) );
  OAI211_X1 U21389 ( .C1(n18322), .C2(n18329), .A(n18321), .B(n18320), .ZN(
        P3_U2852) );
  NAND2_X1 U21390 ( .A1(n18426), .A2(n18323), .ZN(n18327) );
  AOI22_X1 U21391 ( .A1(n18308), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18325), 
        .B2(n18324), .ZN(n18326) );
  OAI221_X1 U21392 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18329), .C1(
        n18328), .C2(n18327), .A(n18326), .ZN(P3_U2853) );
  INV_X1 U21393 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18354) );
  NOR3_X1 U21394 ( .A1(n18354), .A2(n18427), .A3(n18347), .ZN(n18338) );
  AOI21_X1 U21395 ( .B1(n18330), .B2(n18374), .A(n18398), .ZN(n18331) );
  OAI21_X1 U21396 ( .B1(n18332), .B2(n18393), .A(n18331), .ZN(n18356) );
  AOI211_X1 U21397 ( .C1(n18334), .C2(n18333), .A(n18354), .B(n18356), .ZN(
        n18346) );
  OAI21_X1 U21398 ( .B1(n18346), .B2(n18411), .A(n18410), .ZN(n18336) );
  NOR2_X1 U21399 ( .A1(n18426), .A2(n18975), .ZN(n18335) );
  AOI221_X1 U21400 ( .B1(n18338), .B2(n18337), .C1(n18336), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18335), .ZN(n18343) );
  AOI22_X1 U21401 ( .A1(n18425), .A2(n18341), .B1(n18340), .B2(n18339), .ZN(
        n18342) );
  OAI211_X1 U21402 ( .C1(n18345), .C2(n18344), .A(n18343), .B(n18342), .ZN(
        P3_U2854) );
  AOI211_X1 U21403 ( .C1(n18354), .C2(n18347), .A(n18346), .B(n18427), .ZN(
        n18351) );
  OAI22_X1 U21404 ( .A1(n18420), .A2(n18349), .B1(n18385), .B2(n18348), .ZN(
        n18350) );
  NOR2_X1 U21405 ( .A1(n18351), .A2(n18350), .ZN(n18353) );
  NAND2_X1 U21406 ( .A1(n18416), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n18352) );
  OAI211_X1 U21407 ( .C1(n18410), .C2(n18354), .A(n18353), .B(n18352), .ZN(
        P3_U2855) );
  NOR2_X1 U21408 ( .A1(n18426), .A2(n18970), .ZN(n18360) );
  NAND3_X1 U21409 ( .A1(n18409), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18383), .ZN(n18377) );
  NOR2_X1 U21410 ( .A1(n18355), .A2(n18377), .ZN(n18358) );
  OAI21_X1 U21411 ( .B1(n18427), .B2(n18356), .A(n18426), .ZN(n18365) );
  INV_X1 U21412 ( .A(n18365), .ZN(n18357) );
  MUX2_X1 U21413 ( .A(n18358), .B(n18357), .S(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n18359) );
  AOI211_X1 U21414 ( .C1(n18425), .C2(n18361), .A(n18360), .B(n18359), .ZN(
        n18362) );
  OAI21_X1 U21415 ( .B1(n18420), .B2(n18363), .A(n18362), .ZN(P3_U2856) );
  NOR2_X1 U21416 ( .A1(n18377), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18368) );
  INV_X1 U21417 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18366) );
  OAI22_X1 U21418 ( .A1(n18366), .A2(n18365), .B1(n18420), .B2(n18364), .ZN(
        n18367) );
  AOI21_X1 U21419 ( .B1(n18368), .B2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n18367), .ZN(n18370) );
  NAND2_X1 U21420 ( .A1(n18416), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18369) );
  OAI211_X1 U21421 ( .C1(n18371), .C2(n18385), .A(n18370), .B(n18369), .ZN(
        P3_U2857) );
  NAND2_X1 U21422 ( .A1(n18890), .A2(n18372), .ZN(n18399) );
  NAND2_X1 U21423 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18399), .ZN(
        n18373) );
  AOI211_X1 U21424 ( .C1(n18375), .C2(n18374), .A(n18398), .B(n18373), .ZN(
        n18387) );
  OAI21_X1 U21425 ( .B1(n18387), .B2(n18411), .A(n18410), .ZN(n18379) );
  OAI22_X1 U21426 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18377), .B1(
        n18376), .B2(n18385), .ZN(n18378) );
  AOI21_X1 U21427 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18379), .A(
        n18378), .ZN(n18381) );
  NAND2_X1 U21428 ( .A1(n18416), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18380) );
  OAI211_X1 U21429 ( .C1(n18420), .C2(n18382), .A(n18381), .B(n18380), .ZN(
        P3_U2858) );
  OAI21_X1 U21430 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18383), .A(
        n18409), .ZN(n18386) );
  OAI22_X1 U21431 ( .A1(n18387), .A2(n18386), .B1(n18385), .B2(n18384), .ZN(
        n18388) );
  AOI21_X1 U21432 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18404), .A(
        n18388), .ZN(n18390) );
  OAI211_X1 U21433 ( .C1(n18420), .C2(n18391), .A(n18390), .B(n18389), .ZN(
        P3_U2859) );
  NAND2_X1 U21434 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18392) );
  OAI22_X1 U21435 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18392), .ZN(n18397) );
  NOR3_X1 U21436 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19044), .A3(
        n18395), .ZN(n18396) );
  AOI221_X1 U21437 ( .B1(n18398), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18397), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n18396), .ZN(
        n18400) );
  OAI211_X1 U21438 ( .C1(n18402), .C2(n18401), .A(n18400), .B(n18399), .ZN(
        n18403) );
  AOI22_X1 U21439 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18404), .B1(
        n18409), .B2(n18403), .ZN(n18406) );
  OAI211_X1 U21440 ( .C1(n18420), .C2(n18407), .A(n18406), .B(n18405), .ZN(
        P3_U2860) );
  NAND3_X1 U21441 ( .A1(n18409), .A2(n19061), .A3(n18408), .ZN(n18429) );
  AOI21_X1 U21442 ( .B1(n18410), .B2(n18429), .A(n19044), .ZN(n18414) );
  NOR3_X1 U21443 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18412), .A3(
        n18411), .ZN(n18413) );
  AOI211_X1 U21444 ( .C1(n18425), .C2(n18415), .A(n18414), .B(n18413), .ZN(
        n18418) );
  NAND2_X1 U21445 ( .A1(n18416), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18417) );
  OAI211_X1 U21446 ( .C1(n18420), .C2(n18419), .A(n18418), .B(n18417), .ZN(
        P3_U2861) );
  INV_X1 U21447 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19072) );
  NOR2_X1 U21448 ( .A1(n18426), .A2(n19072), .ZN(n18421) );
  AOI221_X1 U21449 ( .B1(n18425), .B2(n18424), .C1(n18423), .C2(n18422), .A(
        n18421), .ZN(n18430) );
  OAI211_X1 U21450 ( .C1(n18878), .C2(n18427), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18426), .ZN(n18428) );
  NAND3_X1 U21451 ( .A1(n18430), .A2(n18429), .A3(n18428), .ZN(P3_U2862) );
  AOI211_X1 U21452 ( .C1(n18432), .C2(n18431), .A(n18931), .B(n19042), .ZN(
        n18924) );
  INV_X1 U21453 ( .A(n18433), .ZN(n18487) );
  OAI21_X1 U21454 ( .B1(n18924), .B2(n18487), .A(n18438), .ZN(n18434) );
  OAI221_X1 U21455 ( .B1(n18903), .B2(n19078), .C1(n18903), .C2(n18438), .A(
        n18434), .ZN(P3_U2863) );
  INV_X1 U21456 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18913) );
  NAND2_X1 U21457 ( .A1(n18910), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18712) );
  INV_X1 U21458 ( .A(n18712), .ZN(n18734) );
  NAND2_X1 U21459 ( .A1(n18913), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18598) );
  INV_X1 U21460 ( .A(n18598), .ZN(n18623) );
  NOR2_X1 U21461 ( .A1(n18734), .A2(n18623), .ZN(n18436) );
  OAI22_X1 U21462 ( .A1(n18437), .A2(n18913), .B1(n18436), .B2(n18435), .ZN(
        P3_U2866) );
  NOR2_X1 U21463 ( .A1(n18914), .A2(n18438), .ZN(P3_U2867) );
  NOR2_X1 U21464 ( .A1(n18440), .A2(n18439), .ZN(n18479) );
  NAND2_X1 U21465 ( .A1(n18479), .A2(n18441), .ZN(n18819) );
  NOR2_X1 U21466 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18554) );
  INV_X1 U21467 ( .A(n18554), .ZN(n18906) );
  NAND2_X1 U21468 ( .A1(n18910), .A2(n18913), .ZN(n18531) );
  NOR2_X2 U21469 ( .A1(n18906), .A2(n18531), .ZN(n18550) );
  INV_X1 U21470 ( .A(n18550), .ZN(n18486) );
  AND2_X1 U21471 ( .A1(n18739), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18810) );
  NOR2_X1 U21472 ( .A1(n18913), .A2(n18621), .ZN(n18813) );
  NAND2_X1 U21473 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18813), .ZN(
        n18865) );
  INV_X1 U21474 ( .A(n18809), .ZN(n18933) );
  AOI21_X1 U21475 ( .B1(n18865), .B2(n18486), .A(n18933), .ZN(n18481) );
  NOR2_X2 U21476 ( .A1(n18442), .A2(n18482), .ZN(n18816) );
  NAND2_X1 U21477 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18444) );
  NOR2_X1 U21478 ( .A1(n18444), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18814) );
  NAND2_X1 U21479 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18814), .ZN(
        n18784) );
  INV_X1 U21480 ( .A(n18784), .ZN(n18856) );
  AOI22_X1 U21481 ( .A1(n18810), .A2(n18481), .B1(n18816), .B2(n18856), .ZN(
        n18447) );
  NAND2_X1 U21482 ( .A1(n18903), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18689) );
  INV_X1 U21483 ( .A(n18689), .ZN(n18445) );
  NOR2_X1 U21484 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18903), .ZN(
        n18666) );
  NOR2_X1 U21485 ( .A1(n18445), .A2(n18666), .ZN(n18737) );
  NOR2_X1 U21486 ( .A1(n18737), .A2(n18444), .ZN(n18788) );
  OAI21_X1 U21487 ( .B1(n19034), .B2(n18903), .A(n18739), .ZN(n18508) );
  AOI21_X1 U21488 ( .B1(n18865), .B2(n18486), .A(n18508), .ZN(n18510) );
  AOI21_X1 U21489 ( .B1(n18815), .B2(n18788), .A(n18510), .ZN(n18483) );
  NOR2_X2 U21490 ( .A1(n18482), .A2(n18443), .ZN(n18811) );
  INV_X1 U21491 ( .A(n18444), .ZN(n18763) );
  NAND2_X1 U21492 ( .A1(n18445), .A2(n18763), .ZN(n18808) );
  INV_X1 U21493 ( .A(n18808), .ZN(n18504) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18483), .B1(
        n18811), .B2(n18504), .ZN(n18446) );
  OAI211_X1 U21495 ( .C1(n18819), .C2(n18486), .A(n18447), .B(n18446), .ZN(
        P3_U2868) );
  NAND2_X1 U21496 ( .A1(n18479), .A2(n18448), .ZN(n18825) );
  NOR2_X2 U21497 ( .A1(n18482), .A2(n18449), .ZN(n18822) );
  AND2_X1 U21498 ( .A1(n18739), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18820) );
  AOI22_X1 U21499 ( .A1(n18822), .A2(n18504), .B1(n18820), .B2(n18481), .ZN(
        n18451) );
  AND2_X1 U21500 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18815), .ZN(n18821) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18483), .B1(
        n18821), .B2(n18856), .ZN(n18450) );
  OAI211_X1 U21502 ( .C1(n18825), .C2(n18486), .A(n18451), .B(n18450), .ZN(
        P3_U2869) );
  NAND2_X1 U21503 ( .A1(n18479), .A2(n18452), .ZN(n18831) );
  INV_X1 U21504 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18453) );
  NOR2_X2 U21505 ( .A1(n18453), .A2(n18482), .ZN(n18827) );
  NOR2_X2 U21506 ( .A1(n18454), .A2(n18488), .ZN(n18826) );
  AOI22_X1 U21507 ( .A1(n18827), .A2(n18504), .B1(n18826), .B2(n18481), .ZN(
        n18456) );
  NOR2_X2 U21508 ( .A1(n19438), .A2(n18482), .ZN(n18828) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18483), .B1(
        n18828), .B2(n18856), .ZN(n18455) );
  OAI211_X1 U21510 ( .C1(n18831), .C2(n18486), .A(n18456), .B(n18455), .ZN(
        P3_U2870) );
  NAND2_X1 U21511 ( .A1(n18479), .A2(n18457), .ZN(n18837) );
  AND2_X1 U21512 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18815), .ZN(n18834) );
  NOR2_X2 U21513 ( .A1(n18458), .A2(n18488), .ZN(n18833) );
  AOI22_X1 U21514 ( .A1(n18834), .A2(n18856), .B1(n18833), .B2(n18481), .ZN(
        n18461) );
  NOR2_X2 U21515 ( .A1(n18459), .A2(n18482), .ZN(n18832) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18483), .B1(
        n18832), .B2(n18504), .ZN(n18460) );
  OAI211_X1 U21517 ( .C1(n18837), .C2(n18486), .A(n18461), .B(n18460), .ZN(
        P3_U2871) );
  NAND2_X1 U21518 ( .A1(n18479), .A2(n18462), .ZN(n18843) );
  NOR2_X2 U21519 ( .A1(n19450), .A2(n18482), .ZN(n18839) );
  NOR2_X2 U21520 ( .A1(n18463), .A2(n18488), .ZN(n18838) );
  AOI22_X1 U21521 ( .A1(n18839), .A2(n18856), .B1(n18838), .B2(n18481), .ZN(
        n18466) );
  NOR2_X2 U21522 ( .A1(n18464), .A2(n18482), .ZN(n18840) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18483), .B1(
        n18840), .B2(n18504), .ZN(n18465) );
  OAI211_X1 U21524 ( .C1(n18843), .C2(n18486), .A(n18466), .B(n18465), .ZN(
        P3_U2872) );
  NAND2_X1 U21525 ( .A1(n18479), .A2(n18467), .ZN(n18849) );
  INV_X1 U21526 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18468) );
  NOR2_X2 U21527 ( .A1(n18468), .A2(n18482), .ZN(n18845) );
  NOR2_X2 U21528 ( .A1(n18469), .A2(n18488), .ZN(n18844) );
  AOI22_X1 U21529 ( .A1(n18845), .A2(n18856), .B1(n18844), .B2(n18481), .ZN(
        n18472) );
  NOR2_X2 U21530 ( .A1(n18470), .A2(n18482), .ZN(n18846) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18483), .B1(
        n18846), .B2(n18504), .ZN(n18471) );
  OAI211_X1 U21532 ( .C1(n18849), .C2(n18486), .A(n18472), .B(n18471), .ZN(
        P3_U2873) );
  NAND2_X1 U21533 ( .A1(n18479), .A2(n18473), .ZN(n18855) );
  AND2_X1 U21534 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18815), .ZN(n18851) );
  NOR2_X2 U21535 ( .A1(n18474), .A2(n18488), .ZN(n18850) );
  AOI22_X1 U21536 ( .A1(n18851), .A2(n18504), .B1(n18850), .B2(n18481), .ZN(
        n18477) );
  INV_X1 U21537 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18475) );
  NOR2_X2 U21538 ( .A1(n18475), .A2(n18482), .ZN(n18852) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18483), .B1(
        n18852), .B2(n18856), .ZN(n18476) );
  OAI211_X1 U21540 ( .C1(n18855), .C2(n18486), .A(n18477), .B(n18476), .ZN(
        P3_U2874) );
  NAND2_X1 U21541 ( .A1(n18479), .A2(n18478), .ZN(n18866) );
  AND2_X1 U21542 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18739), .ZN(n18859) );
  INV_X1 U21543 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18480) );
  NOR2_X2 U21544 ( .A1(n18480), .A2(n18482), .ZN(n18857) );
  AOI22_X1 U21545 ( .A1(n18859), .A2(n18481), .B1(n18857), .B2(n18504), .ZN(
        n18485) );
  NOR2_X2 U21546 ( .A1(n19457), .A2(n18482), .ZN(n18861) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18483), .B1(
        n18861), .B2(n18856), .ZN(n18484) );
  OAI211_X1 U21548 ( .C1(n18866), .C2(n18486), .A(n18485), .B(n18484), .ZN(
        P3_U2875) );
  INV_X1 U21549 ( .A(n18531), .ZN(n18533) );
  NAND2_X1 U21550 ( .A1(n18666), .A2(n18533), .ZN(n18534) );
  INV_X1 U21551 ( .A(n18865), .ZN(n18526) );
  NAND2_X1 U21552 ( .A1(n18905), .A2(n18809), .ZN(n18668) );
  NOR2_X1 U21553 ( .A1(n18531), .A2(n18668), .ZN(n18503) );
  AOI22_X1 U21554 ( .A1(n18811), .A2(n18526), .B1(n18810), .B2(n18503), .ZN(
        n18490) );
  NOR2_X1 U21555 ( .A1(n18488), .A2(n18487), .ZN(n18812) );
  INV_X1 U21556 ( .A(n18812), .ZN(n18532) );
  NOR2_X1 U21557 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18532), .ZN(
        n18762) );
  AOI22_X1 U21558 ( .A1(n18815), .A2(n18813), .B1(n18533), .B2(n18762), .ZN(
        n18505) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18505), .B1(
        n18816), .B2(n18504), .ZN(n18489) );
  OAI211_X1 U21560 ( .C1(n18819), .C2(n18534), .A(n18490), .B(n18489), .ZN(
        P3_U2876) );
  AOI22_X1 U21561 ( .A1(n18822), .A2(n18526), .B1(n18820), .B2(n18503), .ZN(
        n18492) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18505), .B1(
        n18821), .B2(n18504), .ZN(n18491) );
  OAI211_X1 U21563 ( .C1(n18825), .C2(n18534), .A(n18492), .B(n18491), .ZN(
        P3_U2877) );
  AOI22_X1 U21564 ( .A1(n18828), .A2(n18504), .B1(n18826), .B2(n18503), .ZN(
        n18494) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18505), .B1(
        n18827), .B2(n18526), .ZN(n18493) );
  OAI211_X1 U21566 ( .C1(n18831), .C2(n18534), .A(n18494), .B(n18493), .ZN(
        P3_U2878) );
  AOI22_X1 U21567 ( .A1(n18834), .A2(n18504), .B1(n18833), .B2(n18503), .ZN(
        n18496) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18505), .B1(
        n18832), .B2(n18526), .ZN(n18495) );
  OAI211_X1 U21569 ( .C1(n18837), .C2(n18534), .A(n18496), .B(n18495), .ZN(
        P3_U2879) );
  AOI22_X1 U21570 ( .A1(n18840), .A2(n18526), .B1(n18838), .B2(n18503), .ZN(
        n18498) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18505), .B1(
        n18839), .B2(n18504), .ZN(n18497) );
  OAI211_X1 U21572 ( .C1(n18843), .C2(n18534), .A(n18498), .B(n18497), .ZN(
        P3_U2880) );
  AOI22_X1 U21573 ( .A1(n18844), .A2(n18503), .B1(n18846), .B2(n18526), .ZN(
        n18500) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18505), .B1(
        n18845), .B2(n18504), .ZN(n18499) );
  OAI211_X1 U21575 ( .C1(n18849), .C2(n18534), .A(n18500), .B(n18499), .ZN(
        P3_U2881) );
  AOI22_X1 U21576 ( .A1(n18851), .A2(n18526), .B1(n18850), .B2(n18503), .ZN(
        n18502) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18505), .B1(
        n18852), .B2(n18504), .ZN(n18501) );
  OAI211_X1 U21578 ( .C1(n18855), .C2(n18534), .A(n18502), .B(n18501), .ZN(
        P3_U2882) );
  AOI22_X1 U21579 ( .A1(n18861), .A2(n18504), .B1(n18859), .B2(n18503), .ZN(
        n18507) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18505), .B1(
        n18857), .B2(n18526), .ZN(n18506) );
  OAI211_X1 U21581 ( .C1(n18866), .C2(n18534), .A(n18507), .B(n18506), .ZN(
        P3_U2883) );
  NOR2_X2 U21582 ( .A1(n18689), .A2(n18531), .ZN(n18594) );
  INV_X1 U21583 ( .A(n18594), .ZN(n18530) );
  NAND2_X1 U21584 ( .A1(n18534), .A2(n18530), .ZN(n18509) );
  INV_X1 U21585 ( .A(n18509), .ZN(n18556) );
  NOR2_X1 U21586 ( .A1(n18933), .A2(n18556), .ZN(n18525) );
  AOI22_X1 U21587 ( .A1(n18811), .A2(n18550), .B1(n18810), .B2(n18525), .ZN(
        n18512) );
  INV_X1 U21588 ( .A(n18508), .ZN(n18785) );
  AOI22_X1 U21589 ( .A1(n18787), .A2(n18510), .B1(n18785), .B2(n18509), .ZN(
        n18527) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18527), .B1(
        n18816), .B2(n18526), .ZN(n18511) );
  OAI211_X1 U21591 ( .C1(n18819), .C2(n18530), .A(n18512), .B(n18511), .ZN(
        P3_U2884) );
  AOI22_X1 U21592 ( .A1(n18821), .A2(n18526), .B1(n18820), .B2(n18525), .ZN(
        n18514) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18527), .B1(
        n18822), .B2(n18550), .ZN(n18513) );
  OAI211_X1 U21594 ( .C1(n18825), .C2(n18530), .A(n18514), .B(n18513), .ZN(
        P3_U2885) );
  AOI22_X1 U21595 ( .A1(n18827), .A2(n18550), .B1(n18826), .B2(n18525), .ZN(
        n18516) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18527), .B1(
        n18828), .B2(n18526), .ZN(n18515) );
  OAI211_X1 U21597 ( .C1(n18831), .C2(n18530), .A(n18516), .B(n18515), .ZN(
        P3_U2886) );
  AOI22_X1 U21598 ( .A1(n18833), .A2(n18525), .B1(n18832), .B2(n18550), .ZN(
        n18518) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18527), .B1(
        n18834), .B2(n18526), .ZN(n18517) );
  OAI211_X1 U21600 ( .C1(n18837), .C2(n18530), .A(n18518), .B(n18517), .ZN(
        P3_U2887) );
  AOI22_X1 U21601 ( .A1(n18839), .A2(n18526), .B1(n18838), .B2(n18525), .ZN(
        n18520) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18527), .B1(
        n18840), .B2(n18550), .ZN(n18519) );
  OAI211_X1 U21603 ( .C1(n18843), .C2(n18530), .A(n18520), .B(n18519), .ZN(
        P3_U2888) );
  AOI22_X1 U21604 ( .A1(n18844), .A2(n18525), .B1(n18846), .B2(n18550), .ZN(
        n18522) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18527), .B1(
        n18845), .B2(n18526), .ZN(n18521) );
  OAI211_X1 U21606 ( .C1(n18849), .C2(n18530), .A(n18522), .B(n18521), .ZN(
        P3_U2889) );
  AOI22_X1 U21607 ( .A1(n18851), .A2(n18550), .B1(n18850), .B2(n18525), .ZN(
        n18524) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18527), .B1(
        n18852), .B2(n18526), .ZN(n18523) );
  OAI211_X1 U21609 ( .C1(n18855), .C2(n18530), .A(n18524), .B(n18523), .ZN(
        P3_U2890) );
  AOI22_X1 U21610 ( .A1(n18861), .A2(n18526), .B1(n18859), .B2(n18525), .ZN(
        n18529) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18527), .B1(
        n18857), .B2(n18550), .ZN(n18528) );
  OAI211_X1 U21612 ( .C1(n18866), .C2(n18530), .A(n18529), .B(n18528), .ZN(
        P3_U2891) );
  NOR2_X1 U21613 ( .A1(n18905), .A2(n18531), .ZN(n18578) );
  NAND2_X1 U21614 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18578), .ZN(
        n18555) );
  AND2_X1 U21615 ( .A1(n18809), .A2(n18578), .ZN(n18549) );
  AOI22_X1 U21616 ( .A1(n18810), .A2(n18549), .B1(n18816), .B2(n18550), .ZN(
        n18536) );
  AOI21_X1 U21617 ( .B1(n18905), .B2(n18599), .A(n18532), .ZN(n18622) );
  NAND2_X1 U21618 ( .A1(n18533), .A2(n18622), .ZN(n18551) );
  INV_X1 U21619 ( .A(n18534), .ZN(n18573) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18551), .B1(
        n18811), .B2(n18573), .ZN(n18535) );
  OAI211_X1 U21621 ( .C1(n18555), .C2(n18819), .A(n18536), .B(n18535), .ZN(
        P3_U2892) );
  AOI22_X1 U21622 ( .A1(n18821), .A2(n18550), .B1(n18820), .B2(n18549), .ZN(
        n18538) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18551), .B1(
        n18822), .B2(n18573), .ZN(n18537) );
  OAI211_X1 U21624 ( .C1(n18555), .C2(n18825), .A(n18538), .B(n18537), .ZN(
        P3_U2893) );
  AOI22_X1 U21625 ( .A1(n18828), .A2(n18550), .B1(n18826), .B2(n18549), .ZN(
        n18540) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18551), .B1(
        n18827), .B2(n18573), .ZN(n18539) );
  OAI211_X1 U21627 ( .C1(n18555), .C2(n18831), .A(n18540), .B(n18539), .ZN(
        P3_U2894) );
  AOI22_X1 U21628 ( .A1(n18833), .A2(n18549), .B1(n18832), .B2(n18573), .ZN(
        n18542) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18551), .B1(
        n18834), .B2(n18550), .ZN(n18541) );
  OAI211_X1 U21630 ( .C1(n18555), .C2(n18837), .A(n18542), .B(n18541), .ZN(
        P3_U2895) );
  AOI22_X1 U21631 ( .A1(n18839), .A2(n18550), .B1(n18838), .B2(n18549), .ZN(
        n18544) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18551), .B1(
        n18840), .B2(n18573), .ZN(n18543) );
  OAI211_X1 U21633 ( .C1(n18555), .C2(n18843), .A(n18544), .B(n18543), .ZN(
        P3_U2896) );
  AOI22_X1 U21634 ( .A1(n18844), .A2(n18549), .B1(n18846), .B2(n18573), .ZN(
        n18546) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18551), .B1(
        n18845), .B2(n18550), .ZN(n18545) );
  OAI211_X1 U21636 ( .C1(n18555), .C2(n18849), .A(n18546), .B(n18545), .ZN(
        P3_U2897) );
  AOI22_X1 U21637 ( .A1(n18851), .A2(n18573), .B1(n18850), .B2(n18549), .ZN(
        n18548) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18551), .B1(
        n18852), .B2(n18550), .ZN(n18547) );
  OAI211_X1 U21639 ( .C1(n18555), .C2(n18855), .A(n18548), .B(n18547), .ZN(
        P3_U2898) );
  AOI22_X1 U21640 ( .A1(n18861), .A2(n18550), .B1(n18859), .B2(n18549), .ZN(
        n18553) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18551), .B1(
        n18857), .B2(n18573), .ZN(n18552) );
  OAI211_X1 U21642 ( .C1(n18555), .C2(n18866), .A(n18553), .B(n18552), .ZN(
        P3_U2899) );
  NAND2_X1 U21643 ( .A1(n18554), .A2(n18623), .ZN(n18577) );
  INV_X1 U21644 ( .A(n18577), .ZN(n18639) );
  INV_X1 U21645 ( .A(n18555), .ZN(n18617) );
  NOR2_X1 U21646 ( .A1(n18639), .A2(n18617), .ZN(n18600) );
  NOR2_X1 U21647 ( .A1(n18933), .A2(n18600), .ZN(n18572) );
  AOI22_X1 U21648 ( .A1(n18811), .A2(n18594), .B1(n18810), .B2(n18572), .ZN(
        n18559) );
  AOI221_X1 U21649 ( .B1(n18556), .B2(n18555), .C1(n18599), .C2(n18555), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18557) );
  OAI21_X1 U21650 ( .B1(n18639), .B2(n18557), .A(n18739), .ZN(n18574) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18574), .B1(
        n18816), .B2(n18573), .ZN(n18558) );
  OAI211_X1 U21652 ( .C1(n18577), .C2(n18819), .A(n18559), .B(n18558), .ZN(
        P3_U2900) );
  AOI22_X1 U21653 ( .A1(n18821), .A2(n18573), .B1(n18820), .B2(n18572), .ZN(
        n18561) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18574), .B1(
        n18822), .B2(n18594), .ZN(n18560) );
  OAI211_X1 U21655 ( .C1(n18577), .C2(n18825), .A(n18561), .B(n18560), .ZN(
        P3_U2901) );
  AOI22_X1 U21656 ( .A1(n18827), .A2(n18594), .B1(n18826), .B2(n18572), .ZN(
        n18563) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18574), .B1(
        n18828), .B2(n18573), .ZN(n18562) );
  OAI211_X1 U21658 ( .C1(n18577), .C2(n18831), .A(n18563), .B(n18562), .ZN(
        P3_U2902) );
  AOI22_X1 U21659 ( .A1(n18834), .A2(n18573), .B1(n18833), .B2(n18572), .ZN(
        n18565) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18574), .B1(
        n18832), .B2(n18594), .ZN(n18564) );
  OAI211_X1 U21661 ( .C1(n18577), .C2(n18837), .A(n18565), .B(n18564), .ZN(
        P3_U2903) );
  AOI22_X1 U21662 ( .A1(n18839), .A2(n18573), .B1(n18838), .B2(n18572), .ZN(
        n18567) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18574), .B1(
        n18840), .B2(n18594), .ZN(n18566) );
  OAI211_X1 U21664 ( .C1(n18577), .C2(n18843), .A(n18567), .B(n18566), .ZN(
        P3_U2904) );
  AOI22_X1 U21665 ( .A1(n18845), .A2(n18573), .B1(n18844), .B2(n18572), .ZN(
        n18569) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18574), .B1(
        n18846), .B2(n18594), .ZN(n18568) );
  OAI211_X1 U21667 ( .C1(n18577), .C2(n18849), .A(n18569), .B(n18568), .ZN(
        P3_U2905) );
  AOI22_X1 U21668 ( .A1(n18852), .A2(n18573), .B1(n18850), .B2(n18572), .ZN(
        n18571) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18574), .B1(
        n18851), .B2(n18594), .ZN(n18570) );
  OAI211_X1 U21670 ( .C1(n18577), .C2(n18855), .A(n18571), .B(n18570), .ZN(
        P3_U2906) );
  AOI22_X1 U21671 ( .A1(n18859), .A2(n18572), .B1(n18857), .B2(n18594), .ZN(
        n18576) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18574), .B1(
        n18861), .B2(n18573), .ZN(n18575) );
  OAI211_X1 U21673 ( .C1(n18577), .C2(n18866), .A(n18576), .B(n18575), .ZN(
        P3_U2907) );
  NAND2_X1 U21674 ( .A1(n18623), .A2(n18666), .ZN(n18643) );
  NOR2_X1 U21675 ( .A1(n18598), .A2(n18668), .ZN(n18593) );
  AOI22_X1 U21676 ( .A1(n18617), .A2(n18811), .B1(n18810), .B2(n18593), .ZN(
        n18580) );
  AOI22_X1 U21677 ( .A1(n18815), .A2(n18578), .B1(n18623), .B2(n18762), .ZN(
        n18595) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18595), .B1(
        n18816), .B2(n18594), .ZN(n18579) );
  OAI211_X1 U21679 ( .C1(n18643), .C2(n18819), .A(n18580), .B(n18579), .ZN(
        P3_U2908) );
  AOI22_X1 U21680 ( .A1(n18617), .A2(n18822), .B1(n18820), .B2(n18593), .ZN(
        n18582) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18595), .B1(
        n18821), .B2(n18594), .ZN(n18581) );
  OAI211_X1 U21682 ( .C1(n18643), .C2(n18825), .A(n18582), .B(n18581), .ZN(
        P3_U2909) );
  AOI22_X1 U21683 ( .A1(n18617), .A2(n18827), .B1(n18826), .B2(n18593), .ZN(
        n18584) );
  AOI22_X1 U21684 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18595), .B1(
        n18828), .B2(n18594), .ZN(n18583) );
  OAI211_X1 U21685 ( .C1(n18643), .C2(n18831), .A(n18584), .B(n18583), .ZN(
        P3_U2910) );
  AOI22_X1 U21686 ( .A1(n18617), .A2(n18832), .B1(n18833), .B2(n18593), .ZN(
        n18586) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18595), .B1(
        n18834), .B2(n18594), .ZN(n18585) );
  OAI211_X1 U21688 ( .C1(n18643), .C2(n18837), .A(n18586), .B(n18585), .ZN(
        P3_U2911) );
  AOI22_X1 U21689 ( .A1(n18617), .A2(n18840), .B1(n18838), .B2(n18593), .ZN(
        n18588) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18595), .B1(
        n18839), .B2(n18594), .ZN(n18587) );
  OAI211_X1 U21691 ( .C1(n18643), .C2(n18843), .A(n18588), .B(n18587), .ZN(
        P3_U2912) );
  AOI22_X1 U21692 ( .A1(n18845), .A2(n18594), .B1(n18844), .B2(n18593), .ZN(
        n18590) );
  AOI22_X1 U21693 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18595), .B1(
        n18617), .B2(n18846), .ZN(n18589) );
  OAI211_X1 U21694 ( .C1(n18643), .C2(n18849), .A(n18590), .B(n18589), .ZN(
        P3_U2913) );
  AOI22_X1 U21695 ( .A1(n18852), .A2(n18594), .B1(n18850), .B2(n18593), .ZN(
        n18592) );
  AOI22_X1 U21696 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18595), .B1(
        n18617), .B2(n18851), .ZN(n18591) );
  OAI211_X1 U21697 ( .C1(n18643), .C2(n18855), .A(n18592), .B(n18591), .ZN(
        P3_U2914) );
  AOI22_X1 U21698 ( .A1(n18861), .A2(n18594), .B1(n18859), .B2(n18593), .ZN(
        n18597) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18595), .B1(
        n18617), .B2(n18857), .ZN(n18596) );
  OAI211_X1 U21700 ( .C1(n18643), .C2(n18866), .A(n18597), .B(n18596), .ZN(
        P3_U2915) );
  NOR2_X2 U21701 ( .A1(n18689), .A2(n18598), .ZN(n18685) );
  INV_X1 U21702 ( .A(n18685), .ZN(n18644) );
  AOI21_X1 U21703 ( .B1(n18644), .B2(n18643), .A(n18933), .ZN(n18616) );
  AOI22_X1 U21704 ( .A1(n18617), .A2(n18816), .B1(n18810), .B2(n18616), .ZN(
        n18603) );
  AOI221_X1 U21705 ( .B1(n18600), .B2(n18643), .C1(n18599), .C2(n18643), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18601) );
  OAI21_X1 U21706 ( .B1(n18685), .B2(n18601), .A(n18739), .ZN(n18618) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18618), .B1(
        n18639), .B2(n18811), .ZN(n18602) );
  OAI211_X1 U21708 ( .C1(n18644), .C2(n18819), .A(n18603), .B(n18602), .ZN(
        P3_U2916) );
  AOI22_X1 U21709 ( .A1(n18617), .A2(n18821), .B1(n18616), .B2(n18820), .ZN(
        n18605) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18618), .B1(
        n18639), .B2(n18822), .ZN(n18604) );
  OAI211_X1 U21711 ( .C1(n18644), .C2(n18825), .A(n18605), .B(n18604), .ZN(
        P3_U2917) );
  AOI22_X1 U21712 ( .A1(n18617), .A2(n18828), .B1(n18616), .B2(n18826), .ZN(
        n18607) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18618), .B1(
        n18639), .B2(n18827), .ZN(n18606) );
  OAI211_X1 U21714 ( .C1(n18644), .C2(n18831), .A(n18607), .B(n18606), .ZN(
        P3_U2918) );
  AOI22_X1 U21715 ( .A1(n18639), .A2(n18832), .B1(n18616), .B2(n18833), .ZN(
        n18609) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18618), .B1(
        n18617), .B2(n18834), .ZN(n18608) );
  OAI211_X1 U21717 ( .C1(n18644), .C2(n18837), .A(n18609), .B(n18608), .ZN(
        P3_U2919) );
  AOI22_X1 U21718 ( .A1(n18617), .A2(n18839), .B1(n18616), .B2(n18838), .ZN(
        n18611) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18618), .B1(
        n18639), .B2(n18840), .ZN(n18610) );
  OAI211_X1 U21720 ( .C1(n18644), .C2(n18843), .A(n18611), .B(n18610), .ZN(
        P3_U2920) );
  AOI22_X1 U21721 ( .A1(n18639), .A2(n18846), .B1(n18616), .B2(n18844), .ZN(
        n18613) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18618), .B1(
        n18617), .B2(n18845), .ZN(n18612) );
  OAI211_X1 U21723 ( .C1(n18644), .C2(n18849), .A(n18613), .B(n18612), .ZN(
        P3_U2921) );
  AOI22_X1 U21724 ( .A1(n18617), .A2(n18852), .B1(n18616), .B2(n18850), .ZN(
        n18615) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18618), .B1(
        n18639), .B2(n18851), .ZN(n18614) );
  OAI211_X1 U21726 ( .C1(n18644), .C2(n18855), .A(n18615), .B(n18614), .ZN(
        P3_U2922) );
  AOI22_X1 U21727 ( .A1(n18639), .A2(n18857), .B1(n18616), .B2(n18859), .ZN(
        n18620) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18618), .B1(
        n18617), .B2(n18861), .ZN(n18619) );
  OAI211_X1 U21729 ( .C1(n18644), .C2(n18866), .A(n18620), .B(n18619), .ZN(
        P3_U2923) );
  NOR2_X1 U21730 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18621), .ZN(
        n18669) );
  NAND2_X1 U21731 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18669), .ZN(
        n18667) );
  INV_X1 U21732 ( .A(n18643), .ZN(n18662) );
  AOI22_X1 U21733 ( .A1(n18662), .A2(n18811), .B1(n18810), .B2(n18638), .ZN(
        n18625) );
  NAND2_X1 U21734 ( .A1(n18623), .A2(n18622), .ZN(n18640) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18640), .B1(
        n18639), .B2(n18816), .ZN(n18624) );
  OAI211_X1 U21736 ( .C1(n18819), .C2(n18667), .A(n18625), .B(n18624), .ZN(
        P3_U2924) );
  AOI22_X1 U21737 ( .A1(n18662), .A2(n18822), .B1(n18820), .B2(n18638), .ZN(
        n18627) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18640), .B1(
        n18639), .B2(n18821), .ZN(n18626) );
  OAI211_X1 U21739 ( .C1(n18825), .C2(n18667), .A(n18627), .B(n18626), .ZN(
        P3_U2925) );
  AOI22_X1 U21740 ( .A1(n18662), .A2(n18827), .B1(n18826), .B2(n18638), .ZN(
        n18629) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18640), .B1(
        n18639), .B2(n18828), .ZN(n18628) );
  OAI211_X1 U21742 ( .C1(n18831), .C2(n18667), .A(n18629), .B(n18628), .ZN(
        P3_U2926) );
  AOI22_X1 U21743 ( .A1(n18639), .A2(n18834), .B1(n18833), .B2(n18638), .ZN(
        n18631) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18640), .B1(
        n18662), .B2(n18832), .ZN(n18630) );
  OAI211_X1 U21745 ( .C1(n18837), .C2(n18667), .A(n18631), .B(n18630), .ZN(
        P3_U2927) );
  AOI22_X1 U21746 ( .A1(n18662), .A2(n18840), .B1(n18838), .B2(n18638), .ZN(
        n18633) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18640), .B1(
        n18639), .B2(n18839), .ZN(n18632) );
  OAI211_X1 U21748 ( .C1(n18843), .C2(n18667), .A(n18633), .B(n18632), .ZN(
        P3_U2928) );
  AOI22_X1 U21749 ( .A1(n18662), .A2(n18846), .B1(n18844), .B2(n18638), .ZN(
        n18635) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18640), .B1(
        n18639), .B2(n18845), .ZN(n18634) );
  OAI211_X1 U21751 ( .C1(n18849), .C2(n18667), .A(n18635), .B(n18634), .ZN(
        P3_U2929) );
  AOI22_X1 U21752 ( .A1(n18639), .A2(n18852), .B1(n18850), .B2(n18638), .ZN(
        n18637) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18640), .B1(
        n18662), .B2(n18851), .ZN(n18636) );
  OAI211_X1 U21754 ( .C1(n18855), .C2(n18667), .A(n18637), .B(n18636), .ZN(
        P3_U2930) );
  AOI22_X1 U21755 ( .A1(n18662), .A2(n18857), .B1(n18859), .B2(n18638), .ZN(
        n18642) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18640), .B1(
        n18639), .B2(n18861), .ZN(n18641) );
  OAI211_X1 U21757 ( .C1(n18866), .C2(n18667), .A(n18642), .B(n18641), .ZN(
        P3_U2931) );
  NOR2_X2 U21758 ( .A1(n18906), .A2(n18712), .ZN(n18730) );
  INV_X1 U21759 ( .A(n18730), .ZN(n18665) );
  NAND2_X1 U21760 ( .A1(n18667), .A2(n18665), .ZN(n18690) );
  AND2_X1 U21761 ( .A1(n18809), .A2(n18690), .ZN(n18660) );
  AOI22_X1 U21762 ( .A1(n18662), .A2(n18816), .B1(n18810), .B2(n18660), .ZN(
        n18647) );
  NAND2_X1 U21763 ( .A1(n18644), .A2(n18643), .ZN(n18645) );
  OAI221_X1 U21764 ( .B1(n18690), .B2(n18787), .C1(n18690), .C2(n18645), .A(
        n18785), .ZN(n18661) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18661), .B1(
        n18685), .B2(n18811), .ZN(n18646) );
  OAI211_X1 U21766 ( .C1(n18819), .C2(n18665), .A(n18647), .B(n18646), .ZN(
        P3_U2932) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18661), .B1(
        n18820), .B2(n18660), .ZN(n18649) );
  AOI22_X1 U21768 ( .A1(n18685), .A2(n18822), .B1(n18662), .B2(n18821), .ZN(
        n18648) );
  OAI211_X1 U21769 ( .C1(n18825), .C2(n18665), .A(n18649), .B(n18648), .ZN(
        P3_U2933) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18661), .B1(
        n18826), .B2(n18660), .ZN(n18651) );
  AOI22_X1 U21771 ( .A1(n18685), .A2(n18827), .B1(n18662), .B2(n18828), .ZN(
        n18650) );
  OAI211_X1 U21772 ( .C1(n18831), .C2(n18665), .A(n18651), .B(n18650), .ZN(
        P3_U2934) );
  AOI22_X1 U21773 ( .A1(n18662), .A2(n18834), .B1(n18833), .B2(n18660), .ZN(
        n18653) );
  AOI22_X1 U21774 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18661), .B1(
        n18685), .B2(n18832), .ZN(n18652) );
  OAI211_X1 U21775 ( .C1(n18837), .C2(n18665), .A(n18653), .B(n18652), .ZN(
        P3_U2935) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18661), .B1(
        n18838), .B2(n18660), .ZN(n18655) );
  AOI22_X1 U21777 ( .A1(n18685), .A2(n18840), .B1(n18662), .B2(n18839), .ZN(
        n18654) );
  OAI211_X1 U21778 ( .C1(n18843), .C2(n18665), .A(n18655), .B(n18654), .ZN(
        P3_U2936) );
  AOI22_X1 U21779 ( .A1(n18685), .A2(n18846), .B1(n18844), .B2(n18660), .ZN(
        n18657) );
  AOI22_X1 U21780 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18661), .B1(
        n18662), .B2(n18845), .ZN(n18656) );
  OAI211_X1 U21781 ( .C1(n18849), .C2(n18665), .A(n18657), .B(n18656), .ZN(
        P3_U2937) );
  AOI22_X1 U21782 ( .A1(n18685), .A2(n18851), .B1(n18850), .B2(n18660), .ZN(
        n18659) );
  AOI22_X1 U21783 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18661), .B1(
        n18662), .B2(n18852), .ZN(n18658) );
  OAI211_X1 U21784 ( .C1(n18855), .C2(n18665), .A(n18659), .B(n18658), .ZN(
        P3_U2938) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18661), .B1(
        n18859), .B2(n18660), .ZN(n18664) );
  AOI22_X1 U21786 ( .A1(n18685), .A2(n18857), .B1(n18662), .B2(n18861), .ZN(
        n18663) );
  OAI211_X1 U21787 ( .C1(n18866), .C2(n18665), .A(n18664), .B(n18663), .ZN(
        P3_U2939) );
  NAND2_X1 U21788 ( .A1(n18666), .A2(n18734), .ZN(n18714) );
  INV_X1 U21789 ( .A(n18667), .ZN(n18707) );
  NOR2_X1 U21790 ( .A1(n18712), .A2(n18668), .ZN(n18684) );
  AOI22_X1 U21791 ( .A1(n18811), .A2(n18707), .B1(n18810), .B2(n18684), .ZN(
        n18671) );
  NOR2_X1 U21792 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18712), .ZN(
        n18713) );
  AOI22_X1 U21793 ( .A1(n18815), .A2(n18669), .B1(n18812), .B2(n18713), .ZN(
        n18686) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n18816), .ZN(n18670) );
  OAI211_X1 U21795 ( .C1(n18819), .C2(n18714), .A(n18671), .B(n18670), .ZN(
        P3_U2940) );
  AOI22_X1 U21796 ( .A1(n18822), .A2(n18707), .B1(n18820), .B2(n18684), .ZN(
        n18673) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n18821), .ZN(n18672) );
  OAI211_X1 U21798 ( .C1(n18825), .C2(n18714), .A(n18673), .B(n18672), .ZN(
        P3_U2941) );
  AOI22_X1 U21799 ( .A1(n18827), .A2(n18707), .B1(n18826), .B2(n18684), .ZN(
        n18675) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n18828), .ZN(n18674) );
  OAI211_X1 U21801 ( .C1(n18831), .C2(n18714), .A(n18675), .B(n18674), .ZN(
        P3_U2942) );
  AOI22_X1 U21802 ( .A1(n18833), .A2(n18684), .B1(n18832), .B2(n18707), .ZN(
        n18677) );
  AOI22_X1 U21803 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n18834), .ZN(n18676) );
  OAI211_X1 U21804 ( .C1(n18837), .C2(n18714), .A(n18677), .B(n18676), .ZN(
        P3_U2943) );
  AOI22_X1 U21805 ( .A1(n18685), .A2(n18839), .B1(n18838), .B2(n18684), .ZN(
        n18679) );
  AOI22_X1 U21806 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18686), .B1(
        n18840), .B2(n18707), .ZN(n18678) );
  OAI211_X1 U21807 ( .C1(n18843), .C2(n18714), .A(n18679), .B(n18678), .ZN(
        P3_U2944) );
  AOI22_X1 U21808 ( .A1(n18844), .A2(n18684), .B1(n18846), .B2(n18707), .ZN(
        n18681) );
  AOI22_X1 U21809 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n18845), .ZN(n18680) );
  OAI211_X1 U21810 ( .C1(n18849), .C2(n18714), .A(n18681), .B(n18680), .ZN(
        P3_U2945) );
  AOI22_X1 U21811 ( .A1(n18685), .A2(n18852), .B1(n18850), .B2(n18684), .ZN(
        n18683) );
  AOI22_X1 U21812 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18686), .B1(
        n18851), .B2(n18707), .ZN(n18682) );
  OAI211_X1 U21813 ( .C1(n18855), .C2(n18714), .A(n18683), .B(n18682), .ZN(
        P3_U2946) );
  AOI22_X1 U21814 ( .A1(n18859), .A2(n18684), .B1(n18857), .B2(n18707), .ZN(
        n18688) );
  AOI22_X1 U21815 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18686), .B1(
        n18685), .B2(n18861), .ZN(n18687) );
  OAI211_X1 U21816 ( .C1(n18866), .C2(n18714), .A(n18688), .B(n18687), .ZN(
        P3_U2947) );
  NOR2_X2 U21817 ( .A1(n18689), .A2(n18712), .ZN(n18780) );
  INV_X1 U21818 ( .A(n18780), .ZN(n18711) );
  AOI21_X1 U21819 ( .B1(n18714), .B2(n18711), .A(n18933), .ZN(n18706) );
  AOI22_X1 U21820 ( .A1(n18811), .A2(n18730), .B1(n18810), .B2(n18706), .ZN(
        n18693) );
  NAND2_X1 U21821 ( .A1(n18714), .A2(n18711), .ZN(n18691) );
  OAI221_X1 U21822 ( .B1(n18691), .B2(n18787), .C1(n18691), .C2(n18690), .A(
        n18785), .ZN(n18708) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18708), .B1(
        n18816), .B2(n18707), .ZN(n18692) );
  OAI211_X1 U21824 ( .C1(n18819), .C2(n18711), .A(n18693), .B(n18692), .ZN(
        P3_U2948) );
  AOI22_X1 U21825 ( .A1(n18822), .A2(n18730), .B1(n18820), .B2(n18706), .ZN(
        n18695) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18708), .B1(
        n18821), .B2(n18707), .ZN(n18694) );
  OAI211_X1 U21827 ( .C1(n18825), .C2(n18711), .A(n18695), .B(n18694), .ZN(
        P3_U2949) );
  AOI22_X1 U21828 ( .A1(n18828), .A2(n18707), .B1(n18826), .B2(n18706), .ZN(
        n18697) );
  AOI22_X1 U21829 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18708), .B1(
        n18827), .B2(n18730), .ZN(n18696) );
  OAI211_X1 U21830 ( .C1(n18831), .C2(n18711), .A(n18697), .B(n18696), .ZN(
        P3_U2950) );
  AOI22_X1 U21831 ( .A1(n18834), .A2(n18707), .B1(n18833), .B2(n18706), .ZN(
        n18699) );
  AOI22_X1 U21832 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18708), .B1(
        n18832), .B2(n18730), .ZN(n18698) );
  OAI211_X1 U21833 ( .C1(n18837), .C2(n18711), .A(n18699), .B(n18698), .ZN(
        P3_U2951) );
  AOI22_X1 U21834 ( .A1(n18840), .A2(n18730), .B1(n18838), .B2(n18706), .ZN(
        n18701) );
  AOI22_X1 U21835 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18708), .B1(
        n18839), .B2(n18707), .ZN(n18700) );
  OAI211_X1 U21836 ( .C1(n18843), .C2(n18711), .A(n18701), .B(n18700), .ZN(
        P3_U2952) );
  AOI22_X1 U21837 ( .A1(n18845), .A2(n18707), .B1(n18844), .B2(n18706), .ZN(
        n18703) );
  AOI22_X1 U21838 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18708), .B1(
        n18846), .B2(n18730), .ZN(n18702) );
  OAI211_X1 U21839 ( .C1(n18849), .C2(n18711), .A(n18703), .B(n18702), .ZN(
        P3_U2953) );
  AOI22_X1 U21840 ( .A1(n18851), .A2(n18730), .B1(n18850), .B2(n18706), .ZN(
        n18705) );
  AOI22_X1 U21841 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18708), .B1(
        n18852), .B2(n18707), .ZN(n18704) );
  OAI211_X1 U21842 ( .C1(n18855), .C2(n18711), .A(n18705), .B(n18704), .ZN(
        P3_U2954) );
  AOI22_X1 U21843 ( .A1(n18859), .A2(n18706), .B1(n18857), .B2(n18730), .ZN(
        n18710) );
  AOI22_X1 U21844 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18708), .B1(
        n18861), .B2(n18707), .ZN(n18709) );
  OAI211_X1 U21845 ( .C1(n18866), .C2(n18711), .A(n18710), .B(n18709), .ZN(
        P3_U2955) );
  NOR2_X1 U21846 ( .A1(n18905), .A2(n18712), .ZN(n18764) );
  NAND2_X1 U21847 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18764), .ZN(
        n18760) );
  AND2_X1 U21848 ( .A1(n18809), .A2(n18764), .ZN(n18729) );
  AOI22_X1 U21849 ( .A1(n18810), .A2(n18729), .B1(n18816), .B2(n18730), .ZN(
        n18716) );
  AOI22_X1 U21850 ( .A1(n18815), .A2(n18713), .B1(n18812), .B2(n18764), .ZN(
        n18731) );
  INV_X1 U21851 ( .A(n18714), .ZN(n18756) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18731), .B1(
        n18811), .B2(n18756), .ZN(n18715) );
  OAI211_X1 U21853 ( .C1(n18819), .C2(n18760), .A(n18716), .B(n18715), .ZN(
        P3_U2956) );
  AOI22_X1 U21854 ( .A1(n18821), .A2(n18730), .B1(n18820), .B2(n18729), .ZN(
        n18718) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18731), .B1(
        n18822), .B2(n18756), .ZN(n18717) );
  OAI211_X1 U21856 ( .C1(n18825), .C2(n18760), .A(n18718), .B(n18717), .ZN(
        P3_U2957) );
  AOI22_X1 U21857 ( .A1(n18828), .A2(n18730), .B1(n18826), .B2(n18729), .ZN(
        n18720) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18731), .B1(
        n18827), .B2(n18756), .ZN(n18719) );
  OAI211_X1 U21859 ( .C1(n18831), .C2(n18760), .A(n18720), .B(n18719), .ZN(
        P3_U2958) );
  AOI22_X1 U21860 ( .A1(n18834), .A2(n18730), .B1(n18833), .B2(n18729), .ZN(
        n18722) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18731), .B1(
        n18832), .B2(n18756), .ZN(n18721) );
  OAI211_X1 U21862 ( .C1(n18837), .C2(n18760), .A(n18722), .B(n18721), .ZN(
        P3_U2959) );
  AOI22_X1 U21863 ( .A1(n18839), .A2(n18730), .B1(n18838), .B2(n18729), .ZN(
        n18724) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18731), .B1(
        n18840), .B2(n18756), .ZN(n18723) );
  OAI211_X1 U21865 ( .C1(n18843), .C2(n18760), .A(n18724), .B(n18723), .ZN(
        P3_U2960) );
  AOI22_X1 U21866 ( .A1(n18845), .A2(n18730), .B1(n18844), .B2(n18729), .ZN(
        n18726) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18731), .B1(
        n18846), .B2(n18756), .ZN(n18725) );
  OAI211_X1 U21868 ( .C1(n18849), .C2(n18760), .A(n18726), .B(n18725), .ZN(
        P3_U2961) );
  AOI22_X1 U21869 ( .A1(n18851), .A2(n18756), .B1(n18850), .B2(n18729), .ZN(
        n18728) );
  AOI22_X1 U21870 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18731), .B1(
        n18852), .B2(n18730), .ZN(n18727) );
  OAI211_X1 U21871 ( .C1(n18855), .C2(n18760), .A(n18728), .B(n18727), .ZN(
        P3_U2962) );
  AOI22_X1 U21872 ( .A1(n18861), .A2(n18730), .B1(n18859), .B2(n18729), .ZN(
        n18733) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18731), .B1(
        n18857), .B2(n18756), .ZN(n18732) );
  OAI211_X1 U21874 ( .C1(n18866), .C2(n18760), .A(n18733), .B(n18732), .ZN(
        P3_U2963) );
  INV_X1 U21875 ( .A(n18814), .ZN(n18761) );
  NOR2_X2 U21876 ( .A1(n18761), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18860) );
  INV_X1 U21877 ( .A(n18860), .ZN(n18759) );
  NAND2_X1 U21878 ( .A1(n18760), .A2(n18759), .ZN(n18786) );
  INV_X1 U21879 ( .A(n18786), .ZN(n18735) );
  NOR2_X1 U21880 ( .A1(n18933), .A2(n18735), .ZN(n18754) );
  AOI22_X1 U21881 ( .A1(n18810), .A2(n18754), .B1(n18816), .B2(n18756), .ZN(
        n18741) );
  NAND2_X1 U21882 ( .A1(n18787), .A2(n18734), .ZN(n18736) );
  OAI21_X1 U21883 ( .B1(n18737), .B2(n18736), .A(n18735), .ZN(n18738) );
  OAI211_X1 U21884 ( .C1(n18860), .C2(n19034), .A(n18739), .B(n18738), .ZN(
        n18755) );
  AOI22_X1 U21885 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18755), .B1(
        n18811), .B2(n18780), .ZN(n18740) );
  OAI211_X1 U21886 ( .C1(n18819), .C2(n18759), .A(n18741), .B(n18740), .ZN(
        P3_U2964) );
  AOI22_X1 U21887 ( .A1(n18821), .A2(n18756), .B1(n18820), .B2(n18754), .ZN(
        n18743) );
  AOI22_X1 U21888 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18755), .B1(
        n18822), .B2(n18780), .ZN(n18742) );
  OAI211_X1 U21889 ( .C1(n18825), .C2(n18759), .A(n18743), .B(n18742), .ZN(
        P3_U2965) );
  AOI22_X1 U21890 ( .A1(n18828), .A2(n18756), .B1(n18826), .B2(n18754), .ZN(
        n18745) );
  AOI22_X1 U21891 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18755), .B1(
        n18827), .B2(n18780), .ZN(n18744) );
  OAI211_X1 U21892 ( .C1(n18831), .C2(n18759), .A(n18745), .B(n18744), .ZN(
        P3_U2966) );
  AOI22_X1 U21893 ( .A1(n18834), .A2(n18756), .B1(n18833), .B2(n18754), .ZN(
        n18747) );
  AOI22_X1 U21894 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18755), .B1(
        n18832), .B2(n18780), .ZN(n18746) );
  OAI211_X1 U21895 ( .C1(n18837), .C2(n18759), .A(n18747), .B(n18746), .ZN(
        P3_U2967) );
  AOI22_X1 U21896 ( .A1(n18839), .A2(n18756), .B1(n18838), .B2(n18754), .ZN(
        n18749) );
  AOI22_X1 U21897 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18755), .B1(
        n18840), .B2(n18780), .ZN(n18748) );
  OAI211_X1 U21898 ( .C1(n18843), .C2(n18759), .A(n18749), .B(n18748), .ZN(
        P3_U2968) );
  AOI22_X1 U21899 ( .A1(n18845), .A2(n18756), .B1(n18844), .B2(n18754), .ZN(
        n18751) );
  AOI22_X1 U21900 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18755), .B1(
        n18846), .B2(n18780), .ZN(n18750) );
  OAI211_X1 U21901 ( .C1(n18849), .C2(n18759), .A(n18751), .B(n18750), .ZN(
        P3_U2969) );
  AOI22_X1 U21902 ( .A1(n18852), .A2(n18756), .B1(n18850), .B2(n18754), .ZN(
        n18753) );
  AOI22_X1 U21903 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18755), .B1(
        n18851), .B2(n18780), .ZN(n18752) );
  OAI211_X1 U21904 ( .C1(n18855), .C2(n18759), .A(n18753), .B(n18752), .ZN(
        P3_U2970) );
  AOI22_X1 U21905 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18755), .B1(
        n18859), .B2(n18754), .ZN(n18758) );
  AOI22_X1 U21906 ( .A1(n18861), .A2(n18756), .B1(n18857), .B2(n18780), .ZN(
        n18757) );
  OAI211_X1 U21907 ( .C1(n18866), .C2(n18759), .A(n18758), .B(n18757), .ZN(
        P3_U2971) );
  INV_X1 U21908 ( .A(n18760), .ZN(n18804) );
  NOR2_X1 U21909 ( .A1(n18933), .A2(n18761), .ZN(n18779) );
  AOI22_X1 U21910 ( .A1(n18811), .A2(n18804), .B1(n18810), .B2(n18779), .ZN(
        n18766) );
  AOI22_X1 U21911 ( .A1(n18815), .A2(n18764), .B1(n18763), .B2(n18762), .ZN(
        n18781) );
  AOI22_X1 U21912 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18781), .B1(
        n18816), .B2(n18780), .ZN(n18765) );
  OAI211_X1 U21913 ( .C1(n18819), .C2(n18784), .A(n18766), .B(n18765), .ZN(
        P3_U2972) );
  AOI22_X1 U21914 ( .A1(n18822), .A2(n18804), .B1(n18820), .B2(n18779), .ZN(
        n18768) );
  AOI22_X1 U21915 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18781), .B1(
        n18821), .B2(n18780), .ZN(n18767) );
  OAI211_X1 U21916 ( .C1(n18825), .C2(n18784), .A(n18768), .B(n18767), .ZN(
        P3_U2973) );
  AOI22_X1 U21917 ( .A1(n18828), .A2(n18780), .B1(n18826), .B2(n18779), .ZN(
        n18770) );
  AOI22_X1 U21918 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18781), .B1(
        n18827), .B2(n18804), .ZN(n18769) );
  OAI211_X1 U21919 ( .C1(n18831), .C2(n18784), .A(n18770), .B(n18769), .ZN(
        P3_U2974) );
  AOI22_X1 U21920 ( .A1(n18834), .A2(n18780), .B1(n18833), .B2(n18779), .ZN(
        n18772) );
  AOI22_X1 U21921 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18781), .B1(
        n18832), .B2(n18804), .ZN(n18771) );
  OAI211_X1 U21922 ( .C1(n18837), .C2(n18784), .A(n18772), .B(n18771), .ZN(
        P3_U2975) );
  AOI22_X1 U21923 ( .A1(n18840), .A2(n18804), .B1(n18838), .B2(n18779), .ZN(
        n18774) );
  AOI22_X1 U21924 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18781), .B1(
        n18839), .B2(n18780), .ZN(n18773) );
  OAI211_X1 U21925 ( .C1(n18843), .C2(n18784), .A(n18774), .B(n18773), .ZN(
        P3_U2976) );
  AOI22_X1 U21926 ( .A1(n18844), .A2(n18779), .B1(n18846), .B2(n18804), .ZN(
        n18776) );
  AOI22_X1 U21927 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18781), .B1(
        n18845), .B2(n18780), .ZN(n18775) );
  OAI211_X1 U21928 ( .C1(n18849), .C2(n18784), .A(n18776), .B(n18775), .ZN(
        P3_U2977) );
  AOI22_X1 U21929 ( .A1(n18851), .A2(n18804), .B1(n18850), .B2(n18779), .ZN(
        n18778) );
  AOI22_X1 U21930 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18781), .B1(
        n18852), .B2(n18780), .ZN(n18777) );
  OAI211_X1 U21931 ( .C1(n18855), .C2(n18784), .A(n18778), .B(n18777), .ZN(
        P3_U2978) );
  AOI22_X1 U21932 ( .A1(n18859), .A2(n18779), .B1(n18857), .B2(n18804), .ZN(
        n18783) );
  AOI22_X1 U21933 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18781), .B1(
        n18861), .B2(n18780), .ZN(n18782) );
  OAI211_X1 U21934 ( .C1(n18866), .C2(n18784), .A(n18783), .B(n18782), .ZN(
        P3_U2979) );
  AND2_X1 U21935 ( .A1(n18809), .A2(n18788), .ZN(n18803) );
  AOI22_X1 U21936 ( .A1(n18811), .A2(n18860), .B1(n18810), .B2(n18803), .ZN(
        n18790) );
  OAI221_X1 U21937 ( .B1(n18788), .B2(n18787), .C1(n18788), .C2(n18786), .A(
        n18785), .ZN(n18805) );
  AOI22_X1 U21938 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18805), .B1(
        n18816), .B2(n18804), .ZN(n18789) );
  OAI211_X1 U21939 ( .C1(n18819), .C2(n18808), .A(n18790), .B(n18789), .ZN(
        P3_U2980) );
  AOI22_X1 U21940 ( .A1(n18822), .A2(n18860), .B1(n18820), .B2(n18803), .ZN(
        n18792) );
  AOI22_X1 U21941 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18805), .B1(
        n18821), .B2(n18804), .ZN(n18791) );
  OAI211_X1 U21942 ( .C1(n18825), .C2(n18808), .A(n18792), .B(n18791), .ZN(
        P3_U2981) );
  AOI22_X1 U21943 ( .A1(n18827), .A2(n18860), .B1(n18826), .B2(n18803), .ZN(
        n18794) );
  AOI22_X1 U21944 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18805), .B1(
        n18828), .B2(n18804), .ZN(n18793) );
  OAI211_X1 U21945 ( .C1(n18831), .C2(n18808), .A(n18794), .B(n18793), .ZN(
        P3_U2982) );
  AOI22_X1 U21946 ( .A1(n18833), .A2(n18803), .B1(n18832), .B2(n18860), .ZN(
        n18796) );
  AOI22_X1 U21947 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18805), .B1(
        n18834), .B2(n18804), .ZN(n18795) );
  OAI211_X1 U21948 ( .C1(n18837), .C2(n18808), .A(n18796), .B(n18795), .ZN(
        P3_U2983) );
  AOI22_X1 U21949 ( .A1(n18839), .A2(n18804), .B1(n18838), .B2(n18803), .ZN(
        n18798) );
  AOI22_X1 U21950 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18805), .B1(
        n18840), .B2(n18860), .ZN(n18797) );
  OAI211_X1 U21951 ( .C1(n18843), .C2(n18808), .A(n18798), .B(n18797), .ZN(
        P3_U2984) );
  AOI22_X1 U21952 ( .A1(n18845), .A2(n18804), .B1(n18844), .B2(n18803), .ZN(
        n18800) );
  AOI22_X1 U21953 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18805), .B1(
        n18846), .B2(n18860), .ZN(n18799) );
  OAI211_X1 U21954 ( .C1(n18849), .C2(n18808), .A(n18800), .B(n18799), .ZN(
        P3_U2985) );
  AOI22_X1 U21955 ( .A1(n18851), .A2(n18860), .B1(n18850), .B2(n18803), .ZN(
        n18802) );
  AOI22_X1 U21956 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18805), .B1(
        n18852), .B2(n18804), .ZN(n18801) );
  OAI211_X1 U21957 ( .C1(n18855), .C2(n18808), .A(n18802), .B(n18801), .ZN(
        P3_U2986) );
  AOI22_X1 U21958 ( .A1(n18859), .A2(n18803), .B1(n18857), .B2(n18860), .ZN(
        n18807) );
  AOI22_X1 U21959 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18805), .B1(
        n18861), .B2(n18804), .ZN(n18806) );
  OAI211_X1 U21960 ( .C1(n18866), .C2(n18808), .A(n18807), .B(n18806), .ZN(
        P3_U2987) );
  AND2_X1 U21961 ( .A1(n18809), .A2(n18813), .ZN(n18858) );
  AOI22_X1 U21962 ( .A1(n18811), .A2(n18856), .B1(n18810), .B2(n18858), .ZN(
        n18818) );
  AOI22_X1 U21963 ( .A1(n18815), .A2(n18814), .B1(n18813), .B2(n18812), .ZN(
        n18862) );
  AOI22_X1 U21964 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18862), .B1(
        n18816), .B2(n18860), .ZN(n18817) );
  OAI211_X1 U21965 ( .C1(n18819), .C2(n18865), .A(n18818), .B(n18817), .ZN(
        P3_U2988) );
  AOI22_X1 U21966 ( .A1(n18821), .A2(n18860), .B1(n18820), .B2(n18858), .ZN(
        n18824) );
  AOI22_X1 U21967 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18862), .B1(
        n18822), .B2(n18856), .ZN(n18823) );
  OAI211_X1 U21968 ( .C1(n18825), .C2(n18865), .A(n18824), .B(n18823), .ZN(
        P3_U2989) );
  AOI22_X1 U21969 ( .A1(n18827), .A2(n18856), .B1(n18826), .B2(n18858), .ZN(
        n18830) );
  AOI22_X1 U21970 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18862), .B1(
        n18828), .B2(n18860), .ZN(n18829) );
  OAI211_X1 U21971 ( .C1(n18831), .C2(n18865), .A(n18830), .B(n18829), .ZN(
        P3_U2990) );
  AOI22_X1 U21972 ( .A1(n18833), .A2(n18858), .B1(n18832), .B2(n18856), .ZN(
        n18836) );
  AOI22_X1 U21973 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18862), .B1(
        n18834), .B2(n18860), .ZN(n18835) );
  OAI211_X1 U21974 ( .C1(n18837), .C2(n18865), .A(n18836), .B(n18835), .ZN(
        P3_U2991) );
  AOI22_X1 U21975 ( .A1(n18839), .A2(n18860), .B1(n18838), .B2(n18858), .ZN(
        n18842) );
  AOI22_X1 U21976 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18862), .B1(
        n18840), .B2(n18856), .ZN(n18841) );
  OAI211_X1 U21977 ( .C1(n18843), .C2(n18865), .A(n18842), .B(n18841), .ZN(
        P3_U2992) );
  AOI22_X1 U21978 ( .A1(n18845), .A2(n18860), .B1(n18844), .B2(n18858), .ZN(
        n18848) );
  AOI22_X1 U21979 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18862), .B1(
        n18846), .B2(n18856), .ZN(n18847) );
  OAI211_X1 U21980 ( .C1(n18849), .C2(n18865), .A(n18848), .B(n18847), .ZN(
        P3_U2993) );
  AOI22_X1 U21981 ( .A1(n18851), .A2(n18856), .B1(n18850), .B2(n18858), .ZN(
        n18854) );
  AOI22_X1 U21982 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18862), .B1(
        n18852), .B2(n18860), .ZN(n18853) );
  OAI211_X1 U21983 ( .C1(n18855), .C2(n18865), .A(n18854), .B(n18853), .ZN(
        P3_U2994) );
  AOI22_X1 U21984 ( .A1(n18859), .A2(n18858), .B1(n18857), .B2(n18856), .ZN(
        n18864) );
  AOI22_X1 U21985 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18862), .B1(
        n18861), .B2(n18860), .ZN(n18863) );
  OAI211_X1 U21986 ( .C1(n18866), .C2(n18865), .A(n18864), .B(n18863), .ZN(
        P3_U2995) );
  NOR2_X1 U21987 ( .A1(n18890), .A2(n18867), .ZN(n18869) );
  OAI222_X1 U21988 ( .A1(n18873), .A2(n18872), .B1(n18871), .B2(n18870), .C1(
        n18869), .C2(n18868), .ZN(n19077) );
  OAI21_X1 U21989 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18874), .ZN(n18875) );
  OAI211_X1 U21990 ( .C1(n18897), .C2(n18877), .A(n18876), .B(n18875), .ZN(
        n18919) );
  NOR2_X1 U21991 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18878), .ZN(
        n18901) );
  INV_X1 U21992 ( .A(n18901), .ZN(n18879) );
  AOI22_X1 U21993 ( .A1(n18887), .A2(n18879), .B1(n18890), .B2(n18880), .ZN(
        n19035) );
  NOR2_X1 U21994 ( .A1(n18908), .A2(n19035), .ZN(n18884) );
  OAI21_X1 U21995 ( .B1(n18887), .B2(n18900), .A(n18880), .ZN(n18881) );
  AOI21_X1 U21996 ( .B1(n18885), .B2(n18882), .A(n18881), .ZN(n19038) );
  NAND2_X1 U21997 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19038), .ZN(
        n18883) );
  OAI22_X1 U21998 ( .A1(n18884), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18908), .B2(n18883), .ZN(n18917) );
  AOI21_X1 U21999 ( .B1(n19057), .B2(n18891), .A(n18885), .ZN(n18896) );
  NAND2_X1 U22000 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18886), .ZN(
        n18895) );
  AOI21_X1 U22001 ( .B1(n19050), .B2(n19057), .A(n18887), .ZN(n18888) );
  AOI22_X1 U22002 ( .A1(n18890), .A2(n19045), .B1(n18889), .B2(n18888), .ZN(
        n18894) );
  NOR2_X1 U22003 ( .A1(n18898), .A2(n19064), .ZN(n18892) );
  OAI211_X1 U22004 ( .C1(n18892), .C2(n18891), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n19050), .ZN(n18893) );
  OAI211_X1 U22005 ( .C1(n18896), .C2(n18895), .A(n18894), .B(n18893), .ZN(
        n19048) );
  MUX2_X1 U22006 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n19048), .S(
        n18897), .Z(n18912) );
  AND2_X1 U22007 ( .A1(n18899), .A2(n18898), .ZN(n18902) );
  AOI22_X1 U22008 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18900), .B1(
        n18902), .B2(n19064), .ZN(n19059) );
  OAI22_X1 U22009 ( .A1(n18902), .A2(n19051), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18901), .ZN(n19055) );
  OR3_X1 U22010 ( .A1(n19059), .A2(n18905), .A3(n18903), .ZN(n18904) );
  AOI22_X1 U22011 ( .A1(n19059), .A2(n18905), .B1(n19055), .B2(n18904), .ZN(
        n18907) );
  OAI21_X1 U22012 ( .B1(n18908), .B2(n18907), .A(n18906), .ZN(n18911) );
  AND2_X1 U22013 ( .A1(n18912), .A2(n18911), .ZN(n18909) );
  OAI221_X1 U22014 ( .B1(n18912), .B2(n18911), .C1(n18910), .C2(n18909), .A(
        n18914), .ZN(n18916) );
  AOI21_X1 U22015 ( .B1(n18914), .B2(n18913), .A(n18912), .ZN(n18915) );
  AOI222_X1 U22016 ( .A1(n18917), .A2(n18916), .B1(n18917), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18916), .C2(n18915), .ZN(
        n18918) );
  NOR4_X1 U22017 ( .A1(n18920), .A2(n19077), .A3(n18919), .A4(n18918), .ZN(
        n18930) );
  NAND2_X1 U22018 ( .A1(n19042), .A2(n18931), .ZN(n18941) );
  INV_X1 U22019 ( .A(n18941), .ZN(n19087) );
  AOI22_X1 U22020 ( .A1(n18932), .A2(n19081), .B1(n19058), .B2(n19087), .ZN(
        n18921) );
  INV_X1 U22021 ( .A(n18921), .ZN(n18926) );
  OAI211_X1 U22022 ( .C1(n18923), .C2(n18922), .A(n19079), .B(n18930), .ZN(
        n19033) );
  OAI21_X1 U22023 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19085), .A(n19033), 
        .ZN(n18934) );
  NOR2_X1 U22024 ( .A1(n18924), .A2(n18934), .ZN(n18925) );
  MUX2_X1 U22025 ( .A(n18926), .B(n18925), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18928) );
  OAI211_X1 U22026 ( .C1(n18930), .C2(n18929), .A(n18928), .B(n18927), .ZN(
        P3_U2996) );
  NAND2_X1 U22027 ( .A1(n18932), .A2(n19081), .ZN(n18937) );
  NAND4_X1 U22028 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18932), .A4(n18931), .ZN(n18939) );
  OR3_X1 U22029 ( .A1(n18935), .A2(n18934), .A3(n18933), .ZN(n18936) );
  NAND4_X1 U22030 ( .A1(n18938), .A2(n18937), .A3(n18939), .A4(n18936), .ZN(
        P3_U2997) );
  AND4_X1 U22031 ( .A1(n18941), .A2(n18940), .A3(n18939), .A4(n19032), .ZN(
        P3_U2998) );
  AND2_X1 U22032 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18942), .ZN(
        P3_U2999) );
  INV_X1 U22033 ( .A(n19031), .ZN(n18943) );
  AND2_X1 U22034 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18943), .ZN(
        P3_U3000) );
  AND2_X1 U22035 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18942), .ZN(
        P3_U3001) );
  AND2_X1 U22036 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18943), .ZN(
        P3_U3002) );
  AND2_X1 U22037 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18942), .ZN(
        P3_U3003) );
  AND2_X1 U22038 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18942), .ZN(
        P3_U3004) );
  AND2_X1 U22039 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18943), .ZN(
        P3_U3005) );
  AND2_X1 U22040 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18942), .ZN(
        P3_U3006) );
  AND2_X1 U22041 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18942), .ZN(
        P3_U3007) );
  AND2_X1 U22042 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18942), .ZN(
        P3_U3008) );
  AND2_X1 U22043 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18942), .ZN(
        P3_U3009) );
  AND2_X1 U22044 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18943), .ZN(
        P3_U3010) );
  AND2_X1 U22045 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18943), .ZN(
        P3_U3011) );
  AND2_X1 U22046 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18943), .ZN(
        P3_U3012) );
  AND2_X1 U22047 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18943), .ZN(
        P3_U3013) );
  AND2_X1 U22048 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18943), .ZN(
        P3_U3014) );
  AND2_X1 U22049 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18943), .ZN(
        P3_U3015) );
  AND2_X1 U22050 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18942), .ZN(
        P3_U3016) );
  AND2_X1 U22051 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18942), .ZN(
        P3_U3017) );
  AND2_X1 U22052 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18942), .ZN(
        P3_U3018) );
  AND2_X1 U22053 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18942), .ZN(
        P3_U3019) );
  AND2_X1 U22054 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18942), .ZN(
        P3_U3020) );
  AND2_X1 U22055 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18943), .ZN(P3_U3021) );
  AND2_X1 U22056 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18943), .ZN(P3_U3022) );
  AND2_X1 U22057 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18943), .ZN(P3_U3023) );
  AND2_X1 U22058 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18943), .ZN(P3_U3024) );
  AND2_X1 U22059 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18943), .ZN(P3_U3025) );
  AND2_X1 U22060 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18943), .ZN(P3_U3026) );
  AND2_X1 U22061 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18943), .ZN(P3_U3027) );
  AND2_X1 U22062 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18943), .ZN(P3_U3028) );
  NOR2_X1 U22063 ( .A1(n19085), .A2(n18944), .ZN(n18951) );
  INV_X1 U22064 ( .A(n18951), .ZN(n18953) );
  OAI21_X1 U22065 ( .B1(n18945), .B2(n20819), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18947) );
  INV_X1 U22066 ( .A(NA), .ZN(n21056) );
  NOR3_X1 U22067 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .A3(n21056), .ZN(n18946) );
  AOI21_X1 U22068 ( .B1(n19093), .B2(n18947), .A(n18946), .ZN(n18948) );
  OAI221_X1 U22069 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(P3_STATE_REG_0__SCAN_IN), .C1(P3_STATE_REG_2__SCAN_IN), .C2(n18953), .A(n18948), .ZN(P3_U3029) );
  NAND2_X1 U22070 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n18952) );
  AOI22_X1 U22071 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18952), .B1(HOLD), 
        .B2(n18949), .ZN(n18950) );
  OAI211_X1 U22072 ( .C1(n18950), .C2(n18957), .A(n18953), .B(n19082), .ZN(
        P3_U3030) );
  AOI221_X1 U22073 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18957), .C1(n21056), 
        .C2(n18957), .A(n18951), .ZN(n18958) );
  INV_X1 U22074 ( .A(n18952), .ZN(n18955) );
  OAI22_X1 U22075 ( .A1(NA), .A2(n18953), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18954) );
  OAI22_X1 U22076 ( .A1(n18955), .A2(n18954), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18956) );
  OAI22_X1 U22077 ( .A1(n18958), .A2(n18959), .B1(n18957), .B2(n18956), .ZN(
        P3_U3031) );
  INV_X1 U22078 ( .A(n19093), .ZN(n19092) );
  OAI222_X1 U22079 ( .A1(n19066), .A2(n9805), .B1(n18960), .B2(n19092), .C1(
        n18961), .C2(n19022), .ZN(P3_U3032) );
  OAI222_X1 U22080 ( .A1(n19022), .A2(n18964), .B1(n18962), .B2(n19019), .C1(
        n18961), .C2(n9805), .ZN(P3_U3033) );
  OAI222_X1 U22081 ( .A1(n19022), .A2(n18966), .B1(n18965), .B2(n19092), .C1(
        n18964), .C2(n9805), .ZN(P3_U3034) );
  OAI222_X1 U22082 ( .A1(n19022), .A2(n18968), .B1(n18967), .B2(n19019), .C1(
        n18966), .C2(n9805), .ZN(P3_U3035) );
  OAI222_X1 U22083 ( .A1(n19022), .A2(n18970), .B1(n18969), .B2(n19092), .C1(
        n18968), .C2(n9805), .ZN(P3_U3036) );
  OAI222_X1 U22084 ( .A1(n19022), .A2(n18972), .B1(n18971), .B2(n19092), .C1(
        n18970), .C2(n9805), .ZN(P3_U3037) );
  OAI222_X1 U22085 ( .A1(n19022), .A2(n18975), .B1(n18973), .B2(n19026), .C1(
        n18972), .C2(n9805), .ZN(P3_U3038) );
  OAI222_X1 U22086 ( .A1(n18975), .A2(n9805), .B1(n18974), .B2(n19092), .C1(
        n18976), .C2(n19022), .ZN(P3_U3039) );
  INV_X1 U22087 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18978) );
  OAI222_X1 U22088 ( .A1(n19022), .A2(n18978), .B1(n18977), .B2(n19092), .C1(
        n18976), .C2(n9805), .ZN(P3_U3040) );
  OAI222_X1 U22089 ( .A1(n19022), .A2(n18980), .B1(n18979), .B2(n19092), .C1(
        n18978), .C2(n9805), .ZN(P3_U3041) );
  OAI222_X1 U22090 ( .A1(n19022), .A2(n18982), .B1(n18981), .B2(n19092), .C1(
        n18980), .C2(n9805), .ZN(P3_U3042) );
  OAI222_X1 U22091 ( .A1(n19022), .A2(n18984), .B1(n18983), .B2(n19092), .C1(
        n18982), .C2(n9805), .ZN(P3_U3043) );
  OAI222_X1 U22092 ( .A1(n19022), .A2(n18987), .B1(n18985), .B2(n19092), .C1(
        n18984), .C2(n9805), .ZN(P3_U3044) );
  OAI222_X1 U22093 ( .A1(n18987), .A2(n9805), .B1(n18986), .B2(n19092), .C1(
        n18988), .C2(n19022), .ZN(P3_U3045) );
  OAI222_X1 U22094 ( .A1(n19022), .A2(n18990), .B1(n18989), .B2(n19092), .C1(
        n18988), .C2(n9805), .ZN(P3_U3046) );
  OAI222_X1 U22095 ( .A1(n19022), .A2(n18992), .B1(n18991), .B2(n19092), .C1(
        n18990), .C2(n9805), .ZN(P3_U3047) );
  OAI222_X1 U22096 ( .A1(n19022), .A2(n18994), .B1(n18993), .B2(n19092), .C1(
        n18992), .C2(n9805), .ZN(P3_U3048) );
  OAI222_X1 U22097 ( .A1(n19022), .A2(n18996), .B1(n18995), .B2(n19092), .C1(
        n18994), .C2(n9805), .ZN(P3_U3049) );
  INV_X1 U22098 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18999) );
  OAI222_X1 U22099 ( .A1(n19022), .A2(n18999), .B1(n18997), .B2(n19092), .C1(
        n18996), .C2(n9805), .ZN(P3_U3050) );
  OAI222_X1 U22100 ( .A1(n18999), .A2(n9805), .B1(n18998), .B2(n19092), .C1(
        n19000), .C2(n19022), .ZN(P3_U3051) );
  INV_X1 U22101 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19002) );
  OAI222_X1 U22102 ( .A1(n19022), .A2(n19002), .B1(n19001), .B2(n19092), .C1(
        n19000), .C2(n9805), .ZN(P3_U3052) );
  OAI222_X1 U22103 ( .A1(n19022), .A2(n19004), .B1(n19003), .B2(n19092), .C1(
        n19002), .C2(n9805), .ZN(P3_U3053) );
  OAI222_X1 U22104 ( .A1(n19022), .A2(n19006), .B1(n19005), .B2(n19019), .C1(
        n19004), .C2(n9805), .ZN(P3_U3054) );
  OAI222_X1 U22105 ( .A1(n19022), .A2(n19008), .B1(n19007), .B2(n19019), .C1(
        n19006), .C2(n9805), .ZN(P3_U3055) );
  OAI222_X1 U22106 ( .A1(n19022), .A2(n19010), .B1(n19009), .B2(n19019), .C1(
        n19008), .C2(n9805), .ZN(P3_U3056) );
  OAI222_X1 U22107 ( .A1(n19022), .A2(n19013), .B1(n19011), .B2(n19019), .C1(
        n19010), .C2(n9805), .ZN(P3_U3057) );
  OAI222_X1 U22108 ( .A1(n9805), .A2(n19013), .B1(n19012), .B2(n19019), .C1(
        n19014), .C2(n19022), .ZN(P3_U3058) );
  OAI222_X1 U22109 ( .A1(n19022), .A2(n19016), .B1(n19015), .B2(n19019), .C1(
        n19014), .C2(n9805), .ZN(P3_U3059) );
  OAI222_X1 U22110 ( .A1(n19022), .A2(n19018), .B1(n19017), .B2(n19019), .C1(
        n19016), .C2(n9805), .ZN(P3_U3060) );
  INV_X1 U22111 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19020) );
  OAI222_X1 U22112 ( .A1(n19022), .A2(n19021), .B1(n19020), .B2(n19019), .C1(
        n19018), .C2(n9805), .ZN(P3_U3061) );
  OAI22_X1 U22113 ( .A1(n19093), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19092), .ZN(n19023) );
  INV_X1 U22114 ( .A(n19023), .ZN(P3_U3274) );
  OAI22_X1 U22115 ( .A1(n19093), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19092), .ZN(n19024) );
  INV_X1 U22116 ( .A(n19024), .ZN(P3_U3275) );
  OAI22_X1 U22117 ( .A1(n19093), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19092), .ZN(n19025) );
  INV_X1 U22118 ( .A(n19025), .ZN(P3_U3276) );
  OAI22_X1 U22119 ( .A1(n19093), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19026), .ZN(n19027) );
  INV_X1 U22120 ( .A(n19027), .ZN(P3_U3277) );
  OAI21_X1 U22121 ( .B1(n19031), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19029), 
        .ZN(n19028) );
  INV_X1 U22122 ( .A(n19028), .ZN(P3_U3280) );
  OAI21_X1 U22123 ( .B1(n19031), .B2(n19030), .A(n19029), .ZN(P3_U3281) );
  OAI221_X1 U22124 ( .B1(n19034), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19034), 
        .C2(n19033), .A(n19032), .ZN(P3_U3282) );
  NOR3_X1 U22125 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19035), .A3(
        n19095), .ZN(n19036) );
  AOI21_X1 U22126 ( .B1(n19037), .B2(n19058), .A(n19036), .ZN(n19041) );
  OAI21_X1 U22127 ( .B1(n19095), .B2(n19038), .A(n19062), .ZN(n19039) );
  INV_X1 U22128 ( .A(n19039), .ZN(n19040) );
  OAI22_X1 U22129 ( .A1(n19065), .A2(n19041), .B1(n19040), .B2(n17094), .ZN(
        P3_U3285) );
  NOR2_X1 U22130 ( .A1(n19042), .A2(n19061), .ZN(n19052) );
  OAI22_X1 U22131 ( .A1(n19044), .A2(n19043), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19053) );
  INV_X1 U22132 ( .A(n19053), .ZN(n19047) );
  INV_X1 U22133 ( .A(n19045), .ZN(n19046) );
  AOI222_X1 U22134 ( .A1(n19048), .A2(n19060), .B1(n19052), .B2(n19047), .C1(
        n19058), .C2(n19046), .ZN(n19049) );
  AOI22_X1 U22135 ( .A1(n19065), .A2(n19050), .B1(n19049), .B2(n19062), .ZN(
        P3_U3288) );
  INV_X1 U22136 ( .A(n19051), .ZN(n19054) );
  AOI222_X1 U22137 ( .A1(n19055), .A2(n19060), .B1(n19058), .B2(n19054), .C1(
        n19053), .C2(n19052), .ZN(n19056) );
  AOI22_X1 U22138 ( .A1(n19065), .A2(n19057), .B1(n19056), .B2(n19062), .ZN(
        P3_U3289) );
  AOI222_X1 U22139 ( .A1(n19061), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19060), 
        .B2(n19059), .C1(n19064), .C2(n19058), .ZN(n19063) );
  AOI22_X1 U22140 ( .A1(n19065), .A2(n19064), .B1(n19063), .B2(n19062), .ZN(
        P3_U3290) );
  AOI21_X1 U22141 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19067) );
  AOI22_X1 U22142 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19067), .B2(n19066), .ZN(n19069) );
  INV_X1 U22143 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19068) );
  AOI22_X1 U22144 ( .A1(n19070), .A2(n19069), .B1(n19068), .B2(n19073), .ZN(
        P3_U3292) );
  INV_X1 U22145 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19074) );
  NOR2_X1 U22146 ( .A1(n19073), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19071) );
  AOI22_X1 U22147 ( .A1(n19074), .A2(n19073), .B1(n19072), .B2(n19071), .ZN(
        P3_U3293) );
  INV_X1 U22148 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19075) );
  AOI22_X1 U22149 ( .A1(n19092), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19075), 
        .B2(n19093), .ZN(P3_U3294) );
  MUX2_X1 U22150 ( .A(P3_MORE_REG_SCAN_IN), .B(n19077), .S(n19076), .Z(
        P3_U3295) );
  OAI21_X1 U22151 ( .B1(n19079), .B2(n19078), .A(n19097), .ZN(n19080) );
  AOI21_X1 U22152 ( .B1(n19081), .B2(n19085), .A(n19080), .ZN(n19091) );
  AOI21_X1 U22153 ( .B1(n19084), .B2(n19083), .A(n19082), .ZN(n19086) );
  OAI211_X1 U22154 ( .C1(n19096), .C2(n19086), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19085), .ZN(n19088) );
  AOI21_X1 U22155 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19088), .A(n19087), 
        .ZN(n19090) );
  NAND2_X1 U22156 ( .A1(n19091), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19089) );
  OAI21_X1 U22157 ( .B1(n19091), .B2(n19090), .A(n19089), .ZN(P3_U3296) );
  OAI22_X1 U22158 ( .A1(n19093), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19092), .ZN(n19094) );
  INV_X1 U22159 ( .A(n19094), .ZN(P3_U3297) );
  OAI21_X1 U22160 ( .B1(n19095), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n19097), 
        .ZN(n19100) );
  OAI22_X1 U22161 ( .A1(n19100), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19097), 
        .B2(n19096), .ZN(n19098) );
  INV_X1 U22162 ( .A(n19098), .ZN(P3_U3298) );
  OAI21_X1 U22163 ( .B1(n19100), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n19099), 
        .ZN(n19101) );
  INV_X1 U22164 ( .A(n19101), .ZN(P3_U3299) );
  INV_X1 U22165 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19957) );
  NAND2_X1 U22166 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19957), .ZN(n19945) );
  INV_X1 U22167 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19938) );
  AOI22_X1 U22168 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19945), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19938), .ZN(n20028) );
  AOI21_X1 U22169 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20028), .ZN(n19102) );
  INV_X1 U22170 ( .A(n19102), .ZN(P2_U2815) );
  AOI22_X1 U22171 ( .A1(n19104), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n20035), 
        .B2(n19103), .ZN(n19105) );
  INV_X1 U22172 ( .A(n19105), .ZN(P2_U2816) );
  NAND2_X1 U22173 ( .A1(n19938), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20086) );
  INV_X2 U22174 ( .A(n20086), .ZN(n20015) );
  OR2_X1 U22175 ( .A1(n19948), .A2(n20015), .ZN(n19941) );
  AOI21_X1 U22176 ( .B1(n19938), .B2(n19941), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19106) );
  AOI21_X1 U22177 ( .B1(n20015), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n19106), 
        .ZN(P2_U2817) );
  OAI21_X1 U22178 ( .B1(n19948), .B2(BS16), .A(n20028), .ZN(n20026) );
  OAI21_X1 U22179 ( .B1(n20028), .B2(n12350), .A(n20026), .ZN(P2_U2818) );
  NOR4_X1 U22180 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19110) );
  NOR4_X1 U22181 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19109) );
  NOR4_X1 U22182 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19108) );
  NOR4_X1 U22183 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19107) );
  NAND4_X1 U22184 ( .A1(n19110), .A2(n19109), .A3(n19108), .A4(n19107), .ZN(
        n19116) );
  NOR4_X1 U22185 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19114) );
  AOI211_X1 U22186 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19113) );
  NOR4_X1 U22187 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19112) );
  NOR4_X1 U22188 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19111) );
  NAND4_X1 U22189 ( .A1(n19114), .A2(n19113), .A3(n19112), .A4(n19111), .ZN(
        n19115) );
  NOR2_X1 U22190 ( .A1(n19116), .A2(n19115), .ZN(n19127) );
  INV_X1 U22191 ( .A(n19127), .ZN(n19125) );
  NOR2_X1 U22192 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19125), .ZN(n19119) );
  INV_X1 U22193 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19117) );
  AOI22_X1 U22194 ( .A1(n19119), .A2(n19120), .B1(n19125), .B2(n19117), .ZN(
        P2_U2820) );
  OR3_X1 U22195 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19124) );
  INV_X1 U22196 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19118) );
  AOI22_X1 U22197 ( .A1(n19119), .A2(n19124), .B1(n19125), .B2(n19118), .ZN(
        P2_U2821) );
  INV_X1 U22198 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20027) );
  NAND2_X1 U22199 ( .A1(n19119), .A2(n20027), .ZN(n19123) );
  INV_X1 U22200 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19958) );
  OAI21_X1 U22201 ( .B1(n19120), .B2(n19958), .A(n19127), .ZN(n19121) );
  OAI21_X1 U22202 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19127), .A(n19121), 
        .ZN(n19122) );
  OAI221_X1 U22203 ( .B1(n19123), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19123), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19122), .ZN(P2_U2822) );
  INV_X1 U22204 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19126) );
  OAI221_X1 U22205 ( .B1(n19127), .B2(n19126), .C1(n19125), .C2(n19124), .A(
        n19123), .ZN(P2_U2823) );
  OAI21_X1 U22206 ( .B1(n19133), .B2(n19129), .A(n19128), .ZN(n19130) );
  INV_X1 U22207 ( .A(n19130), .ZN(n19131) );
  AOI21_X1 U22208 ( .B1(n19288), .B2(n19132), .A(n19131), .ZN(n19138) );
  INV_X1 U22209 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19996) );
  OAI22_X1 U22210 ( .A1(n19271), .A2(n9973), .B1(n19996), .B2(n19256), .ZN(
        n19135) );
  OAI22_X1 U22211 ( .A1(n15552), .A2(n19264), .B1(n19133), .B2(n19175), .ZN(
        n19134) );
  AOI211_X1 U22212 ( .C1(n19243), .C2(n19136), .A(n19135), .B(n19134), .ZN(
        n19137) );
  OAI211_X1 U22213 ( .C1(n19139), .C2(n19290), .A(n19138), .B(n19137), .ZN(
        P2_U2835) );
  NAND2_X1 U22214 ( .A1(n9797), .A2(n19140), .ZN(n19141) );
  XOR2_X1 U22215 ( .A(n19142), .B(n19141), .Z(n19151) );
  AOI22_X1 U22216 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19298), .B1(
        P2_EBX_REG_19__SCAN_IN), .B2(n19293), .ZN(n19143) );
  OAI21_X1 U22217 ( .B1(n19144), .B2(n19266), .A(n19143), .ZN(n19145) );
  AOI211_X1 U22218 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n19286), .A(n19404), 
        .B(n19145), .ZN(n19150) );
  INV_X1 U22219 ( .A(n19146), .ZN(n19147) );
  AOI22_X1 U22220 ( .A1(n19148), .A2(n19243), .B1(n19147), .B2(n19203), .ZN(
        n19149) );
  OAI211_X1 U22221 ( .C1(n19301), .C2(n19151), .A(n19150), .B(n19149), .ZN(
        P2_U2836) );
  OAI21_X1 U22222 ( .B1(n19992), .B2(n19256), .A(n19254), .ZN(n19154) );
  OAI22_X1 U22223 ( .A1(n19152), .A2(n19266), .B1(n11207), .B2(n19271), .ZN(
        n19153) );
  AOI211_X1 U22224 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19298), .A(
        n19154), .B(n19153), .ZN(n19160) );
  NOR2_X1 U22225 ( .A1(n19277), .A2(n19163), .ZN(n19156) );
  XNOR2_X1 U22226 ( .A(n19156), .B(n19155), .ZN(n19158) );
  AOI22_X1 U22227 ( .A1(n19158), .A2(n19245), .B1(n19157), .B2(n19243), .ZN(
        n19159) );
  OAI211_X1 U22228 ( .C1(n19161), .C2(n19290), .A(n19160), .B(n19159), .ZN(
        P2_U2837) );
  AOI211_X1 U22229 ( .C1(n19165), .C2(n19164), .A(n19163), .B(n19162), .ZN(
        n19169) );
  AOI22_X1 U22230 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19298), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19286), .ZN(n19166) );
  OAI211_X1 U22231 ( .C1(n19167), .C2(n19266), .A(n19166), .B(n19254), .ZN(
        n19168) );
  AOI211_X1 U22232 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19293), .A(n19169), .B(
        n19168), .ZN(n19174) );
  INV_X1 U22233 ( .A(n19170), .ZN(n19171) );
  AOI22_X1 U22234 ( .A1(n19172), .A2(n19243), .B1(n19171), .B2(n19203), .ZN(
        n19173) );
  OAI211_X1 U22235 ( .C1(n19176), .C2(n19175), .A(n19174), .B(n19173), .ZN(
        P2_U2838) );
  OAI21_X1 U22236 ( .B1(n19988), .B2(n19256), .A(n19254), .ZN(n19179) );
  OAI22_X1 U22237 ( .A1(n19177), .A2(n19266), .B1(n10935), .B2(n19271), .ZN(
        n19178) );
  AOI211_X1 U22238 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19298), .A(
        n19179), .B(n19178), .ZN(n19185) );
  XOR2_X1 U22239 ( .A(n19181), .B(n19180), .Z(n19183) );
  AOI22_X1 U22240 ( .A1(n19183), .A2(n19245), .B1(n19182), .B2(n19243), .ZN(
        n19184) );
  OAI211_X1 U22241 ( .C1(n19186), .C2(n19290), .A(n19185), .B(n19184), .ZN(
        P2_U2839) );
  INV_X1 U22242 ( .A(n19187), .ZN(n19189) );
  AOI22_X1 U22243 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19298), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19293), .ZN(n19188) );
  OAI21_X1 U22244 ( .B1(n19189), .B2(n19266), .A(n19188), .ZN(n19190) );
  AOI211_X1 U22245 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19286), .A(n19404), 
        .B(n19190), .ZN(n19196) );
  OR2_X1 U22246 ( .A1(n19277), .A2(n19191), .ZN(n19205) );
  XOR2_X1 U22247 ( .A(n19205), .B(n19192), .Z(n19194) );
  AOI22_X1 U22248 ( .A1(n19194), .A2(n19245), .B1(n19193), .B2(n19243), .ZN(
        n19195) );
  OAI211_X1 U22249 ( .C1(n19313), .C2(n19290), .A(n19196), .B(n19195), .ZN(
        P2_U2841) );
  OAI22_X1 U22250 ( .A1(n19197), .A2(n19264), .B1(n19982), .B2(n19256), .ZN(
        n19198) );
  AOI211_X1 U22251 ( .C1(n19206), .C2(n19199), .A(n19404), .B(n19198), .ZN(
        n19212) );
  AOI22_X1 U22252 ( .A1(n19200), .A2(n19288), .B1(P2_EBX_REG_13__SCAN_IN), 
        .B2(n19293), .ZN(n19211) );
  INV_X1 U22253 ( .A(n19201), .ZN(n19204) );
  AOI22_X1 U22254 ( .A1(n19204), .A2(n19203), .B1(n19243), .B2(n19202), .ZN(
        n19210) );
  AOI211_X1 U22255 ( .C1(n19207), .C2(n19206), .A(n19301), .B(n19205), .ZN(
        n19208) );
  INV_X1 U22256 ( .A(n19208), .ZN(n19209) );
  NAND4_X1 U22257 ( .A1(n19212), .A2(n19211), .A3(n19210), .A4(n19209), .ZN(
        P2_U2842) );
  OAI22_X1 U22258 ( .A1(n19213), .A2(n19266), .B1(n19271), .B2(n13393), .ZN(
        n19214) );
  INV_X1 U22259 ( .A(n19214), .ZN(n19215) );
  OAI211_X1 U22260 ( .C1(n19980), .C2(n19256), .A(n19215), .B(n19254), .ZN(
        n19216) );
  AOI21_X1 U22261 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19298), .A(
        n19216), .ZN(n19223) );
  NOR2_X1 U22262 ( .A1(n19277), .A2(n19217), .ZN(n19219) );
  XNOR2_X1 U22263 ( .A(n19219), .B(n19218), .ZN(n19221) );
  AOI22_X1 U22264 ( .A1(n19221), .A2(n19245), .B1(n19220), .B2(n19243), .ZN(
        n19222) );
  OAI211_X1 U22265 ( .C1(n19224), .C2(n19290), .A(n19223), .B(n19222), .ZN(
        P2_U2843) );
  INV_X1 U22266 ( .A(n19225), .ZN(n19226) );
  AOI22_X1 U22267 ( .A1(n19226), .A2(n19288), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19293), .ZN(n19227) );
  OAI211_X1 U22268 ( .C1(n19976), .C2(n19256), .A(n19227), .B(n19254), .ZN(
        n19228) );
  AOI21_X1 U22269 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19298), .A(
        n19228), .ZN(n19234) );
  NOR2_X1 U22270 ( .A1(n19277), .A2(n19229), .ZN(n19231) );
  XNOR2_X1 U22271 ( .A(n19231), .B(n19230), .ZN(n19232) );
  AOI22_X1 U22272 ( .A1(n19232), .A2(n19245), .B1(n9912), .B2(n19243), .ZN(
        n19233) );
  OAI211_X1 U22273 ( .C1(n19235), .C2(n19290), .A(n19234), .B(n19233), .ZN(
        P2_U2845) );
  AOI22_X1 U22274 ( .A1(n19236), .A2(n19288), .B1(n19293), .B2(
        P2_EBX_REG_8__SCAN_IN), .ZN(n19237) );
  OAI211_X1 U22275 ( .C1(n19972), .C2(n19256), .A(n19237), .B(n19254), .ZN(
        n19238) );
  AOI21_X1 U22276 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19298), .A(
        n19238), .ZN(n19248) );
  NOR2_X1 U22277 ( .A1(n19277), .A2(n19239), .ZN(n19241) );
  XNOR2_X1 U22278 ( .A(n19241), .B(n19240), .ZN(n19246) );
  INV_X1 U22279 ( .A(n19242), .ZN(n19244) );
  AOI22_X1 U22280 ( .A1(n19246), .A2(n19245), .B1(n19244), .B2(n19243), .ZN(
        n19247) );
  OAI211_X1 U22281 ( .C1(n19290), .C2(n19249), .A(n19248), .B(n19247), .ZN(
        P2_U2847) );
  NAND2_X1 U22282 ( .A1(n9797), .A2(n19250), .ZN(n19252) );
  XOR2_X1 U22283 ( .A(n19252), .B(n19251), .Z(n19262) );
  AOI22_X1 U22284 ( .A1(n19288), .A2(n19253), .B1(n19293), .B2(
        P2_EBX_REG_7__SCAN_IN), .ZN(n19255) );
  OAI211_X1 U22285 ( .C1(n19970), .C2(n19256), .A(n19255), .B(n19254), .ZN(
        n19260) );
  OAI22_X1 U22286 ( .A1(n19258), .A2(n19290), .B1(n19257), .B2(n19295), .ZN(
        n19259) );
  AOI211_X1 U22287 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19298), .A(
        n19260), .B(n19259), .ZN(n19261) );
  OAI21_X1 U22288 ( .B1(n19262), .B2(n19301), .A(n19261), .ZN(P2_U2848) );
  OAI22_X1 U22289 ( .A1(n19266), .A2(n19265), .B1(n19264), .B2(n19263), .ZN(
        n19267) );
  INV_X1 U22290 ( .A(n19267), .ZN(n19284) );
  XNOR2_X1 U22291 ( .A(n19269), .B(n19268), .ZN(n19403) );
  OAI22_X1 U22292 ( .A1(n19271), .A2(n19270), .B1(n19290), .B2(n19403), .ZN(
        n19272) );
  AOI211_X1 U22293 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19286), .A(n19404), .B(
        n19272), .ZN(n19283) );
  OAI22_X1 U22294 ( .A1(n19336), .A2(n19273), .B1(n19412), .B2(n19295), .ZN(
        n19274) );
  INV_X1 U22295 ( .A(n19274), .ZN(n19282) );
  INV_X1 U22296 ( .A(n19275), .ZN(n19280) );
  NOR2_X1 U22297 ( .A1(n19277), .A2(n19276), .ZN(n19279) );
  AOI21_X1 U22298 ( .B1(n19280), .B2(n19279), .A(n19301), .ZN(n19278) );
  OAI21_X1 U22299 ( .B1(n19280), .B2(n19279), .A(n19278), .ZN(n19281) );
  NAND4_X1 U22300 ( .A1(n19284), .A2(n19283), .A3(n19282), .A4(n19281), .ZN(
        P2_U2851) );
  INV_X1 U22301 ( .A(n19363), .ZN(n19291) );
  AOI22_X1 U22302 ( .A1(n19288), .A2(n19287), .B1(n19286), .B2(
        P2_REIP_REG_0__SCAN_IN), .ZN(n19289) );
  OAI21_X1 U22303 ( .B1(n19291), .B2(n19290), .A(n19289), .ZN(n19292) );
  AOI21_X1 U22304 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19293), .A(n19292), .ZN(
        n19294) );
  OAI21_X1 U22305 ( .B1(n10384), .B2(n19295), .A(n19294), .ZN(n19296) );
  AOI21_X1 U22306 ( .B1(n19364), .B2(n19297), .A(n19296), .ZN(n19300) );
  NAND2_X1 U22307 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19298), .ZN(
        n19299) );
  OAI211_X1 U22308 ( .C1(n14495), .C2(n19301), .A(n19300), .B(n19299), .ZN(
        P2_U2855) );
  AOI22_X1 U22309 ( .A1(n19303), .A2(n19360), .B1(n19302), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19306) );
  AOI22_X1 U22310 ( .A1(n19304), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19359), .ZN(n19305) );
  NAND2_X1 U22311 ( .A1(n19306), .A2(n19305), .ZN(P2_U2888) );
  AOI22_X1 U22312 ( .A1(n19324), .A2(n19307), .B1(P2_EAX_REG_15__SCAN_IN), 
        .B2(n19359), .ZN(n19308) );
  OAI21_X1 U22313 ( .B1(n19367), .B2(n19309), .A(n19308), .ZN(P2_U2904) );
  INV_X1 U22314 ( .A(n19367), .ZN(n19311) );
  AOI22_X1 U22315 ( .A1(n19311), .A2(n19310), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19359), .ZN(n19312) );
  OAI21_X1 U22316 ( .B1(n19318), .B2(n19313), .A(n19312), .ZN(P2_U2905) );
  AOI22_X1 U22317 ( .A1(n19324), .A2(n19314), .B1(P2_EAX_REG_11__SCAN_IN), 
        .B2(n19359), .ZN(n19315) );
  OAI21_X1 U22318 ( .B1(n19316), .B2(n19367), .A(n19315), .ZN(P2_U2908) );
  INV_X1 U22319 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19317) );
  OAI22_X1 U22320 ( .A1(n19319), .A2(n19318), .B1(n19333), .B2(n19317), .ZN(
        n19320) );
  INV_X1 U22321 ( .A(n19320), .ZN(n19321) );
  OAI21_X1 U22322 ( .B1(n19322), .B2(n19367), .A(n19321), .ZN(P2_U2913) );
  INV_X1 U22323 ( .A(n19323), .ZN(n19325) );
  AOI22_X1 U22324 ( .A1(n19325), .A2(n19324), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19359), .ZN(n19330) );
  XOR2_X1 U22325 ( .A(n20050), .B(n20051), .Z(n19349) );
  XNOR2_X1 U22326 ( .A(n20038), .B(n20062), .ZN(n19354) );
  NAND2_X1 U22327 ( .A1(n19364), .A2(n19363), .ZN(n19362) );
  NAND2_X1 U22328 ( .A1(n19354), .A2(n19362), .ZN(n19353) );
  OAI21_X1 U22329 ( .B1(n20060), .B2(n20062), .A(n19353), .ZN(n19348) );
  NAND2_X1 U22330 ( .A1(n19349), .A2(n19348), .ZN(n19347) );
  OAI21_X1 U22331 ( .B1(n20051), .B2(n20050), .A(n19347), .ZN(n19342) );
  XNOR2_X1 U22332 ( .A(n20039), .B(n20046), .ZN(n19343) );
  NAND2_X1 U22333 ( .A1(n19342), .A2(n19343), .ZN(n19341) );
  OAI21_X1 U22334 ( .B1(n20046), .B2(n19326), .A(n19341), .ZN(n19327) );
  NAND2_X1 U22335 ( .A1(n19327), .A2(n19403), .ZN(n19337) );
  INV_X1 U22336 ( .A(n19336), .ZN(n19328) );
  NAND3_X1 U22337 ( .A1(n19337), .A2(n19328), .A3(n19361), .ZN(n19329) );
  OAI211_X1 U22338 ( .C1(n19331), .C2(n19367), .A(n19330), .B(n19329), .ZN(
        P2_U2914) );
  INV_X1 U22339 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19332) );
  OAI22_X1 U22340 ( .A1(n19403), .A2(n19334), .B1(n19333), .B2(n19332), .ZN(
        n19335) );
  INV_X1 U22341 ( .A(n19335), .ZN(n19340) );
  XNOR2_X1 U22342 ( .A(n19337), .B(n19336), .ZN(n19338) );
  NAND2_X1 U22343 ( .A1(n19338), .A2(n19361), .ZN(n19339) );
  OAI211_X1 U22344 ( .C1(n19452), .C2(n19367), .A(n19340), .B(n19339), .ZN(
        P2_U2915) );
  AOI22_X1 U22345 ( .A1(n20046), .A2(n19360), .B1(n19359), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19346) );
  OAI21_X1 U22346 ( .B1(n19343), .B2(n19342), .A(n19341), .ZN(n19344) );
  NAND2_X1 U22347 ( .A1(n19344), .A2(n19361), .ZN(n19345) );
  OAI211_X1 U22348 ( .C1(n19446), .C2(n19367), .A(n19346), .B(n19345), .ZN(
        P2_U2916) );
  AOI22_X1 U22349 ( .A1(n19360), .A2(n20050), .B1(n19359), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n19352) );
  OAI21_X1 U22350 ( .B1(n19349), .B2(n19348), .A(n19347), .ZN(n19350) );
  NAND2_X1 U22351 ( .A1(n19350), .A2(n19361), .ZN(n19351) );
  OAI211_X1 U22352 ( .C1(n19440), .C2(n19367), .A(n19352), .B(n19351), .ZN(
        P2_U2917) );
  AOI22_X1 U22353 ( .A1(n19360), .A2(n20062), .B1(n19359), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19357) );
  OAI21_X1 U22354 ( .B1(n19354), .B2(n19362), .A(n19353), .ZN(n19355) );
  NAND2_X1 U22355 ( .A1(n19355), .A2(n19361), .ZN(n19356) );
  OAI211_X1 U22356 ( .C1(n19358), .C2(n19367), .A(n19357), .B(n19356), .ZN(
        P2_U2918) );
  AOI22_X1 U22357 ( .A1(n19363), .A2(n19360), .B1(n19359), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19366) );
  OAI211_X1 U22358 ( .C1(n19364), .C2(n19363), .A(n19362), .B(n19361), .ZN(
        n19365) );
  OAI211_X1 U22359 ( .C1(n19368), .C2(n19367), .A(n19366), .B(n19365), .ZN(
        P2_U2919) );
  AND2_X1 U22360 ( .A1(n19384), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  INV_X1 U22361 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19371) );
  AOI22_X1 U22362 ( .A1(n19400), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19370) );
  OAI21_X1 U22363 ( .B1(n19371), .B2(n19402), .A(n19370), .ZN(P2_U2936) );
  AOI22_X1 U22364 ( .A1(n19400), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19372) );
  OAI21_X1 U22365 ( .B1(n19373), .B2(n19402), .A(n19372), .ZN(P2_U2937) );
  AOI22_X1 U22366 ( .A1(n19400), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19374) );
  OAI21_X1 U22367 ( .B1(n19375), .B2(n19402), .A(n19374), .ZN(P2_U2938) );
  AOI22_X1 U22368 ( .A1(n19376), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19377) );
  OAI21_X1 U22369 ( .B1(n19378), .B2(n19402), .A(n19377), .ZN(P2_U2939) );
  INV_X1 U22370 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19380) );
  AOI22_X1 U22371 ( .A1(n19400), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19384), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19379) );
  OAI21_X1 U22372 ( .B1(n19380), .B2(n19402), .A(n19379), .ZN(P2_U2940) );
  AOI22_X1 U22373 ( .A1(n19400), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19384), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19381) );
  OAI21_X1 U22374 ( .B1(n19382), .B2(n19402), .A(n19381), .ZN(P2_U2941) );
  AOI22_X1 U22375 ( .A1(n19400), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19384), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19383) );
  OAI21_X1 U22376 ( .B1(n11320), .B2(n19402), .A(n19383), .ZN(P2_U2942) );
  AOI22_X1 U22377 ( .A1(n19400), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19384), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19385) );
  OAI21_X1 U22378 ( .B1(n19386), .B2(n19402), .A(n19385), .ZN(P2_U2943) );
  AOI22_X1 U22379 ( .A1(n19400), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19387) );
  OAI21_X1 U22380 ( .B1(n19388), .B2(n19402), .A(n19387), .ZN(P2_U2944) );
  AOI22_X1 U22381 ( .A1(n19400), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19389) );
  OAI21_X1 U22382 ( .B1(n19317), .B2(n19402), .A(n19389), .ZN(P2_U2945) );
  INV_X1 U22383 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19391) );
  AOI22_X1 U22384 ( .A1(n19400), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19390) );
  OAI21_X1 U22385 ( .B1(n19391), .B2(n19402), .A(n19390), .ZN(P2_U2946) );
  AOI22_X1 U22386 ( .A1(n19400), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19392) );
  OAI21_X1 U22387 ( .B1(n19332), .B2(n19402), .A(n19392), .ZN(P2_U2947) );
  INV_X1 U22388 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19394) );
  AOI22_X1 U22389 ( .A1(n19400), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19393) );
  OAI21_X1 U22390 ( .B1(n19394), .B2(n19402), .A(n19393), .ZN(P2_U2948) );
  INV_X1 U22391 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19396) );
  AOI22_X1 U22392 ( .A1(n19400), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19395) );
  OAI21_X1 U22393 ( .B1(n19396), .B2(n19402), .A(n19395), .ZN(P2_U2949) );
  INV_X1 U22394 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19398) );
  AOI22_X1 U22395 ( .A1(n19400), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19397) );
  OAI21_X1 U22396 ( .B1(n19398), .B2(n19402), .A(n19397), .ZN(P2_U2950) );
  AOI22_X1 U22397 ( .A1(n19400), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19399), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19401) );
  OAI21_X1 U22398 ( .B1(n11261), .B2(n19402), .A(n19401), .ZN(P2_U2951) );
  INV_X1 U22399 ( .A(n19403), .ZN(n19410) );
  NAND2_X1 U22400 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19404), .ZN(n19405) );
  OAI221_X1 U22401 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19408), .C1(
        n19407), .C2(n19406), .A(n19405), .ZN(n19409) );
  AOI21_X1 U22402 ( .B1(n19420), .B2(n19410), .A(n19409), .ZN(n19417) );
  NOR2_X1 U22403 ( .A1(n19412), .A2(n19411), .ZN(n19413) );
  AOI21_X1 U22404 ( .B1(n19415), .B2(n19414), .A(n19413), .ZN(n19416) );
  OAI211_X1 U22405 ( .C1(n19419), .C2(n19418), .A(n19417), .B(n19416), .ZN(
        P2_U3042) );
  NAND2_X1 U22406 ( .A1(n19420), .A2(n20062), .ZN(n19421) );
  OAI21_X1 U22407 ( .B1(n19423), .B2(n19422), .A(n19421), .ZN(n19424) );
  INV_X1 U22408 ( .A(n19424), .ZN(n19433) );
  NAND2_X1 U22409 ( .A1(n14475), .A2(n19425), .ZN(n19432) );
  OAI211_X1 U22410 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n19427), .B(n19426), .ZN(n19431) );
  NAND2_X1 U22411 ( .A1(n19429), .A2(n19428), .ZN(n19430) );
  AND4_X1 U22412 ( .A1(n19433), .A2(n19432), .A3(n19431), .A4(n19430), .ZN(
        n19435) );
  OAI211_X1 U22413 ( .C1(n19437), .C2(n19436), .A(n19435), .B(n19434), .ZN(
        P2_U3045) );
  INV_X1 U22414 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19444) );
  INV_X1 U22415 ( .A(n19934), .ZN(n19462) );
  NOR2_X2 U22416 ( .A1(n19439), .A2(n19459), .ZN(n19902) );
  AOI22_X1 U22417 ( .A1(n19903), .A2(n19462), .B1(n19461), .B2(n19902), .ZN(
        n19443) );
  AOI22_X1 U22418 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19466), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19465), .ZN(n19906) );
  AOI22_X1 U22419 ( .A1(n19441), .A2(n19467), .B1(n19496), .B2(n19856), .ZN(
        n19442) );
  OAI211_X1 U22420 ( .C1(n19471), .C2(n19444), .A(n19443), .B(n19442), .ZN(
        P2_U3050) );
  AOI22_X1 U22421 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19465), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19466), .ZN(n19817) );
  INV_X1 U22422 ( .A(n19817), .ZN(n19908) );
  NOR2_X2 U22423 ( .A1(n19445), .A2(n19459), .ZN(n19907) );
  AOI22_X1 U22424 ( .A1(n19462), .A2(n19908), .B1(n19461), .B2(n19907), .ZN(
        n19449) );
  AOI22_X1 U22425 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19466), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19465), .ZN(n19911) );
  AOI22_X1 U22426 ( .A1(n19447), .A2(n19467), .B1(n19496), .B2(n19860), .ZN(
        n19448) );
  OAI211_X1 U22427 ( .C1(n19471), .C2(n10661), .A(n19449), .B(n19448), .ZN(
        P2_U3051) );
  NOR2_X2 U22428 ( .A1(n19451), .A2(n19459), .ZN(n19912) );
  AOI22_X1 U22429 ( .A1(n19913), .A2(n19462), .B1(n19461), .B2(n19912), .ZN(
        n19455) );
  AOI22_X1 U22430 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19466), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19465), .ZN(n19916) );
  AOI22_X1 U22431 ( .A1(n19453), .A2(n19467), .B1(n19496), .B2(n19863), .ZN(
        n19454) );
  OAI211_X1 U22432 ( .C1(n19471), .C2(n11780), .A(n19455), .B(n19454), .ZN(
        P2_U3052) );
  NOR2_X2 U22433 ( .A1(n19460), .A2(n19459), .ZN(n19926) );
  AOI22_X1 U22434 ( .A1(n19929), .A2(n19462), .B1(n19461), .B2(n19926), .ZN(
        n19469) );
  AOI22_X1 U22435 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19466), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19465), .ZN(n19935) );
  AOI22_X1 U22436 ( .A1(n19464), .A2(n19467), .B1(n19496), .B2(n19875), .ZN(
        n19468) );
  OAI211_X1 U22437 ( .C1(n19471), .C2(n19470), .A(n19469), .B(n19468), .ZN(
        P2_U3055) );
  NOR2_X1 U22438 ( .A1(n19501), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19479) );
  INV_X1 U22439 ( .A(n19479), .ZN(n19475) );
  INV_X1 U22440 ( .A(n19472), .ZN(n19473) );
  NOR2_X1 U22441 ( .A1(n19698), .A2(n19501), .ZN(n19494) );
  NOR3_X1 U22442 ( .A1(n19473), .A2(n19494), .A3(n20067), .ZN(n19476) );
  AOI211_X2 U22443 ( .C1(n19475), .C2(n20067), .A(n19474), .B(n19476), .ZN(
        n19495) );
  AOI22_X1 U22444 ( .A1(n19495), .A2(n13117), .B1(n19885), .B2(n19494), .ZN(
        n19481) );
  INV_X1 U22445 ( .A(n19494), .ZN(n19477) );
  AOI211_X1 U22446 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19477), .A(n19888), 
        .B(n19476), .ZN(n19478) );
  OAI221_X1 U22447 ( .B1(n19479), .B2(n19699), .C1(n19479), .C2(n19585), .A(
        n19478), .ZN(n19497) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19894), .ZN(n19480) );
  OAI211_X1 U22449 ( .C1(n19897), .C2(n19530), .A(n19481), .B(n19480), .ZN(
        P2_U3056) );
  AOI22_X1 U22450 ( .A1(n19495), .A2(n13681), .B1(n13683), .B2(n19494), .ZN(
        n19483) );
  INV_X1 U22451 ( .A(n19811), .ZN(n19898) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19898), .ZN(n19482) );
  OAI211_X1 U22453 ( .C1(n19901), .C2(n19530), .A(n19483), .B(n19482), .ZN(
        P2_U3057) );
  AOI22_X1 U22454 ( .A1(n19495), .A2(n19441), .B1(n19902), .B2(n19494), .ZN(
        n19485) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19903), .ZN(n19484) );
  OAI211_X1 U22456 ( .C1(n19906), .C2(n19530), .A(n19485), .B(n19484), .ZN(
        P2_U3058) );
  AOI22_X1 U22457 ( .A1(n19495), .A2(n19447), .B1(n19907), .B2(n19494), .ZN(
        n19487) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19908), .ZN(n19486) );
  OAI211_X1 U22459 ( .C1(n19911), .C2(n19530), .A(n19487), .B(n19486), .ZN(
        P2_U3059) );
  AOI22_X1 U22460 ( .A1(n19495), .A2(n19453), .B1(n19912), .B2(n19494), .ZN(
        n19489) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19913), .ZN(n19488) );
  OAI211_X1 U22462 ( .C1(n19916), .C2(n19530), .A(n19489), .B(n19488), .ZN(
        P2_U3060) );
  AOI22_X1 U22463 ( .A1(n19495), .A2(n13305), .B1(n13312), .B2(n19494), .ZN(
        n19491) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19917), .ZN(n19490) );
  OAI211_X1 U22465 ( .C1(n19920), .C2(n19530), .A(n19491), .B(n19490), .ZN(
        P2_U3061) );
  AOI22_X1 U22466 ( .A1(n19495), .A2(n13101), .B1(n19921), .B2(n19494), .ZN(
        n19493) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19922), .ZN(n19492) );
  OAI211_X1 U22468 ( .C1(n19925), .C2(n19530), .A(n19493), .B(n19492), .ZN(
        P2_U3062) );
  AOI22_X1 U22469 ( .A1(n19495), .A2(n19464), .B1(n19926), .B2(n19494), .ZN(
        n19499) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19497), .B1(
        n19496), .B2(n19929), .ZN(n19498) );
  OAI211_X1 U22471 ( .C1(n19935), .C2(n19530), .A(n19499), .B(n19498), .ZN(
        P2_U3063) );
  INV_X1 U22472 ( .A(n19500), .ZN(n19506) );
  NOR2_X1 U22473 ( .A1(n19729), .A2(n19501), .ZN(n19525) );
  OAI21_X1 U22474 ( .B1(n19506), .B2(n19525), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19503) );
  NOR2_X1 U22475 ( .A1(n19732), .A2(n19501), .ZN(n19504) );
  INV_X1 U22476 ( .A(n19504), .ZN(n19502) );
  NAND2_X1 U22477 ( .A1(n19503), .A2(n19502), .ZN(n19526) );
  AOI22_X1 U22478 ( .A1(n19526), .A2(n13117), .B1(n19885), .B2(n19525), .ZN(
        n19511) );
  NAND2_X1 U22479 ( .A1(n19541), .A2(n19530), .ZN(n19505) );
  AOI21_X1 U22480 ( .B1(n19505), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19504), 
        .ZN(n19508) );
  AOI21_X1 U22481 ( .B1(n19506), .B2(n13298), .A(n19525), .ZN(n19507) );
  MUX2_X1 U22482 ( .A(n19508), .B(n19507), .S(n20042), .Z(n19509) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19527), .B1(
        n19547), .B2(n19805), .ZN(n19510) );
  OAI211_X1 U22484 ( .C1(n19808), .C2(n19530), .A(n19511), .B(n19510), .ZN(
        P2_U3064) );
  AOI22_X1 U22485 ( .A1(n19526), .A2(n13681), .B1(n13683), .B2(n19525), .ZN(
        n19513) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19527), .B1(
        n19547), .B2(n19853), .ZN(n19512) );
  OAI211_X1 U22487 ( .C1(n19811), .C2(n19530), .A(n19513), .B(n19512), .ZN(
        P2_U3065) );
  INV_X1 U22488 ( .A(n19903), .ZN(n19814) );
  AOI22_X1 U22489 ( .A1(n19526), .A2(n19441), .B1(n19902), .B2(n19525), .ZN(
        n19515) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19527), .B1(
        n19547), .B2(n19856), .ZN(n19514) );
  OAI211_X1 U22491 ( .C1(n19814), .C2(n19530), .A(n19515), .B(n19514), .ZN(
        P2_U3066) );
  AOI22_X1 U22492 ( .A1(n19526), .A2(n19447), .B1(n19907), .B2(n19525), .ZN(
        n19517) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19527), .B1(
        n19547), .B2(n19860), .ZN(n19516) );
  OAI211_X1 U22494 ( .C1(n19817), .C2(n19530), .A(n19517), .B(n19516), .ZN(
        P2_U3067) );
  AOI22_X1 U22495 ( .A1(n19526), .A2(n19453), .B1(n19912), .B2(n19525), .ZN(
        n19519) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19527), .B1(
        n19547), .B2(n19863), .ZN(n19518) );
  OAI211_X1 U22497 ( .C1(n19820), .C2(n19530), .A(n19519), .B(n19518), .ZN(
        P2_U3068) );
  AOI22_X1 U22498 ( .A1(n19526), .A2(n13305), .B1(n13312), .B2(n19525), .ZN(
        n19521) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19527), .B1(
        n19522), .B2(n19917), .ZN(n19520) );
  OAI211_X1 U22500 ( .C1(n19920), .C2(n19541), .A(n19521), .B(n19520), .ZN(
        P2_U3069) );
  AOI22_X1 U22501 ( .A1(n19526), .A2(n13101), .B1(n19921), .B2(n19525), .ZN(
        n19524) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19527), .B1(
        n19522), .B2(n19922), .ZN(n19523) );
  OAI211_X1 U22503 ( .C1(n19925), .C2(n19541), .A(n19524), .B(n19523), .ZN(
        P2_U3070) );
  AOI22_X1 U22504 ( .A1(n19526), .A2(n19464), .B1(n19926), .B2(n19525), .ZN(
        n19529) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19527), .B1(
        n19547), .B2(n19875), .ZN(n19528) );
  OAI211_X1 U22506 ( .C1(n19833), .C2(n19530), .A(n19529), .B(n19528), .ZN(
        P2_U3071) );
  AOI22_X1 U22507 ( .A1(n19574), .A2(n19805), .B1(n19885), .B2(n19546), .ZN(
        n19532) );
  AOI22_X1 U22508 ( .A1(n13117), .A2(n19548), .B1(n19547), .B2(n19894), .ZN(
        n19531) );
  OAI211_X1 U22509 ( .C1(n19534), .C2(n19533), .A(n19532), .B(n19531), .ZN(
        P2_U3072) );
  AOI22_X1 U22510 ( .A1(n19574), .A2(n19853), .B1(n13683), .B2(n19546), .ZN(
        n19536) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19549), .B1(
        n13681), .B2(n19548), .ZN(n19535) );
  OAI211_X1 U22512 ( .C1(n19811), .C2(n19541), .A(n19536), .B(n19535), .ZN(
        P2_U3073) );
  AOI22_X1 U22513 ( .A1(n19547), .A2(n19903), .B1(n19546), .B2(n19902), .ZN(
        n19538) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19549), .B1(
        n19441), .B2(n19548), .ZN(n19537) );
  OAI211_X1 U22515 ( .C1(n19906), .C2(n19582), .A(n19538), .B(n19537), .ZN(
        P2_U3074) );
  AOI22_X1 U22516 ( .A1(n19574), .A2(n19860), .B1(n19546), .B2(n19907), .ZN(
        n19540) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19549), .B1(
        n19447), .B2(n19548), .ZN(n19539) );
  OAI211_X1 U22518 ( .C1(n19817), .C2(n19541), .A(n19540), .B(n19539), .ZN(
        P2_U3075) );
  AOI22_X1 U22519 ( .A1(n19547), .A2(n19913), .B1(n19546), .B2(n19912), .ZN(
        n19543) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19549), .B1(
        n19453), .B2(n19548), .ZN(n19542) );
  OAI211_X1 U22521 ( .C1(n19916), .C2(n19582), .A(n19543), .B(n19542), .ZN(
        P2_U3076) );
  AOI22_X1 U22522 ( .A1(n19547), .A2(n19922), .B1(n19921), .B2(n19546), .ZN(
        n19545) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19549), .B1(
        n13101), .B2(n19548), .ZN(n19544) );
  OAI211_X1 U22524 ( .C1(n19925), .C2(n19582), .A(n19545), .B(n19544), .ZN(
        P2_U3078) );
  AOI22_X1 U22525 ( .A1(n19547), .A2(n19929), .B1(n19546), .B2(n19926), .ZN(
        n19551) );
  AOI22_X1 U22526 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19549), .B1(
        n19464), .B2(n19548), .ZN(n19550) );
  OAI211_X1 U22527 ( .C1(n19935), .C2(n19582), .A(n19551), .B(n19550), .ZN(
        P2_U3079) );
  NOR2_X1 U22528 ( .A1(n19553), .A2(n19552), .ZN(n19794) );
  NAND2_X1 U22529 ( .A1(n19794), .A2(n20048), .ZN(n19560) );
  OR2_X1 U22530 ( .A1(n19560), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19556) );
  INV_X1 U22531 ( .A(n19554), .ZN(n19555) );
  NAND3_X1 U22532 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20048), .A3(
        n20064), .ZN(n19589) );
  NOR2_X1 U22533 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19589), .ZN(
        n19577) );
  NOR3_X1 U22534 ( .A1(n19555), .A2(n19577), .A3(n20067), .ZN(n19558) );
  AOI21_X1 U22535 ( .B1(n20067), .B2(n19556), .A(n19558), .ZN(n19578) );
  AOI22_X1 U22536 ( .A1(n19578), .A2(n13117), .B1(n19885), .B2(n19577), .ZN(
        n19563) );
  OAI21_X1 U22537 ( .B1(n19574), .B2(n19612), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19559) );
  AOI211_X1 U22538 ( .C1(n19560), .C2(n19559), .A(n19888), .B(n19558), .ZN(
        n19561) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19579), .B1(
        n19612), .B2(n19805), .ZN(n19562) );
  OAI211_X1 U22540 ( .C1(n19808), .C2(n19582), .A(n19563), .B(n19562), .ZN(
        P2_U3080) );
  AOI22_X1 U22541 ( .A1(n19578), .A2(n13681), .B1(n13683), .B2(n19577), .ZN(
        n19565) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19579), .B1(
        n19612), .B2(n19853), .ZN(n19564) );
  OAI211_X1 U22543 ( .C1(n19811), .C2(n19582), .A(n19565), .B(n19564), .ZN(
        P2_U3081) );
  AOI22_X1 U22544 ( .A1(n19578), .A2(n19441), .B1(n19902), .B2(n19577), .ZN(
        n19567) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19579), .B1(
        n19612), .B2(n19856), .ZN(n19566) );
  OAI211_X1 U22546 ( .C1(n19814), .C2(n19582), .A(n19567), .B(n19566), .ZN(
        P2_U3082) );
  AOI22_X1 U22547 ( .A1(n19578), .A2(n19447), .B1(n19907), .B2(n19577), .ZN(
        n19569) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19579), .B1(
        n19612), .B2(n19860), .ZN(n19568) );
  OAI211_X1 U22549 ( .C1(n19817), .C2(n19582), .A(n19569), .B(n19568), .ZN(
        P2_U3083) );
  AOI22_X1 U22550 ( .A1(n19578), .A2(n19453), .B1(n19912), .B2(n19577), .ZN(
        n19571) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19579), .B1(
        n19612), .B2(n19863), .ZN(n19570) );
  OAI211_X1 U22552 ( .C1(n19820), .C2(n19582), .A(n19571), .B(n19570), .ZN(
        P2_U3084) );
  AOI22_X1 U22553 ( .A1(n19578), .A2(n13305), .B1(n13312), .B2(n19577), .ZN(
        n19573) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19579), .B1(
        n19574), .B2(n19917), .ZN(n19572) );
  OAI211_X1 U22555 ( .C1(n19920), .C2(n19619), .A(n19573), .B(n19572), .ZN(
        P2_U3085) );
  AOI22_X1 U22556 ( .A1(n19578), .A2(n13101), .B1(n19921), .B2(n19577), .ZN(
        n19576) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19579), .B1(
        n19574), .B2(n19922), .ZN(n19575) );
  OAI211_X1 U22558 ( .C1(n19925), .C2(n19619), .A(n19576), .B(n19575), .ZN(
        P2_U3086) );
  AOI22_X1 U22559 ( .A1(n19578), .A2(n19464), .B1(n19926), .B2(n19577), .ZN(
        n19581) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19579), .B1(
        n19612), .B2(n19875), .ZN(n19580) );
  OAI211_X1 U22561 ( .C1(n19833), .C2(n19582), .A(n19581), .B(n19580), .ZN(
        P2_U3087) );
  NOR2_X1 U22562 ( .A1(n20074), .A2(n19589), .ZN(n19626) );
  INV_X1 U22563 ( .A(n19626), .ZN(n19583) );
  OAI21_X1 U22564 ( .B1(n19592), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19583), 
        .ZN(n19587) );
  NAND2_X1 U22565 ( .A1(n19585), .A2(n19584), .ZN(n19591) );
  NAND2_X1 U22566 ( .A1(n19591), .A2(n19589), .ZN(n19586) );
  MUX2_X1 U22567 ( .A(n19587), .B(n19586), .S(n20037), .Z(n19588) );
  AND2_X1 U22568 ( .A1(n19588), .A2(n19737), .ZN(n19601) );
  AOI22_X1 U22569 ( .A1(n19612), .A2(n19894), .B1(n19885), .B2(n19626), .ZN(
        n19599) );
  INV_X1 U22570 ( .A(n19589), .ZN(n19590) );
  NAND3_X1 U22571 ( .A1(n19591), .A2(n20037), .A3(n19590), .ZN(n19595) );
  INV_X1 U22572 ( .A(n19592), .ZN(n19593) );
  OAI21_X1 U22573 ( .B1(n19593), .B2(n19626), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19594) );
  NAND2_X1 U22574 ( .A1(n19595), .A2(n19594), .ZN(n19615) );
  AOI22_X1 U22575 ( .A1(n13117), .A2(n19615), .B1(n19646), .B2(n19805), .ZN(
        n19598) );
  OAI211_X1 U22576 ( .C1(n19601), .C2(n19600), .A(n19599), .B(n19598), .ZN(
        P2_U3088) );
  AOI22_X1 U22577 ( .A1(n19646), .A2(n19853), .B1(n13683), .B2(n19626), .ZN(
        n19603) );
  AOI22_X1 U22578 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19616), .B1(
        n13681), .B2(n19615), .ZN(n19602) );
  OAI211_X1 U22579 ( .C1(n19811), .C2(n19619), .A(n19603), .B(n19602), .ZN(
        P2_U3089) );
  AOI22_X1 U22580 ( .A1(n19612), .A2(n19903), .B1(n19626), .B2(n19902), .ZN(
        n19605) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19616), .B1(
        n19441), .B2(n19615), .ZN(n19604) );
  OAI211_X1 U22582 ( .C1(n19906), .C2(n19641), .A(n19605), .B(n19604), .ZN(
        P2_U3090) );
  AOI22_X1 U22583 ( .A1(n19612), .A2(n19908), .B1(n19626), .B2(n19907), .ZN(
        n19607) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19616), .B1(
        n19447), .B2(n19615), .ZN(n19606) );
  OAI211_X1 U22585 ( .C1(n19911), .C2(n19641), .A(n19607), .B(n19606), .ZN(
        P2_U3091) );
  AOI22_X1 U22586 ( .A1(n19646), .A2(n19863), .B1(n19626), .B2(n19912), .ZN(
        n19609) );
  AOI22_X1 U22587 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19616), .B1(
        n19453), .B2(n19615), .ZN(n19608) );
  OAI211_X1 U22588 ( .C1(n19820), .C2(n19619), .A(n19609), .B(n19608), .ZN(
        P2_U3092) );
  AOI22_X1 U22589 ( .A1(n19646), .A2(n19867), .B1(n13312), .B2(n19626), .ZN(
        n19611) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19616), .B1(
        n13305), .B2(n19615), .ZN(n19610) );
  OAI211_X1 U22591 ( .C1(n19823), .C2(n19619), .A(n19611), .B(n19610), .ZN(
        P2_U3093) );
  AOI22_X1 U22592 ( .A1(n19612), .A2(n19922), .B1(n19921), .B2(n19626), .ZN(
        n19614) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19616), .B1(
        n13101), .B2(n19615), .ZN(n19613) );
  OAI211_X1 U22594 ( .C1(n19925), .C2(n19641), .A(n19614), .B(n19613), .ZN(
        P2_U3094) );
  AOI22_X1 U22595 ( .A1(n19646), .A2(n19875), .B1(n19626), .B2(n19926), .ZN(
        n19618) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19616), .B1(
        n19464), .B2(n19615), .ZN(n19617) );
  OAI211_X1 U22597 ( .C1(n19833), .C2(n19619), .A(n19618), .B(n19617), .ZN(
        P2_U3095) );
  NOR2_X1 U22598 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19620), .ZN(
        n19644) );
  NOR2_X1 U22599 ( .A1(n19626), .A2(n19644), .ZN(n19621) );
  OR2_X1 U22600 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19621), .ZN(n19624) );
  INV_X1 U22601 ( .A(n19622), .ZN(n19623) );
  NOR3_X1 U22602 ( .A1(n19623), .A2(n19644), .A3(n20067), .ZN(n19627) );
  AOI21_X1 U22603 ( .B1(n20067), .B2(n19624), .A(n19627), .ZN(n19645) );
  AOI22_X1 U22604 ( .A1(n19645), .A2(n13117), .B1(n19885), .B2(n19644), .ZN(
        n19630) );
  AOI21_X1 U22605 ( .B1(n19641), .B2(n19665), .A(n12350), .ZN(n19625) );
  AOI221_X1 U22606 ( .B1(n13298), .B2(n19626), .C1(n13298), .C2(n19625), .A(
        n19644), .ZN(n19628) );
  AOI22_X1 U22607 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19647), .B1(
        n19658), .B2(n19805), .ZN(n19629) );
  OAI211_X1 U22608 ( .C1(n19808), .C2(n19641), .A(n19630), .B(n19629), .ZN(
        P2_U3096) );
  AOI22_X1 U22609 ( .A1(n19645), .A2(n13681), .B1(n13683), .B2(n19644), .ZN(
        n19632) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19647), .B1(
        n19658), .B2(n19853), .ZN(n19631) );
  OAI211_X1 U22611 ( .C1(n19811), .C2(n19641), .A(n19632), .B(n19631), .ZN(
        P2_U3097) );
  AOI22_X1 U22612 ( .A1(n19645), .A2(n19441), .B1(n19902), .B2(n19644), .ZN(
        n19634) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19647), .B1(
        n19658), .B2(n19856), .ZN(n19633) );
  OAI211_X1 U22614 ( .C1(n19814), .C2(n19641), .A(n19634), .B(n19633), .ZN(
        P2_U3098) );
  AOI22_X1 U22615 ( .A1(n19645), .A2(n19447), .B1(n19907), .B2(n19644), .ZN(
        n19636) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19647), .B1(
        n19658), .B2(n19860), .ZN(n19635) );
  OAI211_X1 U22617 ( .C1(n19817), .C2(n19641), .A(n19636), .B(n19635), .ZN(
        P2_U3099) );
  AOI22_X1 U22618 ( .A1(n19645), .A2(n19453), .B1(n19912), .B2(n19644), .ZN(
        n19638) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19647), .B1(
        n19658), .B2(n19863), .ZN(n19637) );
  OAI211_X1 U22620 ( .C1(n19820), .C2(n19641), .A(n19638), .B(n19637), .ZN(
        P2_U3100) );
  AOI22_X1 U22621 ( .A1(n19645), .A2(n13305), .B1(n13312), .B2(n19644), .ZN(
        n19640) );
  AOI22_X1 U22622 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19647), .B1(
        n19658), .B2(n19867), .ZN(n19639) );
  OAI211_X1 U22623 ( .C1(n19823), .C2(n19641), .A(n19640), .B(n19639), .ZN(
        P2_U3101) );
  AOI22_X1 U22624 ( .A1(n19645), .A2(n13101), .B1(n19921), .B2(n19644), .ZN(
        n19643) );
  AOI22_X1 U22625 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19647), .B1(
        n19646), .B2(n19922), .ZN(n19642) );
  OAI211_X1 U22626 ( .C1(n19925), .C2(n19665), .A(n19643), .B(n19642), .ZN(
        P2_U3102) );
  AOI22_X1 U22627 ( .A1(n19645), .A2(n19464), .B1(n19926), .B2(n19644), .ZN(
        n19649) );
  AOI22_X1 U22628 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19647), .B1(
        n19646), .B2(n19929), .ZN(n19648) );
  OAI211_X1 U22629 ( .C1(n19935), .C2(n19665), .A(n19649), .B(n19648), .ZN(
        P2_U3103) );
  AOI22_X1 U22630 ( .A1(n19661), .A2(n13681), .B1(n19673), .B2(n13683), .ZN(
        n19651) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19662), .B1(
        n19658), .B2(n19898), .ZN(n19650) );
  OAI211_X1 U22632 ( .C1(n19901), .C2(n19697), .A(n19651), .B(n19650), .ZN(
        P2_U3105) );
  AOI22_X1 U22633 ( .A1(n19661), .A2(n19441), .B1(n19673), .B2(n19902), .ZN(
        n19653) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19662), .B1(
        n19658), .B2(n19903), .ZN(n19652) );
  OAI211_X1 U22635 ( .C1(n19906), .C2(n19697), .A(n19653), .B(n19652), .ZN(
        P2_U3106) );
  AOI22_X1 U22636 ( .A1(n19661), .A2(n19447), .B1(n19673), .B2(n19907), .ZN(
        n19655) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19662), .B1(
        n19658), .B2(n19908), .ZN(n19654) );
  OAI211_X1 U22638 ( .C1(n19911), .C2(n19697), .A(n19655), .B(n19654), .ZN(
        P2_U3107) );
  AOI22_X1 U22639 ( .A1(n19661), .A2(n19453), .B1(n19673), .B2(n19912), .ZN(
        n19657) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19662), .B1(
        n19689), .B2(n19863), .ZN(n19656) );
  OAI211_X1 U22641 ( .C1(n19820), .C2(n19665), .A(n19657), .B(n19656), .ZN(
        P2_U3108) );
  AOI22_X1 U22642 ( .A1(n19661), .A2(n13305), .B1(n19673), .B2(n13312), .ZN(
        n19660) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19662), .B1(
        n19658), .B2(n19917), .ZN(n19659) );
  OAI211_X1 U22644 ( .C1(n19920), .C2(n19697), .A(n19660), .B(n19659), .ZN(
        P2_U3109) );
  AOI22_X1 U22645 ( .A1(n19661), .A2(n19464), .B1(n19673), .B2(n19926), .ZN(
        n19664) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19662), .B1(
        n19689), .B2(n19875), .ZN(n19663) );
  OAI211_X1 U22647 ( .C1(n19833), .C2(n19665), .A(n19664), .B(n19663), .ZN(
        P2_U3111) );
  NAND2_X1 U22648 ( .A1(n20056), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19764) );
  OR2_X1 U22649 ( .A1(n19764), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19707) );
  NOR2_X1 U22650 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19707), .ZN(
        n19692) );
  AOI22_X1 U22651 ( .A1(n19724), .A2(n19805), .B1(n19885), .B2(n19692), .ZN(
        n19678) );
  AOI21_X1 U22652 ( .B1(n19697), .B2(n19723), .A(n12350), .ZN(n19667) );
  NOR2_X1 U22653 ( .A1(n19667), .A2(n20042), .ZN(n19672) );
  INV_X1 U22654 ( .A(n19668), .ZN(n19674) );
  OAI21_X1 U22655 ( .B1(n19674), .B2(n20067), .A(n13298), .ZN(n19669) );
  AOI21_X1 U22656 ( .B1(n19672), .B2(n19670), .A(n19669), .ZN(n19671) );
  OAI21_X1 U22657 ( .B1(n19692), .B2(n19671), .A(n19737), .ZN(n19694) );
  OAI21_X1 U22658 ( .B1(n19692), .B2(n19673), .A(n19672), .ZN(n19676) );
  OAI21_X1 U22659 ( .B1(n19674), .B2(n19692), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19675) );
  NAND2_X1 U22660 ( .A1(n19676), .A2(n19675), .ZN(n19693) );
  AOI22_X1 U22661 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19694), .B1(
        n13117), .B2(n19693), .ZN(n19677) );
  OAI211_X1 U22662 ( .C1(n19808), .C2(n19697), .A(n19678), .B(n19677), .ZN(
        P2_U3112) );
  AOI22_X1 U22663 ( .A1(n19724), .A2(n19853), .B1(n13683), .B2(n19692), .ZN(
        n19680) );
  AOI22_X1 U22664 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19694), .B1(
        n13681), .B2(n19693), .ZN(n19679) );
  OAI211_X1 U22665 ( .C1(n19811), .C2(n19697), .A(n19680), .B(n19679), .ZN(
        P2_U3113) );
  AOI22_X1 U22666 ( .A1(n19724), .A2(n19856), .B1(n19902), .B2(n19692), .ZN(
        n19682) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19694), .B1(
        n19441), .B2(n19693), .ZN(n19681) );
  OAI211_X1 U22668 ( .C1(n19814), .C2(n19697), .A(n19682), .B(n19681), .ZN(
        P2_U3114) );
  AOI22_X1 U22669 ( .A1(n19724), .A2(n19860), .B1(n19907), .B2(n19692), .ZN(
        n19684) );
  AOI22_X1 U22670 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19694), .B1(
        n19447), .B2(n19693), .ZN(n19683) );
  OAI211_X1 U22671 ( .C1(n19817), .C2(n19697), .A(n19684), .B(n19683), .ZN(
        P2_U3115) );
  AOI22_X1 U22672 ( .A1(n19724), .A2(n19863), .B1(n19912), .B2(n19692), .ZN(
        n19686) );
  AOI22_X1 U22673 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19694), .B1(
        n19453), .B2(n19693), .ZN(n19685) );
  OAI211_X1 U22674 ( .C1(n19820), .C2(n19697), .A(n19686), .B(n19685), .ZN(
        P2_U3116) );
  AOI22_X1 U22675 ( .A1(n19689), .A2(n19917), .B1(n13312), .B2(n19692), .ZN(
        n19688) );
  AOI22_X1 U22676 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19694), .B1(
        n13305), .B2(n19693), .ZN(n19687) );
  OAI211_X1 U22677 ( .C1(n19920), .C2(n19723), .A(n19688), .B(n19687), .ZN(
        P2_U3117) );
  AOI22_X1 U22678 ( .A1(n19689), .A2(n19922), .B1(n19921), .B2(n19692), .ZN(
        n19691) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19694), .B1(
        n13101), .B2(n19693), .ZN(n19690) );
  OAI211_X1 U22680 ( .C1(n19925), .C2(n19723), .A(n19691), .B(n19690), .ZN(
        P2_U3118) );
  AOI22_X1 U22681 ( .A1(n19724), .A2(n19875), .B1(n19926), .B2(n19692), .ZN(
        n19696) );
  AOI22_X1 U22682 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19694), .B1(
        n19464), .B2(n19693), .ZN(n19695) );
  OAI211_X1 U22683 ( .C1(n19833), .C2(n19697), .A(n19696), .B(n19695), .ZN(
        P2_U3119) );
  NOR2_X1 U22684 ( .A1(n19698), .A2(n19764), .ZN(n19734) );
  AOI22_X1 U22685 ( .A1(n19894), .A2(n19724), .B1(n19885), .B2(n19734), .ZN(
        n19710) );
  AOI21_X1 U22686 ( .B1(n19891), .B2(n19699), .A(n20042), .ZN(n19704) );
  INV_X1 U22687 ( .A(n19734), .ZN(n19700) );
  NAND2_X1 U22688 ( .A1(n19701), .A2(n19700), .ZN(n19705) );
  NOR2_X1 U22689 ( .A1(n19705), .A2(n20067), .ZN(n19702) );
  AOI21_X1 U22690 ( .B1(n19704), .B2(n19707), .A(n19702), .ZN(n19703) );
  OAI211_X1 U22691 ( .C1(n19734), .C2(n13298), .A(n19703), .B(n19737), .ZN(
        n19726) );
  INV_X1 U22692 ( .A(n19704), .ZN(n19708) );
  INV_X1 U22693 ( .A(n19705), .ZN(n19706) );
  OAI22_X1 U22694 ( .A1(n19708), .A2(n19707), .B1(n19706), .B2(n20067), .ZN(
        n19725) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19726), .B1(
        n13117), .B2(n19725), .ZN(n19709) );
  OAI211_X1 U22696 ( .C1(n19897), .C2(n19759), .A(n19710), .B(n19709), .ZN(
        P2_U3120) );
  AOI22_X1 U22697 ( .A1(n19724), .A2(n19898), .B1(n13683), .B2(n19734), .ZN(
        n19712) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19726), .B1(
        n13681), .B2(n19725), .ZN(n19711) );
  OAI211_X1 U22699 ( .C1(n19901), .C2(n19759), .A(n19712), .B(n19711), .ZN(
        P2_U3121) );
  AOI22_X1 U22700 ( .A1(n19751), .A2(n19856), .B1(n19902), .B2(n19734), .ZN(
        n19714) );
  AOI22_X1 U22701 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19726), .B1(
        n19441), .B2(n19725), .ZN(n19713) );
  OAI211_X1 U22702 ( .C1(n19814), .C2(n19723), .A(n19714), .B(n19713), .ZN(
        P2_U3122) );
  AOI22_X1 U22703 ( .A1(n19724), .A2(n19908), .B1(n19907), .B2(n19734), .ZN(
        n19716) );
  AOI22_X1 U22704 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19726), .B1(
        n19447), .B2(n19725), .ZN(n19715) );
  OAI211_X1 U22705 ( .C1(n19911), .C2(n19759), .A(n19716), .B(n19715), .ZN(
        P2_U3123) );
  AOI22_X1 U22706 ( .A1(n19913), .A2(n19724), .B1(n19912), .B2(n19734), .ZN(
        n19718) );
  AOI22_X1 U22707 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19726), .B1(
        n19453), .B2(n19725), .ZN(n19717) );
  OAI211_X1 U22708 ( .C1(n19916), .C2(n19759), .A(n19718), .B(n19717), .ZN(
        P2_U3124) );
  AOI22_X1 U22709 ( .A1(n19724), .A2(n19917), .B1(n13312), .B2(n19734), .ZN(
        n19720) );
  AOI22_X1 U22710 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19726), .B1(
        n13305), .B2(n19725), .ZN(n19719) );
  OAI211_X1 U22711 ( .C1(n19920), .C2(n19759), .A(n19720), .B(n19719), .ZN(
        P2_U3125) );
  AOI22_X1 U22712 ( .A1(n19751), .A2(n19870), .B1(n19921), .B2(n19734), .ZN(
        n19722) );
  AOI22_X1 U22713 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19726), .B1(
        n13101), .B2(n19725), .ZN(n19721) );
  OAI211_X1 U22714 ( .C1(n19826), .C2(n19723), .A(n19722), .B(n19721), .ZN(
        P2_U3126) );
  AOI22_X1 U22715 ( .A1(n19929), .A2(n19724), .B1(n19926), .B2(n19734), .ZN(
        n19728) );
  AOI22_X1 U22716 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19726), .B1(
        n19464), .B2(n19725), .ZN(n19727) );
  OAI211_X1 U22717 ( .C1(n19935), .C2(n19759), .A(n19728), .B(n19727), .ZN(
        P2_U3127) );
  INV_X1 U22718 ( .A(n19736), .ZN(n19730) );
  NOR2_X1 U22719 ( .A1(n19729), .A2(n19764), .ZN(n19754) );
  OAI21_X1 U22720 ( .B1(n19730), .B2(n19754), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19731) );
  OAI21_X1 U22721 ( .B1(n19764), .B2(n19732), .A(n19731), .ZN(n19755) );
  AOI22_X1 U22722 ( .A1(n19755), .A2(n13117), .B1(n19885), .B2(n19754), .ZN(
        n19740) );
  AOI221_X1 U22723 ( .B1(n19783), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19751), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19734), .ZN(n19735) );
  AOI211_X1 U22724 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19736), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19735), .ZN(n19738) );
  OAI21_X1 U22725 ( .B1(n19738), .B2(n19754), .A(n19737), .ZN(n19756) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19756), .B1(
        n19783), .B2(n19805), .ZN(n19739) );
  OAI211_X1 U22727 ( .C1(n19808), .C2(n19759), .A(n19740), .B(n19739), .ZN(
        P2_U3128) );
  AOI22_X1 U22728 ( .A1(n19755), .A2(n13681), .B1(n13683), .B2(n19754), .ZN(
        n19742) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19756), .B1(
        n19783), .B2(n19853), .ZN(n19741) );
  OAI211_X1 U22730 ( .C1(n19811), .C2(n19759), .A(n19742), .B(n19741), .ZN(
        P2_U3129) );
  AOI22_X1 U22731 ( .A1(n19755), .A2(n19441), .B1(n19902), .B2(n19754), .ZN(
        n19744) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19756), .B1(
        n19783), .B2(n19856), .ZN(n19743) );
  OAI211_X1 U22733 ( .C1(n19814), .C2(n19759), .A(n19744), .B(n19743), .ZN(
        P2_U3130) );
  AOI22_X1 U22734 ( .A1(n19755), .A2(n19447), .B1(n19907), .B2(n19754), .ZN(
        n19746) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19756), .B1(
        n19783), .B2(n19860), .ZN(n19745) );
  OAI211_X1 U22736 ( .C1(n19817), .C2(n19759), .A(n19746), .B(n19745), .ZN(
        P2_U3131) );
  AOI22_X1 U22737 ( .A1(n19755), .A2(n19453), .B1(n19912), .B2(n19754), .ZN(
        n19748) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19756), .B1(
        n19783), .B2(n19863), .ZN(n19747) );
  OAI211_X1 U22739 ( .C1(n19820), .C2(n19759), .A(n19748), .B(n19747), .ZN(
        P2_U3132) );
  AOI22_X1 U22740 ( .A1(n19755), .A2(n13305), .B1(n13312), .B2(n19754), .ZN(
        n19750) );
  AOI22_X1 U22741 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19756), .B1(
        n19751), .B2(n19917), .ZN(n19749) );
  OAI211_X1 U22742 ( .C1(n19920), .C2(n19793), .A(n19750), .B(n19749), .ZN(
        P2_U3133) );
  AOI22_X1 U22743 ( .A1(n19755), .A2(n13101), .B1(n19921), .B2(n19754), .ZN(
        n19753) );
  AOI22_X1 U22744 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19756), .B1(
        n19751), .B2(n19922), .ZN(n19752) );
  OAI211_X1 U22745 ( .C1(n19925), .C2(n19793), .A(n19753), .B(n19752), .ZN(
        P2_U3134) );
  AOI22_X1 U22746 ( .A1(n19755), .A2(n19464), .B1(n19926), .B2(n19754), .ZN(
        n19758) );
  AOI22_X1 U22747 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19756), .B1(
        n19783), .B2(n19875), .ZN(n19757) );
  OAI211_X1 U22748 ( .C1(n19833), .C2(n19759), .A(n19758), .B(n19757), .ZN(
        P2_U3135) );
  INV_X1 U22749 ( .A(n19764), .ZN(n19761) );
  NAND2_X1 U22750 ( .A1(n19762), .A2(n19761), .ZN(n19769) );
  NAND3_X1 U22751 ( .A1(n19763), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19769), 
        .ZN(n19767) );
  NOR2_X1 U22752 ( .A1(n20064), .A2(n19764), .ZN(n19772) );
  INV_X1 U22753 ( .A(n19772), .ZN(n19765) );
  OAI21_X1 U22754 ( .B1(n19765), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20067), 
        .ZN(n19766) );
  AND2_X1 U22755 ( .A1(n19767), .A2(n19766), .ZN(n19789) );
  INV_X1 U22756 ( .A(n19769), .ZN(n19788) );
  AOI22_X1 U22757 ( .A1(n19789), .A2(n13117), .B1(n19885), .B2(n19788), .ZN(
        n19774) );
  INV_X1 U22758 ( .A(n19767), .ZN(n19768) );
  AOI211_X1 U22759 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19769), .A(n19888), 
        .B(n19768), .ZN(n19770) );
  OAI221_X1 U22760 ( .B1(n19772), .B2(n19771), .C1(n19772), .C2(n19891), .A(
        n19770), .ZN(n19790) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19790), .B1(
        n19783), .B2(n19894), .ZN(n19773) );
  OAI211_X1 U22762 ( .C1(n19897), .C2(n19832), .A(n19774), .B(n19773), .ZN(
        P2_U3136) );
  AOI22_X1 U22763 ( .A1(n19789), .A2(n13681), .B1(n13683), .B2(n19788), .ZN(
        n19776) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19790), .B1(
        n19800), .B2(n19853), .ZN(n19775) );
  OAI211_X1 U22765 ( .C1(n19811), .C2(n19793), .A(n19776), .B(n19775), .ZN(
        P2_U3137) );
  AOI22_X1 U22766 ( .A1(n19789), .A2(n19441), .B1(n19902), .B2(n19788), .ZN(
        n19778) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19790), .B1(
        n19800), .B2(n19856), .ZN(n19777) );
  OAI211_X1 U22768 ( .C1(n19814), .C2(n19793), .A(n19778), .B(n19777), .ZN(
        P2_U3138) );
  AOI22_X1 U22769 ( .A1(n19789), .A2(n19447), .B1(n19907), .B2(n19788), .ZN(
        n19780) );
  AOI22_X1 U22770 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19790), .B1(
        n19783), .B2(n19908), .ZN(n19779) );
  OAI211_X1 U22771 ( .C1(n19911), .C2(n19832), .A(n19780), .B(n19779), .ZN(
        P2_U3139) );
  AOI22_X1 U22772 ( .A1(n19789), .A2(n19453), .B1(n19912), .B2(n19788), .ZN(
        n19782) );
  AOI22_X1 U22773 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19790), .B1(
        n19783), .B2(n19913), .ZN(n19781) );
  OAI211_X1 U22774 ( .C1(n19916), .C2(n19832), .A(n19782), .B(n19781), .ZN(
        P2_U3140) );
  AOI22_X1 U22775 ( .A1(n19789), .A2(n13305), .B1(n13312), .B2(n19788), .ZN(
        n19785) );
  AOI22_X1 U22776 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19790), .B1(
        n19783), .B2(n19917), .ZN(n19784) );
  OAI211_X1 U22777 ( .C1(n19920), .C2(n19832), .A(n19785), .B(n19784), .ZN(
        P2_U3141) );
  AOI22_X1 U22778 ( .A1(n19789), .A2(n13101), .B1(n19921), .B2(n19788), .ZN(
        n19787) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19790), .B1(
        n19800), .B2(n19870), .ZN(n19786) );
  OAI211_X1 U22780 ( .C1(n19826), .C2(n19793), .A(n19787), .B(n19786), .ZN(
        P2_U3142) );
  AOI22_X1 U22781 ( .A1(n19789), .A2(n19464), .B1(n19926), .B2(n19788), .ZN(
        n19792) );
  AOI22_X1 U22782 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19790), .B1(
        n19800), .B2(n19875), .ZN(n19791) );
  OAI211_X1 U22783 ( .C1(n19833), .C2(n19793), .A(n19792), .B(n19791), .ZN(
        P2_U3143) );
  NAND2_X1 U22784 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19794), .ZN(
        n19802) );
  OR2_X1 U22785 ( .A1(n19802), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19799) );
  INV_X1 U22786 ( .A(n19795), .ZN(n19798) );
  INV_X1 U22787 ( .A(n19796), .ZN(n19797) );
  NOR2_X1 U22788 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19797), .ZN(
        n19827) );
  NOR3_X1 U22789 ( .A1(n19798), .A2(n19827), .A3(n20067), .ZN(n19801) );
  AOI21_X1 U22790 ( .B1(n20067), .B2(n19799), .A(n19801), .ZN(n19828) );
  AOI22_X1 U22791 ( .A1(n19828), .A2(n13117), .B1(n19885), .B2(n19827), .ZN(
        n19807) );
  OAI21_X1 U22792 ( .B1(n19800), .B2(n19848), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19803) );
  AOI211_X1 U22793 ( .C1(n19803), .C2(n19802), .A(n19888), .B(n19801), .ZN(
        n19804) );
  AOI22_X1 U22794 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19829), .B1(
        n19848), .B2(n19805), .ZN(n19806) );
  OAI211_X1 U22795 ( .C1(n19808), .C2(n19832), .A(n19807), .B(n19806), .ZN(
        P2_U3144) );
  AOI22_X1 U22796 ( .A1(n19828), .A2(n13681), .B1(n13683), .B2(n19827), .ZN(
        n19810) );
  AOI22_X1 U22797 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19829), .B1(
        n19848), .B2(n19853), .ZN(n19809) );
  OAI211_X1 U22798 ( .C1(n19811), .C2(n19832), .A(n19810), .B(n19809), .ZN(
        P2_U3145) );
  AOI22_X1 U22799 ( .A1(n19828), .A2(n19441), .B1(n19902), .B2(n19827), .ZN(
        n19813) );
  AOI22_X1 U22800 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19829), .B1(
        n19848), .B2(n19856), .ZN(n19812) );
  OAI211_X1 U22801 ( .C1(n19814), .C2(n19832), .A(n19813), .B(n19812), .ZN(
        P2_U3146) );
  AOI22_X1 U22802 ( .A1(n19828), .A2(n19447), .B1(n19907), .B2(n19827), .ZN(
        n19816) );
  AOI22_X1 U22803 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19829), .B1(
        n19848), .B2(n19860), .ZN(n19815) );
  OAI211_X1 U22804 ( .C1(n19817), .C2(n19832), .A(n19816), .B(n19815), .ZN(
        P2_U3147) );
  AOI22_X1 U22805 ( .A1(n19828), .A2(n19453), .B1(n19912), .B2(n19827), .ZN(
        n19819) );
  AOI22_X1 U22806 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19829), .B1(
        n19848), .B2(n19863), .ZN(n19818) );
  OAI211_X1 U22807 ( .C1(n19820), .C2(n19832), .A(n19819), .B(n19818), .ZN(
        P2_U3148) );
  AOI22_X1 U22808 ( .A1(n19828), .A2(n13305), .B1(n13312), .B2(n19827), .ZN(
        n19822) );
  AOI22_X1 U22809 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19829), .B1(
        n19848), .B2(n19867), .ZN(n19821) );
  OAI211_X1 U22810 ( .C1(n19823), .C2(n19832), .A(n19822), .B(n19821), .ZN(
        P2_U3149) );
  AOI22_X1 U22811 ( .A1(n19828), .A2(n13101), .B1(n19921), .B2(n19827), .ZN(
        n19825) );
  AOI22_X1 U22812 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19829), .B1(
        n19848), .B2(n19870), .ZN(n19824) );
  OAI211_X1 U22813 ( .C1(n19826), .C2(n19832), .A(n19825), .B(n19824), .ZN(
        P2_U3150) );
  AOI22_X1 U22814 ( .A1(n19828), .A2(n19464), .B1(n19926), .B2(n19827), .ZN(
        n19831) );
  AOI22_X1 U22815 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19829), .B1(
        n19848), .B2(n19875), .ZN(n19830) );
  OAI211_X1 U22816 ( .C1(n19833), .C2(n19832), .A(n19831), .B(n19830), .ZN(
        P2_U3151) );
  AOI22_X1 U22817 ( .A1(n19847), .A2(n13681), .B1(n19846), .B2(n13683), .ZN(
        n19835) );
  AOI22_X1 U22818 ( .A1(n19874), .A2(n19853), .B1(n19848), .B2(n19898), .ZN(
        n19834) );
  OAI211_X1 U22819 ( .C1(n19852), .C2(n11908), .A(n19835), .B(n19834), .ZN(
        P2_U3153) );
  AOI22_X1 U22820 ( .A1(n19847), .A2(n19441), .B1(n19846), .B2(n19902), .ZN(
        n19837) );
  AOI22_X1 U22821 ( .A1(n19874), .A2(n19856), .B1(n19848), .B2(n19903), .ZN(
        n19836) );
  OAI211_X1 U22822 ( .C1(n19852), .C2(n11937), .A(n19837), .B(n19836), .ZN(
        P2_U3154) );
  AOI22_X1 U22823 ( .A1(n19847), .A2(n19447), .B1(n19846), .B2(n19907), .ZN(
        n19839) );
  AOI22_X1 U22824 ( .A1(n19874), .A2(n19860), .B1(n19848), .B2(n19908), .ZN(
        n19838) );
  OAI211_X1 U22825 ( .C1(n19852), .C2(n11965), .A(n19839), .B(n19838), .ZN(
        P2_U3155) );
  AOI22_X1 U22826 ( .A1(n19847), .A2(n19453), .B1(n19846), .B2(n19912), .ZN(
        n19841) );
  AOI22_X1 U22827 ( .A1(n19874), .A2(n19863), .B1(n19848), .B2(n19913), .ZN(
        n19840) );
  OAI211_X1 U22828 ( .C1(n19852), .C2(n11991), .A(n19841), .B(n19840), .ZN(
        P2_U3156) );
  AOI22_X1 U22829 ( .A1(n19847), .A2(n13305), .B1(n19846), .B2(n13312), .ZN(
        n19843) );
  AOI22_X1 U22830 ( .A1(n19848), .A2(n19917), .B1(n19874), .B2(n19867), .ZN(
        n19842) );
  OAI211_X1 U22831 ( .C1(n19852), .C2(n12015), .A(n19843), .B(n19842), .ZN(
        P2_U3157) );
  AOI22_X1 U22832 ( .A1(n19847), .A2(n13101), .B1(n19846), .B2(n19921), .ZN(
        n19845) );
  AOI22_X1 U22833 ( .A1(n19848), .A2(n19922), .B1(n19874), .B2(n19870), .ZN(
        n19844) );
  OAI211_X1 U22834 ( .C1(n19852), .C2(n12038), .A(n19845), .B(n19844), .ZN(
        P2_U3158) );
  INV_X1 U22835 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n19851) );
  AOI22_X1 U22836 ( .A1(n19847), .A2(n19464), .B1(n19846), .B2(n19926), .ZN(
        n19850) );
  AOI22_X1 U22837 ( .A1(n19874), .A2(n19875), .B1(n19848), .B2(n19929), .ZN(
        n19849) );
  OAI211_X1 U22838 ( .C1(n19852), .C2(n19851), .A(n19850), .B(n19849), .ZN(
        P2_U3159) );
  AOI22_X1 U22839 ( .A1(n19930), .A2(n19853), .B1(n19873), .B2(n13683), .ZN(
        n19855) );
  AOI22_X1 U22840 ( .A1(n13681), .A2(n19876), .B1(n19874), .B2(n19898), .ZN(
        n19854) );
  OAI211_X1 U22841 ( .C1(n19880), .C2(n10686), .A(n19855), .B(n19854), .ZN(
        P2_U3161) );
  INV_X1 U22842 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19859) );
  AOI22_X1 U22843 ( .A1(n19930), .A2(n19856), .B1(n19873), .B2(n19902), .ZN(
        n19858) );
  AOI22_X1 U22844 ( .A1(n19441), .A2(n19876), .B1(n19874), .B2(n19903), .ZN(
        n19857) );
  OAI211_X1 U22845 ( .C1(n19880), .C2(n19859), .A(n19858), .B(n19857), .ZN(
        P2_U3162) );
  AOI22_X1 U22846 ( .A1(n19874), .A2(n19908), .B1(n19873), .B2(n19907), .ZN(
        n19862) );
  AOI22_X1 U22847 ( .A1(n19447), .A2(n19876), .B1(n19930), .B2(n19860), .ZN(
        n19861) );
  OAI211_X1 U22848 ( .C1(n19880), .C2(n10645), .A(n19862), .B(n19861), .ZN(
        P2_U3163) );
  AOI22_X1 U22849 ( .A1(n19874), .A2(n19913), .B1(n19873), .B2(n19912), .ZN(
        n19865) );
  AOI22_X1 U22850 ( .A1(n19453), .A2(n19876), .B1(n19930), .B2(n19863), .ZN(
        n19864) );
  OAI211_X1 U22851 ( .C1(n19880), .C2(n19866), .A(n19865), .B(n19864), .ZN(
        P2_U3164) );
  AOI22_X1 U22852 ( .A1(n19874), .A2(n19917), .B1(n19873), .B2(n13312), .ZN(
        n19869) );
  AOI22_X1 U22853 ( .A1(n13305), .A2(n19876), .B1(n19930), .B2(n19867), .ZN(
        n19868) );
  OAI211_X1 U22854 ( .C1(n19880), .C2(n10754), .A(n19869), .B(n19868), .ZN(
        P2_U3165) );
  AOI22_X1 U22855 ( .A1(n19874), .A2(n19922), .B1(n19921), .B2(n19873), .ZN(
        n19872) );
  AOI22_X1 U22856 ( .A1(n13101), .A2(n19876), .B1(n19930), .B2(n19870), .ZN(
        n19871) );
  OAI211_X1 U22857 ( .C1(n19880), .C2(n10851), .A(n19872), .B(n19871), .ZN(
        P2_U3166) );
  AOI22_X1 U22858 ( .A1(n19874), .A2(n19929), .B1(n19873), .B2(n19926), .ZN(
        n19878) );
  AOI22_X1 U22859 ( .A1(n19464), .A2(n19876), .B1(n19930), .B2(n19875), .ZN(
        n19877) );
  OAI211_X1 U22860 ( .C1(n19880), .C2(n19879), .A(n19878), .B(n19877), .ZN(
        P2_U3167) );
  NAND3_X1 U22861 ( .A1(n19881), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19889), 
        .ZN(n19886) );
  NOR2_X1 U22862 ( .A1(n20048), .A2(n19882), .ZN(n19893) );
  INV_X1 U22863 ( .A(n19893), .ZN(n19883) );
  OAI21_X1 U22864 ( .B1(n19883), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20067), 
        .ZN(n19884) );
  AND2_X1 U22865 ( .A1(n19886), .A2(n19884), .ZN(n19928) );
  INV_X1 U22866 ( .A(n19889), .ZN(n19927) );
  AOI22_X1 U22867 ( .A1(n19928), .A2(n13117), .B1(n19927), .B2(n19885), .ZN(
        n19896) );
  INV_X1 U22868 ( .A(n19886), .ZN(n19887) );
  AOI211_X1 U22869 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19889), .A(n19888), 
        .B(n19887), .ZN(n19890) );
  OAI221_X1 U22870 ( .B1(n19893), .B2(n19892), .C1(n19893), .C2(n19891), .A(
        n19890), .ZN(n19931) );
  AOI22_X1 U22871 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19931), .B1(
        n19930), .B2(n19894), .ZN(n19895) );
  OAI211_X1 U22872 ( .C1(n19897), .C2(n19934), .A(n19896), .B(n19895), .ZN(
        P2_U3168) );
  AOI22_X1 U22873 ( .A1(n19928), .A2(n13681), .B1(n19927), .B2(n13683), .ZN(
        n19900) );
  AOI22_X1 U22874 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19931), .B1(
        n19930), .B2(n19898), .ZN(n19899) );
  OAI211_X1 U22875 ( .C1(n19901), .C2(n19934), .A(n19900), .B(n19899), .ZN(
        P2_U3169) );
  AOI22_X1 U22876 ( .A1(n19928), .A2(n19441), .B1(n19927), .B2(n19902), .ZN(
        n19905) );
  AOI22_X1 U22877 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19931), .B1(
        n19930), .B2(n19903), .ZN(n19904) );
  OAI211_X1 U22878 ( .C1(n19906), .C2(n19934), .A(n19905), .B(n19904), .ZN(
        P2_U3170) );
  AOI22_X1 U22879 ( .A1(n19928), .A2(n19447), .B1(n19927), .B2(n19907), .ZN(
        n19910) );
  AOI22_X1 U22880 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19931), .B1(
        n19930), .B2(n19908), .ZN(n19909) );
  OAI211_X1 U22881 ( .C1(n19911), .C2(n19934), .A(n19910), .B(n19909), .ZN(
        P2_U3171) );
  AOI22_X1 U22882 ( .A1(n19928), .A2(n19453), .B1(n19927), .B2(n19912), .ZN(
        n19915) );
  AOI22_X1 U22883 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19931), .B1(
        n19930), .B2(n19913), .ZN(n19914) );
  OAI211_X1 U22884 ( .C1(n19916), .C2(n19934), .A(n19915), .B(n19914), .ZN(
        P2_U3172) );
  AOI22_X1 U22885 ( .A1(n19928), .A2(n13305), .B1(n19927), .B2(n13312), .ZN(
        n19919) );
  AOI22_X1 U22886 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19931), .B1(
        n19930), .B2(n19917), .ZN(n19918) );
  OAI211_X1 U22887 ( .C1(n19920), .C2(n19934), .A(n19919), .B(n19918), .ZN(
        P2_U3173) );
  AOI22_X1 U22888 ( .A1(n19928), .A2(n13101), .B1(n19927), .B2(n19921), .ZN(
        n19924) );
  AOI22_X1 U22889 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19931), .B1(
        n19930), .B2(n19922), .ZN(n19923) );
  OAI211_X1 U22890 ( .C1(n19925), .C2(n19934), .A(n19924), .B(n19923), .ZN(
        P2_U3174) );
  AOI22_X1 U22891 ( .A1(n19928), .A2(n19464), .B1(n19927), .B2(n19926), .ZN(
        n19933) );
  AOI22_X1 U22892 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19931), .B1(
        n19930), .B2(n19929), .ZN(n19932) );
  OAI211_X1 U22893 ( .C1(n19935), .C2(n19934), .A(n19933), .B(n19932), .ZN(
        P2_U3175) );
  INV_X1 U22894 ( .A(n20028), .ZN(n19936) );
  AND2_X1 U22895 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19936), .ZN(
        P2_U3179) );
  AND2_X1 U22896 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19936), .ZN(
        P2_U3180) );
  AND2_X1 U22897 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19936), .ZN(
        P2_U3181) );
  AND2_X1 U22898 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19936), .ZN(
        P2_U3182) );
  AND2_X1 U22899 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19936), .ZN(
        P2_U3183) );
  AND2_X1 U22900 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19936), .ZN(
        P2_U3184) );
  AND2_X1 U22901 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19936), .ZN(
        P2_U3185) );
  AND2_X1 U22902 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19936), .ZN(
        P2_U3186) );
  AND2_X1 U22903 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19936), .ZN(
        P2_U3187) );
  AND2_X1 U22904 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19936), .ZN(
        P2_U3188) );
  AND2_X1 U22905 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19936), .ZN(
        P2_U3189) );
  AND2_X1 U22906 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19936), .ZN(
        P2_U3190) );
  AND2_X1 U22907 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19936), .ZN(
        P2_U3191) );
  AND2_X1 U22908 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19936), .ZN(
        P2_U3192) );
  AND2_X1 U22909 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19936), .ZN(
        P2_U3193) );
  AND2_X1 U22910 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19936), .ZN(
        P2_U3194) );
  AND2_X1 U22911 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19936), .ZN(
        P2_U3195) );
  AND2_X1 U22912 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19936), .ZN(
        P2_U3196) );
  AND2_X1 U22913 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19936), .ZN(
        P2_U3197) );
  AND2_X1 U22914 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19936), .ZN(
        P2_U3198) );
  AND2_X1 U22915 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19936), .ZN(
        P2_U3199) );
  AND2_X1 U22916 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19936), .ZN(
        P2_U3200) );
  AND2_X1 U22917 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19936), .ZN(P2_U3201) );
  AND2_X1 U22918 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19936), .ZN(P2_U3202) );
  AND2_X1 U22919 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19936), .ZN(P2_U3203) );
  AND2_X1 U22920 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19936), .ZN(P2_U3204) );
  AND2_X1 U22921 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19936), .ZN(P2_U3205) );
  AND2_X1 U22922 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19936), .ZN(P2_U3206) );
  AND2_X1 U22923 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19936), .ZN(P2_U3207) );
  AND2_X1 U22924 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19936), .ZN(P2_U3208) );
  INV_X1 U22925 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19949) );
  NOR2_X1 U22926 ( .A1(n19937), .A2(n19949), .ZN(n19946) );
  OR3_X1 U22927 ( .A1(n19947), .A2(n19938), .A3(n19946), .ZN(n19939) );
  NOR3_X1 U22928 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21056), .ZN(n19954) );
  AOI21_X1 U22929 ( .B1(n19957), .B2(n19939), .A(n19954), .ZN(n19940) );
  OAI221_X1 U22930 ( .B1(n19941), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n19941), .C2(n20819), .A(n19940), .ZN(P2_U3209) );
  AOI21_X1 U22931 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20819), .A(n19957), 
        .ZN(n19950) );
  NOR3_X1 U22932 ( .A1(n19950), .A2(n19947), .A3(n19938), .ZN(n19942) );
  NOR2_X1 U22933 ( .A1(n19942), .A2(n19946), .ZN(n19944) );
  OAI211_X1 U22934 ( .C1(n20819), .C2(n19945), .A(n19944), .B(n19943), .ZN(
        P2_U3210) );
  AOI22_X1 U22935 ( .A1(n19948), .A2(n19947), .B1(n19946), .B2(n21056), .ZN(
        n19956) );
  OAI21_X1 U22936 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19955) );
  NOR2_X1 U22937 ( .A1(n19949), .A2(n19957), .ZN(n19952) );
  AOI21_X1 U22938 ( .B1(n19952), .B2(n19951), .A(n19950), .ZN(n19953) );
  OAI22_X1 U22939 ( .A1(n19956), .A2(n19955), .B1(n19954), .B2(n19953), .ZN(
        P2_U3211) );
  INV_X1 U22940 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19961) );
  OAI222_X1 U22941 ( .A1(n20021), .A2(n19961), .B1(n19959), .B2(n20015), .C1(
        n19958), .C2(n20017), .ZN(P2_U3212) );
  OAI222_X1 U22942 ( .A1(n20017), .A2(n19961), .B1(n19960), .B2(n20015), .C1(
        n19963), .C2(n20021), .ZN(P2_U3213) );
  OAI222_X1 U22943 ( .A1(n20017), .A2(n19963), .B1(n19962), .B2(n20015), .C1(
        n19964), .C2(n20021), .ZN(P2_U3214) );
  OAI222_X1 U22944 ( .A1(n20021), .A2(n19966), .B1(n19965), .B2(n20015), .C1(
        n19964), .C2(n20017), .ZN(P2_U3215) );
  OAI222_X1 U22945 ( .A1(n20021), .A2(n19968), .B1(n19967), .B2(n20015), .C1(
        n19966), .C2(n20017), .ZN(P2_U3216) );
  OAI222_X1 U22946 ( .A1(n20021), .A2(n19970), .B1(n19969), .B2(n20015), .C1(
        n19968), .C2(n20017), .ZN(P2_U3217) );
  OAI222_X1 U22947 ( .A1(n20021), .A2(n19972), .B1(n19971), .B2(n20015), .C1(
        n19970), .C2(n20017), .ZN(P2_U3218) );
  INV_X1 U22948 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19974) );
  OAI222_X1 U22949 ( .A1(n20021), .A2(n19974), .B1(n19973), .B2(n20015), .C1(
        n19972), .C2(n20017), .ZN(P2_U3219) );
  OAI222_X1 U22950 ( .A1(n20021), .A2(n19976), .B1(n19975), .B2(n20015), .C1(
        n19974), .C2(n20017), .ZN(P2_U3220) );
  INV_X1 U22951 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19978) );
  OAI222_X1 U22952 ( .A1(n20021), .A2(n19978), .B1(n19977), .B2(n20015), .C1(
        n19976), .C2(n20017), .ZN(P2_U3221) );
  OAI222_X1 U22953 ( .A1(n20021), .A2(n19980), .B1(n19979), .B2(n20015), .C1(
        n19978), .C2(n20017), .ZN(P2_U3222) );
  OAI222_X1 U22954 ( .A1(n20021), .A2(n19982), .B1(n19981), .B2(n20015), .C1(
        n19980), .C2(n20017), .ZN(P2_U3223) );
  OAI222_X1 U22955 ( .A1(n20021), .A2(n19984), .B1(n19983), .B2(n20015), .C1(
        n19982), .C2(n20017), .ZN(P2_U3224) );
  INV_X1 U22956 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19986) );
  OAI222_X1 U22957 ( .A1(n20021), .A2(n19986), .B1(n19985), .B2(n20015), .C1(
        n19984), .C2(n20017), .ZN(P2_U3225) );
  OAI222_X1 U22958 ( .A1(n20021), .A2(n19988), .B1(n19987), .B2(n20015), .C1(
        n19986), .C2(n20017), .ZN(P2_U3226) );
  OAI222_X1 U22959 ( .A1(n20021), .A2(n19990), .B1(n19989), .B2(n20015), .C1(
        n19988), .C2(n20017), .ZN(P2_U3227) );
  OAI222_X1 U22960 ( .A1(n20021), .A2(n19992), .B1(n19991), .B2(n20015), .C1(
        n19990), .C2(n20017), .ZN(P2_U3228) );
  INV_X1 U22961 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19994) );
  OAI222_X1 U22962 ( .A1(n20021), .A2(n19994), .B1(n19993), .B2(n20015), .C1(
        n19992), .C2(n20017), .ZN(P2_U3229) );
  OAI222_X1 U22963 ( .A1(n20021), .A2(n19996), .B1(n19995), .B2(n20015), .C1(
        n19994), .C2(n20017), .ZN(P2_U3230) );
  OAI222_X1 U22964 ( .A1(n20021), .A2(n19998), .B1(n19997), .B2(n20015), .C1(
        n19996), .C2(n20017), .ZN(P2_U3231) );
  OAI222_X1 U22965 ( .A1(n20021), .A2(n20000), .B1(n19999), .B2(n20015), .C1(
        n19998), .C2(n20017), .ZN(P2_U3232) );
  INV_X1 U22966 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20002) );
  OAI222_X1 U22967 ( .A1(n20021), .A2(n20002), .B1(n20001), .B2(n20015), .C1(
        n20000), .C2(n20017), .ZN(P2_U3233) );
  OAI222_X1 U22968 ( .A1(n20021), .A2(n20004), .B1(n20003), .B2(n20015), .C1(
        n20002), .C2(n20017), .ZN(P2_U3234) );
  INV_X1 U22969 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20006) );
  OAI222_X1 U22970 ( .A1(n20021), .A2(n20006), .B1(n20005), .B2(n20015), .C1(
        n20004), .C2(n20017), .ZN(P2_U3235) );
  OAI222_X1 U22971 ( .A1(n20021), .A2(n20008), .B1(n20007), .B2(n20015), .C1(
        n20006), .C2(n20017), .ZN(P2_U3236) );
  OAI222_X1 U22972 ( .A1(n20021), .A2(n20011), .B1(n20009), .B2(n20015), .C1(
        n20008), .C2(n20017), .ZN(P2_U3237) );
  INV_X1 U22973 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20012) );
  OAI222_X1 U22974 ( .A1(n20017), .A2(n20011), .B1(n20010), .B2(n20015), .C1(
        n20012), .C2(n20021), .ZN(P2_U3238) );
  OAI222_X1 U22975 ( .A1(n20021), .A2(n20014), .B1(n20013), .B2(n20015), .C1(
        n20012), .C2(n20017), .ZN(P2_U3239) );
  OAI222_X1 U22976 ( .A1(n20021), .A2(n20018), .B1(n20016), .B2(n20015), .C1(
        n20014), .C2(n20017), .ZN(P2_U3240) );
  INV_X1 U22977 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20019) );
  OAI222_X1 U22978 ( .A1(n20021), .A2(n20020), .B1(n20019), .B2(n20015), .C1(
        n20018), .C2(n20017), .ZN(P2_U3241) );
  OAI22_X1 U22979 ( .A1(n20086), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20015), .ZN(n20022) );
  INV_X1 U22980 ( .A(n20022), .ZN(P2_U3585) );
  MUX2_X1 U22981 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20086), .Z(P2_U3586) );
  OAI22_X1 U22982 ( .A1(n20086), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20015), .ZN(n20023) );
  INV_X1 U22983 ( .A(n20023), .ZN(P2_U3587) );
  OAI22_X1 U22984 ( .A1(n20086), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20015), .ZN(n20024) );
  INV_X1 U22985 ( .A(n20024), .ZN(P2_U3588) );
  OAI21_X1 U22986 ( .B1(n20028), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20026), 
        .ZN(n20025) );
  INV_X1 U22987 ( .A(n20025), .ZN(P2_U3591) );
  OAI21_X1 U22988 ( .B1(n20028), .B2(n20027), .A(n20026), .ZN(P2_U3592) );
  OAI22_X1 U22989 ( .A1(n20039), .A2(n20031), .B1(n20030), .B2(n20029), .ZN(
        n20033) );
  MUX2_X1 U22990 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20033), .S(
        n20032), .Z(P2_U3596) );
  NAND2_X1 U22991 ( .A1(n20037), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20059) );
  NOR2_X1 U22992 ( .A1(n20034), .A2(n20059), .ZN(n20053) );
  INV_X1 U22993 ( .A(n20053), .ZN(n20040) );
  AOI211_X1 U22994 ( .C1(n20038), .C2(n20037), .A(n20036), .B(n20035), .ZN(
        n20049) );
  AOI21_X1 U22995 ( .B1(n20040), .B2(n20049), .A(n20039), .ZN(n20045) );
  NOR3_X1 U22996 ( .A1(n20043), .A2(n20042), .A3(n20041), .ZN(n20044) );
  AOI211_X1 U22997 ( .C1(n20046), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20045), 
        .B(n20044), .ZN(n20047) );
  AOI22_X1 U22998 ( .A1(n20072), .A2(n20048), .B1(n20047), .B2(n20073), .ZN(
        P2_U3602) );
  INV_X1 U22999 ( .A(n20049), .ZN(n20052) );
  AOI22_X1 U23000 ( .A1(n20052), .A2(n20051), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20050), .ZN(n20055) );
  NOR2_X1 U23001 ( .A1(n20072), .A2(n20053), .ZN(n20054) );
  AOI22_X1 U23002 ( .A1(n20056), .A2(n20072), .B1(n20055), .B2(n20054), .ZN(
        P2_U3603) );
  NAND3_X1 U23003 ( .A1(n20060), .A2(n20065), .A3(n20057), .ZN(n20058) );
  OAI21_X1 U23004 ( .B1(n20060), .B2(n20059), .A(n20058), .ZN(n20061) );
  AOI21_X1 U23005 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20062), .A(n20061), 
        .ZN(n20063) );
  AOI22_X1 U23006 ( .A1(n20072), .A2(n20064), .B1(n20063), .B2(n20073), .ZN(
        P2_U3604) );
  INV_X1 U23007 ( .A(n20065), .ZN(n20068) );
  OAI22_X1 U23008 ( .A1(n20069), .A2(n20068), .B1(n20067), .B2(n20066), .ZN(
        n20070) );
  AOI21_X1 U23009 ( .B1(n20074), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20070), 
        .ZN(n20071) );
  OAI22_X1 U23010 ( .A1(n20074), .A2(n20073), .B1(n20072), .B2(n20071), .ZN(
        P2_U3605) );
  INV_X1 U23011 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20075) );
  AOI22_X1 U23012 ( .A1(n20015), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20075), 
        .B2(n20086), .ZN(P2_U3608) );
  NAND2_X1 U23013 ( .A1(n20077), .A2(n20076), .ZN(n20078) );
  AOI22_X1 U23014 ( .A1(n20081), .A2(n20080), .B1(n20079), .B2(n20078), .ZN(
        n20082) );
  NAND2_X1 U23015 ( .A1(n20083), .A2(n20082), .ZN(n20085) );
  MUX2_X1 U23016 ( .A(P2_MORE_REG_SCAN_IN), .B(n20085), .S(n20084), .Z(
        P2_U3609) );
  OAI22_X1 U23017 ( .A1(n20086), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20015), .ZN(n20087) );
  INV_X1 U23018 ( .A(n20087), .ZN(P2_U3611) );
  INV_X1 U23019 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20809) );
  AOI21_X1 U23020 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20820), .A(n20809), 
        .ZN(n20810) );
  INV_X1 U23021 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21130) );
  AOI21_X1 U23022 ( .B1(n20810), .B2(n21130), .A(n20912), .ZN(P1_U2802) );
  INV_X1 U23023 ( .A(n20088), .ZN(n20090) );
  OAI21_X1 U23024 ( .B1(n20090), .B2(n20089), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20091) );
  OAI21_X1 U23025 ( .B1(n20092), .B2(n20237), .A(n20091), .ZN(P1_U2803) );
  INV_X2 U23026 ( .A(n20912), .ZN(n20911) );
  NOR2_X1 U23027 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20094) );
  OAI21_X1 U23028 ( .B1(n20094), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20911), .ZN(
        n20093) );
  OAI21_X1 U23029 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20911), .A(n20093), 
        .ZN(P1_U2804) );
  NOR2_X1 U23030 ( .A1(n20810), .A2(n20912), .ZN(n20863) );
  OAI21_X1 U23031 ( .B1(BS16), .B2(n20094), .A(n20863), .ZN(n20861) );
  OAI21_X1 U23032 ( .B1(n20863), .B2(n20703), .A(n20861), .ZN(P1_U2805) );
  OAI21_X1 U23033 ( .B1(n20096), .B2(n21158), .A(n20095), .ZN(P1_U2806) );
  NOR4_X1 U23034 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20100) );
  NOR4_X1 U23035 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20099) );
  NOR4_X1 U23036 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20098) );
  NOR4_X1 U23037 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20097) );
  NAND4_X1 U23038 ( .A1(n20100), .A2(n20099), .A3(n20098), .A4(n20097), .ZN(
        n20106) );
  NOR4_X1 U23039 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20104) );
  AOI211_X1 U23040 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20103) );
  NOR4_X1 U23041 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20102) );
  NOR4_X1 U23042 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20101) );
  NAND4_X1 U23043 ( .A1(n20104), .A2(n20103), .A3(n20102), .A4(n20101), .ZN(
        n20105) );
  NOR2_X1 U23044 ( .A1(n20106), .A2(n20105), .ZN(n20896) );
  INV_X1 U23045 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21199) );
  NOR3_X1 U23046 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20108) );
  OAI21_X1 U23047 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20108), .A(n20896), .ZN(
        n20107) );
  OAI21_X1 U23048 ( .B1(n20896), .B2(n21199), .A(n20107), .ZN(P1_U2807) );
  INV_X1 U23049 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20862) );
  AOI21_X1 U23050 ( .B1(n21013), .B2(n20862), .A(n20108), .ZN(n20109) );
  INV_X1 U23051 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21190) );
  INV_X1 U23052 ( .A(n20896), .ZN(n20898) );
  AOI22_X1 U23053 ( .A1(n20896), .A2(n20109), .B1(n21190), .B2(n20898), .ZN(
        P1_U2808) );
  AOI21_X1 U23054 ( .B1(n20110), .B2(P1_EBX_REG_9__SCAN_IN), .A(n20138), .ZN(
        n20111) );
  OAI21_X1 U23055 ( .B1(n20112), .B2(n20136), .A(n20111), .ZN(n20114) );
  NOR2_X1 U23056 ( .A1(n20170), .A2(n20162), .ZN(n20113) );
  AOI211_X1 U23057 ( .C1(n20115), .C2(n20158), .A(n20114), .B(n20113), .ZN(
        n20119) );
  INV_X1 U23058 ( .A(n20172), .ZN(n20117) );
  AOI22_X1 U23059 ( .A1(n20117), .A2(n20128), .B1(n20121), .B2(n20116), .ZN(
        n20118) );
  OAI211_X1 U23060 ( .C1(n20121), .C2(n20120), .A(n20119), .B(n20118), .ZN(
        P1_U2831) );
  NAND2_X1 U23061 ( .A1(n20110), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n20122) );
  AND2_X1 U23062 ( .A1(n20154), .A2(n20122), .ZN(n20124) );
  NAND2_X1 U23063 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n20123) );
  OAI211_X1 U23064 ( .C1(n20140), .C2(n20125), .A(n20124), .B(n20123), .ZN(
        n20126) );
  AOI21_X1 U23065 ( .B1(n20176), .B2(n20144), .A(n20126), .ZN(n20130) );
  AOI22_X1 U23066 ( .A1(n20177), .A2(n20128), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n20127), .ZN(n20129) );
  OAI211_X1 U23067 ( .C1(P1_REIP_REG_7__SCAN_IN), .C2(n20131), .A(n20130), .B(
        n20129), .ZN(P1_U2833) );
  NAND2_X1 U23068 ( .A1(n9798), .A2(n20132), .ZN(n20168) );
  INV_X1 U23069 ( .A(n20134), .ZN(n20148) );
  NOR2_X1 U23070 ( .A1(n20136), .A2(n20135), .ZN(n20137) );
  AOI211_X1 U23071 ( .C1(n20110), .C2(P1_EBX_REG_5__SCAN_IN), .A(n20138), .B(
        n20137), .ZN(n20139) );
  OAI21_X1 U23072 ( .B1(n20141), .B2(n20140), .A(n20139), .ZN(n20142) );
  AOI21_X1 U23073 ( .B1(n20144), .B2(n20143), .A(n20142), .ZN(n20145) );
  OAI21_X1 U23074 ( .B1(n20146), .B2(P1_REIP_REG_5__SCAN_IN), .A(n20145), .ZN(
        n20147) );
  AOI21_X1 U23075 ( .B1(n20148), .B2(n20165), .A(n20147), .ZN(n20149) );
  OAI21_X1 U23076 ( .B1(n21162), .B2(n20168), .A(n20149), .ZN(P1_U2835) );
  AOI21_X1 U23077 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n20150), .A(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20169) );
  NAND2_X1 U23078 ( .A1(n20152), .A2(n20151), .ZN(n20161) );
  NAND2_X1 U23079 ( .A1(n20153), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20155) );
  OAI211_X1 U23080 ( .C1(n21221), .C2(n20156), .A(n20155), .B(n20154), .ZN(
        n20157) );
  AOI21_X1 U23081 ( .B1(n20159), .B2(n20158), .A(n20157), .ZN(n20160) );
  OAI211_X1 U23082 ( .C1(n20163), .C2(n20162), .A(n20161), .B(n20160), .ZN(
        n20164) );
  AOI21_X1 U23083 ( .B1(n20166), .B2(n20165), .A(n20164), .ZN(n20167) );
  OAI21_X1 U23084 ( .B1(n20169), .B2(n20168), .A(n20167), .ZN(P1_U2836) );
  OAI22_X1 U23085 ( .A1(n20172), .A2(n14803), .B1(n20171), .B2(n20170), .ZN(
        n20173) );
  INV_X1 U23086 ( .A(n20173), .ZN(n20174) );
  OAI21_X1 U23087 ( .B1(n20185), .B2(n20175), .A(n20174), .ZN(P1_U2863) );
  AOI22_X1 U23088 ( .A1(n20177), .A2(n20182), .B1(n20181), .B2(n20176), .ZN(
        n20178) );
  OAI21_X1 U23089 ( .B1(n20185), .B2(n21034), .A(n20178), .ZN(P1_U2865) );
  INV_X1 U23090 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n20995) );
  INV_X1 U23091 ( .A(n20179), .ZN(n20183) );
  AOI22_X1 U23092 ( .A1(n20183), .A2(n20182), .B1(n20181), .B2(n20180), .ZN(
        n20184) );
  OAI21_X1 U23093 ( .B1(n20185), .B2(n20995), .A(n20184), .ZN(P1_U2869) );
  AOI22_X1 U23094 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20189), .B1(n15982), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20186) );
  OAI21_X1 U23095 ( .B1(n20188), .B2(n20187), .A(n20186), .ZN(P1_U2921) );
  INV_X1 U23096 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20191) );
  AOI22_X1 U23097 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20190) );
  OAI21_X1 U23098 ( .B1(n20191), .B2(n20212), .A(n20190), .ZN(P1_U2922) );
  AOI22_X1 U23099 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20192) );
  OAI21_X1 U23100 ( .B1(n14880), .B2(n20212), .A(n20192), .ZN(P1_U2923) );
  INV_X1 U23101 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20194) );
  AOI22_X1 U23102 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20193) );
  OAI21_X1 U23103 ( .B1(n20194), .B2(n20212), .A(n20193), .ZN(P1_U2924) );
  AOI22_X1 U23104 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20195) );
  OAI21_X1 U23105 ( .B1(n13949), .B2(n20212), .A(n20195), .ZN(P1_U2925) );
  AOI22_X1 U23106 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20196) );
  OAI21_X1 U23107 ( .B1(n13900), .B2(n20212), .A(n20196), .ZN(P1_U2926) );
  AOI22_X1 U23108 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20197) );
  OAI21_X1 U23109 ( .B1(n13824), .B2(n20212), .A(n20197), .ZN(P1_U2927) );
  AOI22_X1 U23110 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20198) );
  OAI21_X1 U23111 ( .B1(n20199), .B2(n20212), .A(n20198), .ZN(P1_U2928) );
  AOI22_X1 U23112 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20200) );
  OAI21_X1 U23113 ( .B1(n13590), .B2(n20212), .A(n20200), .ZN(P1_U2929) );
  AOI22_X1 U23114 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20201) );
  OAI21_X1 U23115 ( .B1(n13538), .B2(n20212), .A(n20201), .ZN(P1_U2930) );
  AOI22_X1 U23116 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20202) );
  OAI21_X1 U23117 ( .B1(n13448), .B2(n20212), .A(n20202), .ZN(P1_U2931) );
  AOI22_X1 U23118 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20203) );
  OAI21_X1 U23119 ( .B1(n20204), .B2(n20212), .A(n20203), .ZN(P1_U2932) );
  AOI22_X1 U23120 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20205) );
  OAI21_X1 U23121 ( .B1(n13499), .B2(n20212), .A(n20205), .ZN(P1_U2933) );
  AOI22_X1 U23122 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20206) );
  OAI21_X1 U23123 ( .B1(n20207), .B2(n20212), .A(n20206), .ZN(P1_U2934) );
  AOI22_X1 U23124 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20208) );
  OAI21_X1 U23125 ( .B1(n20209), .B2(n20212), .A(n20208), .ZN(P1_U2935) );
  AOI22_X1 U23126 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20210), .B1(n15982), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20211) );
  OAI21_X1 U23127 ( .B1(n20213), .B2(n20212), .A(n20211), .ZN(P1_U2936) );
  AOI22_X1 U23128 ( .A1(n20225), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20224), .ZN(n20215) );
  NAND2_X1 U23129 ( .A1(n20215), .A2(n20214), .ZN(P1_U2961) );
  AOI22_X1 U23130 ( .A1(n20225), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20224), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20217) );
  NAND2_X1 U23131 ( .A1(n20217), .A2(n20216), .ZN(P1_U2962) );
  AOI22_X1 U23132 ( .A1(n20225), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20224), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20219) );
  NAND2_X1 U23133 ( .A1(n20219), .A2(n20218), .ZN(P1_U2963) );
  AOI22_X1 U23134 ( .A1(n20225), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20224), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20221) );
  NAND2_X1 U23135 ( .A1(n20221), .A2(n20220), .ZN(P1_U2964) );
  AOI22_X1 U23136 ( .A1(n20225), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20224), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20223) );
  NAND2_X1 U23137 ( .A1(n20223), .A2(n20222), .ZN(P1_U2965) );
  AOI22_X1 U23138 ( .A1(n20225), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20224), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20227) );
  NAND2_X1 U23139 ( .A1(n20227), .A2(n20226), .ZN(P1_U2966) );
  NOR2_X1 U23140 ( .A1(n20228), .A2(n20892), .ZN(P1_U3032) );
  INV_X1 U23141 ( .A(DATAI_16_), .ZN(n21145) );
  OAI22_X1 U23142 ( .A1(n21145), .A2(n20291), .B1(n20231), .B2(n20292), .ZN(
        n20753) );
  INV_X1 U23143 ( .A(n20753), .ZN(n20714) );
  INV_X1 U23144 ( .A(n13069), .ZN(n20232) );
  NAND2_X1 U23145 ( .A1(n13069), .A2(n20233), .ZN(n20698) );
  INV_X1 U23146 ( .A(DATAI_24_), .ZN(n21172) );
  OAI22_X1 U23147 ( .A1(n20235), .A2(n20292), .B1(n21172), .B2(n20291), .ZN(
        n20711) );
  NAND3_X1 U23148 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20237), .A3(n20236), 
        .ZN(n20295) );
  NAND2_X1 U23149 ( .A1(n20286), .A2(n20238), .ZN(n20553) );
  NOR3_X1 U23150 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20306) );
  NAND2_X1 U23151 ( .A1(n20670), .A2(n20306), .ZN(n20267) );
  INV_X1 U23152 ( .A(n20267), .ZN(n20296) );
  AOI22_X1 U23153 ( .A1(n20797), .A2(n9941), .B1(n20744), .B2(n20296), .ZN(
        n20251) );
  INV_X1 U23154 ( .A(n20327), .ZN(n20239) );
  OAI21_X1 U23155 ( .B1(n20239), .B2(n20797), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20240) );
  NAND2_X1 U23156 ( .A1(n20240), .A2(n20625), .ZN(n20249) );
  NOR2_X1 U23157 ( .A1(n20359), .A2(n20705), .ZN(n20245) );
  NOR2_X1 U23158 ( .A1(n20246), .A2(n12749), .ZN(n20630) );
  INV_X1 U23159 ( .A(n20497), .ZN(n20242) );
  NAND2_X1 U23160 ( .A1(n20242), .A2(n20699), .ZN(n20392) );
  AOI22_X1 U23161 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20392), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20267), .ZN(n20243) );
  OAI211_X1 U23162 ( .C1(n20249), .C2(n20245), .A(n20559), .B(n20243), .ZN(
        n20299) );
  INV_X1 U23163 ( .A(n20245), .ZN(n20248) );
  INV_X1 U23164 ( .A(n20246), .ZN(n20247) );
  NOR2_X1 U23165 ( .A1(n20247), .A2(n12749), .ZN(n20552) );
  INV_X1 U23166 ( .A(n20552), .ZN(n20498) );
  OAI22_X1 U23167 ( .A1(n20249), .A2(n20248), .B1(n20498), .B2(n20392), .ZN(
        n20298) );
  AOI22_X1 U23168 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20299), .B1(
        n20743), .B2(n20298), .ZN(n20250) );
  OAI211_X1 U23169 ( .C1(n20714), .C2(n20327), .A(n20251), .B(n20250), .ZN(
        P1_U3033) );
  INV_X1 U23170 ( .A(DATAI_17_), .ZN(n21212) );
  OAI22_X1 U23171 ( .A1(n21212), .A2(n20291), .B1(n20252), .B2(n20292), .ZN(
        n20641) );
  INV_X1 U23172 ( .A(n20641), .ZN(n20761) );
  INV_X1 U23173 ( .A(DATAI_25_), .ZN(n21061) );
  OAI22_X2 U23174 ( .A1(n20253), .A2(n20292), .B1(n21061), .B2(n20291), .ZN(
        n20758) );
  NAND2_X1 U23175 ( .A1(n20286), .A2(n20254), .ZN(n20562) );
  AOI22_X1 U23176 ( .A1(n20797), .A2(n20758), .B1(n20757), .B2(n20296), .ZN(
        n20257) );
  AOI22_X1 U23177 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20299), .B1(
        n20756), .B2(n20298), .ZN(n20256) );
  OAI211_X1 U23178 ( .C1(n20761), .C2(n20327), .A(n20257), .B(n20256), .ZN(
        P1_U3034) );
  INV_X1 U23179 ( .A(DATAI_18_), .ZN(n21193) );
  OAI22_X1 U23180 ( .A1(n20258), .A2(n20292), .B1(n21193), .B2(n20291), .ZN(
        n20764) );
  INV_X1 U23181 ( .A(n20764), .ZN(n20720) );
  INV_X1 U23182 ( .A(DATAI_26_), .ZN(n21124) );
  INV_X1 U23183 ( .A(n20717), .ZN(n20767) );
  NAND2_X1 U23184 ( .A1(n20286), .A2(n20260), .ZN(n20566) );
  OAI22_X1 U23185 ( .A1(n20790), .A2(n20767), .B1(n20566), .B2(n20267), .ZN(
        n20261) );
  INV_X1 U23186 ( .A(n20261), .ZN(n20264) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20299), .B1(
        n20762), .B2(n20298), .ZN(n20263) );
  OAI211_X1 U23188 ( .C1(n20720), .C2(n20327), .A(n20264), .B(n20263), .ZN(
        P1_U3035) );
  INV_X1 U23189 ( .A(DATAI_19_), .ZN(n21214) );
  OAI22_X1 U23190 ( .A1(n20265), .A2(n20292), .B1(n21214), .B2(n20291), .ZN(
        n20648) );
  INV_X1 U23191 ( .A(n20648), .ZN(n20773) );
  INV_X1 U23192 ( .A(DATAI_27_), .ZN(n21146) );
  OAI22_X1 U23193 ( .A1(n20266), .A2(n20292), .B1(n21146), .B2(n20291), .ZN(
        n20770) );
  OAI22_X1 U23194 ( .A1(n20790), .A2(n9942), .B1(n20570), .B2(n20267), .ZN(
        n20268) );
  INV_X1 U23195 ( .A(n20268), .ZN(n20271) );
  AOI22_X1 U23196 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20299), .B1(
        n20768), .B2(n20298), .ZN(n20270) );
  OAI211_X1 U23197 ( .C1(n20773), .C2(n20327), .A(n20271), .B(n20270), .ZN(
        P1_U3036) );
  INV_X1 U23198 ( .A(DATAI_20_), .ZN(n20272) );
  OAI22_X1 U23199 ( .A1(n20273), .A2(n20292), .B1(n20272), .B2(n20291), .ZN(
        n20776) );
  INV_X1 U23200 ( .A(n20776), .ZN(n20726) );
  INV_X1 U23201 ( .A(DATAI_28_), .ZN(n21050) );
  OAI22_X1 U23202 ( .A1(n14815), .A2(n20292), .B1(n21050), .B2(n20291), .ZN(
        n20723) );
  NAND2_X1 U23203 ( .A1(n20286), .A2(n13002), .ZN(n20574) );
  AOI22_X1 U23204 ( .A1(n20797), .A2(n9945), .B1(n20775), .B2(n20296), .ZN(
        n20276) );
  AOI22_X1 U23205 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20299), .B1(
        n20774), .B2(n20298), .ZN(n20275) );
  OAI211_X1 U23206 ( .C1(n20726), .C2(n20327), .A(n20276), .B(n20275), .ZN(
        P1_U3037) );
  INV_X1 U23207 ( .A(DATAI_21_), .ZN(n21140) );
  OAI22_X1 U23208 ( .A1(n20277), .A2(n20292), .B1(n21140), .B2(n20291), .ZN(
        n20781) );
  INV_X1 U23209 ( .A(n20781), .ZN(n20730) );
  INV_X1 U23210 ( .A(DATAI_29_), .ZN(n20278) );
  OAI22_X1 U23211 ( .A1(n20279), .A2(n20292), .B1(n20278), .B2(n20291), .ZN(
        n20727) );
  NAND2_X1 U23212 ( .A1(n20286), .A2(n20280), .ZN(n20578) );
  AOI22_X1 U23213 ( .A1(n20797), .A2(n9947), .B1(n20780), .B2(n20296), .ZN(
        n20283) );
  AOI22_X1 U23214 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20299), .B1(
        n20779), .B2(n20298), .ZN(n20282) );
  OAI211_X1 U23215 ( .C1(n20730), .C2(n20327), .A(n20283), .B(n20282), .ZN(
        P1_U3038) );
  INV_X1 U23216 ( .A(DATAI_22_), .ZN(n21001) );
  OAI22_X1 U23217 ( .A1(n20284), .A2(n20292), .B1(n21001), .B2(n20291), .ZN(
        n20658) );
  INV_X1 U23218 ( .A(n20658), .ZN(n20791) );
  INV_X1 U23219 ( .A(DATAI_30_), .ZN(n21287) );
  OAI22_X2 U23220 ( .A1(n14805), .A2(n20292), .B1(n21287), .B2(n20291), .ZN(
        n20786) );
  NAND2_X1 U23221 ( .A1(n20286), .A2(n20285), .ZN(n20583) );
  AOI22_X1 U23222 ( .A1(n20797), .A2(n20786), .B1(n20785), .B2(n20296), .ZN(
        n20289) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20299), .B1(
        n20784), .B2(n20298), .ZN(n20288) );
  OAI211_X1 U23224 ( .C1(n20791), .C2(n20327), .A(n20289), .B(n20288), .ZN(
        P1_U3039) );
  INV_X1 U23225 ( .A(DATAI_23_), .ZN(n21159) );
  OAI22_X1 U23226 ( .A1(n20290), .A2(n20292), .B1(n21159), .B2(n20291), .ZN(
        n20796) );
  INV_X1 U23227 ( .A(DATAI_31_), .ZN(n21002) );
  NOR2_X2 U23228 ( .A1(n20295), .A2(n20294), .ZN(n20793) );
  AOI22_X1 U23229 ( .A1(n20797), .A2(n20735), .B1(n20793), .B2(n20296), .ZN(
        n20301) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20299), .B1(
        n20795), .B2(n20298), .ZN(n20300) );
  OAI211_X1 U23231 ( .C1(n9938), .C2(n20327), .A(n20301), .B(n20300), .ZN(
        P1_U3040) );
  INV_X1 U23232 ( .A(n20306), .ZN(n20303) );
  NOR2_X1 U23233 ( .A1(n20670), .A2(n20303), .ZN(n20322) );
  INV_X1 U23234 ( .A(n20302), .ZN(n20671) );
  AOI21_X1 U23235 ( .B1(n10140), .B2(n20671), .A(n20322), .ZN(n20304) );
  OAI22_X1 U23236 ( .A1(n20304), .A2(n20747), .B1(n20303), .B2(n12749), .ZN(
        n20323) );
  AOI22_X1 U23237 ( .A1(n20744), .A2(n20322), .B1(n20323), .B2(n20743), .ZN(
        n20309) );
  INV_X1 U23238 ( .A(n20360), .ZN(n20363) );
  OAI21_X1 U23239 ( .B1(n20363), .B2(n20703), .A(n20304), .ZN(n20305) );
  OAI221_X1 U23240 ( .B1(n20625), .B2(n20306), .C1(n20747), .C2(n20305), .A(
        n20752), .ZN(n20324) );
  INV_X1 U23241 ( .A(n20669), .ZN(n20307) );
  AOI22_X1 U23242 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20324), .B1(
        n20351), .B2(n20753), .ZN(n20308) );
  OAI211_X1 U23243 ( .C1(n9940), .C2(n20327), .A(n20309), .B(n20308), .ZN(
        P1_U3041) );
  INV_X1 U23244 ( .A(n20758), .ZN(n20607) );
  AOI22_X1 U23245 ( .A1(n20757), .A2(n20322), .B1(n20323), .B2(n20756), .ZN(
        n20311) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20324), .B1(
        n20351), .B2(n20641), .ZN(n20310) );
  OAI211_X1 U23247 ( .C1(n20607), .C2(n20327), .A(n20311), .B(n20310), .ZN(
        P1_U3042) );
  AOI22_X1 U23248 ( .A1(n20763), .A2(n20322), .B1(n20323), .B2(n20762), .ZN(
        n20313) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20324), .B1(
        n20351), .B2(n20764), .ZN(n20312) );
  OAI211_X1 U23250 ( .C1(n20767), .C2(n20327), .A(n20313), .B(n20312), .ZN(
        P1_U3043) );
  AOI22_X1 U23251 ( .A1(n20769), .A2(n20322), .B1(n20323), .B2(n20768), .ZN(
        n20315) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20324), .B1(
        n20351), .B2(n20648), .ZN(n20314) );
  OAI211_X1 U23253 ( .C1(n9942), .C2(n20327), .A(n20315), .B(n20314), .ZN(
        P1_U3044) );
  AOI22_X1 U23254 ( .A1(n20775), .A2(n20322), .B1(n20323), .B2(n20774), .ZN(
        n20317) );
  AOI22_X1 U23255 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20324), .B1(
        n20351), .B2(n20776), .ZN(n20316) );
  OAI211_X1 U23256 ( .C1(n9944), .C2(n20327), .A(n20317), .B(n20316), .ZN(
        P1_U3045) );
  AOI22_X1 U23257 ( .A1(n20780), .A2(n20322), .B1(n20323), .B2(n20779), .ZN(
        n20319) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20324), .B1(
        n20351), .B2(n20781), .ZN(n20318) );
  OAI211_X1 U23259 ( .C1(n9946), .C2(n20327), .A(n20319), .B(n20318), .ZN(
        P1_U3046) );
  INV_X1 U23260 ( .A(n20786), .ZN(n20618) );
  AOI22_X1 U23261 ( .A1(n20785), .A2(n20322), .B1(n20323), .B2(n20784), .ZN(
        n20321) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20324), .B1(
        n20351), .B2(n20658), .ZN(n20320) );
  OAI211_X1 U23263 ( .C1(n20618), .C2(n20327), .A(n20321), .B(n20320), .ZN(
        P1_U3047) );
  INV_X1 U23264 ( .A(n20735), .ZN(n20802) );
  AOI22_X1 U23265 ( .A1(n20323), .A2(n20795), .B1(n20793), .B2(n20322), .ZN(
        n20326) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20324), .B1(
        n20351), .B2(n9939), .ZN(n20325) );
  OAI211_X1 U23267 ( .C1(n20802), .C2(n20327), .A(n20326), .B(n20325), .ZN(
        P1_U3048) );
  INV_X1 U23268 ( .A(n20351), .ZN(n20328) );
  NAND2_X1 U23269 ( .A1(n20328), .A2(n20625), .ZN(n20330) );
  OAI21_X1 U23270 ( .B1(n20330), .B2(n20384), .A(n20882), .ZN(n20331) );
  NOR2_X1 U23271 ( .A1(n20359), .A2(n20702), .ZN(n20334) );
  INV_X1 U23272 ( .A(n20743), .ZN(n20640) );
  NOR3_X1 U23273 ( .A1(n20631), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20364) );
  NAND2_X1 U23274 ( .A1(n20670), .A2(n20364), .ZN(n20332) );
  INV_X1 U23275 ( .A(n20332), .ZN(n20350) );
  AOI22_X1 U23276 ( .A1(n20351), .A2(n9941), .B1(n20744), .B2(n20350), .ZN(
        n20337) );
  INV_X1 U23277 ( .A(n20331), .ZN(n20335) );
  NOR2_X1 U23278 ( .A1(n9933), .A2(n12749), .ZN(n20445) );
  AOI21_X1 U23279 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20332), .A(n20445), 
        .ZN(n20333) );
  AOI22_X1 U23280 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20352), .B1(
        n20384), .B2(n20753), .ZN(n20336) );
  OAI211_X1 U23281 ( .C1(n20355), .C2(n20640), .A(n20337), .B(n20336), .ZN(
        P1_U3049) );
  INV_X1 U23282 ( .A(n20756), .ZN(n20644) );
  AOI22_X1 U23283 ( .A1(n20351), .A2(n20758), .B1(n20757), .B2(n20350), .ZN(
        n20339) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20352), .B1(
        n20384), .B2(n20641), .ZN(n20338) );
  OAI211_X1 U23285 ( .C1(n20355), .C2(n20644), .A(n20339), .B(n20338), .ZN(
        P1_U3050) );
  INV_X1 U23286 ( .A(n20762), .ZN(n20647) );
  AOI22_X1 U23287 ( .A1(n20384), .A2(n20764), .B1(n20763), .B2(n20350), .ZN(
        n20341) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20352), .B1(
        n20351), .B2(n20717), .ZN(n20340) );
  OAI211_X1 U23289 ( .C1(n20355), .C2(n20647), .A(n20341), .B(n20340), .ZN(
        P1_U3051) );
  INV_X1 U23290 ( .A(n20768), .ZN(n20651) );
  AOI22_X1 U23291 ( .A1(n20384), .A2(n20648), .B1(n20769), .B2(n20350), .ZN(
        n20343) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20352), .B1(
        n20351), .B2(n9943), .ZN(n20342) );
  OAI211_X1 U23293 ( .C1(n20355), .C2(n20651), .A(n20343), .B(n20342), .ZN(
        P1_U3052) );
  INV_X1 U23294 ( .A(n20774), .ZN(n20654) );
  AOI22_X1 U23295 ( .A1(n20351), .A2(n9945), .B1(n20775), .B2(n20350), .ZN(
        n20345) );
  AOI22_X1 U23296 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20352), .B1(
        n20384), .B2(n20776), .ZN(n20344) );
  OAI211_X1 U23297 ( .C1(n20355), .C2(n20654), .A(n20345), .B(n20344), .ZN(
        P1_U3053) );
  INV_X1 U23298 ( .A(n20779), .ZN(n20657) );
  AOI22_X1 U23299 ( .A1(n20384), .A2(n20781), .B1(n20780), .B2(n20350), .ZN(
        n20347) );
  AOI22_X1 U23300 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20352), .B1(
        n20351), .B2(n9947), .ZN(n20346) );
  OAI211_X1 U23301 ( .C1(n20355), .C2(n20657), .A(n20347), .B(n20346), .ZN(
        P1_U3054) );
  INV_X1 U23302 ( .A(n20784), .ZN(n20661) );
  AOI22_X1 U23303 ( .A1(n20384), .A2(n20658), .B1(n20785), .B2(n20350), .ZN(
        n20349) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20352), .B1(
        n20351), .B2(n20786), .ZN(n20348) );
  OAI211_X1 U23305 ( .C1(n20355), .C2(n20661), .A(n20349), .B(n20348), .ZN(
        P1_U3055) );
  INV_X1 U23306 ( .A(n20795), .ZN(n20667) );
  AOI22_X1 U23307 ( .A1(n20351), .A2(n20735), .B1(n20793), .B2(n20350), .ZN(
        n20354) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20352), .B1(
        n20384), .B2(n9939), .ZN(n20353) );
  OAI211_X1 U23309 ( .C1(n20355), .C2(n20667), .A(n20354), .B(n20353), .ZN(
        P1_U3056) );
  AND2_X1 U23310 ( .A1(n20356), .A2(n12646), .ZN(n20741) );
  INV_X1 U23311 ( .A(n20741), .ZN(n20358) );
  NOR2_X1 U23312 ( .A1(n20595), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20383) );
  INV_X1 U23313 ( .A(n20383), .ZN(n20357) );
  OAI21_X1 U23314 ( .B1(n20359), .B2(n20358), .A(n20357), .ZN(n20367) );
  OR2_X1 U23315 ( .A1(n20360), .A2(n20747), .ZN(n20361) );
  AND2_X1 U23316 ( .A1(n20361), .A2(n20745), .ZN(n20368) );
  INV_X1 U23317 ( .A(n20368), .ZN(n20362) );
  AOI22_X1 U23318 ( .A1(n20414), .A2(n20753), .B1(n20744), .B2(n20383), .ZN(
        n20370) );
  INV_X1 U23319 ( .A(n20364), .ZN(n20365) );
  INV_X1 U23320 ( .A(n20752), .ZN(n20674) );
  AOI21_X1 U23321 ( .B1(n20747), .B2(n20365), .A(n20674), .ZN(n20366) );
  OAI21_X1 U23322 ( .B1(n20368), .B2(n20367), .A(n20366), .ZN(n20385) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n9941), .ZN(n20369) );
  OAI211_X1 U23324 ( .C1(n20388), .C2(n20640), .A(n20370), .B(n20369), .ZN(
        P1_U3057) );
  AOI22_X1 U23325 ( .A1(n20414), .A2(n20641), .B1(n20757), .B2(n20383), .ZN(
        n20372) );
  AOI22_X1 U23326 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20758), .ZN(n20371) );
  OAI211_X1 U23327 ( .C1(n20388), .C2(n20644), .A(n20372), .B(n20371), .ZN(
        P1_U3058) );
  AOI22_X1 U23328 ( .A1(n20414), .A2(n20764), .B1(n20763), .B2(n20383), .ZN(
        n20374) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20717), .ZN(n20373) );
  OAI211_X1 U23330 ( .C1(n20388), .C2(n20647), .A(n20374), .B(n20373), .ZN(
        P1_U3059) );
  AOI22_X1 U23331 ( .A1(n20384), .A2(n9943), .B1(n20769), .B2(n20383), .ZN(
        n20376) );
  AOI22_X1 U23332 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20385), .B1(
        n20414), .B2(n20648), .ZN(n20375) );
  OAI211_X1 U23333 ( .C1(n20388), .C2(n20651), .A(n20376), .B(n20375), .ZN(
        P1_U3060) );
  AOI22_X1 U23334 ( .A1(n20414), .A2(n20776), .B1(n20775), .B2(n20383), .ZN(
        n20378) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n9945), .ZN(n20377) );
  OAI211_X1 U23336 ( .C1(n20388), .C2(n20654), .A(n20378), .B(n20377), .ZN(
        P1_U3061) );
  AOI22_X1 U23337 ( .A1(n20384), .A2(n9947), .B1(n20780), .B2(n20383), .ZN(
        n20380) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20385), .B1(
        n20414), .B2(n20781), .ZN(n20379) );
  OAI211_X1 U23339 ( .C1(n20388), .C2(n20657), .A(n20380), .B(n20379), .ZN(
        P1_U3062) );
  AOI22_X1 U23340 ( .A1(n20414), .A2(n20658), .B1(n20785), .B2(n20383), .ZN(
        n20382) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20786), .ZN(n20381) );
  OAI211_X1 U23342 ( .C1(n20388), .C2(n20661), .A(n20382), .B(n20381), .ZN(
        P1_U3063) );
  AOI22_X1 U23343 ( .A1(n20414), .A2(n9939), .B1(n20793), .B2(n20383), .ZN(
        n20387) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20735), .ZN(n20386) );
  OAI211_X1 U23345 ( .C1(n20388), .C2(n20667), .A(n20387), .B(n20386), .ZN(
        P1_U3064) );
  NOR3_X1 U23346 ( .A1(n12471), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20421) );
  INV_X1 U23347 ( .A(n20421), .ZN(n20418) );
  NOR2_X1 U23348 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20418), .ZN(
        n20412) );
  INV_X1 U23349 ( .A(n20630), .ZN(n20700) );
  NOR2_X1 U23350 ( .A1(n13189), .A2(n20390), .ZN(n20470) );
  NAND3_X1 U23351 ( .A1(n20470), .A2(n20625), .A3(n20702), .ZN(n20391) );
  OAI21_X1 U23352 ( .B1(n20392), .B2(n20700), .A(n20391), .ZN(n20413) );
  AOI22_X1 U23353 ( .A1(n20744), .A2(n20412), .B1(n20743), .B2(n20413), .ZN(
        n20399) );
  INV_X1 U23354 ( .A(n20414), .ZN(n20393) );
  AOI21_X1 U23355 ( .B1(n20393), .B2(n20441), .A(n20703), .ZN(n20394) );
  AOI21_X1 U23356 ( .B1(n20470), .B2(n20702), .A(n20394), .ZN(n20395) );
  NOR2_X1 U23357 ( .A1(n20395), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20397) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n9941), .ZN(n20398) );
  OAI211_X1 U23359 ( .C1(n20714), .C2(n20441), .A(n20399), .B(n20398), .ZN(
        P1_U3065) );
  AOI22_X1 U23360 ( .A1(n20757), .A2(n20412), .B1(n20756), .B2(n20413), .ZN(
        n20401) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n20758), .ZN(n20400) );
  OAI211_X1 U23362 ( .C1(n20761), .C2(n20441), .A(n20401), .B(n20400), .ZN(
        P1_U3066) );
  AOI22_X1 U23363 ( .A1(n20763), .A2(n20412), .B1(n20762), .B2(n20413), .ZN(
        n20403) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n20717), .ZN(n20402) );
  OAI211_X1 U23365 ( .C1(n20720), .C2(n20441), .A(n20403), .B(n20402), .ZN(
        P1_U3067) );
  AOI22_X1 U23366 ( .A1(n20769), .A2(n20412), .B1(n20768), .B2(n20413), .ZN(
        n20405) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n9943), .ZN(n20404) );
  OAI211_X1 U23368 ( .C1(n20773), .C2(n20441), .A(n20405), .B(n20404), .ZN(
        P1_U3068) );
  AOI22_X1 U23369 ( .A1(n20775), .A2(n20412), .B1(n20774), .B2(n20413), .ZN(
        n20407) );
  AOI22_X1 U23370 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n9945), .ZN(n20406) );
  OAI211_X1 U23371 ( .C1(n20726), .C2(n20441), .A(n20407), .B(n20406), .ZN(
        P1_U3069) );
  AOI22_X1 U23372 ( .A1(n20780), .A2(n20412), .B1(n20779), .B2(n20413), .ZN(
        n20409) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n9947), .ZN(n20408) );
  OAI211_X1 U23374 ( .C1(n20730), .C2(n20441), .A(n20409), .B(n20408), .ZN(
        P1_U3070) );
  AOI22_X1 U23375 ( .A1(n20785), .A2(n20412), .B1(n20784), .B2(n20413), .ZN(
        n20411) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n20786), .ZN(n20410) );
  OAI211_X1 U23377 ( .C1(n20791), .C2(n20441), .A(n20411), .B(n20410), .ZN(
        P1_U3071) );
  AOI22_X1 U23378 ( .A1(n20795), .A2(n20413), .B1(n20793), .B2(n20412), .ZN(
        n20417) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20415), .B1(
        n20414), .B2(n20735), .ZN(n20416) );
  OAI211_X1 U23380 ( .C1(n9938), .C2(n20441), .A(n20417), .B(n20416), .ZN(
        P1_U3072) );
  NOR2_X1 U23381 ( .A1(n20670), .A2(n20418), .ZN(n20436) );
  AOI21_X1 U23382 ( .B1(n20470), .B2(n20671), .A(n20436), .ZN(n20419) );
  OAI22_X1 U23383 ( .A1(n20419), .A2(n20747), .B1(n20418), .B2(n12749), .ZN(
        n20437) );
  AOI22_X1 U23384 ( .A1(n20744), .A2(n20436), .B1(n20743), .B2(n20437), .ZN(
        n20423) );
  OAI21_X1 U23385 ( .B1(n20473), .B2(n20703), .A(n20419), .ZN(n20420) );
  OAI221_X1 U23386 ( .B1(n20625), .B2(n20421), .C1(n20747), .C2(n20420), .A(
        n20752), .ZN(n20438) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20438), .B1(
        n20464), .B2(n20753), .ZN(n20422) );
  OAI211_X1 U23388 ( .C1(n9940), .C2(n20441), .A(n20423), .B(n20422), .ZN(
        P1_U3073) );
  AOI22_X1 U23389 ( .A1(n20757), .A2(n20436), .B1(n20756), .B2(n20437), .ZN(
        n20425) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20438), .B1(
        n20464), .B2(n20641), .ZN(n20424) );
  OAI211_X1 U23391 ( .C1(n20607), .C2(n20441), .A(n20425), .B(n20424), .ZN(
        P1_U3074) );
  AOI22_X1 U23392 ( .A1(n20763), .A2(n20436), .B1(n20762), .B2(n20437), .ZN(
        n20427) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20438), .B1(
        n20464), .B2(n20764), .ZN(n20426) );
  OAI211_X1 U23394 ( .C1(n20767), .C2(n20441), .A(n20427), .B(n20426), .ZN(
        P1_U3075) );
  AOI22_X1 U23395 ( .A1(n20769), .A2(n20436), .B1(n20768), .B2(n20437), .ZN(
        n20429) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20438), .B1(
        n20464), .B2(n20648), .ZN(n20428) );
  OAI211_X1 U23397 ( .C1(n9942), .C2(n20441), .A(n20429), .B(n20428), .ZN(
        P1_U3076) );
  AOI22_X1 U23398 ( .A1(n20775), .A2(n20436), .B1(n20774), .B2(n20437), .ZN(
        n20431) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20438), .B1(
        n20464), .B2(n20776), .ZN(n20430) );
  OAI211_X1 U23400 ( .C1(n9944), .C2(n20441), .A(n20431), .B(n20430), .ZN(
        P1_U3077) );
  AOI22_X1 U23401 ( .A1(n20780), .A2(n20436), .B1(n20779), .B2(n20437), .ZN(
        n20433) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20438), .B1(
        n20464), .B2(n20781), .ZN(n20432) );
  OAI211_X1 U23403 ( .C1(n9946), .C2(n20441), .A(n20433), .B(n20432), .ZN(
        P1_U3078) );
  AOI22_X1 U23404 ( .A1(n20785), .A2(n20436), .B1(n20784), .B2(n20437), .ZN(
        n20435) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20438), .B1(
        n20464), .B2(n20658), .ZN(n20434) );
  OAI211_X1 U23406 ( .C1(n20618), .C2(n20441), .A(n20435), .B(n20434), .ZN(
        P1_U3079) );
  AOI22_X1 U23407 ( .A1(n20795), .A2(n20437), .B1(n20793), .B2(n20436), .ZN(
        n20440) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20438), .B1(
        n20464), .B2(n9939), .ZN(n20439) );
  OAI211_X1 U23409 ( .C1(n20802), .C2(n20441), .A(n20440), .B(n20439), .ZN(
        P1_U3080) );
  INV_X1 U23410 ( .A(n20464), .ZN(n20442) );
  NAND2_X1 U23411 ( .A1(n20442), .A2(n20625), .ZN(n20443) );
  OAI21_X1 U23412 ( .B1(n20443), .B2(n20492), .A(n20882), .ZN(n20447) );
  AND2_X1 U23413 ( .A1(n20470), .A2(n20705), .ZN(n20444) );
  NOR2_X1 U23414 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20471), .ZN(
        n20463) );
  AOI22_X1 U23415 ( .A1(n20492), .A2(n20753), .B1(n20463), .B2(n20744), .ZN(
        n20450) );
  INV_X1 U23416 ( .A(n20444), .ZN(n20446) );
  AOI21_X1 U23417 ( .B1(n20447), .B2(n20446), .A(n20445), .ZN(n20448) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n9941), .ZN(n20449) );
  OAI211_X1 U23419 ( .C1(n20468), .C2(n20640), .A(n20450), .B(n20449), .ZN(
        P1_U3081) );
  AOI22_X1 U23420 ( .A1(n20492), .A2(n20641), .B1(n20463), .B2(n20757), .ZN(
        n20452) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20758), .ZN(n20451) );
  OAI211_X1 U23422 ( .C1(n20468), .C2(n20644), .A(n20452), .B(n20451), .ZN(
        P1_U3082) );
  AOI22_X1 U23423 ( .A1(n20492), .A2(n20764), .B1(n20463), .B2(n20763), .ZN(
        n20454) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20717), .ZN(n20453) );
  OAI211_X1 U23425 ( .C1(n20468), .C2(n20647), .A(n20454), .B(n20453), .ZN(
        P1_U3083) );
  AOI22_X1 U23426 ( .A1(n20464), .A2(n9943), .B1(n20769), .B2(n20463), .ZN(
        n20456) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20465), .B1(
        n20492), .B2(n20648), .ZN(n20455) );
  OAI211_X1 U23428 ( .C1(n20468), .C2(n20651), .A(n20456), .B(n20455), .ZN(
        P1_U3084) );
  AOI22_X1 U23429 ( .A1(n20492), .A2(n20776), .B1(n20463), .B2(n20775), .ZN(
        n20458) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n9945), .ZN(n20457) );
  OAI211_X1 U23431 ( .C1(n20468), .C2(n20654), .A(n20458), .B(n20457), .ZN(
        P1_U3085) );
  AOI22_X1 U23432 ( .A1(n20492), .A2(n20781), .B1(n20463), .B2(n20780), .ZN(
        n20460) );
  AOI22_X1 U23433 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n9947), .ZN(n20459) );
  OAI211_X1 U23434 ( .C1(n20468), .C2(n20657), .A(n20460), .B(n20459), .ZN(
        P1_U3086) );
  AOI22_X1 U23435 ( .A1(n20464), .A2(n20786), .B1(n20463), .B2(n20785), .ZN(
        n20462) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20465), .B1(
        n20492), .B2(n20658), .ZN(n20461) );
  OAI211_X1 U23437 ( .C1(n20468), .C2(n20661), .A(n20462), .B(n20461), .ZN(
        P1_U3087) );
  AOI22_X1 U23438 ( .A1(n20492), .A2(n9939), .B1(n20463), .B2(n20793), .ZN(
        n20467) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20735), .ZN(n20466) );
  OAI211_X1 U23440 ( .C1(n20468), .C2(n20667), .A(n20467), .B(n20466), .ZN(
        P1_U3088) );
  INV_X1 U23441 ( .A(n20469), .ZN(n20490) );
  AOI21_X1 U23442 ( .B1(n20470), .B2(n20741), .A(n20490), .ZN(n20472) );
  OAI22_X1 U23443 ( .A1(n20472), .A2(n20747), .B1(n20471), .B2(n12749), .ZN(
        n20491) );
  AOI22_X1 U23444 ( .A1(n20744), .A2(n20490), .B1(n20743), .B2(n20491), .ZN(
        n20477) );
  OR2_X1 U23445 ( .A1(n20473), .A2(n20599), .ZN(n20887) );
  INV_X1 U23446 ( .A(n20887), .ZN(n20475) );
  OAI21_X1 U23447 ( .B1(n20475), .B2(n20474), .A(n20752), .ZN(n20493) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20493), .B1(
        n20492), .B2(n9941), .ZN(n20476) );
  OAI211_X1 U23449 ( .C1(n20714), .C2(n20499), .A(n20477), .B(n20476), .ZN(
        P1_U3089) );
  AOI22_X1 U23450 ( .A1(n20757), .A2(n20490), .B1(n20756), .B2(n20491), .ZN(
        n20479) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20493), .B1(
        n20492), .B2(n20758), .ZN(n20478) );
  OAI211_X1 U23452 ( .C1(n20761), .C2(n20499), .A(n20479), .B(n20478), .ZN(
        P1_U3090) );
  AOI22_X1 U23453 ( .A1(n20763), .A2(n20490), .B1(n20762), .B2(n20491), .ZN(
        n20481) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20493), .B1(
        n20492), .B2(n20717), .ZN(n20480) );
  OAI211_X1 U23455 ( .C1(n20720), .C2(n20499), .A(n20481), .B(n20480), .ZN(
        P1_U3091) );
  AOI22_X1 U23456 ( .A1(n20769), .A2(n20490), .B1(n20768), .B2(n20491), .ZN(
        n20483) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20493), .B1(
        n20492), .B2(n9943), .ZN(n20482) );
  OAI211_X1 U23458 ( .C1(n20773), .C2(n20499), .A(n20483), .B(n20482), .ZN(
        P1_U3092) );
  AOI22_X1 U23459 ( .A1(n20775), .A2(n20490), .B1(n20774), .B2(n20491), .ZN(
        n20485) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20493), .B1(
        n20492), .B2(n9945), .ZN(n20484) );
  OAI211_X1 U23461 ( .C1(n20726), .C2(n20499), .A(n20485), .B(n20484), .ZN(
        P1_U3093) );
  AOI22_X1 U23462 ( .A1(n20780), .A2(n20490), .B1(n20779), .B2(n20491), .ZN(
        n20487) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20493), .B1(
        n20492), .B2(n9947), .ZN(n20486) );
  OAI211_X1 U23464 ( .C1(n20730), .C2(n20499), .A(n20487), .B(n20486), .ZN(
        P1_U3094) );
  AOI22_X1 U23465 ( .A1(n20785), .A2(n20490), .B1(n20784), .B2(n20491), .ZN(
        n20489) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20493), .B1(
        n20492), .B2(n20786), .ZN(n20488) );
  OAI211_X1 U23467 ( .C1(n20791), .C2(n20499), .A(n20489), .B(n20488), .ZN(
        P1_U3095) );
  AOI22_X1 U23468 ( .A1(n20795), .A2(n20491), .B1(n20793), .B2(n20490), .ZN(
        n20495) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20493), .B1(
        n20492), .B2(n20735), .ZN(n20494) );
  OAI211_X1 U23470 ( .C1(n9938), .C2(n20499), .A(n20495), .B(n20494), .ZN(
        P1_U3096) );
  NOR3_X1 U23471 ( .A1(n20594), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20527) );
  INV_X1 U23472 ( .A(n20527), .ZN(n20524) );
  NOR2_X1 U23473 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20524), .ZN(
        n20518) );
  AOI21_X1 U23474 ( .B1(n20596), .B2(n20702), .A(n20518), .ZN(n20501) );
  AND2_X1 U23475 ( .A1(n20497), .A2(n20699), .ZN(n20629) );
  INV_X1 U23476 ( .A(n20629), .ZN(n20633) );
  OAI22_X1 U23477 ( .A1(n20501), .A2(n20747), .B1(n20633), .B2(n20498), .ZN(
        n20519) );
  AOI22_X1 U23478 ( .A1(n20744), .A2(n20518), .B1(n20519), .B2(n20743), .ZN(
        n20505) );
  INV_X1 U23479 ( .A(n20547), .ZN(n20500) );
  OAI21_X1 U23480 ( .B1(n20500), .B2(n20520), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20502) );
  NAND2_X1 U23481 ( .A1(n20502), .A2(n20501), .ZN(n20503) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n9941), .ZN(n20504) );
  OAI211_X1 U23483 ( .C1(n20714), .C2(n20547), .A(n20505), .B(n20504), .ZN(
        P1_U3097) );
  AOI22_X1 U23484 ( .A1(n20757), .A2(n20518), .B1(n20519), .B2(n20756), .ZN(
        n20507) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20758), .ZN(n20506) );
  OAI211_X1 U23486 ( .C1(n20761), .C2(n20547), .A(n20507), .B(n20506), .ZN(
        P1_U3098) );
  AOI22_X1 U23487 ( .A1(n20763), .A2(n20518), .B1(n20762), .B2(n20519), .ZN(
        n20509) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20717), .ZN(n20508) );
  OAI211_X1 U23489 ( .C1(n20720), .C2(n20547), .A(n20509), .B(n20508), .ZN(
        P1_U3099) );
  AOI22_X1 U23490 ( .A1(n20769), .A2(n20518), .B1(n20768), .B2(n20519), .ZN(
        n20511) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n9943), .ZN(n20510) );
  OAI211_X1 U23492 ( .C1(n20773), .C2(n20547), .A(n20511), .B(n20510), .ZN(
        P1_U3100) );
  AOI22_X1 U23493 ( .A1(n20775), .A2(n20518), .B1(n20774), .B2(n20519), .ZN(
        n20513) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n9945), .ZN(n20512) );
  OAI211_X1 U23495 ( .C1(n20726), .C2(n20547), .A(n20513), .B(n20512), .ZN(
        P1_U3101) );
  AOI22_X1 U23496 ( .A1(n20780), .A2(n20518), .B1(n20779), .B2(n20519), .ZN(
        n20515) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n9947), .ZN(n20514) );
  OAI211_X1 U23498 ( .C1(n20730), .C2(n20547), .A(n20515), .B(n20514), .ZN(
        P1_U3102) );
  AOI22_X1 U23499 ( .A1(n20785), .A2(n20518), .B1(n20784), .B2(n20519), .ZN(
        n20517) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20786), .ZN(n20516) );
  OAI211_X1 U23501 ( .C1(n20791), .C2(n20547), .A(n20517), .B(n20516), .ZN(
        P1_U3103) );
  AOI22_X1 U23502 ( .A1(n20795), .A2(n20519), .B1(n20793), .B2(n20518), .ZN(
        n20523) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20735), .ZN(n20522) );
  OAI211_X1 U23504 ( .C1(n9938), .C2(n20547), .A(n20523), .B(n20522), .ZN(
        P1_U3104) );
  NOR2_X1 U23505 ( .A1(n20670), .A2(n20524), .ZN(n20542) );
  AOI21_X1 U23506 ( .B1(n20596), .B2(n20671), .A(n20542), .ZN(n20525) );
  OAI22_X1 U23507 ( .A1(n20525), .A2(n20747), .B1(n20524), .B2(n12749), .ZN(
        n20543) );
  AOI22_X1 U23508 ( .A1(n20744), .A2(n20542), .B1(n20543), .B2(n20743), .ZN(
        n20529) );
  OAI21_X1 U23509 ( .B1(n20602), .B2(n20703), .A(n20525), .ZN(n20526) );
  OAI221_X1 U23510 ( .B1(n20625), .B2(n20527), .C1(n20747), .C2(n20526), .A(
        n20752), .ZN(n20544) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20544), .B1(
        n20588), .B2(n20753), .ZN(n20528) );
  OAI211_X1 U23512 ( .C1(n9940), .C2(n20547), .A(n20529), .B(n20528), .ZN(
        P1_U3105) );
  AOI22_X1 U23513 ( .A1(n20757), .A2(n20542), .B1(n20543), .B2(n20756), .ZN(
        n20531) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20544), .B1(
        n20588), .B2(n20641), .ZN(n20530) );
  OAI211_X1 U23515 ( .C1(n20607), .C2(n20547), .A(n20531), .B(n20530), .ZN(
        P1_U3106) );
  AOI22_X1 U23516 ( .A1(n20763), .A2(n20542), .B1(n20762), .B2(n20543), .ZN(
        n20533) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20544), .B1(
        n20588), .B2(n20764), .ZN(n20532) );
  OAI211_X1 U23518 ( .C1(n20767), .C2(n20547), .A(n20533), .B(n20532), .ZN(
        P1_U3107) );
  AOI22_X1 U23519 ( .A1(n20769), .A2(n20542), .B1(n20768), .B2(n20543), .ZN(
        n20535) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20544), .B1(
        n20588), .B2(n20648), .ZN(n20534) );
  OAI211_X1 U23521 ( .C1(n9942), .C2(n20547), .A(n20535), .B(n20534), .ZN(
        P1_U3108) );
  AOI22_X1 U23522 ( .A1(n20775), .A2(n20542), .B1(n20774), .B2(n20543), .ZN(
        n20537) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20544), .B1(
        n20588), .B2(n20776), .ZN(n20536) );
  OAI211_X1 U23524 ( .C1(n9944), .C2(n20547), .A(n20537), .B(n20536), .ZN(
        P1_U3109) );
  AOI22_X1 U23525 ( .A1(n20780), .A2(n20542), .B1(n20779), .B2(n20543), .ZN(
        n20539) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20544), .B1(
        n20588), .B2(n20781), .ZN(n20538) );
  OAI211_X1 U23527 ( .C1(n9946), .C2(n20547), .A(n20539), .B(n20538), .ZN(
        P1_U3110) );
  AOI22_X1 U23528 ( .A1(n20785), .A2(n20542), .B1(n20784), .B2(n20543), .ZN(
        n20541) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20544), .B1(
        n20588), .B2(n20658), .ZN(n20540) );
  OAI211_X1 U23530 ( .C1(n20618), .C2(n20547), .A(n20541), .B(n20540), .ZN(
        P1_U3111) );
  AOI22_X1 U23531 ( .A1(n20795), .A2(n20543), .B1(n20793), .B2(n20542), .ZN(
        n20546) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20544), .B1(
        n20588), .B2(n9939), .ZN(n20545) );
  OAI211_X1 U23533 ( .C1(n20802), .C2(n20547), .A(n20546), .B(n20545), .ZN(
        P1_U3112) );
  INV_X1 U23534 ( .A(n20588), .ZN(n20549) );
  NAND3_X1 U23535 ( .A1(n20549), .A2(n20625), .A3(n20624), .ZN(n20550) );
  NAND2_X1 U23536 ( .A1(n20550), .A2(n20882), .ZN(n20557) );
  AND2_X1 U23537 ( .A1(n20596), .A2(n20705), .ZN(n20555) );
  NOR2_X1 U23538 ( .A1(n20699), .A2(n20594), .ZN(n20551) );
  NAND3_X1 U23539 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n12471), .ZN(n20598) );
  NOR2_X1 U23540 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20598), .ZN(
        n20587) );
  INV_X1 U23541 ( .A(n20587), .ZN(n20582) );
  OAI22_X1 U23542 ( .A1(n20624), .A2(n20714), .B1(n20553), .B2(n20582), .ZN(
        n20554) );
  INV_X1 U23543 ( .A(n20554), .ZN(n20561) );
  INV_X1 U23544 ( .A(n20555), .ZN(n20556) );
  AOI22_X1 U23545 ( .A1(n20557), .A2(n20556), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20582), .ZN(n20558) );
  OAI21_X1 U23546 ( .B1(n20594), .B2(n20699), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20707) );
  NAND3_X1 U23547 ( .A1(n20559), .A2(n20558), .A3(n20707), .ZN(n20590) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20590), .B1(
        n20588), .B2(n9941), .ZN(n20560) );
  OAI211_X1 U23549 ( .C1(n20593), .C2(n20640), .A(n20561), .B(n20560), .ZN(
        P1_U3113) );
  OAI22_X1 U23550 ( .A1(n20624), .A2(n20761), .B1(n20562), .B2(n20582), .ZN(
        n20563) );
  INV_X1 U23551 ( .A(n20563), .ZN(n20565) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20590), .B1(
        n20588), .B2(n20758), .ZN(n20564) );
  OAI211_X1 U23553 ( .C1(n20593), .C2(n20644), .A(n20565), .B(n20564), .ZN(
        P1_U3114) );
  OAI22_X1 U23554 ( .A1(n20624), .A2(n20720), .B1(n20566), .B2(n20582), .ZN(
        n20567) );
  INV_X1 U23555 ( .A(n20567), .ZN(n20569) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20590), .B1(
        n20588), .B2(n20717), .ZN(n20568) );
  OAI211_X1 U23557 ( .C1(n20593), .C2(n20647), .A(n20569), .B(n20568), .ZN(
        P1_U3115) );
  OAI22_X1 U23558 ( .A1(n20624), .A2(n20773), .B1(n20570), .B2(n20582), .ZN(
        n20571) );
  INV_X1 U23559 ( .A(n20571), .ZN(n20573) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20590), .B1(
        n20588), .B2(n9943), .ZN(n20572) );
  OAI211_X1 U23561 ( .C1(n20593), .C2(n20651), .A(n20573), .B(n20572), .ZN(
        P1_U3116) );
  OAI22_X1 U23562 ( .A1(n20624), .A2(n20726), .B1(n20574), .B2(n20582), .ZN(
        n20575) );
  INV_X1 U23563 ( .A(n20575), .ZN(n20577) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20590), .B1(
        n20588), .B2(n9945), .ZN(n20576) );
  OAI211_X1 U23565 ( .C1(n20593), .C2(n20654), .A(n20577), .B(n20576), .ZN(
        P1_U3117) );
  OAI22_X1 U23566 ( .A1(n20624), .A2(n20730), .B1(n20578), .B2(n20582), .ZN(
        n20579) );
  INV_X1 U23567 ( .A(n20579), .ZN(n20581) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20590), .B1(
        n20588), .B2(n9947), .ZN(n20580) );
  OAI211_X1 U23569 ( .C1(n20593), .C2(n20657), .A(n20581), .B(n20580), .ZN(
        P1_U3118) );
  OAI22_X1 U23570 ( .A1(n20624), .A2(n20791), .B1(n20583), .B2(n20582), .ZN(
        n20584) );
  INV_X1 U23571 ( .A(n20584), .ZN(n20586) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20590), .B1(
        n20588), .B2(n20786), .ZN(n20585) );
  OAI211_X1 U23573 ( .C1(n20593), .C2(n20661), .A(n20586), .B(n20585), .ZN(
        P1_U3119) );
  AOI22_X1 U23574 ( .A1(n20588), .A2(n20735), .B1(n20793), .B2(n20587), .ZN(
        n20592) );
  INV_X1 U23575 ( .A(n20624), .ZN(n20589) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n9939), .ZN(n20591) );
  OAI211_X1 U23577 ( .C1(n20593), .C2(n20667), .A(n20592), .B(n20591), .ZN(
        P1_U3120) );
  NOR2_X1 U23578 ( .A1(n20595), .A2(n20594), .ZN(n20619) );
  AOI21_X1 U23579 ( .B1(n20596), .B2(n20741), .A(n20619), .ZN(n20597) );
  OAI22_X1 U23580 ( .A1(n20597), .A2(n20747), .B1(n20598), .B2(n12749), .ZN(
        n20620) );
  AOI22_X1 U23581 ( .A1(n20744), .A2(n20619), .B1(n20743), .B2(n20620), .ZN(
        n20604) );
  OAI21_X1 U23582 ( .B1(n20602), .B2(n20599), .A(n20598), .ZN(n20600) );
  NAND2_X1 U23583 ( .A1(n20600), .A2(n20752), .ZN(n20621) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20621), .B1(
        n20663), .B2(n20753), .ZN(n20603) );
  OAI211_X1 U23585 ( .C1(n9940), .C2(n20624), .A(n20604), .B(n20603), .ZN(
        P1_U3121) );
  AOI22_X1 U23586 ( .A1(n20757), .A2(n20619), .B1(n20756), .B2(n20620), .ZN(
        n20606) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20621), .B1(
        n20663), .B2(n20641), .ZN(n20605) );
  OAI211_X1 U23588 ( .C1(n20607), .C2(n20624), .A(n20606), .B(n20605), .ZN(
        P1_U3122) );
  AOI22_X1 U23589 ( .A1(n20763), .A2(n20619), .B1(n20762), .B2(n20620), .ZN(
        n20609) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20621), .B1(
        n20663), .B2(n20764), .ZN(n20608) );
  OAI211_X1 U23591 ( .C1(n20767), .C2(n20624), .A(n20609), .B(n20608), .ZN(
        P1_U3123) );
  AOI22_X1 U23592 ( .A1(n20769), .A2(n20619), .B1(n20768), .B2(n20620), .ZN(
        n20611) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20621), .B1(
        n20663), .B2(n20648), .ZN(n20610) );
  OAI211_X1 U23594 ( .C1(n9942), .C2(n20624), .A(n20611), .B(n20610), .ZN(
        P1_U3124) );
  AOI22_X1 U23595 ( .A1(n20775), .A2(n20619), .B1(n20774), .B2(n20620), .ZN(
        n20613) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20621), .B1(
        n20663), .B2(n20776), .ZN(n20612) );
  OAI211_X1 U23597 ( .C1(n9944), .C2(n20624), .A(n20613), .B(n20612), .ZN(
        P1_U3125) );
  AOI22_X1 U23598 ( .A1(n20780), .A2(n20619), .B1(n20779), .B2(n20620), .ZN(
        n20615) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20621), .B1(
        n20663), .B2(n20781), .ZN(n20614) );
  OAI211_X1 U23600 ( .C1(n9946), .C2(n20624), .A(n20615), .B(n20614), .ZN(
        P1_U3126) );
  AOI22_X1 U23601 ( .A1(n20785), .A2(n20619), .B1(n20784), .B2(n20620), .ZN(
        n20617) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20621), .B1(
        n20663), .B2(n20658), .ZN(n20616) );
  OAI211_X1 U23603 ( .C1(n20618), .C2(n20624), .A(n20617), .B(n20616), .ZN(
        P1_U3127) );
  AOI22_X1 U23604 ( .A1(n20795), .A2(n20620), .B1(n20793), .B2(n20619), .ZN(
        n20623) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20621), .B1(
        n20663), .B2(n9939), .ZN(n20622) );
  OAI211_X1 U23606 ( .C1(n20802), .C2(n20624), .A(n20623), .B(n20622), .ZN(
        P1_U3128) );
  INV_X1 U23607 ( .A(n20663), .ZN(n20626) );
  NAND2_X1 U23608 ( .A1(n20626), .A2(n20625), .ZN(n20628) );
  NOR2_X2 U23609 ( .A1(n20698), .A2(n20627), .ZN(n20693) );
  OAI21_X1 U23610 ( .B1(n20628), .B2(n20693), .A(n20882), .ZN(n20635) );
  NOR2_X1 U23611 ( .A1(n13189), .A2(n10142), .ZN(n20742) );
  AND2_X1 U23612 ( .A1(n20742), .A2(n20702), .ZN(n20632) );
  NAND3_X1 U23613 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20631), .ZN(n20675) );
  NOR2_X1 U23614 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20675), .ZN(
        n20662) );
  AOI22_X1 U23615 ( .A1(n20693), .A2(n20753), .B1(n20744), .B2(n20662), .ZN(
        n20639) );
  INV_X1 U23616 ( .A(n20632), .ZN(n20634) );
  AOI22_X1 U23617 ( .A1(n20635), .A2(n20634), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20633), .ZN(n20636) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20664), .B1(
        n20663), .B2(n9941), .ZN(n20638) );
  OAI211_X1 U23619 ( .C1(n20668), .C2(n20640), .A(n20639), .B(n20638), .ZN(
        P1_U3129) );
  AOI22_X1 U23620 ( .A1(n20693), .A2(n20641), .B1(n20757), .B2(n20662), .ZN(
        n20643) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20664), .B1(
        n20663), .B2(n20758), .ZN(n20642) );
  OAI211_X1 U23622 ( .C1(n20668), .C2(n20644), .A(n20643), .B(n20642), .ZN(
        P1_U3130) );
  AOI22_X1 U23623 ( .A1(n20693), .A2(n20764), .B1(n20763), .B2(n20662), .ZN(
        n20646) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20664), .B1(
        n20663), .B2(n20717), .ZN(n20645) );
  OAI211_X1 U23625 ( .C1(n20668), .C2(n20647), .A(n20646), .B(n20645), .ZN(
        P1_U3131) );
  AOI22_X1 U23626 ( .A1(n20693), .A2(n20648), .B1(n20769), .B2(n20662), .ZN(
        n20650) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20664), .B1(
        n20663), .B2(n9943), .ZN(n20649) );
  OAI211_X1 U23628 ( .C1(n20668), .C2(n20651), .A(n20650), .B(n20649), .ZN(
        P1_U3132) );
  AOI22_X1 U23629 ( .A1(n20693), .A2(n20776), .B1(n20775), .B2(n20662), .ZN(
        n20653) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20664), .B1(
        n20663), .B2(n9945), .ZN(n20652) );
  OAI211_X1 U23631 ( .C1(n20668), .C2(n20654), .A(n20653), .B(n20652), .ZN(
        P1_U3133) );
  AOI22_X1 U23632 ( .A1(n20693), .A2(n20781), .B1(n20780), .B2(n20662), .ZN(
        n20656) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20664), .B1(
        n20663), .B2(n9947), .ZN(n20655) );
  OAI211_X1 U23634 ( .C1(n20668), .C2(n20657), .A(n20656), .B(n20655), .ZN(
        P1_U3134) );
  AOI22_X1 U23635 ( .A1(n20693), .A2(n20658), .B1(n20785), .B2(n20662), .ZN(
        n20660) );
  AOI22_X1 U23636 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20664), .B1(
        n20663), .B2(n20786), .ZN(n20659) );
  OAI211_X1 U23637 ( .C1(n20668), .C2(n20661), .A(n20660), .B(n20659), .ZN(
        P1_U3135) );
  AOI22_X1 U23638 ( .A1(n20693), .A2(n9939), .B1(n20793), .B2(n20662), .ZN(
        n20666) );
  AOI22_X1 U23639 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20664), .B1(
        n20663), .B2(n20735), .ZN(n20665) );
  OAI211_X1 U23640 ( .C1(n20668), .C2(n20667), .A(n20666), .B(n20665), .ZN(
        P1_U3136) );
  NOR2_X1 U23641 ( .A1(n20670), .A2(n20675), .ZN(n20691) );
  AOI21_X1 U23642 ( .B1(n20742), .B2(n20671), .A(n20691), .ZN(n20672) );
  OAI22_X1 U23643 ( .A1(n20672), .A2(n20747), .B1(n20675), .B2(n12749), .ZN(
        n20692) );
  AOI22_X1 U23644 ( .A1(n20744), .A2(n20691), .B1(n20743), .B2(n20692), .ZN(
        n20678) );
  INV_X1 U23645 ( .A(n20698), .ZN(n20746) );
  INV_X1 U23646 ( .A(n9811), .ZN(n20673) );
  NAND3_X1 U23647 ( .A1(n20746), .A2(n20673), .A3(n20885), .ZN(n20888) );
  AOI21_X1 U23648 ( .B1(n20675), .B2(n20888), .A(n20674), .ZN(n20676) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n9941), .ZN(n20677) );
  OAI211_X1 U23650 ( .C1(n20714), .C2(n20710), .A(n20678), .B(n20677), .ZN(
        P1_U3137) );
  AOI22_X1 U23651 ( .A1(n20757), .A2(n20691), .B1(n20756), .B2(n20692), .ZN(
        n20680) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n20758), .ZN(n20679) );
  OAI211_X1 U23653 ( .C1(n20761), .C2(n20710), .A(n20680), .B(n20679), .ZN(
        P1_U3138) );
  AOI22_X1 U23654 ( .A1(n20763), .A2(n20691), .B1(n20762), .B2(n20692), .ZN(
        n20682) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n20717), .ZN(n20681) );
  OAI211_X1 U23656 ( .C1(n20720), .C2(n20710), .A(n20682), .B(n20681), .ZN(
        P1_U3139) );
  AOI22_X1 U23657 ( .A1(n20769), .A2(n20691), .B1(n20768), .B2(n20692), .ZN(
        n20684) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n9943), .ZN(n20683) );
  OAI211_X1 U23659 ( .C1(n20773), .C2(n20710), .A(n20684), .B(n20683), .ZN(
        P1_U3140) );
  AOI22_X1 U23660 ( .A1(n20775), .A2(n20691), .B1(n20774), .B2(n20692), .ZN(
        n20686) );
  AOI22_X1 U23661 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n9945), .ZN(n20685) );
  OAI211_X1 U23662 ( .C1(n20726), .C2(n20710), .A(n20686), .B(n20685), .ZN(
        P1_U3141) );
  AOI22_X1 U23663 ( .A1(n20780), .A2(n20691), .B1(n20779), .B2(n20692), .ZN(
        n20688) );
  AOI22_X1 U23664 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n9947), .ZN(n20687) );
  OAI211_X1 U23665 ( .C1(n20730), .C2(n20710), .A(n20688), .B(n20687), .ZN(
        P1_U3142) );
  AOI22_X1 U23666 ( .A1(n20785), .A2(n20691), .B1(n20784), .B2(n20692), .ZN(
        n20690) );
  AOI22_X1 U23667 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n20786), .ZN(n20689) );
  OAI211_X1 U23668 ( .C1(n20791), .C2(n20710), .A(n20690), .B(n20689), .ZN(
        P1_U3143) );
  AOI22_X1 U23669 ( .A1(n20795), .A2(n20692), .B1(n20793), .B2(n20691), .ZN(
        n20696) );
  AOI22_X1 U23670 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20694), .B1(
        n20693), .B2(n20735), .ZN(n20695) );
  OAI211_X1 U23671 ( .C1(n9938), .C2(n20710), .A(n20696), .B(n20695), .ZN(
        P1_U3144) );
  INV_X1 U23672 ( .A(n20742), .ZN(n20701) );
  OAI33_X1 U23673 ( .A1(n20747), .A2(n20702), .A3(n20701), .B1(n20700), .B2(
        n20699), .B3(n20594), .ZN(n20734) );
  NOR2_X1 U23674 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20748), .ZN(
        n20733) );
  AOI22_X1 U23675 ( .A1(n9949), .A2(n20743), .B1(n20744), .B2(n20733), .ZN(
        n20713) );
  AOI21_X1 U23676 ( .B1(n20801), .B2(n20710), .A(n20703), .ZN(n20704) );
  AOI21_X1 U23677 ( .B1(n20742), .B2(n20705), .A(n20704), .ZN(n20706) );
  NOR2_X1 U23678 ( .A1(n20706), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20709) );
  AOI22_X1 U23679 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20737), .B1(
        n20736), .B2(n9941), .ZN(n20712) );
  OAI211_X1 U23680 ( .C1(n20714), .C2(n20801), .A(n20713), .B(n20712), .ZN(
        P1_U3145) );
  AOI22_X1 U23681 ( .A1(n9949), .A2(n20756), .B1(n20757), .B2(n20733), .ZN(
        n20716) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20737), .B1(
        n20736), .B2(n20758), .ZN(n20715) );
  OAI211_X1 U23683 ( .C1(n20761), .C2(n20801), .A(n20716), .B(n20715), .ZN(
        P1_U3146) );
  AOI22_X1 U23684 ( .A1(n9949), .A2(n20762), .B1(n20763), .B2(n20733), .ZN(
        n20719) );
  AOI22_X1 U23685 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20737), .B1(
        n20736), .B2(n20717), .ZN(n20718) );
  OAI211_X1 U23686 ( .C1(n20720), .C2(n20801), .A(n20719), .B(n20718), .ZN(
        P1_U3147) );
  AOI22_X1 U23687 ( .A1(n9949), .A2(n20768), .B1(n20769), .B2(n20733), .ZN(
        n20722) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20737), .B1(
        n20736), .B2(n9943), .ZN(n20721) );
  OAI211_X1 U23689 ( .C1(n20773), .C2(n20801), .A(n20722), .B(n20721), .ZN(
        P1_U3148) );
  AOI22_X1 U23690 ( .A1(n9949), .A2(n20774), .B1(n20775), .B2(n20733), .ZN(
        n20725) );
  AOI22_X1 U23691 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20737), .B1(
        n20736), .B2(n9945), .ZN(n20724) );
  OAI211_X1 U23692 ( .C1(n20726), .C2(n20801), .A(n20725), .B(n20724), .ZN(
        P1_U3149) );
  AOI22_X1 U23693 ( .A1(n9949), .A2(n20779), .B1(n20780), .B2(n20733), .ZN(
        n20729) );
  AOI22_X1 U23694 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20737), .B1(
        n20736), .B2(n9947), .ZN(n20728) );
  OAI211_X1 U23695 ( .C1(n20730), .C2(n20801), .A(n20729), .B(n20728), .ZN(
        P1_U3150) );
  AOI22_X1 U23696 ( .A1(n9949), .A2(n20784), .B1(n20785), .B2(n20733), .ZN(
        n20732) );
  AOI22_X1 U23697 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20737), .B1(
        n20736), .B2(n20786), .ZN(n20731) );
  OAI211_X1 U23698 ( .C1(n20791), .C2(n20801), .A(n20732), .B(n20731), .ZN(
        P1_U3151) );
  AOI22_X1 U23699 ( .A1(n9949), .A2(n20795), .B1(n20793), .B2(n20733), .ZN(
        n20739) );
  AOI22_X1 U23700 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20737), .B1(
        n20736), .B2(n20735), .ZN(n20738) );
  OAI211_X1 U23701 ( .C1(n9938), .C2(n20801), .A(n20739), .B(n20738), .ZN(
        P1_U3152) );
  INV_X1 U23702 ( .A(n20740), .ZN(n20792) );
  AOI21_X1 U23703 ( .B1(n20742), .B2(n20741), .A(n20792), .ZN(n20750) );
  OAI22_X1 U23704 ( .A1(n20750), .A2(n20747), .B1(n20748), .B2(n12749), .ZN(
        n20794) );
  AOI22_X1 U23705 ( .A1(n20744), .A2(n20792), .B1(n20743), .B2(n20794), .ZN(
        n20755) );
  OAI21_X1 U23706 ( .B1(n20746), .B2(n20747), .A(n20745), .ZN(n20749) );
  AOI22_X1 U23707 ( .A1(n20750), .A2(n20749), .B1(n20748), .B2(n20747), .ZN(
        n20751) );
  NAND2_X1 U23708 ( .A1(n20752), .A2(n20751), .ZN(n20798) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n20753), .ZN(n20754) );
  OAI211_X1 U23710 ( .C1(n9940), .C2(n20801), .A(n20755), .B(n20754), .ZN(
        P1_U3153) );
  AOI22_X1 U23711 ( .A1(n20757), .A2(n20792), .B1(n20756), .B2(n20794), .ZN(
        n20760) );
  INV_X1 U23712 ( .A(n20801), .ZN(n20787) );
  AOI22_X1 U23713 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20798), .B1(
        n20787), .B2(n20758), .ZN(n20759) );
  OAI211_X1 U23714 ( .C1(n20761), .C2(n20790), .A(n20760), .B(n20759), .ZN(
        P1_U3154) );
  AOI22_X1 U23715 ( .A1(n20763), .A2(n20792), .B1(n20762), .B2(n20794), .ZN(
        n20766) );
  AOI22_X1 U23716 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n20764), .ZN(n20765) );
  OAI211_X1 U23717 ( .C1(n20767), .C2(n20801), .A(n20766), .B(n20765), .ZN(
        P1_U3155) );
  AOI22_X1 U23718 ( .A1(n20769), .A2(n20792), .B1(n20768), .B2(n20794), .ZN(
        n20772) );
  AOI22_X1 U23719 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20798), .B1(
        n20787), .B2(n9943), .ZN(n20771) );
  OAI211_X1 U23720 ( .C1(n20773), .C2(n20790), .A(n20772), .B(n20771), .ZN(
        P1_U3156) );
  AOI22_X1 U23721 ( .A1(n20775), .A2(n20792), .B1(n20774), .B2(n20794), .ZN(
        n20778) );
  AOI22_X1 U23722 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n20776), .ZN(n20777) );
  OAI211_X1 U23723 ( .C1(n9944), .C2(n20801), .A(n20778), .B(n20777), .ZN(
        P1_U3157) );
  AOI22_X1 U23724 ( .A1(n20780), .A2(n20792), .B1(n20779), .B2(n20794), .ZN(
        n20783) );
  AOI22_X1 U23725 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n20781), .ZN(n20782) );
  OAI211_X1 U23726 ( .C1(n9946), .C2(n20801), .A(n20783), .B(n20782), .ZN(
        P1_U3158) );
  AOI22_X1 U23727 ( .A1(n20785), .A2(n20792), .B1(n20784), .B2(n20794), .ZN(
        n20789) );
  AOI22_X1 U23728 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20798), .B1(
        n20787), .B2(n20786), .ZN(n20788) );
  OAI211_X1 U23729 ( .C1(n20791), .C2(n20790), .A(n20789), .B(n20788), .ZN(
        P1_U3159) );
  AOI22_X1 U23730 ( .A1(n20795), .A2(n20794), .B1(n20793), .B2(n20792), .ZN(
        n20800) );
  AOI22_X1 U23731 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20798), .B1(
        n20797), .B2(n9939), .ZN(n20799) );
  OAI211_X1 U23732 ( .C1(n20802), .C2(n20801), .A(n20800), .B(n20799), .ZN(
        P1_U3160) );
  MUX2_X1 U23733 ( .A(n20804), .B(n20803), .S(n12749), .Z(P1_U3163) );
  AND2_X1 U23734 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20805), .ZN(
        P1_U3164) );
  AND2_X1 U23735 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20805), .ZN(
        P1_U3165) );
  AND2_X1 U23736 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20805), .ZN(
        P1_U3166) );
  AND2_X1 U23737 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20805), .ZN(
        P1_U3167) );
  AND2_X1 U23738 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20805), .ZN(
        P1_U3168) );
  AND2_X1 U23739 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20805), .ZN(
        P1_U3169) );
  AND2_X1 U23740 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20805), .ZN(
        P1_U3170) );
  AND2_X1 U23741 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20805), .ZN(
        P1_U3171) );
  AND2_X1 U23742 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20805), .ZN(
        P1_U3172) );
  AND2_X1 U23743 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20805), .ZN(
        P1_U3173) );
  AND2_X1 U23744 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20805), .ZN(
        P1_U3174) );
  AND2_X1 U23745 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20805), .ZN(
        P1_U3175) );
  AND2_X1 U23746 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20805), .ZN(
        P1_U3176) );
  AND2_X1 U23747 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20805), .ZN(
        P1_U3177) );
  AND2_X1 U23748 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20805), .ZN(
        P1_U3178) );
  AND2_X1 U23749 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20805), .ZN(
        P1_U3179) );
  AND2_X1 U23750 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20805), .ZN(
        P1_U3180) );
  AND2_X1 U23751 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20805), .ZN(
        P1_U3181) );
  AND2_X1 U23752 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20805), .ZN(
        P1_U3182) );
  AND2_X1 U23753 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20805), .ZN(
        P1_U3183) );
  AND2_X1 U23754 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20805), .ZN(
        P1_U3184) );
  AND2_X1 U23755 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20805), .ZN(
        P1_U3185) );
  AND2_X1 U23756 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20805), .ZN(P1_U3186) );
  AND2_X1 U23757 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20805), .ZN(P1_U3187) );
  AND2_X1 U23758 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20805), .ZN(P1_U3188) );
  AND2_X1 U23759 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20805), .ZN(P1_U3189) );
  AND2_X1 U23760 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20805), .ZN(P1_U3190) );
  AND2_X1 U23761 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20805), .ZN(P1_U3191) );
  AND2_X1 U23762 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20805), .ZN(P1_U3192) );
  AND2_X1 U23763 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20805), .ZN(P1_U3193) );
  AOI21_X1 U23764 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20811), .A(n20809), 
        .ZN(n20816) );
  NOR2_X1 U23765 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20806) );
  OAI22_X1 U23766 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21056), .B1(n20806), 
        .B2(n20819), .ZN(n20807) );
  NOR2_X1 U23767 ( .A1(n20999), .A2(n20807), .ZN(n20808) );
  OAI22_X1 U23768 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20816), .B1(n20912), 
        .B2(n20808), .ZN(P1_U3194) );
  NOR2_X1 U23769 ( .A1(NA), .A2(n20809), .ZN(n20812) );
  AOI21_X1 U23770 ( .B1(n20812), .B2(n20811), .A(n20810), .ZN(n20818) );
  AOI21_X1 U23771 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20812), .A(
        P1_STATE_REG_2__SCAN_IN), .ZN(n20815) );
  AND2_X1 U23772 ( .A1(n20813), .A2(NA), .ZN(n20814) );
  OAI33_X1 U23773 ( .A1(n20819), .A2(n20818), .A3(n20817), .B1(n20816), .B2(
        n20815), .B3(n20814), .ZN(P1_U3196) );
  OR2_X1 U23774 ( .A1(n20911), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20843) );
  NOR2_X1 U23775 ( .A1(n20820), .A2(n20911), .ZN(n20854) );
  INV_X1 U23776 ( .A(n20854), .ZN(n20841) );
  INV_X1 U23777 ( .A(n20841), .ZN(n20849) );
  AOI222_X1 U23778 ( .A1(n9806), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20849), .ZN(n20821) );
  INV_X1 U23779 ( .A(n20821), .ZN(P1_U3197) );
  AOI222_X1 U23780 ( .A1(n20854), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n9806), .ZN(n20822) );
  INV_X1 U23781 ( .A(n20822), .ZN(P1_U3198) );
  OAI222_X1 U23782 ( .A1(n20841), .A2(n13415), .B1(n20824), .B2(n20912), .C1(
        n20823), .C2(n20843), .ZN(P1_U3199) );
  AOI222_X1 U23783 ( .A1(n20849), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n9806), .ZN(n20825) );
  INV_X1 U23784 ( .A(n20825), .ZN(P1_U3200) );
  AOI222_X1 U23785 ( .A1(n20854), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n9806), .ZN(n20826) );
  INV_X1 U23786 ( .A(n20826), .ZN(P1_U3201) );
  AOI222_X1 U23787 ( .A1(n9806), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20849), .ZN(n20827) );
  INV_X1 U23788 ( .A(n20827), .ZN(P1_U3202) );
  AOI222_X1 U23789 ( .A1(n9806), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20849), .ZN(n20828) );
  INV_X1 U23790 ( .A(n20828), .ZN(P1_U3203) );
  AOI222_X1 U23791 ( .A1(n20849), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n9806), .ZN(n20829) );
  INV_X1 U23792 ( .A(n20829), .ZN(P1_U3204) );
  AOI222_X1 U23793 ( .A1(n20854), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n9806), .ZN(n20830) );
  INV_X1 U23794 ( .A(n20830), .ZN(P1_U3205) );
  AOI222_X1 U23795 ( .A1(n20849), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n9806), .ZN(n20831) );
  INV_X1 U23796 ( .A(n20831), .ZN(P1_U3206) );
  AOI222_X1 U23797 ( .A1(n20849), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n9806), .ZN(n20832) );
  INV_X1 U23798 ( .A(n20832), .ZN(P1_U3207) );
  AOI222_X1 U23799 ( .A1(n9806), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20849), .ZN(n20833) );
  INV_X1 U23800 ( .A(n20833), .ZN(P1_U3208) );
  AOI222_X1 U23801 ( .A1(n9806), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20849), .ZN(n20834) );
  INV_X1 U23802 ( .A(n20834), .ZN(P1_U3209) );
  AOI222_X1 U23803 ( .A1(n9806), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20849), .ZN(n20835) );
  INV_X1 U23804 ( .A(n20835), .ZN(P1_U3210) );
  AOI222_X1 U23805 ( .A1(n9806), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20849), .ZN(n20836) );
  INV_X1 U23806 ( .A(n20836), .ZN(P1_U3211) );
  AOI222_X1 U23807 ( .A1(n20849), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n9806), .ZN(n20837) );
  INV_X1 U23808 ( .A(n20837), .ZN(P1_U3212) );
  AOI222_X1 U23809 ( .A1(n9806), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20849), .ZN(n20838) );
  INV_X1 U23810 ( .A(n20838), .ZN(P1_U3213) );
  AOI222_X1 U23811 ( .A1(n20849), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n9806), .ZN(n20839) );
  INV_X1 U23812 ( .A(n20839), .ZN(P1_U3214) );
  AOI22_X1 U23813 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20911), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n9806), .ZN(n20840) );
  OAI21_X1 U23814 ( .B1(n21024), .B2(n20841), .A(n20840), .ZN(P1_U3215) );
  AOI22_X1 U23815 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20911), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20854), .ZN(n20842) );
  OAI21_X1 U23816 ( .B1(n21288), .B2(n20843), .A(n20842), .ZN(P1_U3216) );
  AOI222_X1 U23817 ( .A1(n9806), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20849), .ZN(n20844) );
  INV_X1 U23818 ( .A(n20844), .ZN(P1_U3217) );
  AOI222_X1 U23819 ( .A1(n20849), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n9806), .ZN(n20845) );
  INV_X1 U23820 ( .A(n20845), .ZN(P1_U3218) );
  AOI222_X1 U23821 ( .A1(n9806), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20849), .ZN(n20846) );
  INV_X1 U23822 ( .A(n20846), .ZN(P1_U3219) );
  AOI222_X1 U23823 ( .A1(n9806), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20854), .ZN(n20847) );
  INV_X1 U23824 ( .A(n20847), .ZN(P1_U3220) );
  AOI222_X1 U23825 ( .A1(n20854), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n9806), .ZN(n20848) );
  INV_X1 U23826 ( .A(n20848), .ZN(P1_U3221) );
  AOI222_X1 U23827 ( .A1(n9806), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20849), .ZN(n20850) );
  INV_X1 U23828 ( .A(n20850), .ZN(P1_U3222) );
  AOI222_X1 U23829 ( .A1(n20854), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n9806), .ZN(n20851) );
  INV_X1 U23830 ( .A(n20851), .ZN(P1_U3223) );
  AOI222_X1 U23831 ( .A1(n9806), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20854), .ZN(n20852) );
  INV_X1 U23832 ( .A(n20852), .ZN(P1_U3224) );
  AOI222_X1 U23833 ( .A1(n9806), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20854), .ZN(n20853) );
  INV_X1 U23834 ( .A(n20853), .ZN(P1_U3225) );
  AOI222_X1 U23835 ( .A1(n20854), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20911), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n9806), .ZN(n20855) );
  INV_X1 U23836 ( .A(n20855), .ZN(P1_U3226) );
  OAI22_X1 U23837 ( .A1(n20911), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20912), .ZN(n20856) );
  INV_X1 U23838 ( .A(n20856), .ZN(P1_U3458) );
  OAI22_X1 U23839 ( .A1(n20911), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20912), .ZN(n20857) );
  INV_X1 U23840 ( .A(n20857), .ZN(P1_U3459) );
  OAI22_X1 U23841 ( .A1(n20911), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20912), .ZN(n20858) );
  INV_X1 U23842 ( .A(n20858), .ZN(P1_U3460) );
  OAI22_X1 U23843 ( .A1(n20911), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20912), .ZN(n20859) );
  INV_X1 U23844 ( .A(n20859), .ZN(P1_U3461) );
  OAI21_X1 U23845 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20863), .A(n20861), 
        .ZN(n20860) );
  INV_X1 U23846 ( .A(n20860), .ZN(P1_U3464) );
  OAI21_X1 U23847 ( .B1(n20863), .B2(n20862), .A(n20861), .ZN(P1_U3465) );
  INV_X1 U23848 ( .A(n20864), .ZN(n20866) );
  OAI22_X1 U23849 ( .A1(n20866), .A2(n20871), .B1(n20865), .B2(n20875), .ZN(
        n20867) );
  MUX2_X1 U23850 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20867), .S(
        n20878), .Z(P1_U3469) );
  INV_X1 U23851 ( .A(n20868), .ZN(n20873) );
  INV_X1 U23852 ( .A(n20869), .ZN(n20870) );
  OAI222_X1 U23853 ( .A1(n20875), .A2(n20874), .B1(n20873), .B2(n20872), .C1(
        n20871), .C2(n20870), .ZN(n20877) );
  OAI22_X1 U23854 ( .A1(n20878), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20877), .B2(n20876), .ZN(n20879) );
  INV_X1 U23855 ( .A(n20879), .ZN(P1_U3472) );
  OAI22_X1 U23856 ( .A1(n20883), .A2(n20882), .B1(n20881), .B2(n20880), .ZN(
        n20884) );
  AOI21_X1 U23857 ( .B1(n20886), .B2(n20885), .A(n20884), .ZN(n20889) );
  NAND3_X1 U23858 ( .A1(n20889), .A2(n20888), .A3(n20887), .ZN(n20890) );
  NAND2_X1 U23859 ( .A1(n20892), .A2(n20890), .ZN(n20891) );
  OAI21_X1 U23860 ( .B1(n20892), .B2(n20594), .A(n20891), .ZN(P1_U3475) );
  AOI21_X1 U23861 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20893) );
  AOI22_X1 U23862 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20893), .B2(n21013), .ZN(n20895) );
  INV_X1 U23863 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20894) );
  AOI22_X1 U23864 ( .A1(n20896), .A2(n20895), .B1(n20894), .B2(n20898), .ZN(
        P1_U3481) );
  INV_X1 U23865 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20899) );
  NOR2_X1 U23866 ( .A1(n20898), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20897) );
  AOI22_X1 U23867 ( .A1(n20899), .A2(n20898), .B1(n21207), .B2(n20897), .ZN(
        P1_U3482) );
  AOI22_X1 U23868 ( .A1(n20912), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21178), 
        .B2(n20911), .ZN(P1_U3483) );
  AOI211_X1 U23869 ( .C1(n20210), .C2(n20902), .A(n20901), .B(n20900), .ZN(
        n20910) );
  INV_X1 U23870 ( .A(n20903), .ZN(n20904) );
  OAI211_X1 U23871 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20905), .A(n20904), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20907) );
  AOI21_X1 U23872 ( .B1(n20907), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20906), 
        .ZN(n20909) );
  NAND2_X1 U23873 ( .A1(n20910), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20908) );
  OAI21_X1 U23874 ( .B1(n20910), .B2(n20909), .A(n20908), .ZN(P1_U3485) );
  AOI22_X1 U23875 ( .A1(n20912), .A2(n21225), .B1(n21282), .B2(n20911), .ZN(
        P1_U3486) );
  AOI22_X1 U23876 ( .A1(n16743), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16745), .ZN(n21303) );
  OAI22_X1 U23877 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(keyinput_g100), .B1(
        keyinput_g15), .B2(DATAI_17_), .ZN(n20913) );
  AOI221_X1 U23878 ( .B1(P1_EBX_REG_15__SCAN_IN), .B2(keyinput_g100), .C1(
        DATAI_17_), .C2(keyinput_g15), .A(n20913), .ZN(n20920) );
  OAI22_X1 U23879 ( .A1(DATAI_21_), .A2(keyinput_g11), .B1(keyinput_g33), .B2(
        HOLD), .ZN(n20914) );
  AOI221_X1 U23880 ( .B1(DATAI_21_), .B2(keyinput_g11), .C1(HOLD), .C2(
        keyinput_g33), .A(n20914), .ZN(n20919) );
  OAI22_X1 U23881 ( .A1(P1_EBX_REG_24__SCAN_IN), .A2(keyinput_g91), .B1(
        DATAI_3_), .B2(keyinput_g29), .ZN(n20915) );
  AOI221_X1 U23882 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(keyinput_g91), .C1(
        keyinput_g29), .C2(DATAI_3_), .A(n20915), .ZN(n20918) );
  OAI22_X1 U23883 ( .A1(DATAI_18_), .A2(keyinput_g14), .B1(DATAI_2_), .B2(
        keyinput_g30), .ZN(n20916) );
  AOI221_X1 U23884 ( .B1(DATAI_18_), .B2(keyinput_g14), .C1(keyinput_g30), 
        .C2(DATAI_2_), .A(n20916), .ZN(n20917) );
  NAND4_X1 U23885 ( .A1(n20920), .A2(n20919), .A3(n20918), .A4(n20917), .ZN(
        n20948) );
  OAI22_X1 U23886 ( .A1(READY1), .A2(keyinput_g36), .B1(P1_EBX_REG_21__SCAN_IN), .B2(keyinput_g94), .ZN(n20921) );
  AOI221_X1 U23887 ( .B1(READY1), .B2(keyinput_g36), .C1(keyinput_g94), .C2(
        P1_EBX_REG_21__SCAN_IN), .A(n20921), .ZN(n20928) );
  OAI22_X1 U23888 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(keyinput_g55), .B1(
        keyinput_g3), .B2(DATAI_29_), .ZN(n20922) );
  AOI221_X1 U23889 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_g55), .C1(
        DATAI_29_), .C2(keyinput_g3), .A(n20922), .ZN(n20927) );
  OAI22_X1 U23890 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(keyinput_g106), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .ZN(n20923) );
  AOI221_X1 U23891 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(keyinput_g106), .C1(
        keyinput_g63), .C2(P1_REIP_REG_20__SCAN_IN), .A(n20923), .ZN(n20926)
         );
  OAI22_X1 U23892 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput_g75), .B1(
        keyinput_g60), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n20924) );
  AOI221_X1 U23893 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput_g75), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_g60), .A(n20924), .ZN(n20925)
         );
  NAND4_X1 U23894 ( .A1(n20928), .A2(n20927), .A3(n20926), .A4(n20925), .ZN(
        n20947) );
  OAI22_X1 U23895 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_g123), .B1(
        keyinput_g118), .B2(P1_EAX_REG_29__SCAN_IN), .ZN(n20929) );
  AOI221_X1 U23896 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_g123), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput_g118), .A(n20929), .ZN(n20936)
         );
  OAI22_X1 U23897 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_g65), .B1(
        keyinput_g49), .B2(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20930) );
  AOI221_X1 U23898 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(keyinput_g65), .C1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_g49), .A(n20930), .ZN(
        n20935) );
  OAI22_X1 U23899 ( .A1(P1_EAX_REG_23__SCAN_IN), .A2(keyinput_g124), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_g58), .ZN(n20931) );
  AOI221_X1 U23900 ( .B1(P1_EAX_REG_23__SCAN_IN), .B2(keyinput_g124), .C1(
        keyinput_g58), .C2(P1_REIP_REG_25__SCAN_IN), .A(n20931), .ZN(n20934)
         );
  OAI22_X1 U23901 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(keyinput_g79), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_g61), .ZN(n20932) );
  AOI221_X1 U23902 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(keyinput_g79), .C1(
        keyinput_g61), .C2(P1_REIP_REG_22__SCAN_IN), .A(n20932), .ZN(n20933)
         );
  NAND4_X1 U23903 ( .A1(n20936), .A2(n20935), .A3(n20934), .A4(n20933), .ZN(
        n20946) );
  OAI22_X1 U23904 ( .A1(P1_EBX_REG_29__SCAN_IN), .A2(keyinput_g86), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(keyinput_g70), .ZN(n20937) );
  AOI221_X1 U23905 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(keyinput_g86), .C1(
        keyinput_g70), .C2(P1_REIP_REG_13__SCAN_IN), .A(n20937), .ZN(n20944)
         );
  OAI22_X1 U23906 ( .A1(P1_EBX_REG_4__SCAN_IN), .A2(keyinput_g111), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .ZN(n20938) );
  AOI221_X1 U23907 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(keyinput_g111), .C1(
        keyinput_g57), .C2(P1_REIP_REG_26__SCAN_IN), .A(n20938), .ZN(n20943)
         );
  OAI22_X1 U23908 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(keyinput_g96), .B1(
        keyinput_g76), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n20939) );
  AOI221_X1 U23909 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(keyinput_g96), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(keyinput_g76), .A(n20939), .ZN(n20942) );
  OAI22_X1 U23910 ( .A1(DATAI_0_), .A2(keyinput_g32), .B1(
        P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_g40), .ZN(n20940) );
  AOI221_X1 U23911 ( .B1(DATAI_0_), .B2(keyinput_g32), .C1(keyinput_g40), .C2(
        P1_CODEFETCH_REG_SCAN_IN), .A(n20940), .ZN(n20941) );
  NAND4_X1 U23912 ( .A1(n20944), .A2(n20943), .A3(n20942), .A4(n20941), .ZN(
        n20945) );
  NOR4_X1 U23913 ( .A1(n20948), .A2(n20947), .A3(n20946), .A4(n20945), .ZN(
        n21087) );
  OAI22_X1 U23914 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(keyinput_g101), .B1(
        DATAI_4_), .B2(keyinput_g28), .ZN(n20949) );
  AOI221_X1 U23915 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(keyinput_g101), .C1(
        keyinput_g28), .C2(DATAI_4_), .A(n20949), .ZN(n20956) );
  OAI22_X1 U23916 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(keyinput_g104), .B1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g48), .ZN(n20950) );
  AOI221_X1 U23917 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput_g104), .C1(
        keyinput_g48), .C2(P1_BYTEENABLE_REG_0__SCAN_IN), .A(n20950), .ZN(
        n20955) );
  OAI22_X1 U23918 ( .A1(P1_EAX_REG_25__SCAN_IN), .A2(keyinput_g122), .B1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g50), .ZN(n20951) );
  AOI221_X1 U23919 ( .B1(P1_EAX_REG_25__SCAN_IN), .B2(keyinput_g122), .C1(
        keyinput_g50), .C2(P1_BYTEENABLE_REG_2__SCAN_IN), .A(n20951), .ZN(
        n20954) );
  OAI22_X1 U23920 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(keyinput_g113), .B1(
        DATAI_30_), .B2(keyinput_g2), .ZN(n20952) );
  AOI221_X1 U23921 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(keyinput_g113), .C1(
        keyinput_g2), .C2(DATAI_30_), .A(n20952), .ZN(n20953) );
  NAND4_X1 U23922 ( .A1(n20956), .A2(n20955), .A3(n20954), .A4(n20953), .ZN(
        n21085) );
  OAI22_X1 U23923 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(keyinput_g116), .B1(
        keyinput_g13), .B2(DATAI_19_), .ZN(n20957) );
  AOI221_X1 U23924 ( .B1(P1_EAX_REG_31__SCAN_IN), .B2(keyinput_g116), .C1(
        DATAI_19_), .C2(keyinput_g13), .A(n20957), .ZN(n20983) );
  OAI22_X1 U23925 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(keyinput_g114), .B1(
        keyinput_g16), .B2(DATAI_16_), .ZN(n20958) );
  AOI221_X1 U23926 ( .B1(P1_EBX_REG_1__SCAN_IN), .B2(keyinput_g114), .C1(
        DATAI_16_), .C2(keyinput_g16), .A(n20958), .ZN(n20961) );
  OAI22_X1 U23927 ( .A1(P1_EAX_REG_30__SCAN_IN), .A2(keyinput_g117), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(keyinput_g53), .ZN(n20959) );
  AOI221_X1 U23928 ( .B1(P1_EAX_REG_30__SCAN_IN), .B2(keyinput_g117), .C1(
        keyinput_g53), .C2(P1_REIP_REG_30__SCAN_IN), .A(n20959), .ZN(n20960)
         );
  OAI211_X1 U23929 ( .C1(n20963), .C2(keyinput_g69), .A(n20961), .B(n20960), 
        .ZN(n20962) );
  AOI21_X1 U23930 ( .B1(n20963), .B2(keyinput_g69), .A(n20962), .ZN(n20982) );
  AOI22_X1 U23931 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput_g38), .B1(
        DATAI_12_), .B2(keyinput_g20), .ZN(n20964) );
  OAI221_X1 U23932 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_g38), .C1(
        DATAI_12_), .C2(keyinput_g20), .A(n20964), .ZN(n20971) );
  AOI22_X1 U23933 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput_g67), .B1(
        P1_EBX_REG_22__SCAN_IN), .B2(keyinput_g93), .ZN(n20965) );
  OAI221_X1 U23934 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(keyinput_g67), .C1(
        P1_EBX_REG_22__SCAN_IN), .C2(keyinput_g93), .A(n20965), .ZN(n20970) );
  AOI22_X1 U23935 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P1_FLUSH_REG_SCAN_IN), .B2(keyinput_g46), .ZN(n20966) );
  OAI221_X1 U23936 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P1_FLUSH_REG_SCAN_IN), .C2(keyinput_g46), .A(n20966), .ZN(n20969) );
  AOI22_X1 U23937 ( .A1(P1_EBX_REG_30__SCAN_IN), .A2(keyinput_g85), .B1(
        P1_EBX_REG_23__SCAN_IN), .B2(keyinput_g92), .ZN(n20967) );
  OAI221_X1 U23938 ( .B1(P1_EBX_REG_30__SCAN_IN), .B2(keyinput_g85), .C1(
        P1_EBX_REG_23__SCAN_IN), .C2(keyinput_g92), .A(n20967), .ZN(n20968) );
  NOR4_X1 U23939 ( .A1(n20971), .A2(n20970), .A3(n20969), .A4(n20968), .ZN(
        n20981) );
  AOI22_X1 U23940 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(keyinput_g56), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(keyinput_g74), .ZN(n20972) );
  OAI221_X1 U23941 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(keyinput_g56), .C1(
        P1_REIP_REG_9__SCAN_IN), .C2(keyinput_g74), .A(n20972), .ZN(n20979) );
  AOI22_X1 U23942 ( .A1(DATAI_7_), .A2(keyinput_g25), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(keyinput_g71), .ZN(n20973) );
  OAI221_X1 U23943 ( .B1(DATAI_7_), .B2(keyinput_g25), .C1(
        P1_REIP_REG_12__SCAN_IN), .C2(keyinput_g71), .A(n20973), .ZN(n20978)
         );
  AOI22_X1 U23944 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(keyinput_g99), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(keyinput_g126), .ZN(n20974) );
  OAI221_X1 U23945 ( .B1(P1_EBX_REG_16__SCAN_IN), .B2(keyinput_g99), .C1(
        P1_EAX_REG_21__SCAN_IN), .C2(keyinput_g126), .A(n20974), .ZN(n20977)
         );
  AOI22_X1 U23946 ( .A1(READY2), .A2(keyinput_g37), .B1(P1_REIP_REG_2__SCAN_IN), .B2(keyinput_g81), .ZN(n20975) );
  OAI221_X1 U23947 ( .B1(READY2), .B2(keyinput_g37), .C1(
        P1_REIP_REG_2__SCAN_IN), .C2(keyinput_g81), .A(n20975), .ZN(n20976) );
  NOR4_X1 U23948 ( .A1(n20979), .A2(n20978), .A3(n20977), .A4(n20976), .ZN(
        n20980) );
  NAND4_X1 U23949 ( .A1(n20983), .A2(n20982), .A3(n20981), .A4(n20980), .ZN(
        n21084) );
  AOI22_X1 U23950 ( .A1(DATAI_10_), .A2(keyinput_g22), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(keyinput_g121), .ZN(n20984) );
  OAI221_X1 U23951 ( .B1(DATAI_10_), .B2(keyinput_g22), .C1(
        P1_EAX_REG_26__SCAN_IN), .C2(keyinput_g121), .A(n20984), .ZN(n20993)
         );
  AOI22_X1 U23952 ( .A1(DATAI_20_), .A2(keyinput_g12), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_g44), .ZN(n20985) );
  OAI221_X1 U23953 ( .B1(DATAI_20_), .B2(keyinput_g12), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_g44), .A(n20985), .ZN(n20992)
         );
  AOI22_X1 U23954 ( .A1(DATAI_23_), .A2(keyinput_g9), .B1(
        P1_EBX_REG_12__SCAN_IN), .B2(keyinput_g103), .ZN(n20986) );
  OAI221_X1 U23955 ( .B1(DATAI_23_), .B2(keyinput_g9), .C1(
        P1_EBX_REG_12__SCAN_IN), .C2(keyinput_g103), .A(n20986), .ZN(n20991)
         );
  AOI22_X1 U23956 ( .A1(n20989), .A2(keyinput_g18), .B1(n20988), .B2(
        keyinput_g54), .ZN(n20987) );
  OAI221_X1 U23957 ( .B1(n20989), .B2(keyinput_g18), .C1(n20988), .C2(
        keyinput_g54), .A(n20987), .ZN(n20990) );
  NOR4_X1 U23958 ( .A1(n20993), .A2(n20992), .A3(n20991), .A4(n20990), .ZN(
        n21032) );
  AOI22_X1 U23959 ( .A1(n21196), .A2(keyinput_g23), .B1(n20995), .B2(
        keyinput_g112), .ZN(n20994) );
  OAI221_X1 U23960 ( .B1(n21196), .B2(keyinput_g23), .C1(n20995), .C2(
        keyinput_g112), .A(n20994), .ZN(n21006) );
  AOI22_X1 U23961 ( .A1(n20997), .A2(keyinput_g115), .B1(keyinput_g80), .B2(
        n13415), .ZN(n20996) );
  OAI221_X1 U23962 ( .B1(n20997), .B2(keyinput_g115), .C1(n13415), .C2(
        keyinput_g80), .A(n20996), .ZN(n21005) );
  AOI22_X1 U23963 ( .A1(n21165), .A2(keyinput_g97), .B1(keyinput_g43), .B2(
        n20999), .ZN(n20998) );
  OAI221_X1 U23964 ( .B1(n21165), .B2(keyinput_g97), .C1(n20999), .C2(
        keyinput_g43), .A(n20998), .ZN(n21004) );
  AOI22_X1 U23965 ( .A1(n21002), .A2(keyinput_g1), .B1(keyinput_g10), .B2(
        n21001), .ZN(n21000) );
  OAI221_X1 U23966 ( .B1(n21002), .B2(keyinput_g1), .C1(n21001), .C2(
        keyinput_g10), .A(n21000), .ZN(n21003) );
  NOR4_X1 U23967 ( .A1(n21006), .A2(n21005), .A3(n21004), .A4(n21003), .ZN(
        n21031) );
  INV_X1 U23968 ( .A(DATAI_1_), .ZN(n21156) );
  AOI22_X1 U23969 ( .A1(n21175), .A2(keyinput_g88), .B1(keyinput_g31), .B2(
        n21156), .ZN(n21007) );
  OAI221_X1 U23970 ( .B1(n21175), .B2(keyinput_g88), .C1(n21156), .C2(
        keyinput_g31), .A(n21007), .ZN(n21017) );
  AOI22_X1 U23971 ( .A1(n21009), .A2(keyinput_g87), .B1(keyinput_g27), .B2(
        n12538), .ZN(n21008) );
  OAI221_X1 U23972 ( .B1(n21009), .B2(keyinput_g87), .C1(n12538), .C2(
        keyinput_g27), .A(n21008), .ZN(n21016) );
  INV_X1 U23973 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21011) );
  AOI22_X1 U23974 ( .A1(n21146), .A2(keyinput_g5), .B1(n21011), .B2(
        keyinput_g109), .ZN(n21010) );
  OAI221_X1 U23975 ( .B1(n21146), .B2(keyinput_g5), .C1(n21011), .C2(
        keyinput_g109), .A(n21010), .ZN(n21015) );
  AOI22_X1 U23976 ( .A1(n21013), .A2(keyinput_g82), .B1(n21239), .B2(
        keyinput_g107), .ZN(n21012) );
  OAI221_X1 U23977 ( .B1(n21013), .B2(keyinput_g82), .C1(n21239), .C2(
        keyinput_g107), .A(n21012), .ZN(n21014) );
  NOR4_X1 U23978 ( .A1(n21017), .A2(n21016), .A3(n21015), .A4(n21014), .ZN(
        n21030) );
  AOI22_X1 U23979 ( .A1(n21177), .A2(keyinput_g59), .B1(keyinput_g83), .B2(
        n21207), .ZN(n21018) );
  OAI221_X1 U23980 ( .B1(n21177), .B2(keyinput_g59), .C1(n21207), .C2(
        keyinput_g83), .A(n21018), .ZN(n21028) );
  AOI22_X1 U23981 ( .A1(n21235), .A2(keyinput_g90), .B1(keyinput_g39), .B2(
        n21130), .ZN(n21019) );
  OAI221_X1 U23982 ( .B1(n21235), .B2(keyinput_g90), .C1(n21130), .C2(
        keyinput_g39), .A(n21019), .ZN(n21027) );
  AOI22_X1 U23983 ( .A1(n21162), .A2(keyinput_g78), .B1(keyinput_g19), .B2(
        n21021), .ZN(n21020) );
  OAI221_X1 U23984 ( .B1(n21162), .B2(keyinput_g78), .C1(n21021), .C2(
        keyinput_g19), .A(n21020), .ZN(n21026) );
  AOI22_X1 U23985 ( .A1(n21024), .A2(keyinput_g64), .B1(n21023), .B2(
        keyinput_g120), .ZN(n21022) );
  OAI221_X1 U23986 ( .B1(n21024), .B2(keyinput_g64), .C1(n21023), .C2(
        keyinput_g120), .A(n21022), .ZN(n21025) );
  NOR4_X1 U23987 ( .A1(n21028), .A2(n21027), .A3(n21026), .A4(n21025), .ZN(
        n21029) );
  NAND4_X1 U23988 ( .A1(n21032), .A2(n21031), .A3(n21030), .A4(n21029), .ZN(
        n21083) );
  AOI22_X1 U23989 ( .A1(n21034), .A2(keyinput_g108), .B1(keyinput_g26), .B2(
        n12523), .ZN(n21033) );
  OAI221_X1 U23990 ( .B1(n21034), .B2(keyinput_g108), .C1(n12523), .C2(
        keyinput_g26), .A(n21033), .ZN(n21044) );
  AOI22_X1 U23991 ( .A1(n21242), .A2(keyinput_g45), .B1(n21172), .B2(
        keyinput_g8), .ZN(n21035) );
  OAI221_X1 U23992 ( .B1(n21242), .B2(keyinput_g45), .C1(n21172), .C2(
        keyinput_g8), .A(n21035), .ZN(n21043) );
  AOI22_X1 U23993 ( .A1(n21037), .A2(keyinput_g84), .B1(keyinput_g6), .B2(
        n21124), .ZN(n21036) );
  OAI221_X1 U23994 ( .B1(n21037), .B2(keyinput_g84), .C1(n21124), .C2(
        keyinput_g6), .A(n21036), .ZN(n21042) );
  AOI22_X1 U23995 ( .A1(n21040), .A2(keyinput_g72), .B1(n21039), .B2(
        keyinput_g105), .ZN(n21038) );
  OAI221_X1 U23996 ( .B1(n21040), .B2(keyinput_g72), .C1(n21039), .C2(
        keyinput_g105), .A(n21038), .ZN(n21041) );
  NOR4_X1 U23997 ( .A1(n21044), .A2(n21043), .A3(n21042), .A4(n21041), .ZN(
        n21081) );
  AOI22_X1 U23998 ( .A1(n12622), .A2(keyinput_g17), .B1(n21215), .B2(
        keyinput_g77), .ZN(n21045) );
  OAI221_X1 U23999 ( .B1(n12622), .B2(keyinput_g17), .C1(n21215), .C2(
        keyinput_g77), .A(n21045), .ZN(n21054) );
  AOI22_X1 U24000 ( .A1(n21243), .A2(keyinput_g21), .B1(keyinput_g51), .B2(
        n21190), .ZN(n21046) );
  OAI221_X1 U24001 ( .B1(n21243), .B2(keyinput_g21), .C1(n21190), .C2(
        keyinput_g51), .A(n21046), .ZN(n21053) );
  AOI22_X1 U24002 ( .A1(n21191), .A2(keyinput_g125), .B1(keyinput_g73), .B2(
        n21048), .ZN(n21047) );
  OAI221_X1 U24003 ( .B1(n21191), .B2(keyinput_g125), .C1(n21048), .C2(
        keyinput_g73), .A(n21047), .ZN(n21052) );
  INV_X1 U24004 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n21143) );
  AOI22_X1 U24005 ( .A1(n21050), .A2(keyinput_g4), .B1(n21143), .B2(
        keyinput_g102), .ZN(n21049) );
  OAI221_X1 U24006 ( .B1(n21050), .B2(keyinput_g4), .C1(n21143), .C2(
        keyinput_g102), .A(n21049), .ZN(n21051) );
  NOR4_X1 U24007 ( .A1(n21054), .A2(n21053), .A3(n21052), .A4(n21051), .ZN(
        n21080) );
  AOI22_X1 U24008 ( .A1(n21194), .A2(keyinput_g24), .B1(keyinput_g34), .B2(
        n21056), .ZN(n21055) );
  OAI221_X1 U24009 ( .B1(n21194), .B2(keyinput_g24), .C1(n21056), .C2(
        keyinput_g34), .A(n21055), .ZN(n21066) );
  AOI22_X1 U24010 ( .A1(n21058), .A2(keyinput_g68), .B1(keyinput_g41), .B2(
        n21282), .ZN(n21057) );
  OAI221_X1 U24011 ( .B1(n21058), .B2(keyinput_g68), .C1(n21282), .C2(
        keyinput_g41), .A(n21057), .ZN(n21065) );
  INV_X1 U24012 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n21060) );
  AOI22_X1 U24013 ( .A1(n21061), .A2(keyinput_g7), .B1(n21060), .B2(
        keyinput_g110), .ZN(n21059) );
  OAI221_X1 U24014 ( .B1(n21061), .B2(keyinput_g7), .C1(n21060), .C2(
        keyinput_g110), .A(n21059), .ZN(n21064) );
  AOI22_X1 U24015 ( .A1(n21222), .A2(keyinput_g98), .B1(keyinput_g47), .B2(
        n21178), .ZN(n21062) );
  OAI221_X1 U24016 ( .B1(n21222), .B2(keyinput_g98), .C1(n21178), .C2(
        keyinput_g47), .A(n21062), .ZN(n21063) );
  NOR4_X1 U24017 ( .A1(n21066), .A2(n21065), .A3(n21064), .A4(n21063), .ZN(
        n21079) );
  AOI22_X1 U24018 ( .A1(n21180), .A2(keyinput_g95), .B1(n21068), .B2(
        keyinput_g119), .ZN(n21067) );
  OAI221_X1 U24019 ( .B1(n21180), .B2(keyinput_g95), .C1(n21068), .C2(
        keyinput_g119), .A(n21067), .ZN(n21077) );
  INV_X1 U24020 ( .A(BS16), .ZN(n21070) );
  AOI22_X1 U24021 ( .A1(n21070), .A2(keyinput_g35), .B1(n21210), .B2(
        keyinput_g66), .ZN(n21069) );
  OAI221_X1 U24022 ( .B1(n21070), .B2(keyinput_g35), .C1(n21210), .C2(
        keyinput_g66), .A(n21069), .ZN(n21076) );
  AOI22_X1 U24023 ( .A1(n21072), .A2(keyinput_g89), .B1(n21155), .B2(
        keyinput_g127), .ZN(n21071) );
  OAI221_X1 U24024 ( .B1(n21072), .B2(keyinput_g89), .C1(n21155), .C2(
        keyinput_g127), .A(n21071), .ZN(n21075) );
  AOI22_X1 U24025 ( .A1(n21288), .A2(keyinput_g62), .B1(n21285), .B2(
        keyinput_g52), .ZN(n21073) );
  OAI221_X1 U24026 ( .B1(n21288), .B2(keyinput_g62), .C1(n21285), .C2(
        keyinput_g52), .A(n21073), .ZN(n21074) );
  NOR4_X1 U24027 ( .A1(n21077), .A2(n21076), .A3(n21075), .A4(n21074), .ZN(
        n21078) );
  NAND4_X1 U24028 ( .A1(n21081), .A2(n21080), .A3(n21079), .A4(n21078), .ZN(
        n21082) );
  NOR4_X1 U24029 ( .A1(n21085), .A2(n21084), .A3(n21083), .A4(n21082), .ZN(
        n21086) );
  AOI22_X1 U24030 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_g42), .B1(n21087), 
        .B2(n21086), .ZN(n21301) );
  OAI22_X1 U24031 ( .A1(P1_EBX_REG_28__SCAN_IN), .A2(keyinput_f87), .B1(
        keyinput_f113), .B2(P1_EBX_REG_2__SCAN_IN), .ZN(n21088) );
  AOI221_X1 U24032 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(keyinput_f87), .C1(
        P1_EBX_REG_2__SCAN_IN), .C2(keyinput_f113), .A(n21088), .ZN(n21095) );
  OAI22_X1 U24033 ( .A1(DATAI_31_), .A2(keyinput_f1), .B1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_f50), .ZN(n21089) );
  AOI221_X1 U24034 ( .B1(DATAI_31_), .B2(keyinput_f1), .C1(keyinput_f50), .C2(
        P1_BYTEENABLE_REG_2__SCAN_IN), .A(n21089), .ZN(n21094) );
  OAI22_X1 U24035 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(keyinput_f109), .B1(HOLD), 
        .B2(keyinput_f33), .ZN(n21090) );
  AOI221_X1 U24036 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(keyinput_f109), .C1(
        keyinput_f33), .C2(HOLD), .A(n21090), .ZN(n21093) );
  OAI22_X1 U24037 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_f123), .B1(
        keyinput_f70), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n21091) );
  AOI221_X1 U24038 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_f123), .C1(
        P1_REIP_REG_13__SCAN_IN), .C2(keyinput_f70), .A(n21091), .ZN(n21092)
         );
  NAND4_X1 U24039 ( .A1(n21095), .A2(n21094), .A3(n21093), .A4(n21092), .ZN(
        n21255) );
  OAI22_X1 U24040 ( .A1(P1_EBX_REG_29__SCAN_IN), .A2(keyinput_f86), .B1(
        keyinput_f82), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n21096) );
  AOI221_X1 U24041 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(keyinput_f86), .C1(
        P1_REIP_REG_1__SCAN_IN), .C2(keyinput_f82), .A(n21096), .ZN(n21122) );
  OAI22_X1 U24042 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(keyinput_f96), .B1(
        keyinput_f25), .B2(DATAI_7_), .ZN(n21097) );
  AOI221_X1 U24043 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(keyinput_f96), .C1(
        DATAI_7_), .C2(keyinput_f25), .A(n21097), .ZN(n21100) );
  OAI22_X1 U24044 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(keyinput_f94), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(keyinput_f68), .ZN(n21098) );
  AOI221_X1 U24045 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(keyinput_f94), .C1(
        keyinput_f68), .C2(P1_REIP_REG_15__SCAN_IN), .A(n21098), .ZN(n21099)
         );
  OAI211_X1 U24046 ( .C1(n21102), .C2(keyinput_f56), .A(n21100), .B(n21099), 
        .ZN(n21101) );
  AOI21_X1 U24047 ( .B1(n21102), .B2(keyinput_f56), .A(n21101), .ZN(n21121) );
  AOI22_X1 U24048 ( .A1(DATAI_25_), .A2(keyinput_f7), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(keyinput_f119), .ZN(n21103) );
  OAI221_X1 U24049 ( .B1(DATAI_25_), .B2(keyinput_f7), .C1(
        P1_EAX_REG_28__SCAN_IN), .C2(keyinput_f119), .A(n21103), .ZN(n21110)
         );
  AOI22_X1 U24050 ( .A1(DATAI_3_), .A2(keyinput_f29), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(keyinput_f79), .ZN(n21104) );
  OAI221_X1 U24051 ( .B1(DATAI_3_), .B2(keyinput_f29), .C1(
        P1_REIP_REG_4__SCAN_IN), .C2(keyinput_f79), .A(n21104), .ZN(n21109) );
  AOI22_X1 U24052 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(keyinput_f73), .B1(
        P1_EBX_REG_10__SCAN_IN), .B2(keyinput_f105), .ZN(n21105) );
  OAI221_X1 U24053 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(keyinput_f73), .C1(
        P1_EBX_REG_10__SCAN_IN), .C2(keyinput_f105), .A(n21105), .ZN(n21108)
         );
  AOI22_X1 U24054 ( .A1(DATAI_28_), .A2(keyinput_f4), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(keyinput_f74), .ZN(n21106) );
  OAI221_X1 U24055 ( .B1(DATAI_28_), .B2(keyinput_f4), .C1(
        P1_REIP_REG_9__SCAN_IN), .C2(keyinput_f74), .A(n21106), .ZN(n21107) );
  NOR4_X1 U24056 ( .A1(n21110), .A2(n21109), .A3(n21108), .A4(n21107), .ZN(
        n21120) );
  AOI22_X1 U24057 ( .A1(keyinput_f48), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_EBX_REG_11__SCAN_IN), .B2(keyinput_f104), .ZN(n21111) );
  OAI221_X1 U24058 ( .B1(keyinput_f48), .B2(P1_BYTEENABLE_REG_0__SCAN_IN), 
        .C1(P1_EBX_REG_11__SCAN_IN), .C2(keyinput_f104), .A(n21111), .ZN(
        n21118) );
  AOI22_X1 U24059 ( .A1(READY1), .A2(keyinput_f36), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n21112) );
  OAI221_X1 U24060 ( .B1(READY1), .B2(keyinput_f36), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_f44), .A(n21112), .ZN(n21117)
         );
  AOI22_X1 U24061 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(keyinput_f81), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(keyinput_f85), .ZN(n21113) );
  OAI221_X1 U24062 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(keyinput_f81), .C1(
        P1_EBX_REG_30__SCAN_IN), .C2(keyinput_f85), .A(n21113), .ZN(n21116) );
  AOI22_X1 U24063 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(keyinput_f106), .B1(
        P1_EBX_REG_0__SCAN_IN), .B2(keyinput_f115), .ZN(n21114) );
  OAI221_X1 U24064 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(keyinput_f106), .C1(
        P1_EBX_REG_0__SCAN_IN), .C2(keyinput_f115), .A(n21114), .ZN(n21115) );
  NOR4_X1 U24065 ( .A1(n21118), .A2(n21117), .A3(n21116), .A4(n21115), .ZN(
        n21119) );
  NAND4_X1 U24066 ( .A1(n21122), .A2(n21121), .A3(n21120), .A4(n21119), .ZN(
        n21254) );
  AOI22_X1 U24067 ( .A1(n21125), .A2(keyinput_f103), .B1(keyinput_f6), .B2(
        n21124), .ZN(n21123) );
  OAI221_X1 U24068 ( .B1(n21125), .B2(keyinput_f103), .C1(n21124), .C2(
        keyinput_f6), .A(n21123), .ZN(n21137) );
  AOI22_X1 U24069 ( .A1(n21128), .A2(keyinput_f114), .B1(n21127), .B2(
        keyinput_f101), .ZN(n21126) );
  OAI221_X1 U24070 ( .B1(n21128), .B2(keyinput_f114), .C1(n21127), .C2(
        keyinput_f101), .A(n21126), .ZN(n21136) );
  AOI22_X1 U24071 ( .A1(n21130), .A2(keyinput_f39), .B1(n12523), .B2(
        keyinput_f26), .ZN(n21129) );
  OAI221_X1 U24072 ( .B1(n21130), .B2(keyinput_f39), .C1(n12523), .C2(
        keyinput_f26), .A(n21129), .ZN(n21135) );
  INV_X1 U24073 ( .A(DATAI_0_), .ZN(n21133) );
  AOI22_X1 U24074 ( .A1(n21133), .A2(keyinput_f32), .B1(n21132), .B2(
        keyinput_f126), .ZN(n21131) );
  OAI221_X1 U24075 ( .B1(n21133), .B2(keyinput_f32), .C1(n21132), .C2(
        keyinput_f126), .A(n21131), .ZN(n21134) );
  NOR4_X1 U24076 ( .A1(n21137), .A2(n21136), .A3(n21135), .A4(n21134), .ZN(
        n21188) );
  AOI22_X1 U24077 ( .A1(n21140), .A2(keyinput_f11), .B1(n21139), .B2(
        keyinput_f57), .ZN(n21138) );
  OAI221_X1 U24078 ( .B1(n21140), .B2(keyinput_f11), .C1(n21139), .C2(
        keyinput_f57), .A(n21138), .ZN(n21153) );
  INV_X1 U24079 ( .A(READY2), .ZN(n21142) );
  AOI22_X1 U24080 ( .A1(n21143), .A2(keyinput_f102), .B1(keyinput_f37), .B2(
        n21142), .ZN(n21141) );
  OAI221_X1 U24081 ( .B1(n21143), .B2(keyinput_f102), .C1(n21142), .C2(
        keyinput_f37), .A(n21141), .ZN(n21152) );
  AOI22_X1 U24082 ( .A1(n21146), .A2(keyinput_f5), .B1(keyinput_f16), .B2(
        n21145), .ZN(n21144) );
  OAI221_X1 U24083 ( .B1(n21146), .B2(keyinput_f5), .C1(n21145), .C2(
        keyinput_f16), .A(n21144), .ZN(n21151) );
  AOI22_X1 U24084 ( .A1(n21149), .A2(keyinput_f118), .B1(keyinput_f60), .B2(
        n21148), .ZN(n21147) );
  OAI221_X1 U24085 ( .B1(n21149), .B2(keyinput_f118), .C1(n21148), .C2(
        keyinput_f60), .A(n21147), .ZN(n21150) );
  NOR4_X1 U24086 ( .A1(n21153), .A2(n21152), .A3(n21151), .A4(n21150), .ZN(
        n21187) );
  AOI22_X1 U24087 ( .A1(n21156), .A2(keyinput_f31), .B1(n21155), .B2(
        keyinput_f127), .ZN(n21154) );
  OAI221_X1 U24088 ( .B1(n21156), .B2(keyinput_f31), .C1(n21155), .C2(
        keyinput_f127), .A(n21154), .ZN(n21169) );
  AOI22_X1 U24089 ( .A1(n21159), .A2(keyinput_f9), .B1(keyinput_f46), .B2(
        n21158), .ZN(n21157) );
  OAI221_X1 U24090 ( .B1(n21159), .B2(keyinput_f9), .C1(n21158), .C2(
        keyinput_f46), .A(n21157), .ZN(n21168) );
  AOI22_X1 U24091 ( .A1(n21162), .A2(keyinput_f78), .B1(n21161), .B2(
        keyinput_f100), .ZN(n21160) );
  OAI221_X1 U24092 ( .B1(n21162), .B2(keyinput_f78), .C1(n21161), .C2(
        keyinput_f100), .A(n21160), .ZN(n21167) );
  AOI22_X1 U24093 ( .A1(n21165), .A2(keyinput_f97), .B1(keyinput_f99), .B2(
        n21164), .ZN(n21163) );
  OAI221_X1 U24094 ( .B1(n21165), .B2(keyinput_f97), .C1(n21164), .C2(
        keyinput_f99), .A(n21163), .ZN(n21166) );
  NOR4_X1 U24095 ( .A1(n21169), .A2(n21168), .A3(n21167), .A4(n21166), .ZN(
        n21186) );
  INV_X1 U24096 ( .A(keyinput_f35), .ZN(n21171) );
  AOI22_X1 U24097 ( .A1(n21172), .A2(keyinput_f8), .B1(BS16), .B2(n21171), 
        .ZN(n21170) );
  OAI221_X1 U24098 ( .B1(n21172), .B2(keyinput_f8), .C1(n21171), .C2(BS16), 
        .A(n21170), .ZN(n21184) );
  INV_X1 U24099 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21174) );
  AOI22_X1 U24100 ( .A1(n21175), .A2(keyinput_f88), .B1(keyinput_f38), .B2(
        n21174), .ZN(n21173) );
  OAI221_X1 U24101 ( .B1(n21175), .B2(keyinput_f88), .C1(n21174), .C2(
        keyinput_f38), .A(n21173), .ZN(n21183) );
  AOI22_X1 U24102 ( .A1(n21178), .A2(keyinput_f47), .B1(n21177), .B2(
        keyinput_f59), .ZN(n21176) );
  OAI221_X1 U24103 ( .B1(n21178), .B2(keyinput_f47), .C1(n21177), .C2(
        keyinput_f59), .A(n21176), .ZN(n21182) );
  AOI22_X1 U24104 ( .A1(n12622), .A2(keyinput_f17), .B1(n21180), .B2(
        keyinput_f95), .ZN(n21179) );
  OAI221_X1 U24105 ( .B1(n12622), .B2(keyinput_f17), .C1(n21180), .C2(
        keyinput_f95), .A(n21179), .ZN(n21181) );
  NOR4_X1 U24106 ( .A1(n21184), .A2(n21183), .A3(n21182), .A4(n21181), .ZN(
        n21185) );
  NAND4_X1 U24107 ( .A1(n21188), .A2(n21187), .A3(n21186), .A4(n21185), .ZN(
        n21253) );
  AOI22_X1 U24108 ( .A1(n21191), .A2(keyinput_f125), .B1(keyinput_f51), .B2(
        n21190), .ZN(n21189) );
  OAI221_X1 U24109 ( .B1(n21191), .B2(keyinput_f125), .C1(n21190), .C2(
        keyinput_f51), .A(n21189), .ZN(n21204) );
  AOI22_X1 U24110 ( .A1(n21194), .A2(keyinput_f24), .B1(keyinput_f14), .B2(
        n21193), .ZN(n21192) );
  OAI221_X1 U24111 ( .B1(n21194), .B2(keyinput_f24), .C1(n21193), .C2(
        keyinput_f14), .A(n21192), .ZN(n21203) );
  AOI22_X1 U24112 ( .A1(n21197), .A2(keyinput_f122), .B1(keyinput_f23), .B2(
        n21196), .ZN(n21195) );
  OAI221_X1 U24113 ( .B1(n21197), .B2(keyinput_f122), .C1(n21196), .C2(
        keyinput_f23), .A(n21195), .ZN(n21202) );
  AOI22_X1 U24114 ( .A1(n21200), .A2(keyinput_f71), .B1(keyinput_f49), .B2(
        n21199), .ZN(n21198) );
  OAI221_X1 U24115 ( .B1(n21200), .B2(keyinput_f71), .C1(n21199), .C2(
        keyinput_f49), .A(n21198), .ZN(n21201) );
  NOR4_X1 U24116 ( .A1(n21204), .A2(n21203), .A3(n21202), .A4(n21201), .ZN(
        n21251) );
  AOI22_X1 U24117 ( .A1(n21207), .A2(keyinput_f83), .B1(n21206), .B2(
        keyinput_f121), .ZN(n21205) );
  OAI221_X1 U24118 ( .B1(n21207), .B2(keyinput_f83), .C1(n21206), .C2(
        keyinput_f121), .A(n21205), .ZN(n21219) );
  AOI22_X1 U24119 ( .A1(n21210), .A2(keyinput_f66), .B1(keyinput_f61), .B2(
        n21209), .ZN(n21208) );
  OAI221_X1 U24120 ( .B1(n21210), .B2(keyinput_f66), .C1(n21209), .C2(
        keyinput_f61), .A(n21208), .ZN(n21218) );
  AOI22_X1 U24121 ( .A1(n14928), .A2(keyinput_f58), .B1(keyinput_f15), .B2(
        n21212), .ZN(n21211) );
  OAI221_X1 U24122 ( .B1(n14928), .B2(keyinput_f58), .C1(n21212), .C2(
        keyinput_f15), .A(n21211), .ZN(n21217) );
  AOI22_X1 U24123 ( .A1(n21215), .A2(keyinput_f77), .B1(keyinput_f13), .B2(
        n21214), .ZN(n21213) );
  OAI221_X1 U24124 ( .B1(n21215), .B2(keyinput_f77), .C1(n21214), .C2(
        keyinput_f13), .A(n21213), .ZN(n21216) );
  NOR4_X1 U24125 ( .A1(n21219), .A2(n21218), .A3(n21217), .A4(n21216), .ZN(
        n21250) );
  AOI22_X1 U24126 ( .A1(n21222), .A2(keyinput_f98), .B1(keyinput_f111), .B2(
        n21221), .ZN(n21220) );
  OAI221_X1 U24127 ( .B1(n21222), .B2(keyinput_f98), .C1(n21221), .C2(
        keyinput_f111), .A(n21220), .ZN(n21232) );
  AOI22_X1 U24128 ( .A1(n21225), .A2(keyinput_f0), .B1(n21224), .B2(
        keyinput_f92), .ZN(n21223) );
  OAI221_X1 U24129 ( .B1(n21225), .B2(keyinput_f0), .C1(n21224), .C2(
        keyinput_f92), .A(n21223), .ZN(n21231) );
  INV_X1 U24130 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21227) );
  AOI22_X1 U24131 ( .A1(n21227), .A2(keyinput_f40), .B1(n12543), .B2(
        keyinput_f28), .ZN(n21226) );
  OAI221_X1 U24132 ( .B1(n21227), .B2(keyinput_f40), .C1(n12543), .C2(
        keyinput_f28), .A(n21226), .ZN(n21230) );
  AOI22_X1 U24133 ( .A1(n13790), .A2(keyinput_f75), .B1(n13415), .B2(
        keyinput_f80), .ZN(n21228) );
  OAI221_X1 U24134 ( .B1(n13790), .B2(keyinput_f75), .C1(n13415), .C2(
        keyinput_f80), .A(n21228), .ZN(n21229) );
  NOR4_X1 U24135 ( .A1(n21232), .A2(n21231), .A3(n21230), .A4(n21229), .ZN(
        n21249) );
  AOI22_X1 U24136 ( .A1(n21235), .A2(keyinput_f90), .B1(keyinput_f22), .B2(
        n21234), .ZN(n21233) );
  OAI221_X1 U24137 ( .B1(n21235), .B2(keyinput_f90), .C1(n21234), .C2(
        keyinput_f22), .A(n21233), .ZN(n21247) );
  AOI22_X1 U24138 ( .A1(n21237), .A2(keyinput_f65), .B1(keyinput_f27), .B2(
        n12538), .ZN(n21236) );
  OAI221_X1 U24139 ( .B1(n21237), .B2(keyinput_f65), .C1(n12538), .C2(
        keyinput_f27), .A(n21236), .ZN(n21246) );
  INV_X1 U24140 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n21240) );
  AOI22_X1 U24141 ( .A1(n21240), .A2(keyinput_f116), .B1(keyinput_f107), .B2(
        n21239), .ZN(n21238) );
  OAI221_X1 U24142 ( .B1(n21240), .B2(keyinput_f116), .C1(n21239), .C2(
        keyinput_f107), .A(n21238), .ZN(n21245) );
  AOI22_X1 U24143 ( .A1(n21243), .A2(keyinput_f21), .B1(keyinput_f45), .B2(
        n21242), .ZN(n21241) );
  OAI221_X1 U24144 ( .B1(n21243), .B2(keyinput_f21), .C1(n21242), .C2(
        keyinput_f45), .A(n21241), .ZN(n21244) );
  NOR4_X1 U24145 ( .A1(n21247), .A2(n21246), .A3(n21245), .A4(n21244), .ZN(
        n21248) );
  NAND4_X1 U24146 ( .A1(n21251), .A2(n21250), .A3(n21249), .A4(n21248), .ZN(
        n21252) );
  NOR4_X1 U24147 ( .A1(n21255), .A2(n21254), .A3(n21253), .A4(n21252), .ZN(
        n21298) );
  OAI22_X1 U24148 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(keyinput_f76), .B1(
        keyinput_f63), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n21256) );
  AOI221_X1 U24149 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(keyinput_f76), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_f63), .A(n21256), .ZN(n21263)
         );
  OAI22_X1 U24150 ( .A1(P1_EBX_REG_22__SCAN_IN), .A2(keyinput_f93), .B1(
        keyinput_f54), .B2(P1_REIP_REG_29__SCAN_IN), .ZN(n21257) );
  AOI221_X1 U24151 ( .B1(P1_EBX_REG_22__SCAN_IN), .B2(keyinput_f93), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_f54), .A(n21257), .ZN(n21262)
         );
  OAI22_X1 U24152 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(keyinput_f108), .B1(
        DATAI_13_), .B2(keyinput_f19), .ZN(n21258) );
  AOI221_X1 U24153 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(keyinput_f108), .C1(
        keyinput_f19), .C2(DATAI_13_), .A(n21258), .ZN(n21261) );
  OAI22_X1 U24154 ( .A1(P1_EAX_REG_27__SCAN_IN), .A2(keyinput_f120), .B1(
        P1_EBX_REG_3__SCAN_IN), .B2(keyinput_f112), .ZN(n21259) );
  AOI221_X1 U24155 ( .B1(P1_EAX_REG_27__SCAN_IN), .B2(keyinput_f120), .C1(
        keyinput_f112), .C2(P1_EBX_REG_3__SCAN_IN), .A(n21259), .ZN(n21260) );
  NAND4_X1 U24156 ( .A1(n21263), .A2(n21262), .A3(n21261), .A4(n21260), .ZN(
        n21296) );
  OAI22_X1 U24157 ( .A1(P1_EAX_REG_30__SCAN_IN), .A2(keyinput_f117), .B1(
        P1_EBX_REG_24__SCAN_IN), .B2(keyinput_f91), .ZN(n21264) );
  AOI221_X1 U24158 ( .B1(P1_EAX_REG_30__SCAN_IN), .B2(keyinput_f117), .C1(
        keyinput_f91), .C2(P1_EBX_REG_24__SCAN_IN), .A(n21264), .ZN(n21271) );
  OAI22_X1 U24159 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput_f67), .B1(
        DATAI_2_), .B2(keyinput_f30), .ZN(n21265) );
  AOI221_X1 U24160 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(keyinput_f67), .C1(
        keyinput_f30), .C2(DATAI_2_), .A(n21265), .ZN(n21270) );
  OAI22_X1 U24161 ( .A1(DATAI_12_), .A2(keyinput_f20), .B1(keyinput_f43), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21266) );
  AOI221_X1 U24162 ( .B1(DATAI_12_), .B2(keyinput_f20), .C1(
        P1_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_f43), .A(n21266), .ZN(
        n21269) );
  OAI22_X1 U24163 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(keyinput_f84), .B1(
        keyinput_f3), .B2(DATAI_29_), .ZN(n21267) );
  AOI221_X1 U24164 ( .B1(P1_EBX_REG_31__SCAN_IN), .B2(keyinput_f84), .C1(
        DATAI_29_), .C2(keyinput_f3), .A(n21267), .ZN(n21268) );
  NAND4_X1 U24165 ( .A1(n21271), .A2(n21270), .A3(n21269), .A4(n21268), .ZN(
        n21295) );
  OAI22_X1 U24166 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(keyinput_f55), .B1(
        keyinput_f34), .B2(NA), .ZN(n21272) );
  AOI221_X1 U24167 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_f55), .C1(NA), 
        .C2(keyinput_f34), .A(n21272), .ZN(n21279) );
  OAI22_X1 U24168 ( .A1(P1_EBX_REG_5__SCAN_IN), .A2(keyinput_f110), .B1(
        keyinput_f10), .B2(DATAI_22_), .ZN(n21273) );
  AOI221_X1 U24169 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(keyinput_f110), .C1(
        DATAI_22_), .C2(keyinput_f10), .A(n21273), .ZN(n21278) );
  OAI22_X1 U24170 ( .A1(P1_EBX_REG_26__SCAN_IN), .A2(keyinput_f89), .B1(
        DATAI_14_), .B2(keyinput_f18), .ZN(n21274) );
  AOI221_X1 U24171 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(keyinput_f89), .C1(
        keyinput_f18), .C2(DATAI_14_), .A(n21274), .ZN(n21277) );
  OAI22_X1 U24172 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(keyinput_f72), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(keyinput_f69), .ZN(n21275) );
  AOI221_X1 U24173 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(keyinput_f72), .C1(
        keyinput_f69), .C2(P1_REIP_REG_14__SCAN_IN), .A(n21275), .ZN(n21276)
         );
  NAND4_X1 U24174 ( .A1(n21279), .A2(n21278), .A3(n21277), .A4(n21276), .ZN(
        n21294) );
  OAI22_X1 U24175 ( .A1(P1_EAX_REG_23__SCAN_IN), .A2(keyinput_f124), .B1(
        keyinput_f12), .B2(DATAI_20_), .ZN(n21280) );
  AOI221_X1 U24176 ( .B1(P1_EAX_REG_23__SCAN_IN), .B2(keyinput_f124), .C1(
        DATAI_20_), .C2(keyinput_f12), .A(n21280), .ZN(n21292) );
  OAI22_X1 U24177 ( .A1(n21282), .A2(keyinput_f41), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(keyinput_f64), .ZN(n21281) );
  AOI221_X1 U24178 ( .B1(n21282), .B2(keyinput_f41), .C1(keyinput_f64), .C2(
        P1_REIP_REG_19__SCAN_IN), .A(n21281), .ZN(n21291) );
  INV_X1 U24179 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21284) );
  OAI22_X1 U24180 ( .A1(n21285), .A2(keyinput_f52), .B1(n21284), .B2(
        keyinput_f53), .ZN(n21283) );
  AOI221_X1 U24181 ( .B1(n21285), .B2(keyinput_f52), .C1(keyinput_f53), .C2(
        n21284), .A(n21283), .ZN(n21290) );
  OAI22_X1 U24182 ( .A1(n21288), .A2(keyinput_f62), .B1(n21287), .B2(
        keyinput_f2), .ZN(n21286) );
  AOI221_X1 U24183 ( .B1(n21288), .B2(keyinput_f62), .C1(keyinput_f2), .C2(
        n21287), .A(n21286), .ZN(n21289) );
  NAND4_X1 U24184 ( .A1(n21292), .A2(n21291), .A3(n21290), .A4(n21289), .ZN(
        n21293) );
  NOR4_X1 U24185 ( .A1(n21296), .A2(n21295), .A3(n21294), .A4(n21293), .ZN(
        n21297) );
  AOI22_X1 U24186 ( .A1(n21298), .A2(n21297), .B1(P1_D_C_N_REG_SCAN_IN), .B2(
        keyinput_f42), .ZN(n21299) );
  OAI21_X1 U24187 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_f42), .A(n21299), 
        .ZN(n21300) );
  OAI211_X1 U24188 ( .C1(P1_D_C_N_REG_SCAN_IN), .C2(keyinput_g42), .A(n21301), 
        .B(n21300), .ZN(n21302) );
  XOR2_X1 U24189 ( .A(n21303), .B(n21302), .Z(U355) );
  AND2_X1 U15433 ( .A1(n13176), .A2(n15173), .ZN(n14394) );
  INV_X1 U11274 ( .A(n9926), .ZN(n17417) );
  INV_X1 U11271 ( .A(n12096), .ZN(n19460) );
  NOR2_X1 U11269 ( .A1(n20260), .A2(n10136), .ZN(n13168) );
  INV_X1 U11257 ( .A(n11251), .ZN(n14459) );
  CLKBUF_X1 U11256 ( .A(n12256), .Z(n14331) );
  CLKBUF_X1 U11299 ( .A(n12449), .Z(n12450) );
  CLKBUF_X1 U11332 ( .A(n12665), .Z(n14223) );
  CLKBUF_X1 U11488 ( .A(n12475), .Z(n12478) );
  OR2_X1 U11656 ( .A1(n12954), .A2(n12953), .ZN(n12955) );
  CLKBUF_X1 U12270 ( .A(n11168), .Z(n11169) );
  CLKBUF_X1 U12441 ( .A(n11477), .Z(n17261) );
  INV_X1 U12540 ( .A(n20254), .ZN(n12508) );
  CLKBUF_X1 U12675 ( .A(n13211), .Z(n9811) );
  CLKBUF_X1 U12730 ( .A(n11491), .Z(n17453) );
  CLKBUF_X1 U13068 ( .A(n20133), .Z(n9798) );
  CLKBUF_X1 U13085 ( .A(n14671), .Z(n14672) );
  OR2_X1 U13113 ( .A1(n13052), .A2(n10248), .ZN(n15222) );
  CLKBUF_X1 U16027 ( .A(n19384), .Z(n19399) );
  INV_X1 U16331 ( .A(n13682), .ZN(n11259) );
  CLKBUF_X1 U18117 ( .A(n17744), .Z(n17747) );
endmodule

