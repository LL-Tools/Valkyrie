

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906;

  OR2_X2 U3418 ( .A1(n5219), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3820) );
  INV_X1 U3419 ( .A(n5662), .ZN(n5760) );
  INV_X1 U3420 ( .A(n3190), .ZN(n3201) );
  INV_X4 U3421 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5165) );
  CLKBUF_X2 U3422 ( .A(n4320), .Z(n4748) );
  CLKBUF_X3 U3423 ( .A(n3468), .Z(n4343) );
  INV_X1 U3424 ( .A(n4344), .ZN(n4296) );
  INV_X1 U3425 ( .A(n3426), .ZN(n4595) );
  BUF_X2 U3426 ( .A(n4317), .Z(n4350) );
  CLKBUF_X3 U3427 ( .A(n3474), .Z(n4353) );
  AND4_X2 U3428 ( .A1(n3303), .A2(n3301), .A3(n3302), .A4(n3300), .ZN(n4599)
         );
  AND4_X1 U3429 ( .A1(n3299), .A2(n3298), .A3(n3297), .A4(n3296), .ZN(n3300)
         );
  AND4_X1 U3430 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3384)
         );
  AND2_X1 U3431 ( .A1(n4744), .A2(n3158), .ZN(n3403) );
  AND2_X2 U3432 ( .A1(n3163), .A2(n4745), .ZN(n3476) );
  AND2_X2 U3433 ( .A1(n5194), .A2(n4742), .ZN(n3386) );
  NAND2_X1 U3434 ( .A1(n3462), .A2(n5479), .ZN(n3554) );
  NAND2_X1 U3435 ( .A1(n3536), .A2(n3535), .ZN(n3593) );
  AND4_X1 U3436 ( .A1(n3381), .A2(n3380), .A3(n3379), .A4(n3378), .ZN(n3382)
         );
  NOR2_X1 U3437 ( .A1(n3765), .A2(n3105), .ZN(n3104) );
  INV_X1 U3438 ( .A(n4599), .ZN(n3453) );
  NAND3_X1 U3439 ( .A1(n3434), .A2(n3524), .A3(n3433), .ZN(n3531) );
  AND2_X2 U3440 ( .A1(n3152), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4745)
         );
  AND2_X2 U3441 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4742) );
  AND2_X1 U3444 ( .A1(n3400), .A2(n3421), .ZN(n5479) );
  NAND2_X1 U34450 ( .A1(n4588), .A2(n3426), .ZN(n3431) );
  OR3_X1 U34460 ( .A1(n6725), .A2(n6368), .A3(n3831), .ZN(n6197) );
  NAND2_X1 U34470 ( .A1(n5452), .A2(n2996), .ZN(n5419) );
  INV_X2 U34480 ( .A(n5179), .ZN(n3941) );
  OAI21_X2 U3449 ( .B1(n3514), .B2(n3513), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3520) );
  INV_X2 U34510 ( .A(n5662), .ZN(n5757) );
  OR2_X1 U34520 ( .A1(n4397), .A2(n6015), .ZN(n4398) );
  NAND2_X1 U34530 ( .A1(n3017), .A2(n3768), .ZN(n5653) );
  NAND2_X1 U3454 ( .A1(n3585), .A2(n3584), .ZN(n3589) );
  AND2_X1 U34550 ( .A1(n5554), .A2(n3113), .ZN(n5471) );
  OAI21_X1 U34560 ( .B1(n3531), .B2(n3422), .A(n3556), .ZN(n3519) );
  NAND2_X1 U3457 ( .A1(n3555), .A2(n3507), .ZN(n3784) );
  NAND2_X1 U3458 ( .A1(n3530), .A2(n3422), .ZN(n6711) );
  NAND2_X1 U34590 ( .A1(n3862), .A2(n3453), .ZN(n3430) );
  INV_X2 U34610 ( .A(n3421), .ZN(n2971) );
  CLKBUF_X3 U34620 ( .A(n4027), .Z(n4197) );
  CLKBUF_X3 U34630 ( .A(n3412), .Z(n4352) );
  AND2_X1 U34650 ( .A1(n4432), .A2(n4430), .ZN(n3047) );
  AOI21_X1 U3466 ( .B1(n5622), .B2(n5804), .A(n5621), .ZN(n5623) );
  AND2_X1 U3467 ( .A1(n3056), .A2(n3055), .ZN(n5639) );
  AND2_X1 U34680 ( .A1(n4404), .A2(n4403), .ZN(n5622) );
  XNOR2_X1 U34690 ( .A(n4373), .B(n4372), .ZN(n5215) );
  OR2_X1 U34700 ( .A1(n5272), .A2(n5259), .ZN(n3055) );
  OR2_X1 U34710 ( .A1(n4397), .A2(n6101), .ZN(n3011) );
  OAI21_X1 U34720 ( .B1(n5247), .B2(n5248), .A(n4401), .ZN(n5626) );
  OR2_X1 U34730 ( .A1(n5688), .A2(n2998), .ZN(n3145) );
  NAND2_X1 U34740 ( .A1(n3016), .A2(n3015), .ZN(n5616) );
  INV_X1 U3475 ( .A(n5653), .ZN(n3016) );
  NAND2_X1 U3476 ( .A1(n3040), .A2(n3043), .ZN(n5651) );
  NAND2_X1 U3477 ( .A1(n5705), .A2(n3767), .ZN(n3017) );
  NAND2_X1 U3478 ( .A1(n3101), .A2(n3102), .ZN(n5705) );
  INV_X1 U3479 ( .A(n5416), .ZN(n3128) );
  NAND2_X1 U3480 ( .A1(n5736), .A2(n3104), .ZN(n3101) );
  NAND2_X1 U3481 ( .A1(n3079), .A2(n2981), .ZN(n5745) );
  AND2_X1 U3482 ( .A1(n2993), .A2(n3097), .ZN(n3096) );
  NAND2_X1 U3483 ( .A1(n5798), .A2(n5799), .ZN(n3107) );
  NOR2_X1 U3484 ( .A1(n5778), .A2(n3078), .ZN(n3077) );
  INV_X1 U3485 ( .A(n3104), .ZN(n3099) );
  NOR2_X1 U3486 ( .A1(n5662), .A2(n3770), .ZN(n3015) );
  XNOR2_X1 U3487 ( .A(n3728), .B(n3727), .ZN(n5054) );
  OAI21_X1 U3488 ( .B1(n3912), .B2(n3726), .A(n3725), .ZN(n3728) );
  INV_X2 U3489 ( .A(n3753), .ZN(n5662) );
  NAND2_X1 U3490 ( .A1(n3741), .A2(n3744), .ZN(n3753) );
  NAND2_X1 U3491 ( .A1(n3741), .A2(n3723), .ZN(n3912) );
  AND2_X1 U3492 ( .A1(n3675), .A2(n3696), .ZN(n3895) );
  CLKBUF_X1 U3493 ( .A(n5288), .Z(n5306) );
  AND2_X1 U3494 ( .A1(n5288), .A2(n5289), .ZN(n5279) );
  NAND2_X2 U3495 ( .A1(n3650), .A2(n3649), .ZN(n4627) );
  NAND2_X1 U3496 ( .A1(n3623), .A2(n3624), .ZN(n3657) );
  CLKBUF_X1 U3497 ( .A(n5370), .Z(n5406) );
  NAND2_X2 U3498 ( .A1(n3589), .A2(n3588), .ZN(n4587) );
  CLKBUF_X1 U3499 ( .A(n5559), .Z(n5598) );
  NAND2_X1 U3500 ( .A1(n4580), .A2(n6722), .ZN(n3650) );
  NOR2_X1 U3501 ( .A1(n6295), .A2(n6018), .ZN(n6577) );
  OR2_X2 U3502 ( .A1(n6329), .A2(n4518), .ZN(n6341) );
  NAND2_X1 U3503 ( .A1(n3867), .A2(n3866), .ZN(n4517) );
  OAI211_X1 U3504 ( .C1(n4534), .C2(n4529), .A(n4528), .B(n6324), .ZN(n5213)
         );
  AND2_X2 U3505 ( .A1(n6101), .A2(n4380), .ZN(n6329) );
  AND2_X1 U3506 ( .A1(n3581), .A2(n3580), .ZN(n2974) );
  AOI21_X1 U3507 ( .B1(n4557), .B2(n4558), .A(n3197), .ZN(n4856) );
  NAND2_X1 U3508 ( .A1(n3499), .A2(n3498), .ZN(n3586) );
  MUX2_X1 U3509 ( .A(n3537), .B(n3743), .S(n3590), .Z(n3587) );
  NAND2_X1 U3510 ( .A1(n3517), .A2(n3431), .ZN(n3518) );
  INV_X1 U3511 ( .A(n3857), .ZN(n5216) );
  AND2_X1 U3512 ( .A1(n4409), .A2(n3501), .ZN(n3537) );
  AND2_X2 U3513 ( .A1(n3329), .A2(n3453), .ZN(n3517) );
  CLKBUF_X1 U3514 ( .A(n3509), .Z(n4469) );
  OR2_X2 U3515 ( .A1(n3461), .A2(n3530), .ZN(n3274) );
  INV_X1 U3516 ( .A(n3461), .ZN(n4603) );
  CLKBUF_X2 U3517 ( .A(n3432), .Z(n4405) );
  CLKBUF_X1 U3518 ( .A(n3427), .Z(n4530) );
  NAND2_X1 U3519 ( .A1(n2980), .A2(n3189), .ZN(n3461) );
  NOR2_X1 U3520 ( .A1(n3480), .A2(n3479), .ZN(n3484) );
  NAND2_X1 U3521 ( .A1(n3144), .A2(n3417), .ZN(n3432) );
  AND4_X2 U3522 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3421)
         );
  AND4_X1 U3523 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(n3417)
         );
  AND4_X1 U3524 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3303)
         );
  AND4_X1 U3525 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(n3170)
         );
  AND4_X1 U3526 ( .A1(n3156), .A2(n3155), .A3(n3154), .A4(n3153), .ZN(n3171)
         );
  AND4_X1 U3527 ( .A1(n3295), .A2(n3294), .A3(n3293), .A4(n3292), .ZN(n3301)
         );
  AND4_X1 U3528 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3302)
         );
  INV_X2 U3529 ( .A(n6099), .ZN(n6673) );
  INV_X2 U3530 ( .A(n3409), .ZN(n3387) );
  BUF_X2 U3531 ( .A(n4345), .Z(n4278) );
  AND2_X1 U3532 ( .A1(n3157), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3164)
         );
  AND2_X1 U3533 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4744) );
  INV_X2 U3534 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3146) );
  NOR2_X2 U3535 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6437) );
  NAND2_X1 U3536 ( .A1(n4550), .A2(n3592), .ZN(n6331) );
  AND2_X2 U3537 ( .A1(n5187), .A2(n3164), .ZN(n3392) );
  XNOR2_X2 U3538 ( .A(n3655), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4661)
         );
  NOR2_X4 U3539 ( .A1(n5271), .A2(n5273), .ZN(n5260) );
  NAND2_X2 U3540 ( .A1(n3107), .A2(n3106), .ZN(n3079) );
  AND2_X2 U3541 ( .A1(n5260), .A2(n3139), .ZN(n4425) );
  NAND2_X2 U3542 ( .A1(n3128), .A2(n2978), .ZN(n5367) );
  NAND2_X2 U3543 ( .A1(n4521), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6380)
         );
  NOR2_X1 U3544 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3908) );
  OR2_X1 U3545 ( .A1(n4759), .A2(n6722), .ZN(n4334) );
  NAND2_X1 U3547 ( .A1(n3026), .A2(n3030), .ZN(n4534) );
  INV_X1 U3548 ( .A(n3031), .ZN(n3030) );
  NAND2_X1 U3549 ( .A1(n3028), .A2(n3027), .ZN(n3026) );
  OAI21_X1 U3550 ( .B1(n3034), .B2(n3032), .A(n5208), .ZN(n3031) );
  INV_X1 U3551 ( .A(n3657), .ZN(n3010) );
  AOI21_X1 U3552 ( .B1(n3349), .B2(n3348), .A(n3347), .ZN(n3354) );
  AND2_X1 U3553 ( .A1(n6519), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3347)
         );
  NAND2_X1 U3554 ( .A1(n3517), .A2(n3742), .ZN(n3351) );
  NOR2_X1 U3555 ( .A1(n6395), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3357)
         );
  AND2_X1 U3556 ( .A1(n3718), .A2(n3717), .ZN(n3721) );
  NAND2_X1 U3557 ( .A1(n3674), .A2(n3133), .ZN(n3722) );
  NOR2_X1 U3558 ( .A1(n3672), .A2(n3134), .ZN(n3133) );
  INV_X1 U3559 ( .A(n3671), .ZN(n3674) );
  OAI211_X1 U3560 ( .C1(n4456), .C2(n3560), .A(n3559), .B(n3558), .ZN(n3567)
         );
  INV_X1 U3561 ( .A(n3573), .ZN(n3418) );
  NAND2_X1 U3562 ( .A1(n3862), .A2(n3506), .ZN(n3452) );
  INV_X1 U3563 ( .A(n3517), .ZN(n3731) );
  NOR2_X1 U3564 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3158) );
  INV_X1 U3565 ( .A(n5551), .ZN(n3940) );
  AND2_X2 U3566 ( .A1(n3423), .A2(n3427), .ZN(n3862) );
  AND2_X1 U3567 ( .A1(n5652), .A2(n3044), .ZN(n3043) );
  NAND2_X1 U3568 ( .A1(n3768), .A2(n3045), .ZN(n3044) );
  INV_X1 U3569 ( .A(n3767), .ZN(n3045) );
  AND2_X1 U3570 ( .A1(n3461), .A2(n3422), .ZN(n3507) );
  NAND2_X1 U3571 ( .A1(n3098), .A2(n3104), .ZN(n3097) );
  INV_X1 U3572 ( .A(n3759), .ZN(n3098) );
  AND2_X1 U3573 ( .A1(n3743), .A2(n3742), .ZN(n3744) );
  AND2_X1 U3574 ( .A1(n3422), .A2(n3426), .ZN(n3742) );
  AND2_X1 U3575 ( .A1(n5165), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4370) );
  MUX2_X1 U3576 ( .A(n4312), .B(n5628), .S(n4369), .Z(n5248) );
  NAND2_X1 U3577 ( .A1(n4275), .A2(n3065), .ZN(n4313) );
  INV_X1 U3578 ( .A(n4111), .ZN(n4112) );
  NAND2_X1 U3579 ( .A1(n4112), .A2(n3072), .ZN(n4148) );
  NOR2_X1 U3580 ( .A1(n5425), .A2(n4022), .ZN(n3071) );
  INV_X1 U3581 ( .A(n4060), .ZN(n4061) );
  NAND2_X1 U3582 ( .A1(n3986), .A2(n3066), .ZN(n4060) );
  AND2_X1 U3583 ( .A1(n2976), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3066)
         );
  NOR3_X1 U3584 ( .A1(n5261), .A2(n5262), .A3(n5249), .ZN(n5250) );
  OR2_X1 U3585 ( .A1(n3775), .A2(n4524), .ZN(n4529) );
  AND2_X1 U3586 ( .A1(n3460), .A2(n3459), .ZN(n3792) );
  OR3_X1 U3587 ( .A1(n4534), .A2(n3458), .A3(n4405), .ZN(n3459) );
  NAND2_X1 U3588 ( .A1(n3029), .A2(n3363), .ZN(n4492) );
  NAND2_X1 U3589 ( .A1(n3035), .A2(n3034), .ZN(n3029) );
  NAND2_X1 U3590 ( .A1(n3028), .A2(n3025), .ZN(n3035) );
  INV_X1 U3591 ( .A(n3033), .ZN(n3025) );
  AND2_X1 U3592 ( .A1(n4673), .A2(n4672), .ZN(n4953) );
  OR2_X1 U3593 ( .A1(n5811), .A2(n5557), .ZN(n4421) );
  BUF_X1 U3594 ( .A(n3387), .Z(n4319) );
  NAND2_X1 U3595 ( .A1(n4599), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3500) );
  INV_X1 U3596 ( .A(n3351), .ZN(n3362) );
  NAND2_X1 U3597 ( .A1(n3412), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3368)
         );
  AND2_X1 U3598 ( .A1(n6395), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3355)
         );
  NOR2_X1 U3599 ( .A1(n3231), .A2(n3123), .ZN(n3122) );
  INV_X1 U3600 ( .A(n5453), .ZN(n3123) );
  INV_X1 U3601 ( .A(n3500), .ZN(n4409) );
  NOR2_X1 U3602 ( .A1(n4184), .A2(n5682), .ZN(n3076) );
  AND2_X1 U3603 ( .A1(n5315), .A2(n4181), .ZN(n3132) );
  INV_X1 U3604 ( .A(n5328), .ZN(n4181) );
  AND2_X1 U3605 ( .A1(n3940), .A2(n3058), .ZN(n3057) );
  INV_X1 U3606 ( .A(n5467), .ZN(n3058) );
  NOR2_X1 U3607 ( .A1(n3033), .A2(n3032), .ZN(n3027) );
  AND2_X1 U3608 ( .A1(n3857), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3881) );
  INV_X1 U3609 ( .A(n3768), .ZN(n3046) );
  NOR2_X1 U3610 ( .A1(n5303), .A2(n5304), .ZN(n5288) );
  AND2_X1 U3611 ( .A1(n5336), .A2(n5345), .ZN(n3126) );
  AOI21_X1 U3612 ( .B1(n3104), .B2(n3762), .A(n3103), .ZN(n3102) );
  INV_X1 U3613 ( .A(n3764), .ZN(n3103) );
  AND2_X1 U3614 ( .A1(n5744), .A2(n3755), .ZN(n3756) );
  INV_X1 U3615 ( .A(n3751), .ZN(n3078) );
  INV_X1 U3616 ( .A(n3204), .ZN(n3271) );
  NOR2_X1 U3617 ( .A1(n5548), .A2(n3116), .ZN(n3115) );
  INV_X1 U3618 ( .A(n5553), .ZN(n3116) );
  NOR2_X1 U3619 ( .A1(n3190), .A2(n4410), .ZN(n3266) );
  OAI21_X1 U3620 ( .B1(n3898), .B2(n3726), .A(n3703), .ZN(n3704) );
  NOR2_X1 U3621 ( .A1(n4489), .A2(n3789), .ZN(n3791) );
  INV_X1 U3622 ( .A(n3742), .ZN(n3726) );
  OR2_X1 U3623 ( .A1(n3565), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3566)
         );
  INV_X1 U3624 ( .A(n3328), .ZN(n3329) );
  NAND2_X1 U3625 ( .A1(n3515), .A2(n3500), .ZN(n3729) );
  AND2_X1 U3626 ( .A1(n3127), .A2(n3597), .ZN(n3623) );
  INV_X1 U3627 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4948) );
  AOI22_X1 U3628 ( .A1(n4320), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3180) );
  AND4_X1 U3629 ( .A1(n3188), .A2(n3187), .A3(n3186), .A4(n3185), .ZN(n3189)
         );
  AND2_X1 U3630 ( .A1(n4581), .A2(n5498), .ZN(n4951) );
  AND2_X1 U3631 ( .A1(n4459), .A2(n3829), .ZN(n4449) );
  AOI21_X1 U3632 ( .B1(n5238), .B2(n4369), .A(n4368), .ZN(n4424) );
  AOI22_X1 U3633 ( .A1(n4320), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3309) );
  NAND2_X1 U3634 ( .A1(n4516), .A2(n3869), .ZN(n4732) );
  NAND2_X1 U3635 ( .A1(n4731), .A2(n4732), .ZN(n4733) );
  INV_X1 U3636 ( .A(n5479), .ZN(n4524) );
  NOR2_X1 U3637 ( .A1(n4498), .A2(n4477), .ZN(n4527) );
  OR2_X1 U3638 ( .A1(n4315), .A2(n4314), .ZN(n4374) );
  INV_X1 U3639 ( .A(n3140), .ZN(n3138) );
  INV_X1 U3640 ( .A(n4129), .ZN(n5368) );
  NAND2_X1 U3641 ( .A1(n4061), .A2(n3003), .ZN(n4111) );
  INV_X1 U3642 ( .A(n4057), .ZN(n4058) );
  NOR2_X1 U3643 ( .A1(n6144), .A2(n3068), .ZN(n3067) );
  INV_X1 U3644 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3068) );
  AND2_X1 U3645 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n3982), .ZN(n3986)
         );
  AND2_X1 U3646 ( .A1(n3956), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3982)
         );
  NOR2_X1 U3647 ( .A1(n3923), .A2(n6755), .ZN(n3956) );
  AND3_X1 U3648 ( .A1(n3939), .A2(n3938), .A3(n3937), .ZN(n5551) );
  AND2_X1 U3649 ( .A1(n5908), .A2(n3819), .ZN(n5845) );
  NAND2_X1 U3650 ( .A1(n3089), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3082) );
  OR2_X1 U3651 ( .A1(n3090), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3087)
         );
  NAND2_X1 U3652 ( .A1(n5991), .A2(n3798), .ZN(n3020) );
  NOR2_X1 U3653 ( .A1(n5992), .A2(n3797), .ZN(n5931) );
  AND2_X1 U3654 ( .A1(n3141), .A2(n3750), .ZN(n3106) );
  INV_X1 U3655 ( .A(n6372), .ZN(n4664) );
  OR2_X1 U3656 ( .A1(n3775), .A2(n3506), .ZN(n4790) );
  NAND2_X1 U3657 ( .A1(n4459), .A2(n3422), .ZN(n4761) );
  INV_X1 U3658 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U3659 ( .A1(n3637), .A2(n3636), .ZN(n4674) );
  NAND2_X1 U3660 ( .A1(n4579), .A2(n6722), .ZN(n6018) );
  AND2_X1 U3661 ( .A1(n6021), .A2(n4587), .ZN(n6042) );
  AND2_X1 U3662 ( .A1(n6437), .A2(n6435), .ZN(n6582) );
  AND2_X1 U3663 ( .A1(n4949), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4676)
         );
  NOR2_X1 U3664 ( .A1(n6024), .A2(n4586), .ZN(n4673) );
  AOI21_X1 U3665 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6574), .A(n6018), .ZN(
        n6400) );
  AND2_X1 U3666 ( .A1(n4786), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3561) );
  NAND2_X1 U3667 ( .A1(n5225), .A2(n5223), .ZN(n5481) );
  INV_X1 U3668 ( .A(n5481), .ZN(n6890) );
  NAND2_X1 U3669 ( .A1(n6197), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6186) );
  AND2_X1 U3670 ( .A1(n5484), .A2(n5234), .ZN(n6895) );
  AND2_X1 U3671 ( .A1(n5484), .A2(n3833), .ZN(n6220) );
  INV_X1 U3672 ( .A(n6895), .ZN(n6229) );
  NOR2_X2 U3673 ( .A1(n5225), .A2(n5224), .ZN(n6889) );
  NAND2_X2 U3674 ( .A1(n5552), .A2(n5558), .ZN(n5557) );
  INV_X1 U3675 ( .A(n5639), .ZN(n5570) );
  INV_X2 U3676 ( .A(n5213), .ZN(n5612) );
  AND2_X1 U3677 ( .A1(n5213), .A2(n4532), .ZN(n5613) );
  XNOR2_X1 U3678 ( .A(n3070), .B(n4383), .ZN(n5225) );
  NOR2_X1 U3679 ( .A1(n4374), .A2(n5235), .ZN(n3070) );
  NAND2_X1 U3680 ( .A1(n4275), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4276)
         );
  NAND2_X1 U3681 ( .A1(n4183), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4185)
         );
  NAND2_X1 U3682 ( .A1(n4061), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4089)
         );
  INV_X1 U3683 ( .A(n6341), .ZN(n5787) );
  OR2_X2 U3684 ( .A1(n4534), .A2(n4790), .ZN(n6101) );
  INV_X1 U3685 ( .A(n6329), .ZN(n5784) );
  OR2_X1 U3686 ( .A1(n6641), .A2(n6578), .ZN(n5797) );
  XNOR2_X1 U3687 ( .A(n4388), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4397)
         );
  XNOR2_X1 U3688 ( .A(n3828), .B(n3827), .ZN(n5504) );
  NAND2_X1 U3689 ( .A1(n3825), .A2(n2987), .ZN(n3828) );
  OR2_X1 U3690 ( .A1(n5813), .A2(n3807), .ZN(n4396) );
  XNOR2_X1 U3691 ( .A(n3080), .B(n3808), .ZN(n4431) );
  NAND2_X1 U3692 ( .A1(n3772), .A2(n3771), .ZN(n3080) );
  NAND2_X1 U3693 ( .A1(n5617), .A2(n5807), .ZN(n3772) );
  NAND2_X1 U3694 ( .A1(n5616), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3771) );
  OR2_X1 U3695 ( .A1(n4418), .A2(n4417), .ZN(n5811) );
  NAND2_X1 U3696 ( .A1(n3018), .A2(n2986), .ZN(n5867) );
  INV_X1 U3697 ( .A(n5885), .ZN(n3018) );
  OR2_X1 U3698 ( .A1(n3792), .A2(n3465), .ZN(n6387) );
  CLKBUF_X1 U3699 ( .A(n4582), .Z(n4583) );
  NAND2_X1 U3701 ( .A1(n3610), .A2(n4496), .ZN(n4503) );
  NAND2_X1 U3702 ( .A1(n3431), .A2(n3461), .ZN(n3524) );
  NAND2_X1 U3703 ( .A1(n3478), .A2(n3477), .ZN(n3479) );
  INV_X1 U3704 ( .A(n3475), .ZN(n3480) );
  AOI21_X1 U3705 ( .B1(n3431), .B2(n3453), .A(n4603), .ZN(n3527) );
  AND2_X1 U3706 ( .A1(n6574), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3317)
         );
  AOI22_X1 U3707 ( .A1(n4027), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3396) );
  NAND2_X1 U3708 ( .A1(n3010), .A2(n4627), .ZN(n3671) );
  NAND2_X1 U3709 ( .A1(n3009), .A2(n3010), .ZN(n3696) );
  AND2_X1 U3710 ( .A1(n4627), .A2(n3673), .ZN(n3009) );
  INV_X1 U3711 ( .A(n3722), .ZN(n3720) );
  OR2_X1 U3712 ( .A1(n3693), .A2(n3692), .ZN(n3701) );
  OR2_X1 U3713 ( .A1(n3668), .A2(n3667), .ZN(n3698) );
  NAND2_X1 U3714 ( .A1(n3526), .A2(n3418), .ZN(n3513) );
  OR2_X1 U3715 ( .A1(n3547), .A2(n3546), .ZN(n3572) );
  NAND2_X1 U3716 ( .A1(n2971), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3328) );
  AOI21_X1 U3717 ( .B1(INSTQUEUE_REG_14__0__SCAN_IN), .B2(n3386), .A(n3151), 
        .ZN(n3172) );
  OR2_X1 U3718 ( .A1(n3409), .A2(n3147), .ZN(n3148) );
  AOI22_X1 U3719 ( .A1(n3466), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U3720 ( .A1(n4351), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3185) );
  INV_X1 U3721 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6789) );
  AOI22_X1 U3722 ( .A1(n3466), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U3723 ( .A1(n3412), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U3724 ( .A1(n4027), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U3725 ( .A1(n3387), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        INSTQUEUE_REG_4__5__SCAN_IN), .B2(n3474), .ZN(n3308) );
  AOI22_X1 U3726 ( .A1(n4351), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3311) );
  NOR2_X1 U3727 ( .A1(n4402), .A2(n3140), .ZN(n3139) );
  NAND2_X1 U3728 ( .A1(n5248), .A2(n5259), .ZN(n3140) );
  NOR2_X1 U3729 ( .A1(n5264), .A2(n4267), .ZN(n3065) );
  OR2_X1 U3730 ( .A1(n4266), .A2(n4265), .ZN(n4289) );
  NAND2_X1 U3731 ( .A1(n3131), .A2(n3060), .ZN(n3059) );
  AND2_X1 U3732 ( .A1(n3132), .A2(n5302), .ZN(n3131) );
  INV_X1 U3733 ( .A(n3061), .ZN(n3060) );
  NAND2_X1 U3734 ( .A1(n3062), .A2(n4166), .ZN(n3061) );
  INV_X1 U3735 ( .A(n3063), .ZN(n3062) );
  INV_X1 U3736 ( .A(n4334), .ZN(n4366) );
  NOR2_X1 U3737 ( .A1(n4113), .A2(n3073), .ZN(n3072) );
  NAND2_X1 U3738 ( .A1(n5401), .A2(n3130), .ZN(n3129) );
  CLKBUF_X1 U3739 ( .A(n5434), .Z(n5435) );
  INV_X1 U3740 ( .A(n3908), .ZN(n4339) );
  INV_X1 U3741 ( .A(n3363), .ZN(n3032) );
  NAND2_X1 U3742 ( .A1(n5745), .A2(n3756), .ZN(n3760) );
  INV_X1 U3743 ( .A(n3761), .ZN(n3105) );
  INV_X1 U3744 ( .A(n5404), .ZN(n3245) );
  AND2_X1 U3745 ( .A1(n3122), .A2(n3121), .ZN(n3120) );
  INV_X1 U3746 ( .A(n5527), .ZN(n3121) );
  INV_X1 U3747 ( .A(n3274), .ZN(n3232) );
  NAND2_X1 U3748 ( .A1(n3204), .A2(n6230), .ZN(n3194) );
  OAI21_X1 U3749 ( .B1(n3345), .B2(n3344), .A(n2997), .ZN(n3033) );
  AND2_X1 U3750 ( .A1(n3361), .A2(n3360), .ZN(n3034) );
  AOI21_X1 U3751 ( .B1(n3362), .B2(n3353), .A(n3352), .ZN(n3361) );
  NAND2_X1 U3752 ( .A1(n2992), .A2(n3036), .ZN(n3028) );
  AOI21_X1 U3753 ( .B1(n3634), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3605), 
        .ZN(n3609) );
  INV_X1 U3754 ( .A(n3604), .ZN(n3605) );
  XNOR2_X1 U3755 ( .A(n4496), .B(n4674), .ZN(n4580) );
  OR2_X1 U3756 ( .A1(n4858), .A2(n4859), .ZN(n6398) );
  BUF_X1 U3757 ( .A(n3550), .Z(n3634) );
  AND4_X2 U3758 ( .A1(n3385), .A2(n3384), .A3(n3383), .A4(n3382), .ZN(n3423)
         );
  NOR2_X1 U3759 ( .A1(n3377), .A2(n3376), .ZN(n3383) );
  INV_X1 U3760 ( .A(n3561), .ZN(n4795) );
  INV_X1 U3761 ( .A(n4469), .ZN(n6713) );
  AND2_X1 U3762 ( .A1(n3557), .A2(n3435), .ZN(n4459) );
  AND2_X1 U3763 ( .A1(n3447), .A2(n3446), .ZN(n4458) );
  NAND2_X1 U3764 ( .A1(n3552), .A2(n2971), .ZN(n4456) );
  AND2_X1 U3765 ( .A1(n5295), .A2(n3838), .ZN(n5254) );
  OR3_X1 U3766 ( .A1(n5352), .A2(n6682), .A3(n5691), .ZN(n5319) );
  INV_X1 U3767 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6755) );
  INV_X1 U3768 ( .A(n5250), .ZN(n3822) );
  AND2_X1 U3769 ( .A1(n3230), .A2(n3229), .ZN(n5970) );
  NAND2_X1 U3770 ( .A1(n5452), .A2(n3122), .ZN(n5973) );
  NOR2_X1 U3771 ( .A1(n3137), .A2(n3136), .ZN(n3135) );
  INV_X1 U3772 ( .A(n3139), .ZN(n3137) );
  INV_X1 U3773 ( .A(n4424), .ZN(n3136) );
  CLKBUF_X1 U3774 ( .A(n4877), .Z(n4878) );
  AOI21_X1 U3775 ( .B1(n3905), .B2(n4018), .A(n3904), .ZN(n4852) );
  INV_X1 U3776 ( .A(n3903), .ZN(n3904) );
  INV_X1 U3777 ( .A(n3898), .ZN(n3905) );
  CLKBUF_X1 U3778 ( .A(n4850), .Z(n4851) );
  NAND2_X1 U3779 ( .A1(n4858), .A2(n4018), .ZN(n3887) );
  INV_X1 U3780 ( .A(n4274), .ZN(n4275) );
  AND2_X1 U3781 ( .A1(n3076), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3075)
         );
  INV_X1 U3782 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5292) );
  OR2_X1 U3783 ( .A1(n4247), .A2(n5292), .ZN(n4274) );
  CLKBUF_X1 U3784 ( .A(n5284), .Z(n5285) );
  INV_X1 U3785 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4184) );
  INV_X1 U3786 ( .A(n4182), .ZN(n4183) );
  NAND2_X1 U3787 ( .A1(n4183), .A2(n3076), .ZN(n4246) );
  OR2_X1 U3788 ( .A1(n4149), .A2(n6788), .ZN(n4182) );
  INV_X1 U3789 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6788) );
  OR2_X1 U3790 ( .A1(n3064), .A2(n5368), .ZN(n3063) );
  INV_X1 U3791 ( .A(n5360), .ZN(n3064) );
  AND3_X1 U3792 ( .A1(n3955), .A2(n3954), .A3(n3953), .ZN(n5467) );
  OR2_X1 U3793 ( .A1(n3915), .A2(n3914), .ZN(n3923) );
  NAND2_X1 U3794 ( .A1(n3906), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3915)
         );
  NOR2_X1 U3795 ( .A1(n3899), .A2(n6185), .ZN(n3906) );
  AND2_X1 U3796 ( .A1(n3891), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3892)
         );
  NAND2_X1 U3797 ( .A1(n3892), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3899)
         );
  CLKBUF_X1 U3798 ( .A(n4547), .Z(n4548) );
  AND2_X1 U3799 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3891) );
  NAND2_X1 U3800 ( .A1(n3049), .A2(n4225), .ZN(n4546) );
  AND2_X1 U3801 ( .A1(n3627), .A2(n4018), .ZN(n3050) );
  OAI22_X1 U3802 ( .A1(n3823), .A2(n3190), .B1(n5261), .B2(n3109), .ZN(n4418)
         );
  NAND2_X1 U3803 ( .A1(n3111), .A2(n3110), .ZN(n3109) );
  NOR2_X1 U3804 ( .A1(n5249), .A2(n4414), .ZN(n3110) );
  INV_X1 U3805 ( .A(n5262), .ZN(n3111) );
  NAND2_X1 U3806 ( .A1(n3042), .A2(n3041), .ZN(n5643) );
  AOI21_X1 U3807 ( .B1(n3043), .B2(n3046), .A(n2989), .ZN(n3041) );
  AND2_X1 U3808 ( .A1(n3265), .A2(n3264), .ZN(n5304) );
  AND2_X1 U3809 ( .A1(n3126), .A2(n3125), .ZN(n3124) );
  INV_X1 U3810 ( .A(n5317), .ZN(n3125) );
  NAND2_X1 U3811 ( .A1(n3091), .A2(n5680), .ZN(n3090) );
  INV_X1 U3812 ( .A(n5689), .ZN(n3091) );
  NAND2_X1 U3813 ( .A1(n5346), .A2(n3126), .ZN(n5338) );
  AND2_X1 U3814 ( .A1(n3257), .A2(n3256), .ZN(n5345) );
  AND2_X1 U3815 ( .A1(n5346), .A2(n5345), .ZN(n5348) );
  AND2_X1 U3816 ( .A1(n3239), .A2(n3238), .ZN(n5444) );
  AND2_X1 U3817 ( .A1(n5452), .A2(n3120), .ZN(n5528) );
  INV_X1 U3818 ( .A(n3013), .ZN(n3012) );
  INV_X1 U3819 ( .A(n3756), .ZN(n3014) );
  NOR2_X1 U3820 ( .A1(n3114), .A2(n5472), .ZN(n3113) );
  INV_X1 U3821 ( .A(n3115), .ZN(n3114) );
  NAND2_X1 U3822 ( .A1(n4664), .A2(n3023), .ZN(n5992) );
  NOR2_X1 U3823 ( .A1(n3024), .A2(n3796), .ZN(n3023) );
  NOR2_X1 U3824 ( .A1(n3118), .A2(n4847), .ZN(n3117) );
  INV_X1 U3825 ( .A(n3143), .ZN(n3118) );
  INV_X1 U3826 ( .A(n3039), .ZN(n3038) );
  AND2_X1 U3827 ( .A1(n3633), .A2(n6874), .ZN(n3037) );
  NAND2_X1 U3828 ( .A1(n6392), .A2(n3800), .ZN(n5936) );
  OR2_X1 U3829 ( .A1(n3551), .A2(n6713), .ZN(n4798) );
  NAND2_X1 U3830 ( .A1(n3201), .A2(n3274), .ZN(n4872) );
  CLKBUF_X1 U3831 ( .A(n3863), .Z(n5498) );
  OR2_X1 U3832 ( .A1(n6024), .A2(n4627), .ZN(n4695) );
  NAND2_X1 U3833 ( .A1(n3399), .A2(n3426), .ZN(n4759) );
  INV_X1 U3834 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4747) );
  NAND2_X1 U3835 ( .A1(n4485), .A2(n4484), .ZN(n4782) );
  NOR2_X1 U3836 ( .A1(n6398), .A2(n6021), .ZN(n5015) );
  AND2_X1 U3837 ( .A1(n3635), .A2(n4619), .ZN(n6476) );
  CLKBUF_X1 U3838 ( .A(n4580), .Z(n4581) );
  INV_X1 U3839 ( .A(n6398), .ZN(n6396) );
  AND3_X1 U3840 ( .A1(n6519), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4802) );
  INV_X1 U3841 ( .A(n4695), .ZN(n4630) );
  NAND2_X1 U3842 ( .A1(n4858), .A2(n6024), .ZN(n6514) );
  OR2_X1 U3843 ( .A1(n6018), .A2(n6050), .ZN(n4618) );
  NOR2_X1 U3844 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n4577) );
  AND2_X1 U3845 ( .A1(n6722), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4377) );
  INV_X1 U3846 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6435) );
  NAND2_X1 U3847 ( .A1(n3986), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4019)
         );
  INV_X1 U3848 ( .A(n6896), .ZN(n6188) );
  NAND2_X1 U3849 ( .A1(n5484), .A2(n3836), .ZN(n6206) );
  INV_X1 U3850 ( .A(n6889), .ZN(n6223) );
  INV_X1 U3851 ( .A(n6186), .ZN(n6894) );
  NAND2_X1 U3852 ( .A1(n6206), .A2(n6197), .ZN(n6170) );
  OR2_X1 U3853 ( .A1(n5251), .A2(n5250), .ZN(n5508) );
  OR2_X1 U3854 ( .A1(n5552), .A2(n5511), .ZN(n3053) );
  INV_X1 U3855 ( .A(n5557), .ZN(n6232) );
  OR2_X1 U3856 ( .A1(n4525), .A2(n4410), .ZN(n4411) );
  OR3_X1 U3857 ( .A1(n4492), .A2(n4455), .A3(n4506), .ZN(n4412) );
  CLKBUF_X1 U3858 ( .A(n4733), .Z(n4734) );
  AOI21_X1 U3859 ( .B1(n4527), .B2(n5208), .A(n4526), .ZN(n4528) );
  INV_X1 U3860 ( .A(n5613), .ZN(n5180) );
  OR3_X1 U3861 ( .A1(n4534), .A2(n4533), .A3(n6716), .ZN(n6269) );
  AND2_X1 U3862 ( .A1(n4761), .A2(n4798), .ZN(n4533) );
  OR3_X2 U3863 ( .A1(n4534), .A2(READY_N), .A3(n4473), .ZN(n6324) );
  OR2_X1 U3864 ( .A1(n4534), .A2(n4798), .ZN(n6327) );
  INV_X1 U3865 ( .A(n6327), .ZN(n6322) );
  INV_X1 U3866 ( .A(n5247), .ZN(n3056) );
  OR2_X1 U3867 ( .A1(n5301), .A2(n5316), .ZN(n5673) );
  NAND2_X1 U3868 ( .A1(n4112), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4114)
         );
  NAND2_X1 U3869 ( .A1(n4061), .A2(n3071), .ZN(n4090) );
  NAND2_X1 U3870 ( .A1(n3986), .A2(n3067), .ZN(n4021) );
  INV_X1 U3871 ( .A(n3820), .ZN(n6368) );
  INV_X1 U3872 ( .A(n6101), .ZN(n6336) );
  OR2_X1 U3873 ( .A1(n4393), .A2(n4392), .ZN(n4394) );
  AND2_X1 U3874 ( .A1(n5845), .A2(n5836), .ZN(n5829) );
  NOR2_X1 U3875 ( .A1(n5867), .A2(n3803), .ZN(n5855) );
  NAND2_X1 U3876 ( .A1(n3086), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3083) );
  OR2_X1 U3877 ( .A1(n5688), .A2(n3082), .ZN(n3081) );
  OAI211_X1 U3878 ( .C1(n5688), .C2(n3088), .A(n3085), .B(n6853), .ZN(n3084)
         );
  NAND2_X1 U3879 ( .A1(n3021), .A2(n3019), .ZN(n5885) );
  OR2_X1 U3880 ( .A1(n5991), .A2(n3795), .ZN(n3021) );
  AOI21_X1 U3881 ( .B1(n3020), .B2(n3005), .A(n5890), .ZN(n3019) );
  AND2_X1 U3882 ( .A1(n5928), .A2(n3817), .ZN(n5908) );
  OR2_X1 U3883 ( .A1(n6348), .A2(n5935), .ZN(n5945) );
  NAND2_X1 U3884 ( .A1(n3079), .A2(n3751), .ZN(n5780) );
  NAND2_X1 U3885 ( .A1(n3107), .A2(n3750), .ZN(n5791) );
  NAND2_X1 U3886 ( .A1(n3094), .A2(n3705), .ZN(n5055) );
  NAND2_X1 U3887 ( .A1(n4664), .A2(n5056), .ZN(n4841) );
  AND2_X1 U3888 ( .A1(n5995), .A2(n4553), .ZN(n6367) );
  OR2_X1 U3889 ( .A1(n3792), .A2(n4506), .ZN(n6372) );
  INV_X1 U3890 ( .A(n6387), .ZN(n6359) );
  OR2_X1 U3891 ( .A1(n3792), .A2(n4761), .ZN(n6392) );
  AND2_X2 U3892 ( .A1(n4472), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5194)
         );
  AND2_X2 U3893 ( .A1(n3146), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5187)
         );
  INV_X1 U3894 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4768) );
  NAND2_X1 U3895 ( .A1(n4492), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6036) );
  INV_X1 U3896 ( .A(n5045), .ZN(n4943) );
  INV_X1 U3897 ( .A(n4918), .ZN(n4946) );
  INV_X1 U3898 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5022) );
  INV_X1 U3899 ( .A(n6436), .ZN(n6460) );
  NAND2_X1 U3900 ( .A1(n4700), .A2(n5014), .ZN(n6468) );
  NAND2_X1 U3901 ( .A1(n4630), .A2(n6042), .ZN(n6474) );
  INV_X1 U3902 ( .A(n6507), .ZN(n6479) );
  INV_X1 U3903 ( .A(n6083), .ZN(n6091) );
  NOR2_X2 U3904 ( .A1(n4885), .A2(n5014), .ZN(n6503) );
  INV_X1 U3905 ( .A(n6529), .ZN(n6593) );
  INV_X1 U3906 ( .A(n6534), .ZN(n6599) );
  INV_X1 U3907 ( .A(n6539), .ZN(n6605) );
  INV_X1 U3908 ( .A(n6544), .ZN(n6611) );
  INV_X1 U3909 ( .A(n6549), .ZN(n6617) );
  OAI22_X1 U3910 ( .A1(n4959), .A2(n4958), .B1(n5165), .B2(n4957), .ZN(n4990)
         );
  AND2_X1 U3911 ( .A1(n4953), .A2(n4587), .ZN(n6633) );
  NOR2_X1 U3912 ( .A1(n4678), .A2(n4677), .ZN(n5075) );
  NAND2_X1 U3913 ( .A1(n4953), .A2(n5014), .ZN(n5100) );
  OR2_X1 U3914 ( .A1(n4618), .A2(n4603), .ZN(n6539) );
  NAND2_X1 U3915 ( .A1(n4673), .A2(n6508), .ZN(n4941) );
  OR2_X1 U3916 ( .A1(n4618), .A2(n5558), .ZN(n6560) );
  INV_X1 U3917 ( .A(n4941), .ZN(n4868) );
  OAI211_X1 U3918 ( .C1(n4676), .C2(n6437), .A(n4592), .B(n6400), .ZN(n4616)
         );
  NOR2_X1 U3919 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5164) );
  AND2_X1 U3920 ( .A1(n6673), .A2(n4446), .ZN(n6702) );
  AND2_X1 U3921 ( .A1(n6645), .A2(STATE_REG_1__SCAN_IN), .ZN(n6099) );
  OR2_X1 U3922 ( .A1(n3854), .A2(n3853), .ZN(n3855) );
  OR2_X1 U3923 ( .A1(n5562), .A2(n5481), .ZN(n5240) );
  AND2_X1 U3924 ( .A1(n4421), .A2(n4420), .ZN(n4422) );
  NAND2_X1 U3925 ( .A1(n3054), .A2(n3051), .ZN(U2832) );
  INV_X1 U3926 ( .A(n3052), .ZN(n3051) );
  NAND2_X1 U3927 ( .A1(n5639), .A2(n6233), .ZN(n3054) );
  OAI21_X1 U3928 ( .B1(n5510), .B2(n5557), .A(n3053), .ZN(n3052) );
  NAND2_X1 U3929 ( .A1(n3011), .A2(n2984), .ZN(U2955) );
  OAI21_X1 U3930 ( .B1(n4431), .B2(n6101), .A(n3047), .ZN(U2956) );
  INV_X1 U3931 ( .A(n4429), .ZN(n4430) );
  AOI21_X1 U3932 ( .B1(n5630), .B2(n5804), .A(n5629), .ZN(n5631) );
  OAI211_X1 U3933 ( .C1(n4431), .C2(n6015), .A(n3022), .B(n2975), .ZN(U2988)
         );
  OR2_X1 U3934 ( .A1(n3809), .A2(n3808), .ZN(n3022) );
  INV_X1 U3935 ( .A(n4396), .ZN(n3809) );
  AND2_X1 U3936 ( .A1(n4667), .A2(n4669), .ZN(n3119) );
  INV_X1 U3937 ( .A(n3422), .ZN(n3400) );
  INV_X2 U3938 ( .A(n3466), .ZN(n3467) );
  NAND2_X1 U3939 ( .A1(n2983), .A2(n5450), .ZN(n5449) );
  NOR2_X1 U3940 ( .A1(n5367), .A2(n3061), .ZN(n5327) );
  AND4_X1 U3941 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n2973)
         );
  NOR3_X1 U3942 ( .A1(n5261), .A2(n5262), .A3(n3001), .ZN(n3108) );
  NOR2_X1 U3943 ( .A1(n2994), .A2(n3821), .ZN(n2975) );
  AND2_X1 U3944 ( .A1(n3670), .A2(n3669), .ZN(n3672) );
  NAND2_X1 U3945 ( .A1(n3119), .A2(n3143), .ZN(n4689) );
  AOI21_X1 U3946 ( .B1(n4587), .B2(n3862), .A(n5165), .ZN(n4515) );
  AND2_X1 U3947 ( .A1(n3067), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n2976)
         );
  AND2_X1 U3948 ( .A1(n3057), .A2(n5542), .ZN(n2977) );
  INV_X1 U3949 ( .A(n3119), .ZN(n4668) );
  NOR2_X1 U3950 ( .A1(n5389), .A2(n3129), .ZN(n2978) );
  NAND2_X1 U3951 ( .A1(n3720), .A2(n3719), .ZN(n3741) );
  INV_X1 U3952 ( .A(n3431), .ZN(n3516) );
  NOR2_X1 U3953 ( .A1(n5367), .A2(n5368), .ZN(n5359) );
  AND2_X1 U3954 ( .A1(n5327), .A2(n3132), .ZN(n5301) );
  OR2_X1 U3955 ( .A1(n5416), .A2(n3129), .ZN(n5387) );
  AND2_X1 U3956 ( .A1(n5327), .A2(n4181), .ZN(n5314) );
  AND2_X1 U3957 ( .A1(n3941), .A2(n3057), .ZN(n2979) );
  AND4_X1 U3958 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .ZN(n2980)
         );
  NAND2_X1 U3959 ( .A1(n3941), .A2(n3940), .ZN(n5466) );
  OAI21_X1 U3960 ( .B1(n5736), .B2(n3762), .A(n3761), .ZN(n5711) );
  AND2_X1 U3961 ( .A1(n3077), .A2(n3752), .ZN(n2981) );
  OR2_X1 U3962 ( .A1(n5261), .A2(n5262), .ZN(n2982) );
  AND2_X1 U3963 ( .A1(n3941), .A2(n2977), .ZN(n2983) );
  OR2_X1 U3964 ( .A1(n5367), .A2(n3063), .ZN(n5342) );
  NAND2_X1 U3965 ( .A1(n3452), .A2(n3402), .ZN(n3526) );
  XNOR2_X1 U3966 ( .A(n3741), .B(n3732), .ZN(n3920) );
  AND2_X1 U3967 ( .A1(n4390), .A2(n4389), .ZN(n2984) );
  AND2_X1 U3968 ( .A1(n3728), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n2985)
         );
  NAND2_X1 U3969 ( .A1(n5936), .A2(n5873), .ZN(n2986) );
  NAND2_X1 U3970 ( .A1(n3823), .A2(n3201), .ZN(n2987) );
  NAND2_X1 U3971 ( .A1(n5760), .A2(n5907), .ZN(n2988) );
  NOR2_X1 U3972 ( .A1(n3422), .A2(n3421), .ZN(n3509) );
  NOR2_X1 U3973 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n2989)
         );
  AND4_X1 U3974 ( .A1(n3473), .A2(n3472), .A3(n3471), .A4(n3470), .ZN(n2990)
         );
  NAND2_X1 U3975 ( .A1(n3079), .A2(n3077), .ZN(n2991) );
  NOR2_X1 U3976 ( .A1(n3332), .A2(n3331), .ZN(n2992) );
  INV_X1 U3977 ( .A(n3086), .ZN(n3085) );
  NOR2_X1 U3978 ( .A1(n5690), .A2(n3087), .ZN(n3086) );
  AND2_X1 U3979 ( .A1(n3102), .A2(n2988), .ZN(n2993) );
  NOR2_X1 U3980 ( .A1(n5507), .A2(n6387), .ZN(n2994) );
  AND2_X1 U3981 ( .A1(n3784), .A2(n3510), .ZN(n2995) );
  AND2_X1 U3982 ( .A1(n3120), .A2(n5444), .ZN(n2996) );
  NAND2_X1 U3983 ( .A1(n3731), .A2(n3350), .ZN(n2997) );
  BUF_X1 U3984 ( .A(n3423), .Z(n4588) );
  NAND2_X1 U3985 ( .A1(n5452), .A2(n5453), .ZN(n5451) );
  NAND2_X1 U3986 ( .A1(n3880), .A2(n3879), .ZN(n4544) );
  NAND2_X1 U3987 ( .A1(n5554), .A2(n3115), .ZN(n5470) );
  INV_X1 U3988 ( .A(n5249), .ZN(n3112) );
  AND2_X1 U3989 ( .A1(n3277), .A2(n3276), .ZN(n5249) );
  NAND2_X1 U3990 ( .A1(n5554), .A2(n5553), .ZN(n5547) );
  NOR2_X1 U3991 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n2998)
         );
  NAND2_X1 U3992 ( .A1(n3008), .A2(n3740), .ZN(n5798) );
  AND2_X1 U3993 ( .A1(n3986), .A2(n2976), .ZN(n2999) );
  AND2_X1 U3994 ( .A1(n4003), .A2(n5450), .ZN(n3000) );
  OAI21_X1 U3995 ( .B1(n3912), .B2(n4052), .A(n3911), .ZN(n4876) );
  OAI21_X1 U3996 ( .B1(n3731), .B2(n4945), .A(n3694), .ZN(n3695) );
  INV_X1 U3997 ( .A(n3695), .ZN(n3134) );
  NAND2_X1 U3998 ( .A1(n4733), .A2(n3876), .ZN(n4543) );
  INV_X1 U3999 ( .A(n4166), .ZN(n5344) );
  NAND2_X1 U4000 ( .A1(n3112), .A2(n4413), .ZN(n3001) );
  INV_X1 U4001 ( .A(n3089), .ZN(n3088) );
  NOR2_X1 U4002 ( .A1(n5663), .A2(n2998), .ZN(n3089) );
  INV_X1 U4003 ( .A(n4018), .ZN(n4052) );
  NOR2_X1 U4004 ( .A1(n3401), .A2(n5165), .ZN(n4018) );
  NAND2_X1 U4005 ( .A1(n3861), .A2(n3860), .ZN(n4731) );
  AND2_X1 U4006 ( .A1(n2977), .A2(n3000), .ZN(n3002) );
  INV_X1 U4007 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6722) );
  INV_X2 U4008 ( .A(n5797), .ZN(n5804) );
  AND2_X1 U4009 ( .A1(n4856), .A2(n4855), .ZN(n4667) );
  AND2_X1 U4010 ( .A1(n3071), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3003)
         );
  INV_X1 U4011 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6131) );
  AND2_X1 U4012 ( .A1(n3072), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3004)
         );
  OR2_X1 U4013 ( .A1(n3816), .A2(n5872), .ZN(n3005) );
  INV_X1 U4014 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3073) );
  AND2_X1 U4015 ( .A1(n3065), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3006)
         );
  INV_X1 U4016 ( .A(n5056), .ZN(n3024) );
  INV_X1 U4017 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3074) );
  INV_X1 U4018 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3069) );
  CLKBUF_X1 U4019 ( .A(n6459), .Z(n3007) );
  AND2_X2 U4020 ( .A1(n4745), .A2(n4502), .ZN(n3412) );
  NAND2_X1 U4021 ( .A1(n5182), .A2(n5183), .ZN(n3008) );
  NAND2_X1 U4022 ( .A1(n3092), .A2(n3093), .ZN(n5182) );
  NAND3_X1 U4023 ( .A1(n3784), .A2(n3510), .A3(n3512), .ZN(n3514) );
  OAI21_X1 U4024 ( .B1(n2981), .B2(n3014), .A(n3759), .ZN(n3013) );
  OAI21_X2 U4025 ( .B1(n3079), .B2(n3014), .A(n3012), .ZN(n5736) );
  NAND2_X2 U4026 ( .A1(n3426), .A2(n4599), .ZN(n3506) );
  OAI211_X1 U4027 ( .C1(n3426), .C2(n3423), .A(n4599), .B(n3427), .ZN(n3508)
         );
  NAND2_X1 U4028 ( .A1(n5931), .A2(n3799), .ZN(n5888) );
  INV_X1 U4029 ( .A(n3344), .ZN(n3036) );
  AOI21_X1 U4030 ( .B1(n6024), .B2(n3633), .A(n3038), .ZN(n6332) );
  OAI21_X1 U4031 ( .B1(n6024), .B2(n3726), .A(n3037), .ZN(n6333) );
  AOI21_X1 U4032 ( .B1(n3633), .B2(n3726), .A(n6874), .ZN(n3039) );
  OR2_X1 U4033 ( .A1(n5705), .A2(n3046), .ZN(n3040) );
  NAND2_X1 U4034 ( .A1(n5705), .A2(n3043), .ZN(n3042) );
  NAND2_X1 U4035 ( .A1(n3048), .A2(n3622), .ZN(n3624) );
  NAND3_X1 U4036 ( .A1(n3610), .A2(n4496), .A3(n6722), .ZN(n3048) );
  NAND2_X1 U4037 ( .A1(n3657), .A2(n3627), .ZN(n6024) );
  NAND2_X1 U4038 ( .A1(n3050), .A2(n3657), .ZN(n3049) );
  NAND2_X1 U4039 ( .A1(n3941), .A2(n3002), .ZN(n5434) );
  OR2_X2 U4040 ( .A1(n5367), .A2(n3059), .ZN(n5284) );
  NAND2_X1 U4041 ( .A1(n4275), .A2(n3006), .ZN(n4315) );
  NAND2_X1 U4042 ( .A1(n4112), .A2(n3004), .ZN(n4149) );
  NAND2_X1 U4043 ( .A1(n4183), .A2(n3075), .ZN(n4247) );
  NAND3_X1 U4044 ( .A1(n3084), .A2(n3083), .A3(n3081), .ZN(n5861) );
  OR2_X2 U4045 ( .A1(n5690), .A2(n3090), .ZN(n5670) );
  NOR2_X2 U4046 ( .A1(n5690), .A2(n5689), .ZN(n5688) );
  NAND3_X1 U4047 ( .A1(n4837), .A2(n4838), .A3(n5054), .ZN(n3092) );
  AOI21_X1 U4048 ( .B1(n5054), .B2(n3095), .A(n2985), .ZN(n3093) );
  NAND2_X1 U4049 ( .A1(n4837), .A2(n4838), .ZN(n3094) );
  INV_X1 U4050 ( .A(n3705), .ZN(n3095) );
  OAI21_X2 U4051 ( .B1(n3760), .B2(n3099), .A(n3096), .ZN(n3100) );
  INV_X1 U4052 ( .A(n3100), .ZN(n5660) );
  XNOR2_X2 U4053 ( .A(n4627), .B(n3657), .ZN(n4858) );
  INV_X1 U4054 ( .A(n2970), .ZN(n3823) );
  NAND2_X1 U4055 ( .A1(n3117), .A2(n3119), .ZN(n4996) );
  NAND2_X1 U4056 ( .A1(n5346), .A2(n3124), .ZN(n5303) );
  INV_X2 U4057 ( .A(n4558), .ZN(n4410) );
  AND2_X2 U4058 ( .A1(n3190), .A2(n4558), .ZN(n3204) );
  AND2_X2 U4059 ( .A1(n2971), .A2(n3422), .ZN(n4558) );
  XNOR2_X1 U4060 ( .A(n3570), .B(n3127), .ZN(n3856) );
  OAI21_X1 U4061 ( .B1(n4582), .B2(STATE2_REG_0__SCAN_IN), .A(n3569), .ZN(
        n3127) );
  INV_X1 U4062 ( .A(n5434), .ZN(n4059) );
  NOR2_X1 U4063 ( .A1(n5416), .A2(n5417), .ZN(n5400) );
  INV_X1 U4064 ( .A(n5417), .ZN(n3130) );
  INV_X1 U4065 ( .A(n5284), .ZN(n4251) );
  NAND2_X1 U4066 ( .A1(n5260), .A2(n3135), .ZN(n4373) );
  AND2_X1 U4067 ( .A1(n5260), .A2(n5259), .ZN(n5247) );
  NAND2_X1 U4068 ( .A1(n5260), .A2(n3138), .ZN(n4401) );
  NAND2_X1 U4069 ( .A1(n5403), .A2(n3245), .ZN(n5370) );
  OAI22_X2 U4070 ( .A1(n4662), .A2(n4661), .B1(n3656), .B2(n4666), .ZN(n4688)
         );
  OAI211_X1 U4071 ( .C1(n3822), .C2(n2970), .A(n3824), .B(n2987), .ZN(n3281)
         );
  NOR2_X2 U4072 ( .A1(n5419), .A2(n5422), .ZN(n5403) );
  NAND2_X1 U4073 ( .A1(n4426), .A2(n5804), .ZN(n4432) );
  INV_X1 U4074 ( .A(n4625), .ZN(n3896) );
  NAND2_X2 U4075 ( .A1(n5213), .A2(n4531), .ZN(n5591) );
  OR2_X1 U4076 ( .A1(n5760), .A2(n6841), .ZN(n3141) );
  INV_X1 U4077 ( .A(n4587), .ZN(n5014) );
  AND4_X1 U4078 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3142)
         );
  OR2_X1 U4079 ( .A1(n3207), .A2(n3206), .ZN(n3143) );
  NAND2_X1 U4080 ( .A1(n4617), .A2(n3461), .ZN(n3573) );
  AND2_X1 U4081 ( .A1(n5552), .A2(n4530), .ZN(n6233) );
  INV_X1 U4082 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4784) );
  INV_X1 U4083 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3914) );
  INV_X1 U4084 ( .A(n5552), .ZN(n5518) );
  NAND2_X2 U4085 ( .A1(n4412), .A2(n4411), .ZN(n5552) );
  AND4_X1 U4086 ( .A1(n3407), .A2(n3406), .A3(n3405), .A4(n3404), .ZN(n3144)
         );
  CLKBUF_X3 U4087 ( .A(n4351), .Z(n4198) );
  CLKBUF_X3 U4088 ( .A(n3507), .Z(n3190) );
  INV_X1 U4089 ( .A(n5327), .ZN(n5343) );
  AND2_X1 U4090 ( .A1(n3442), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3324) );
  INV_X1 U4091 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3147) );
  NAND2_X1 U4092 ( .A1(n3341), .A2(n3340), .ZN(n3349) );
  OR2_X1 U4093 ( .A1(n3408), .A2(n5022), .ZN(n3150) );
  OR2_X1 U4094 ( .A1(n4233), .A2(n4232), .ZN(n4252) );
  INV_X1 U4095 ( .A(n3721), .ZN(n3719) );
  OR2_X1 U4096 ( .A1(n3621), .A2(n3620), .ZN(n3628) );
  AOI22_X1 U4097 ( .A1(n3386), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4098 ( .A1(n3412), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U4099 ( .A1(n4351), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3295) );
  INV_X1 U4100 ( .A(n3672), .ZN(n3673) );
  INV_X1 U4101 ( .A(n5534), .ZN(n4003) );
  OR2_X1 U4102 ( .A1(n3716), .A2(n3715), .ZN(n3734) );
  OR2_X1 U4103 ( .A1(n3356), .A2(n3355), .ZN(n3359) );
  AND4_X1 U4104 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n3169)
         );
  OR2_X1 U4105 ( .A1(n4224), .A2(n4223), .ZN(n4231) );
  INV_X1 U4106 ( .A(n3452), .ZN(n3454) );
  INV_X1 U4107 ( .A(n3913), .ZN(n3882) );
  OR2_X1 U4108 ( .A1(n3648), .A2(n3647), .ZN(n3652) );
  AND2_X1 U4109 ( .A1(n3359), .A2(n3358), .ZN(n3440) );
  INV_X1 U4110 ( .A(n3609), .ZN(n3606) );
  INV_X1 U4111 ( .A(n3551), .ZN(n3552) );
  INV_X1 U4112 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4113) );
  INV_X1 U4113 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6776) );
  INV_X1 U4114 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6144) );
  INV_X1 U4115 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3808) );
  NAND2_X1 U4116 ( .A1(n3362), .A2(n3440), .ZN(n3363) );
  INV_X1 U4117 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4769) );
  OR2_X1 U4118 ( .A1(n5395), .A2(n3841), .ZN(n5352) );
  INV_X1 U4119 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6185) );
  AND2_X1 U4120 ( .A1(n6197), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5484) );
  INV_X1 U4121 ( .A(n5403), .ZN(n5420) );
  INV_X1 U4123 ( .A(n4250), .ZN(n5287) );
  AND2_X1 U4124 ( .A1(n3241), .A2(n3240), .ZN(n5422) );
  INV_X1 U4125 ( .A(n5662), .ZN(n5789) );
  NAND2_X1 U4126 ( .A1(n6036), .A2(n4578), .ZN(n4579) );
  OR2_X1 U4127 ( .A1(n4581), .A2(n6481), .ZN(n5006) );
  OR2_X1 U4128 ( .A1(n4581), .A2(n6046), .ZN(n6399) );
  NOR2_X1 U4129 ( .A1(n4695), .A2(n6021), .ZN(n4700) );
  INV_X1 U4130 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6519) );
  OR2_X1 U4131 ( .A1(n6514), .A2(n6021), .ZN(n4885) );
  OR2_X1 U4132 ( .A1(n4503), .A2(n6218), .ZN(n6580) );
  INV_X1 U4133 ( .A(n6580), .ZN(n4950) );
  INV_X1 U4134 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6050) );
  OR2_X1 U4135 ( .A1(n4618), .A2(n4595), .ZN(n6549) );
  INV_X1 U4136 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4786) );
  OR2_X1 U4137 ( .A1(n4534), .A2(n4456), .ZN(n4465) );
  INV_X1 U4138 ( .A(n4378), .ZN(n6724) );
  AND2_X1 U4139 ( .A1(n6197), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5223) );
  OR2_X1 U4140 ( .A1(n5552), .A2(n4419), .ZN(n4420) );
  AND2_X1 U4141 ( .A1(n3248), .A2(n3247), .ZN(n5374) );
  NOR2_X2 U4142 ( .A1(n4996), .A2(n4995), .ZN(n5554) );
  NOR2_X2 U4143 ( .A1(n5612), .A2(n5216), .ZN(n5597) );
  NOR2_X1 U4144 ( .A1(n6269), .A2(n3530), .ZN(n6239) );
  INV_X1 U4145 ( .A(n6269), .ZN(n6251) );
  INV_X2 U4146 ( .A(n6253), .ZN(n6266) );
  INV_X1 U4147 ( .A(n6273), .ZN(n6320) );
  OR2_X1 U4148 ( .A1(n3551), .A2(n4410), .ZN(n4473) );
  NOR2_X1 U4149 ( .A1(n5945), .A2(n3815), .ZN(n5928) );
  INV_X1 U4150 ( .A(n6015), .ZN(n6381) );
  INV_X1 U4151 ( .A(n6437), .ZN(n6578) );
  INV_X1 U4152 ( .A(n5120), .ZN(n5154) );
  OAI21_X1 U4153 ( .B1(n6405), .B2(n6404), .A(n6403), .ZN(n6428) );
  OAI211_X1 U4154 ( .C1(n6443), .C2(n6442), .A(n6441), .B(n6440), .ZN(n6461)
         );
  OAI211_X1 U4155 ( .C1(n6437), .C2(n6434), .A(n4704), .B(n6400), .ZN(n4727)
         );
  INV_X1 U4156 ( .A(n6474), .ZN(n4834) );
  OAI211_X1 U4157 ( .C1(n4802), .C2(n6437), .A(n4634), .B(n6400), .ZN(n4657)
         );
  AND2_X1 U4158 ( .A1(n6021), .A2(n5014), .ZN(n6508) );
  OAI211_X1 U4159 ( .C1(n6437), .C2(n4890), .A(n4889), .B(n6400), .ZN(n5001)
         );
  NOR2_X1 U4160 ( .A1(n4885), .A2(n4587), .ZN(n6083) );
  OAI22_X1 U4161 ( .A1(n6057), .A2(n6516), .B1(n6056), .B2(n6055), .ZN(n6095)
         );
  OAI21_X1 U4162 ( .B1(n6525), .B2(n6524), .A(n6523), .ZN(n6563) );
  INV_X1 U4163 ( .A(n6511), .ZN(n6576) );
  INV_X1 U4164 ( .A(n6560), .ZN(n6630) );
  INV_X1 U4165 ( .A(n5075), .ZN(n5103) );
  INV_X1 U4166 ( .A(n6530), .ZN(n6595) );
  INV_X1 U4167 ( .A(n6553), .ZN(n6619) );
  INV_X1 U4168 ( .A(n6561), .ZN(n6634) );
  AND2_X1 U4169 ( .A1(n3561), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5208) );
  INV_X1 U4170 ( .A(READY_N), .ZN(n6712) );
  INV_X1 U4171 ( .A(n6698), .ZN(n6692) );
  NAND2_X1 U4172 ( .A1(n4465), .A2(n4466), .ZN(n6725) );
  INV_X1 U4173 ( .A(n6220), .ZN(n6899) );
  INV_X1 U4174 ( .A(n6239), .ZN(n4575) );
  OR2_X1 U4175 ( .A1(n6251), .A2(n6267), .ZN(n6253) );
  INV_X1 U4176 ( .A(n4470), .ZN(n6273) );
  OR2_X1 U4177 ( .A1(n5369), .A2(n5359), .ZN(n5710) );
  NOR2_X1 U4178 ( .A1(n5958), .A2(n3814), .ZN(n6348) );
  OR2_X2 U4179 ( .A1(n3792), .A2(n3777), .ZN(n6015) );
  INV_X1 U4180 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6395) );
  AND2_X1 U4181 ( .A1(n4500), .A2(n4487), .ZN(n6040) );
  NAND2_X1 U4182 ( .A1(n5015), .A2(n4587), .ZN(n5045) );
  AOI21_X1 U4183 ( .B1(n5010), .B2(n5012), .A(n5009), .ZN(n5050) );
  AOI21_X1 U4184 ( .B1(n5116), .B2(n5125), .A(n5115), .ZN(n5156) );
  NAND2_X1 U4185 ( .A1(n6396), .A2(n6042), .ZN(n6432) );
  NAND2_X1 U4186 ( .A1(n6396), .A2(n6508), .ZN(n6464) );
  AOI22_X1 U4187 ( .A1(n4703), .A2(n4699), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6434), .ZN(n4730) );
  AOI21_X1 U4188 ( .B1(n4805), .B2(n4804), .A(n4803), .ZN(n6467) );
  AOI22_X1 U4189 ( .A1(n4633), .A2(n4629), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4802), .ZN(n4660) );
  NAND2_X1 U4190 ( .A1(n4630), .A2(n6508), .ZN(n6507) );
  AOI22_X1 U4191 ( .A1(n4888), .A2(n4884), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4890), .ZN(n5005) );
  AOI21_X1 U4192 ( .B1(n6052), .B2(n6516), .A(n6051), .ZN(n6098) );
  OR2_X1 U4193 ( .A1(n6514), .A2(n6043), .ZN(n6567) );
  OR2_X1 U4194 ( .A1(n6514), .A2(n6509), .ZN(n6638) );
  AOI21_X1 U4195 ( .B1(n4956), .B2(n4958), .A(n4952), .ZN(n4994) );
  NAND2_X1 U4196 ( .A1(n4673), .A2(n6042), .ZN(n5096) );
  NOR2_X1 U4197 ( .A1(n4799), .A2(n5168), .ZN(n5201) );
  INV_X1 U4198 ( .A(n6702), .ZN(n6644) );
  OR2_X1 U4199 ( .A1(n3511), .A2(STATE_REG_0__SCAN_IN), .ZN(n6716) );
  NAND2_X1 U4200 ( .A1(n6099), .A2(STATE_REG_2__SCAN_IN), .ZN(n6694) );
  NAND2_X1 U4201 ( .A1(n4423), .A2(n4422), .ZN(U2830) );
  NOR2_X4 U4202 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4741) );
  NAND2_X2 U4203 ( .A1(n5187), .A2(n4741), .ZN(n3408) );
  AND2_X2 U4204 ( .A1(n5194), .A2(n4741), .ZN(n3468) );
  NAND2_X1 U4205 ( .A1(n3468), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3149) );
  NOR2_X4 U4206 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3163) );
  NAND2_X2 U4207 ( .A1(n3163), .A2(n4742), .ZN(n3409) );
  NAND3_X1 U4208 ( .A1(n3150), .A2(n3149), .A3(n3148), .ZN(n3151) );
  AND2_X2 U4209 ( .A1(n3163), .A2(n4741), .ZN(n3486) );
  NAND2_X1 U4210 ( .A1(n3486), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3156) );
  INV_X1 U4211 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U4212 ( .A1(n3476), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3155) );
  AND2_X4 U4213 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4502) );
  NAND2_X1 U4214 ( .A1(n3412), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3154)
         );
  AND2_X2 U4215 ( .A1(n4742), .A2(n4502), .ZN(n4345) );
  NAND2_X1 U4216 ( .A1(n4345), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3153)
         );
  INV_X1 U4217 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U4218 ( .A1(n3392), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3162) );
  AND2_X4 U4219 ( .A1(n4745), .A2(n5194), .ZN(n4027) );
  NAND2_X1 U4220 ( .A1(n4027), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3161)
         );
  AND2_X4 U4221 ( .A1(n5187), .A2(n4742), .ZN(n4317) );
  NAND2_X1 U4222 ( .A1(n4317), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3160)
         );
  NAND2_X1 U4223 ( .A1(n3403), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3159) );
  AND2_X2 U4224 ( .A1(n3164), .A2(n3163), .ZN(n3474) );
  NAND2_X1 U4225 ( .A1(n3474), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3168) );
  AND2_X4 U4226 ( .A1(n3164), .A2(n4502), .ZN(n4320) );
  NAND2_X1 U4227 ( .A1(n4320), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3167) );
  AND2_X4 U4228 ( .A1(n5187), .A2(n4745), .ZN(n4351) );
  NAND2_X1 U4229 ( .A1(n4351), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3166) );
  AND2_X2 U4230 ( .A1(n4741), .A2(n4502), .ZN(n3469) );
  NAND2_X1 U4231 ( .A1(n3469), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3165) );
  INV_X2 U4232 ( .A(n3408), .ZN(n3466) );
  AOI22_X1 U4233 ( .A1(n3387), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U4234 ( .A1(n4317), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4235 ( .A1(n3486), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4236 ( .A1(n4351), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3178) );
  NAND2_X2 U4237 ( .A1(n3142), .A2(n2973), .ZN(n3422) );
  AOI22_X1 U4238 ( .A1(n3466), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4239 ( .A1(n3412), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4240 ( .A1(n3476), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3486), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4241 ( .A1(n4317), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4242 ( .A1(n3386), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4243 ( .A1(n3387), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4244 ( .A1(n3468), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3186) );
  INV_X1 U4245 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6230) );
  INV_X1 U4246 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4554) );
  NAND2_X1 U4247 ( .A1(n3274), .A2(n4554), .ZN(n3192) );
  NAND2_X1 U4248 ( .A1(n4558), .A2(n6230), .ZN(n3191) );
  NAND3_X1 U4249 ( .A1(n3192), .A2(n3201), .A3(n3191), .ZN(n3193) );
  NAND2_X1 U4250 ( .A1(n3194), .A2(n3193), .ZN(n3196) );
  NAND2_X1 U4251 ( .A1(n3274), .A2(EBX_REG_0__SCAN_IN), .ZN(n3195) );
  OAI21_X1 U4252 ( .B1(n3190), .B2(EBX_REG_0__SCAN_IN), .A(n3195), .ZN(n4871)
         );
  XNOR2_X1 U4253 ( .A(n3196), .B(n4871), .ZN(n4557) );
  INV_X1 U4254 ( .A(n3196), .ZN(n3197) );
  MUX2_X1 U4255 ( .A(n3271), .B(n3274), .S(EBX_REG_2__SCAN_IN), .Z(n3200) );
  NAND2_X1 U4256 ( .A1(n3232), .A2(n4410), .ZN(n3234) );
  NAND2_X1 U4257 ( .A1(n4410), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3198)
         );
  AND2_X1 U4258 ( .A1(n3234), .A2(n3198), .ZN(n3199) );
  NAND2_X1 U4259 ( .A1(n3200), .A2(n3199), .ZN(n4855) );
  MUX2_X1 U4260 ( .A(n3266), .B(n3190), .S(EBX_REG_3__SCAN_IN), .Z(n3203) );
  NOR2_X1 U4261 ( .A1(n4872), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3202)
         );
  NOR2_X1 U4262 ( .A1(n3203), .A2(n3202), .ZN(n4669) );
  MUX2_X1 U4263 ( .A(n3204), .B(n3232), .S(EBX_REG_4__SCAN_IN), .Z(n3207) );
  NAND2_X1 U4264 ( .A1(n4410), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3205)
         );
  NAND2_X1 U4265 ( .A1(n3234), .A2(n3205), .ZN(n3206) );
  INV_X1 U4266 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6839) );
  NAND2_X1 U4267 ( .A1(n3266), .A2(n6839), .ZN(n3210) );
  INV_X1 U4268 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U4269 ( .A1(n4558), .A2(n6839), .ZN(n3208) );
  OAI211_X1 U4270 ( .C1(n3190), .C2(n4842), .A(n3208), .B(n3274), .ZN(n3209)
         );
  NAND2_X1 U4271 ( .A1(n3210), .A2(n3209), .ZN(n4847) );
  MUX2_X1 U4272 ( .A(n3204), .B(n3232), .S(EBX_REG_6__SCAN_IN), .Z(n3213) );
  NAND2_X1 U4273 ( .A1(n4410), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3211)
         );
  NAND2_X1 U4274 ( .A1(n3234), .A2(n3211), .ZN(n3212) );
  NOR2_X1 U4275 ( .A1(n3213), .A2(n3212), .ZN(n4995) );
  MUX2_X1 U4276 ( .A(n3266), .B(n3190), .S(EBX_REG_7__SCAN_IN), .Z(n3215) );
  NOR2_X1 U4277 ( .A1(n4872), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3214)
         );
  NOR2_X1 U4278 ( .A1(n3215), .A2(n3214), .ZN(n5553) );
  MUX2_X1 U4279 ( .A(n3204), .B(n3232), .S(EBX_REG_8__SCAN_IN), .Z(n3217) );
  INV_X1 U4280 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6006) );
  OAI21_X1 U4281 ( .B1(n4558), .B2(n6006), .A(n3234), .ZN(n3216) );
  NOR2_X1 U4282 ( .A1(n3217), .A2(n3216), .ZN(n5548) );
  INV_X1 U4283 ( .A(n3266), .ZN(n3272) );
  MUX2_X1 U4284 ( .A(n3272), .B(n3201), .S(EBX_REG_9__SCAN_IN), .Z(n3218) );
  OAI21_X1 U4285 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n4872), .A(n3218), 
        .ZN(n5472) );
  MUX2_X1 U4286 ( .A(n3271), .B(n3274), .S(EBX_REG_10__SCAN_IN), .Z(n3221) );
  NAND2_X1 U4287 ( .A1(n4410), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3219) );
  AND2_X1 U4288 ( .A1(n3234), .A2(n3219), .ZN(n3220) );
  NAND2_X1 U4289 ( .A1(n3221), .A2(n3220), .ZN(n5540) );
  AND2_X2 U4290 ( .A1(n5471), .A2(n5540), .ZN(n5452) );
  INV_X1 U4291 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U4292 ( .A1(n3266), .A2(n5537), .ZN(n3224) );
  INV_X1 U4293 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U4294 ( .A1(n4558), .A2(n5537), .ZN(n3222) );
  OAI211_X1 U4295 ( .C1(n3190), .C2(n5983), .A(n3222), .B(n3274), .ZN(n3223)
         );
  AND2_X1 U4296 ( .A1(n3224), .A2(n3223), .ZN(n5453) );
  MUX2_X1 U4297 ( .A(n3271), .B(n3274), .S(EBX_REG_12__SCAN_IN), .Z(n3227) );
  NAND2_X1 U4298 ( .A1(n4410), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3225) );
  AND2_X1 U4299 ( .A1(n3234), .A2(n3225), .ZN(n3226) );
  NAND2_X1 U4300 ( .A1(n3227), .A2(n3226), .ZN(n5535) );
  INV_X1 U4301 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U4302 ( .A1(n3266), .A2(n6236), .ZN(n3230) );
  INV_X1 U4303 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3757) );
  NAND2_X1 U4304 ( .A1(n4558), .A2(n6236), .ZN(n3228) );
  OAI211_X1 U4305 ( .C1(n3190), .C2(n3757), .A(n3228), .B(n3274), .ZN(n3229)
         );
  NAND2_X1 U4306 ( .A1(n5535), .A2(n5970), .ZN(n3231) );
  MUX2_X1 U4307 ( .A(n3204), .B(n3232), .S(EBX_REG_14__SCAN_IN), .Z(n3236) );
  NAND2_X1 U4308 ( .A1(n4410), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3233) );
  NAND2_X1 U4309 ( .A1(n3234), .A2(n3233), .ZN(n3235) );
  NOR2_X1 U4310 ( .A1(n3236), .A2(n3235), .ZN(n5527) );
  INV_X1 U4311 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U4312 ( .A1(n3266), .A2(n5526), .ZN(n3239) );
  INV_X1 U4313 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U4314 ( .A1(n4558), .A2(n5526), .ZN(n3237) );
  OAI211_X1 U4315 ( .C1(n3190), .C2(n5950), .A(n3237), .B(n3274), .ZN(n3238)
         );
  MUX2_X1 U4316 ( .A(n3271), .B(n3274), .S(EBX_REG_16__SCAN_IN), .Z(n3241) );
  NAND2_X1 U4317 ( .A1(n4410), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3240) );
  INV_X1 U4318 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U4319 ( .A1(n3266), .A2(n5524), .ZN(n3244) );
  INV_X1 U4320 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U4321 ( .A1(n4558), .A2(n5524), .ZN(n3242) );
  OAI211_X1 U4322 ( .C1(n3190), .C2(n5927), .A(n3242), .B(n3274), .ZN(n3243)
         );
  NAND2_X1 U4323 ( .A1(n3244), .A2(n3243), .ZN(n5404) );
  INV_X1 U4324 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U4325 ( .A1(n3204), .A2(n5521), .ZN(n3248) );
  INV_X1 U4326 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U4327 ( .A1(n3274), .A2(n5907), .ZN(n3246) );
  OAI211_X1 U4328 ( .C1(EBX_REG_19__SCAN_IN), .C2(n4410), .A(n3246), .B(n3201), 
        .ZN(n3247) );
  NOR2_X2 U4329 ( .A1(n5370), .A2(n5374), .ZN(n5356) );
  INV_X1 U4330 ( .A(n4872), .ZN(n3279) );
  INV_X1 U4331 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5917) );
  NOR2_X1 U4332 ( .A1(n4410), .A2(EBX_REG_18__SCAN_IN), .ZN(n5371) );
  AOI21_X1 U4333 ( .B1(n3279), .B2(n5917), .A(n5371), .ZN(n5372) );
  OAI22_X1 U4334 ( .A1(n4872), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4410), .ZN(n5358) );
  NAND2_X1 U4335 ( .A1(n5372), .A2(n5358), .ZN(n3250) );
  NAND2_X1 U4336 ( .A1(n3190), .A2(EBX_REG_20__SCAN_IN), .ZN(n3249) );
  OAI211_X1 U4337 ( .C1(n5372), .C2(n3190), .A(n3250), .B(n3249), .ZN(n3251)
         );
  INV_X1 U4338 ( .A(n3251), .ZN(n3252) );
  AND2_X2 U4339 ( .A1(n5356), .A2(n3252), .ZN(n5346) );
  INV_X1 U4340 ( .A(EBX_REG_21__SCAN_IN), .ZN(n3253) );
  NAND2_X1 U4341 ( .A1(n3266), .A2(n3253), .ZN(n3257) );
  INV_X1 U4342 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3255) );
  NAND2_X1 U4343 ( .A1(n4558), .A2(n3253), .ZN(n3254) );
  OAI211_X1 U4344 ( .C1(n3190), .C2(n3255), .A(n3254), .B(n3274), .ZN(n3256)
         );
  MUX2_X1 U4345 ( .A(n3271), .B(n3274), .S(EBX_REG_22__SCAN_IN), .Z(n3259) );
  NAND2_X1 U4346 ( .A1(n4410), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3258) );
  NAND2_X1 U4347 ( .A1(n3259), .A2(n3258), .ZN(n5336) );
  INV_X1 U4348 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U4349 ( .A1(n3266), .A2(n5516), .ZN(n3263) );
  INV_X1 U4350 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U4351 ( .A1(n4558), .A2(n5516), .ZN(n3260) );
  OAI211_X1 U4352 ( .C1(n3190), .C2(n3261), .A(n3260), .B(n3274), .ZN(n3262)
         );
  NAND2_X1 U4353 ( .A1(n3263), .A2(n3262), .ZN(n5317) );
  MUX2_X1 U4354 ( .A(n3271), .B(n3274), .S(EBX_REG_24__SCAN_IN), .Z(n3265) );
  NAND2_X1 U4355 ( .A1(n4410), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3264) );
  MUX2_X1 U4356 ( .A(n3266), .B(n3190), .S(EBX_REG_25__SCAN_IN), .Z(n3268) );
  NOR2_X1 U4357 ( .A1(n4872), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3267)
         );
  NOR2_X1 U4358 ( .A1(n3268), .A2(n3267), .ZN(n5289) );
  INV_X1 U4359 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U4360 ( .A1(n3274), .A2(n5641), .ZN(n3269) );
  OAI211_X1 U4361 ( .C1(EBX_REG_26__SCAN_IN), .C2(n4410), .A(n3269), .B(n3201), 
        .ZN(n3270) );
  OAI21_X1 U4362 ( .B1(n3271), .B2(EBX_REG_26__SCAN_IN), .A(n3270), .ZN(n5280)
         );
  NAND2_X1 U4363 ( .A1(n5279), .A2(n5280), .ZN(n5261) );
  MUX2_X1 U4364 ( .A(n3272), .B(n3201), .S(EBX_REG_27__SCAN_IN), .Z(n3273) );
  OAI21_X1 U4365 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4872), .A(n3273), 
        .ZN(n5262) );
  INV_X1 U4366 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U4367 ( .A1(n3204), .A2(n5509), .ZN(n3277) );
  INV_X1 U4368 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3769) );
  NAND2_X1 U4369 ( .A1(n3274), .A2(n3769), .ZN(n3275) );
  OAI211_X1 U4370 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4410), .A(n3275), .B(n3201), 
        .ZN(n3276) );
  INV_X1 U4371 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5807) );
  NOR2_X1 U4372 ( .A1(n4410), .A2(EBX_REG_29__SCAN_IN), .ZN(n3278) );
  AOI21_X1 U4373 ( .B1(n3279), .B2(n5807), .A(n3278), .ZN(n4413) );
  AND2_X1 U4374 ( .A1(n4410), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3280)
         );
  AOI21_X1 U4375 ( .B1(n4872), .B2(EBX_REG_30__SCAN_IN), .A(n3280), .ZN(n3824)
         );
  INV_X1 U4376 ( .A(n3281), .ZN(n3283) );
  AOI211_X1 U4377 ( .C1(n3190), .C2(n3822), .A(n3824), .B(n2970), .ZN(n3282)
         );
  NOR2_X1 U4378 ( .A1(n3283), .A2(n3282), .ZN(n5507) );
  NAND2_X1 U4379 ( .A1(n3530), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3515) );
  NAND2_X1 U4380 ( .A1(n3386), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3287)
         );
  NAND2_X1 U4381 ( .A1(n3466), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3286) );
  NAND2_X1 U4382 ( .A1(n3412), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3285)
         );
  NAND2_X1 U4383 ( .A1(n3468), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3284) );
  NAND2_X1 U4384 ( .A1(n3392), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3291) );
  NAND2_X1 U4385 ( .A1(n4027), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3290)
         );
  NAND2_X1 U4386 ( .A1(n4317), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3289)
         );
  NAND2_X1 U4387 ( .A1(n3403), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U4388 ( .A1(n3474), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3294) );
  NAND2_X1 U4389 ( .A1(n3469), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3293) );
  NAND2_X1 U4390 ( .A1(n3387), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3292)
         );
  NAND2_X1 U4391 ( .A1(n3476), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3299) );
  NAND2_X1 U4392 ( .A1(n4320), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3298) );
  NAND2_X1 U4393 ( .A1(n3486), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3297) );
  NAND2_X1 U4394 ( .A1(n4345), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3296)
         );
  NAND2_X1 U4395 ( .A1(n3729), .A2(n3422), .ZN(n3314) );
  AOI22_X1 U4396 ( .A1(n3486), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3304) );
  AND4_X2 U4397 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n3313)
         );
  AOI22_X1 U4398 ( .A1(n3468), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3310) );
  NAND2_X1 U4401 ( .A1(n3314), .A2(n3426), .ZN(n3323) );
  XNOR2_X1 U4402 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3318) );
  INV_X1 U4403 ( .A(n3318), .ZN(n3316) );
  INV_X1 U4404 ( .A(n3317), .ZN(n3315) );
  NAND2_X1 U4405 ( .A1(n3316), .A2(n3315), .ZN(n3319) );
  NAND2_X1 U4406 ( .A1(n3318), .A2(n3317), .ZN(n3334) );
  AND2_X1 U4407 ( .A1(n3319), .A2(n3334), .ZN(n3442) );
  XNOR2_X1 U4408 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3322) );
  AOI21_X1 U4409 ( .B1(n3506), .B2(n3322), .A(n3328), .ZN(n3321) );
  NAND2_X1 U4410 ( .A1(n2972), .A2(n3426), .ZN(n3320) );
  NAND2_X1 U4411 ( .A1(n4524), .A2(n3320), .ZN(n3342) );
  OAI22_X1 U4412 ( .A1(n3323), .A2(n3324), .B1(n3321), .B2(n3342), .ZN(n3330)
         );
  NAND2_X1 U4413 ( .A1(n3729), .A2(n3322), .ZN(n3327) );
  INV_X1 U4414 ( .A(n3323), .ZN(n3326) );
  INV_X1 U4415 ( .A(n3324), .ZN(n3325) );
  OAI22_X1 U4416 ( .A1(n3330), .A2(n3327), .B1(n3326), .B2(n3325), .ZN(n3332)
         );
  AOI21_X1 U4417 ( .B1(n3330), .B2(n3442), .A(n3351), .ZN(n3331) );
  NAND2_X1 U4418 ( .A1(n4948), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U4419 ( .A1(n3334), .A2(n3333), .ZN(n3339) );
  XNOR2_X1 U4420 ( .A(n4768), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3337)
         );
  XNOR2_X1 U4421 ( .A(n3339), .B(n3337), .ZN(n3441) );
  NAND2_X1 U4422 ( .A1(n3729), .A2(n3441), .ZN(n3336) );
  INV_X1 U4423 ( .A(n3342), .ZN(n3335) );
  OAI211_X1 U4424 ( .C1(n3441), .C2(n3731), .A(n3336), .B(n3335), .ZN(n3345)
         );
  INV_X1 U4425 ( .A(n3337), .ZN(n3338) );
  NAND2_X1 U4426 ( .A1(n3339), .A2(n3338), .ZN(n3341) );
  NAND2_X1 U4427 ( .A1(n4769), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3340) );
  XNOR2_X1 U4428 ( .A(n4747), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3346)
         );
  XNOR2_X1 U4429 ( .A(n3349), .B(n3346), .ZN(n3443) );
  NAND3_X1 U4430 ( .A1(n3342), .A2(n3729), .A3(n3441), .ZN(n3343) );
  OAI21_X1 U4431 ( .B1(n3443), .B2(n3726), .A(n3343), .ZN(n3344) );
  INV_X1 U4432 ( .A(n3346), .ZN(n3348) );
  AND2_X1 U4433 ( .A1(n3354), .A2(n3357), .ZN(n3353) );
  INV_X1 U4434 ( .A(n3353), .ZN(n3446) );
  NAND2_X1 U4435 ( .A1(n3446), .A2(n3443), .ZN(n3350) );
  NOR2_X1 U4436 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4784), .ZN(n3352) );
  INV_X1 U4437 ( .A(n3354), .ZN(n3356) );
  INV_X1 U4438 ( .A(n3357), .ZN(n3358) );
  NAND2_X1 U4439 ( .A1(n3729), .A2(n3440), .ZN(n3360) );
  NAND2_X1 U4440 ( .A1(n3466), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3367) );
  NAND2_X1 U4441 ( .A1(n3392), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3366) );
  NAND2_X1 U4442 ( .A1(n4320), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3365) );
  NAND2_X1 U4443 ( .A1(n3387), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3364)
         );
  AND4_X2 U4444 ( .A1(n3367), .A2(n3366), .A3(n3365), .A4(n3364), .ZN(n3385)
         );
  NAND2_X1 U4445 ( .A1(n3476), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3371) );
  NAND2_X1 U4446 ( .A1(n3468), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3370) );
  NAND2_X1 U4447 ( .A1(n3386), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3369)
         );
  NAND2_X1 U4448 ( .A1(n4345), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3373)
         );
  NAND2_X1 U4449 ( .A1(n3474), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3372) );
  NAND2_X1 U4450 ( .A1(n3373), .A2(n3372), .ZN(n3377) );
  NAND2_X1 U4451 ( .A1(n4351), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3375) );
  NAND2_X1 U4452 ( .A1(n3486), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3374) );
  NAND2_X1 U4453 ( .A1(n3375), .A2(n3374), .ZN(n3376) );
  NAND2_X1 U4454 ( .A1(n4317), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3381)
         );
  NAND2_X1 U4455 ( .A1(n4027), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3380)
         );
  NAND2_X1 U4456 ( .A1(n3403), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3379) );
  NAND2_X1 U4457 ( .A1(n3469), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4458 ( .A1(n3412), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4459 ( .A1(n3468), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4460 ( .A1(n3466), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3387), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4461 ( .A1(n3486), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3388) );
  NAND4_X1 U4462 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3398)
         );
  AOI22_X1 U4463 ( .A1(n4351), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4464 ( .A1(n4320), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4465 ( .A1(n3392), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3393) );
  NAND4_X1 U4466 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3397)
         );
  OR2_X2 U4467 ( .A1(n3398), .A2(n3397), .ZN(n3427) );
  INV_X1 U4468 ( .A(n3430), .ZN(n3399) );
  NOR2_X1 U4469 ( .A1(n4759), .A2(n2972), .ZN(n3790) );
  INV_X1 U4470 ( .A(n3790), .ZN(n3450) );
  INV_X1 U4471 ( .A(n3423), .ZN(n3401) );
  AND2_X2 U4472 ( .A1(n3401), .A2(n3427), .ZN(n3455) );
  NAND2_X1 U4473 ( .A1(n3455), .A2(n3426), .ZN(n3402) );
  AOI22_X1 U4474 ( .A1(n4027), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4475 ( .A1(n4351), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3474), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4476 ( .A1(n4320), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3469), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4477 ( .A1(n3392), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3403), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4478 ( .A1(n3386), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3468), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3416) );
  INV_X1 U4479 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5030) );
  BUF_X4 U4480 ( .A(n3409), .Z(n4297) );
  INV_X1 U4481 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3410) );
  OAI22_X1 U4482 ( .A1(n3408), .A2(n5030), .B1(n4297), .B2(n3410), .ZN(n3411)
         );
  INV_X1 U4483 ( .A(n3411), .ZN(n3415) );
  AOI22_X1 U4484 ( .A1(n3486), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4485 ( .A1(n3412), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3476), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3413) );
  INV_X2 U4486 ( .A(n3432), .ZN(n4617) );
  INV_X1 U4487 ( .A(n3513), .ZN(n3420) );
  NAND2_X1 U4488 ( .A1(n4759), .A2(n3530), .ZN(n3419) );
  NAND2_X1 U4489 ( .A1(n3420), .A2(n3419), .ZN(n3775) );
  INV_X1 U4490 ( .A(n3775), .ZN(n3425) );
  NAND2_X1 U4491 ( .A1(n3508), .A2(n2971), .ZN(n3424) );
  MUX2_X1 U4492 ( .A(n3424), .B(n6713), .S(n3516), .Z(n3781) );
  NAND2_X1 U4493 ( .A1(n3425), .A2(n3781), .ZN(n3437) );
  NAND2_X1 U4494 ( .A1(n3455), .A2(n4595), .ZN(n3429) );
  NAND2_X1 U4495 ( .A1(n3432), .A2(n3427), .ZN(n3428) );
  NAND3_X1 U4496 ( .A1(n3430), .A2(n3429), .A3(n3428), .ZN(n3434) );
  NAND2_X1 U4497 ( .A1(n3862), .A2(n4405), .ZN(n3433) );
  INV_X1 U4498 ( .A(n3531), .ZN(n3557) );
  OR2_X1 U4499 ( .A1(n3506), .A2(n2971), .ZN(n3532) );
  INV_X1 U4500 ( .A(n3532), .ZN(n3435) );
  INV_X1 U4501 ( .A(n4459), .ZN(n3436) );
  NAND2_X1 U4502 ( .A1(n3437), .A2(n3436), .ZN(n4480) );
  INV_X1 U4503 ( .A(STATE_REG_1__SCAN_IN), .ZN(n3438) );
  INV_X1 U4504 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4440) );
  NAND2_X1 U4505 ( .A1(n3438), .A2(n4440), .ZN(n4437) );
  NAND2_X1 U4506 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n3439) );
  NAND2_X1 U4507 ( .A1(n4437), .A2(n3439), .ZN(n3511) );
  NAND2_X1 U4508 ( .A1(n3422), .A2(n6716), .ZN(n3448) );
  INV_X1 U4509 ( .A(n3440), .ZN(n3445) );
  NAND3_X1 U4510 ( .A1(n3443), .A2(n3442), .A3(n3441), .ZN(n3444) );
  NAND2_X1 U4511 ( .A1(n3445), .A2(n3444), .ZN(n3447) );
  NOR2_X1 U4512 ( .A1(n4458), .A2(READY_N), .ZN(n4476) );
  NAND3_X1 U4513 ( .A1(n3448), .A2(n4476), .A3(n4405), .ZN(n3449) );
  OAI211_X1 U4514 ( .C1(n4492), .C2(n3450), .A(n4480), .B(n3449), .ZN(n3451)
         );
  NAND2_X1 U4515 ( .A1(n3451), .A2(n5208), .ZN(n3460) );
  NAND3_X1 U4516 ( .A1(n3418), .A2(n3454), .A3(n4599), .ZN(n3551) );
  NAND2_X1 U4517 ( .A1(n2972), .A2(n6716), .ZN(n3834) );
  NAND2_X1 U4518 ( .A1(n3834), .A2(n6712), .ZN(n3456) );
  OAI211_X1 U4519 ( .C1(n3551), .C2(n3456), .A(n2971), .B(n5216), .ZN(n3457)
         );
  INV_X1 U4520 ( .A(n3457), .ZN(n3458) );
  AND3_X1 U4521 ( .A1(n4603), .A2(n4617), .A3(n4595), .ZN(n3462) );
  NAND2_X1 U4522 ( .A1(n3857), .A2(n4599), .ZN(n3463) );
  OAI21_X1 U4523 ( .B1(n3554), .B2(n3463), .A(n4798), .ZN(n3464) );
  INV_X1 U4524 ( .A(n3464), .ZN(n3465) );
  NAND2_X1 U4525 ( .A1(n3517), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3499) );
  INV_X2 U4526 ( .A(n3467), .ZN(n4342) );
  AOI22_X1 U4527 ( .A1(n4342), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3473) );
  CLKBUF_X3 U4528 ( .A(n3486), .Z(n4325) );
  AOI22_X1 U4529 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4352), .B1(n4325), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3472) );
  CLKBUF_X3 U4530 ( .A(n3392), .Z(n4355) );
  CLKBUF_X3 U4531 ( .A(n3469), .Z(n4199) );
  AOI22_X1 U4532 ( .A1(n4355), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3471) );
  CLKBUF_X3 U4533 ( .A(n3403), .Z(n4354) );
  AOI22_X1 U4534 ( .A1(n4748), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4535 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n4198), .B1(n4353), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4536 ( .A1(n4197), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3478) );
  CLKBUF_X3 U4537 ( .A(n3476), .Z(n4318) );
  AOI22_X1 U4538 ( .A1(n4318), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3477) );
  CLKBUF_X3 U4539 ( .A(n3386), .Z(n4344) );
  INV_X1 U4540 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3481) );
  INV_X1 U4541 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4970) );
  OAI22_X1 U4542 ( .A1(n4296), .A2(n3481), .B1(n4297), .B2(n4970), .ZN(n3482)
         );
  INV_X1 U4543 ( .A(n3482), .ZN(n3483) );
  NAND3_X1 U4544 ( .A1(n2990), .A2(n3484), .A3(n3483), .ZN(n3571) );
  INV_X1 U4545 ( .A(n3571), .ZN(n3590) );
  AOI22_X1 U4546 ( .A1(n4344), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U4547 ( .A1(n4352), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3489) );
  INV_X1 U4548 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6749) );
  INV_X1 U4549 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4962) );
  OAI22_X1 U4550 ( .A1(n3467), .A2(n6749), .B1(n4297), .B2(n4962), .ZN(n3485)
         );
  INV_X1 U4551 ( .A(n3485), .ZN(n3488) );
  AOI22_X1 U4552 ( .A1(n4325), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3487) );
  NAND4_X1 U4553 ( .A1(n3490), .A2(n3489), .A3(n3488), .A4(n3487), .ZN(n3496)
         );
  AOI22_X1 U4554 ( .A1(n4197), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4555 ( .A1(n4198), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4556 ( .A1(n4748), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4557 ( .A1(n4355), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3491) );
  NAND4_X1 U4558 ( .A1(n3494), .A2(n3493), .A3(n3492), .A4(n3491), .ZN(n3495)
         );
  OR2_X2 U4559 ( .A1(n3496), .A2(n3495), .ZN(n3745) );
  NAND2_X1 U4560 ( .A1(n3745), .A2(n4599), .ZN(n3502) );
  OAI211_X1 U4561 ( .C1(n3590), .C2(n2971), .A(n3502), .B(
        STATE2_REG_0__SCAN_IN), .ZN(n3497) );
  INV_X1 U4562 ( .A(n3497), .ZN(n3498) );
  INV_X1 U4563 ( .A(n3586), .ZN(n3505) );
  INV_X1 U4564 ( .A(n3745), .ZN(n3501) );
  NOR2_X2 U4565 ( .A1(n3502), .A2(n6722), .ZN(n3743) );
  INV_X1 U4566 ( .A(n3587), .ZN(n3584) );
  INV_X1 U4567 ( .A(n3743), .ZN(n3503) );
  AND2_X1 U4568 ( .A1(n3584), .A2(n3503), .ZN(n3504) );
  OR2_X2 U4569 ( .A1(n3505), .A2(n3504), .ZN(n3536) );
  INV_X1 U4570 ( .A(n3506), .ZN(n3555) );
  NAND2_X1 U4571 ( .A1(n3509), .A2(n3508), .ZN(n3510) );
  NAND2_X1 U4572 ( .A1(n3400), .A2(n3511), .ZN(n3553) );
  NAND2_X1 U4573 ( .A1(n3553), .A2(n4595), .ZN(n3512) );
  INV_X1 U4574 ( .A(n3515), .ZN(n3556) );
  NAND3_X1 U4575 ( .A1(n3520), .A2(n3519), .A3(n3518), .ZN(n3550) );
  NAND2_X1 U4576 ( .A1(n3550), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3522) );
  NAND2_X1 U4577 ( .A1(n5164), .A2(n6722), .ZN(n4378) );
  MUX2_X1 U4578 ( .A(n3561), .B(n4378), .S(n6574), .Z(n3521) );
  NAND2_X1 U4579 ( .A1(n3522), .A2(n3521), .ZN(n3578) );
  NAND3_X1 U4580 ( .A1(n3530), .A2(n4617), .A3(n4603), .ZN(n3787) );
  NAND2_X1 U4581 ( .A1(n5164), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3523) );
  AOI21_X1 U4582 ( .B1(n3524), .B2(n3509), .A(n3523), .ZN(n3525) );
  OAI211_X1 U4583 ( .C1(n3430), .C2(n3787), .A(n2995), .B(n3525), .ZN(n3529)
         );
  AOI21_X1 U4584 ( .B1(n3526), .B2(n3527), .A(n2972), .ZN(n3528) );
  NOR2_X1 U4585 ( .A1(n3529), .A2(n3528), .ZN(n3534) );
  NAND2_X1 U4586 ( .A1(n6711), .A2(n4617), .ZN(n3533) );
  AOI22_X1 U4587 ( .A1(n3533), .A2(n3532), .B1(n3531), .B2(n5479), .ZN(n3783)
         );
  NAND2_X1 U4588 ( .A1(n3534), .A2(n3783), .ZN(n3579) );
  NAND2_X2 U4589 ( .A1(n3578), .A2(n3579), .ZN(n3599) );
  NAND2_X1 U4590 ( .A1(n3599), .A2(n6722), .ZN(n3535) );
  INV_X1 U4591 ( .A(n3537), .ZN(n3549) );
  AOI22_X1 U4592 ( .A1(n4198), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4593 ( .A1(n4343), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4594 ( .A1(n4344), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4595 ( .A1(n4325), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3538) );
  NAND4_X1 U4596 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3547)
         );
  AOI22_X1 U4597 ( .A1(n4319), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4598 ( .A1(n4342), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4599 ( .A1(n4748), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4600 ( .A1(n4355), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3542) );
  NAND4_X1 U4601 ( .A1(n3545), .A2(n3544), .A3(n3543), .A4(n3542), .ZN(n3546)
         );
  NAND2_X1 U4602 ( .A1(n3556), .A2(n3572), .ZN(n3548) );
  OAI211_X1 U4603 ( .C1(n3731), .C2(n6825), .A(n3549), .B(n3548), .ZN(n3594)
         );
  XNOR2_X1 U4604 ( .A(n3593), .B(n3594), .ZN(n3570) );
  NAND2_X1 U4605 ( .A1(n3550), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3563) );
  NAND2_X1 U4606 ( .A1(n3553), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3560) );
  NOR2_X2 U4607 ( .A1(n3554), .A2(n5216), .ZN(n3773) );
  NAND2_X1 U4608 ( .A1(n3773), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3559) );
  NAND4_X1 U4609 ( .A1(n3557), .A2(n3556), .A3(n2972), .A4(n3555), .ZN(n3558)
         );
  INV_X1 U4610 ( .A(n3567), .ZN(n3562) );
  XNOR2_X1 U4611 ( .A(n6574), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6433)
         );
  AOI22_X1 U4612 ( .A1(n6724), .A2(n6433), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n4795), .ZN(n3564) );
  NAND3_X1 U4613 ( .A1(n3563), .A2(n3562), .A3(n3564), .ZN(n3600) );
  INV_X1 U4614 ( .A(n3564), .ZN(n3565) );
  NAND2_X1 U4615 ( .A1(n3567), .A2(n3566), .ZN(n3598) );
  NAND2_X1 U4616 ( .A1(n3600), .A2(n3598), .ZN(n3568) );
  XNOR2_X1 U4617 ( .A(n3568), .B(n3599), .ZN(n4582) );
  NAND2_X1 U4618 ( .A1(n4409), .A2(n3572), .ZN(n3569) );
  NAND2_X1 U4619 ( .A1(n3856), .A2(n3742), .ZN(n3577) );
  NAND2_X1 U4620 ( .A1(n3572), .A2(n3571), .ZN(n3629) );
  OAI211_X1 U4621 ( .C1(n3572), .C2(n3571), .A(n4469), .B(n3629), .ZN(n3575)
         );
  NOR2_X1 U4622 ( .A1(n3573), .A2(n4595), .ZN(n3574) );
  AND2_X1 U4623 ( .A1(n3575), .A2(n3574), .ZN(n3576) );
  NAND2_X1 U4624 ( .A1(n3577), .A2(n3576), .ZN(n4551) );
  INV_X1 U4625 ( .A(n3599), .ZN(n3582) );
  INV_X1 U4626 ( .A(n3578), .ZN(n3581) );
  INV_X1 U4627 ( .A(n3579), .ZN(n3580) );
  NOR2_X1 U4628 ( .A1(n3582), .A2(n2974), .ZN(n3863) );
  NAND2_X1 U4629 ( .A1(n3863), .A2(n6722), .ZN(n3583) );
  NAND2_X1 U4630 ( .A1(n3583), .A2(n3586), .ZN(n3585) );
  NAND2_X1 U4631 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  AND2_X1 U4632 ( .A1(n3530), .A2(n3461), .ZN(n3631) );
  AOI21_X1 U4633 ( .B1(n3590), .B2(n4469), .A(n3631), .ZN(n3591) );
  OAI21_X1 U4634 ( .B1(n4587), .B2(n3726), .A(n3591), .ZN(n4521) );
  XNOR2_X1 U4635 ( .A(n6380), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4552)
         );
  NAND2_X1 U4636 ( .A1(n4551), .A2(n4552), .ZN(n4550) );
  OR2_X1 U4637 ( .A1(n6380), .A2(n4554), .ZN(n3592) );
  INV_X1 U4638 ( .A(n3593), .ZN(n3596) );
  INV_X1 U4639 ( .A(n3594), .ZN(n3595) );
  NAND2_X1 U4640 ( .A1(n3596), .A2(n3595), .ZN(n3597) );
  NAND2_X1 U4641 ( .A1(n3599), .A2(n3598), .ZN(n3601) );
  NAND2_X1 U4642 ( .A1(n3601), .A2(n3600), .ZN(n3608) );
  INV_X1 U4643 ( .A(n3608), .ZN(n3607) );
  AND2_X1 U4644 ( .A1(n4769), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6522)
         );
  NAND2_X1 U4645 ( .A1(n6522), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U4646 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3602) );
  NAND2_X1 U4647 ( .A1(n3602), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3603) );
  NAND2_X1 U4648 ( .A1(n6510), .A2(n3603), .ZN(n4679) );
  AOI22_X1 U4649 ( .A1(n4679), .A2(n6724), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n4795), .ZN(n3604) );
  NAND2_X2 U4650 ( .A1(n3607), .A2(n3606), .ZN(n4496) );
  NAND2_X1 U4651 ( .A1(n3608), .A2(n3609), .ZN(n3610) );
  AOI22_X1 U4652 ( .A1(n4344), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4653 ( .A1(n4352), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3614) );
  INV_X1 U4654 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5145) );
  INV_X1 U4655 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4974) );
  OAI22_X1 U4656 ( .A1(n3467), .A2(n5145), .B1(n4297), .B2(n4974), .ZN(n3611)
         );
  INV_X1 U4657 ( .A(n3611), .ZN(n3613) );
  AOI22_X1 U4658 ( .A1(n4325), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3612) );
  NAND4_X1 U4659 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3621)
         );
  AOI22_X1 U4660 ( .A1(n4197), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4661 ( .A1(n4198), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4662 ( .A1(n4748), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3617) );
  INV_X1 U4663 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6739) );
  AOI22_X1 U4664 ( .A1(n4355), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3616) );
  NAND4_X1 U4665 ( .A1(n3619), .A2(n3618), .A3(n3617), .A4(n3616), .ZN(n3620)
         );
  AOI22_X1 U4666 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n3517), .B1(n3729), 
        .B2(n3628), .ZN(n3622) );
  INV_X1 U4667 ( .A(n3623), .ZN(n3626) );
  INV_X1 U4668 ( .A(n3624), .ZN(n3625) );
  NAND2_X1 U4669 ( .A1(n3626), .A2(n3625), .ZN(n3627) );
  INV_X1 U4670 ( .A(n3628), .ZN(n3630) );
  NAND2_X1 U4671 ( .A1(n3629), .A2(n3630), .ZN(n3651) );
  OAI21_X1 U4672 ( .B1(n3630), .B2(n3629), .A(n3651), .ZN(n3632) );
  AOI21_X1 U4673 ( .B1(n3632), .B2(n4469), .A(n3631), .ZN(n3633) );
  OAI21_X1 U4674 ( .B1(n6331), .B2(n6332), .A(n6333), .ZN(n4662) );
  NAND2_X1 U4675 ( .A1(n3634), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4676 ( .A1(n4802), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4655) );
  NAND2_X1 U4677 ( .A1(n4655), .A2(n6519), .ZN(n3635) );
  AND2_X1 U4678 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4949) );
  NAND2_X1 U4679 ( .A1(n4676), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4619) );
  AOI22_X1 U4680 ( .A1(n6476), .A2(n6724), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4795), .ZN(n3636) );
  AOI22_X1 U4681 ( .A1(n4344), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4682 ( .A1(n4352), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3641) );
  INV_X1 U4683 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5137) );
  INV_X1 U4684 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4983) );
  OAI22_X1 U4685 ( .A1(n3467), .A2(n5137), .B1(n4297), .B2(n4983), .ZN(n3638)
         );
  INV_X1 U4686 ( .A(n3638), .ZN(n3640) );
  AOI22_X1 U4687 ( .A1(n4325), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3639) );
  NAND4_X1 U4688 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n3648)
         );
  AOI22_X1 U4689 ( .A1(n4197), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4690 ( .A1(n4198), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4691 ( .A1(n4748), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4692 ( .A1(n4355), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3643) );
  NAND4_X1 U4693 ( .A1(n3646), .A2(n3645), .A3(n3644), .A4(n3643), .ZN(n3647)
         );
  AOI22_X1 U4694 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n3517), .B1(n3729), 
        .B2(n3652), .ZN(n3649) );
  NAND2_X1 U4695 ( .A1(n4858), .A2(n3742), .ZN(n3654) );
  NAND2_X1 U4696 ( .A1(n3651), .A2(n3652), .ZN(n3700) );
  OAI211_X1 U4697 ( .C1(n3652), .C2(n3651), .A(n3700), .B(n4469), .ZN(n3653)
         );
  NAND2_X1 U4698 ( .A1(n3654), .A2(n3653), .ZN(n3655) );
  INV_X1 U4699 ( .A(n3655), .ZN(n3656) );
  INV_X1 U4700 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4666) );
  NAND2_X1 U4701 ( .A1(n3517), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4702 ( .A1(n4344), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4703 ( .A1(n4352), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3661) );
  INV_X1 U4704 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5129) );
  INV_X1 U4705 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4987) );
  OAI22_X1 U4706 ( .A1(n3467), .A2(n5129), .B1(n4297), .B2(n4987), .ZN(n3658)
         );
  INV_X1 U4707 ( .A(n3658), .ZN(n3660) );
  AOI22_X1 U4708 ( .A1(n4325), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3659) );
  NAND4_X1 U4709 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(n3668)
         );
  AOI22_X1 U4710 ( .A1(n4197), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3666) );
  INV_X1 U4711 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6770) );
  AOI22_X1 U4712 ( .A1(n4198), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4713 ( .A1(n4748), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4714 ( .A1(n4355), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3663) );
  NAND4_X1 U4715 ( .A1(n3666), .A2(n3665), .A3(n3664), .A4(n3663), .ZN(n3667)
         );
  NAND2_X1 U4716 ( .A1(n3729), .A2(n3698), .ZN(n3669) );
  NAND2_X1 U4717 ( .A1(n3671), .A2(n3672), .ZN(n3675) );
  NAND2_X1 U4718 ( .A1(n3895), .A2(n3742), .ZN(n3678) );
  XNOR2_X1 U4719 ( .A(n3700), .B(n3698), .ZN(n3676) );
  NAND2_X1 U4720 ( .A1(n3676), .A2(n4469), .ZN(n3677) );
  NAND2_X1 U4721 ( .A1(n3678), .A2(n3677), .ZN(n3680) );
  INV_X1 U4722 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3679) );
  XNOR2_X1 U4723 ( .A(n3680), .B(n3679), .ZN(n4687) );
  NAND2_X1 U4724 ( .A1(n4688), .A2(n4687), .ZN(n3682) );
  NAND2_X1 U4725 ( .A1(n3680), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3681)
         );
  NAND2_X1 U4726 ( .A1(n3682), .A2(n3681), .ZN(n4837) );
  INV_X1 U4727 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U4728 ( .A1(n4344), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4729 ( .A1(n4352), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3686) );
  INV_X1 U4730 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4966) );
  OAI22_X1 U4731 ( .A1(n3467), .A2(n6842), .B1(n4297), .B2(n4966), .ZN(n3683)
         );
  INV_X1 U4732 ( .A(n3683), .ZN(n3685) );
  AOI22_X1 U4733 ( .A1(n4325), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4734 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3693)
         );
  AOI22_X1 U4735 ( .A1(n4197), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4736 ( .A1(n4198), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4737 ( .A1(n4748), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4738 ( .A1(n4355), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3688) );
  NAND4_X1 U4739 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3692)
         );
  NAND2_X1 U4740 ( .A1(n3729), .A2(n3701), .ZN(n3694) );
  NAND2_X1 U4741 ( .A1(n3696), .A2(n3134), .ZN(n3697) );
  NAND2_X1 U4742 ( .A1(n3722), .A2(n3697), .ZN(n3898) );
  INV_X1 U4743 ( .A(n3698), .ZN(n3699) );
  NOR2_X1 U4744 ( .A1(n3700), .A2(n3699), .ZN(n3702) );
  NAND2_X1 U4745 ( .A1(n3702), .A2(n3701), .ZN(n3733) );
  OAI211_X1 U4746 ( .C1(n3702), .C2(n3701), .A(n3733), .B(n4469), .ZN(n3703)
         );
  XNOR2_X1 U4747 ( .A(n3704), .B(n4842), .ZN(n4838) );
  NAND2_X1 U4748 ( .A1(n3704), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3705)
         );
  NAND2_X1 U4749 ( .A1(n3517), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4750 ( .A1(n4344), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4751 ( .A1(n4352), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3709) );
  INV_X1 U4752 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5124) );
  INV_X1 U4753 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4979) );
  OAI22_X1 U4754 ( .A1(n3467), .A2(n5124), .B1(n4297), .B2(n4979), .ZN(n3706)
         );
  INV_X1 U4755 ( .A(n3706), .ZN(n3708) );
  INV_X1 U4756 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6869) );
  AOI22_X1 U4757 ( .A1(n4325), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3707) );
  NAND4_X1 U4758 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3716)
         );
  AOI22_X1 U4759 ( .A1(n4197), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4760 ( .A1(n4198), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4761 ( .A1(n4748), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4762 ( .A1(n4355), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3711) );
  NAND4_X1 U4763 ( .A1(n3714), .A2(n3713), .A3(n3712), .A4(n3711), .ZN(n3715)
         );
  NAND2_X1 U4764 ( .A1(n3729), .A2(n3734), .ZN(n3717) );
  NAND2_X1 U4765 ( .A1(n3722), .A2(n3721), .ZN(n3723) );
  XNOR2_X1 U4766 ( .A(n3733), .B(n3734), .ZN(n3724) );
  NAND2_X1 U4767 ( .A1(n3724), .A2(n4469), .ZN(n3725) );
  INV_X1 U4768 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3727) );
  INV_X1 U4769 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U4770 ( .A1(n3729), .A2(n3745), .ZN(n3730) );
  OAI21_X1 U4771 ( .B1(n4937), .B2(n3731), .A(n3730), .ZN(n3732) );
  NAND2_X1 U4772 ( .A1(n3920), .A2(n3742), .ZN(n3738) );
  INV_X1 U4773 ( .A(n3733), .ZN(n3735) );
  NAND2_X1 U4774 ( .A1(n3735), .A2(n3734), .ZN(n3747) );
  XNOR2_X1 U4775 ( .A(n3747), .B(n3745), .ZN(n3736) );
  NAND2_X1 U4776 ( .A1(n3736), .A2(n4469), .ZN(n3737) );
  NAND2_X1 U4777 ( .A1(n3738), .A2(n3737), .ZN(n3739) );
  INV_X1 U4778 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6365) );
  XNOR2_X1 U4779 ( .A(n3739), .B(n6365), .ZN(n5183) );
  NAND2_X1 U4780 ( .A1(n3739), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3740)
         );
  NAND2_X1 U4781 ( .A1(n4469), .A2(n3745), .ZN(n3746) );
  OR2_X1 U4782 ( .A1(n3747), .A2(n3746), .ZN(n3748) );
  NAND2_X1 U4783 ( .A1(n3753), .A2(n3748), .ZN(n3749) );
  XNOR2_X1 U4784 ( .A(n3749), .B(n6006), .ZN(n5799) );
  NAND2_X1 U4785 ( .A1(n3749), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3750)
         );
  INV_X1 U4786 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U4787 ( .A1(n5760), .A2(n6841), .ZN(n3751) );
  INV_X1 U4788 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6000) );
  AND2_X1 U4789 ( .A1(n5760), .A2(n6000), .ZN(n5778) );
  NAND2_X1 U4790 ( .A1(n5757), .A2(n5983), .ZN(n5767) );
  INV_X1 U4791 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U4792 ( .A1(n5757), .A2(n5759), .ZN(n5758) );
  AND2_X1 U4793 ( .A1(n5767), .A2(n5758), .ZN(n3752) );
  NAND2_X1 U4794 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5777) );
  OAI21_X1 U4795 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A(n5662), .ZN(n3754) );
  AND2_X1 U4796 ( .A1(n5777), .A2(n3754), .ZN(n5744) );
  OAI21_X1 U4797 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .A(n5662), .ZN(n3755) );
  NAND2_X1 U4798 ( .A1(n5757), .A2(n3757), .ZN(n5746) );
  INV_X1 U4799 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U4800 ( .A1(n5757), .A2(n5967), .ZN(n3758) );
  AND2_X1 U4801 ( .A1(n5746), .A2(n3758), .ZN(n3759) );
  AND2_X1 U4802 ( .A1(n5760), .A2(n5950), .ZN(n3762) );
  NAND2_X1 U4803 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3761) );
  INV_X1 U4804 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5944) );
  AND3_X1 U4805 ( .A1(n5927), .A2(n5917), .A3(n5944), .ZN(n3763) );
  NOR2_X1 U4806 ( .A1(n5757), .A2(n3763), .ZN(n3765) );
  NAND2_X1 U4807 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3816) );
  OAI21_X1 U4808 ( .B1(n3816), .B2(n5944), .A(n5757), .ZN(n3764) );
  NOR2_X1 U4809 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5856) );
  NOR2_X1 U4810 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5874) );
  NOR2_X1 U4811 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5896) );
  NAND3_X1 U4812 ( .A1(n5856), .A2(n5874), .A3(n5896), .ZN(n3766) );
  NAND2_X1 U4813 ( .A1(n5662), .A2(n3766), .ZN(n3767) );
  NAND2_X1 U4814 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U4815 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5873) );
  NOR2_X1 U4816 ( .A1(n5872), .A2(n5873), .ZN(n5854) );
  AND2_X1 U4817 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3801) );
  NAND2_X1 U4818 ( .A1(n5854), .A2(n3801), .ZN(n3818) );
  NAND2_X1 U4819 ( .A1(n5757), .A2(n3818), .ZN(n3768) );
  XNOR2_X1 U4820 ( .A(n5789), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5652)
         );
  INV_X1 U4821 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U4822 ( .A1(n5828), .A2(n3769), .ZN(n5817) );
  NOR3_X1 U4823 ( .A1(n5757), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5817), 
        .ZN(n4385) );
  NAND2_X1 U4824 ( .A1(n5643), .A2(n4385), .ZN(n5617) );
  AND2_X1 U4825 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5836) );
  AND2_X1 U4826 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U4827 ( .A1(n5836), .A2(n5808), .ZN(n3770) );
  NAND2_X1 U4828 ( .A1(n4459), .A2(n2972), .ZN(n4498) );
  NAND2_X1 U4829 ( .A1(n3773), .A2(n3453), .ZN(n3774) );
  AND2_X1 U4830 ( .A1(n4473), .A2(n3774), .ZN(n3776) );
  AND4_X1 U4831 ( .A1(n4498), .A2(n3776), .A3(n4790), .A4(n4529), .ZN(n3777)
         );
  NOR2_X1 U4832 ( .A1(n6711), .A2(n4405), .ZN(n4478) );
  OAI21_X1 U4833 ( .B1(n4478), .B2(n4872), .A(n3573), .ZN(n3779) );
  NAND2_X1 U4834 ( .A1(n5216), .A2(n4405), .ZN(n3778) );
  OAI211_X1 U4835 ( .C1(n3201), .C2(n3526), .A(n3779), .B(n3778), .ZN(n3780)
         );
  INV_X1 U4836 ( .A(n3780), .ZN(n3782) );
  NAND3_X1 U4837 ( .A1(n3783), .A2(n3782), .A3(n3781), .ZN(n4489) );
  INV_X1 U4838 ( .A(n3862), .ZN(n3785) );
  OAI22_X1 U4839 ( .A1(n3554), .A2(n3785), .B1(n3784), .B2(n2971), .ZN(n3786)
         );
  INV_X1 U4840 ( .A(n3786), .ZN(n3788) );
  OR2_X1 U4841 ( .A1(n4759), .A2(n3787), .ZN(n4750) );
  NAND2_X1 U4842 ( .A1(n3788), .A2(n4750), .ZN(n3789) );
  NAND2_X1 U4843 ( .A1(n3791), .A2(n3790), .ZN(n4506) );
  NAND2_X1 U4844 ( .A1(n6437), .A2(n4786), .ZN(n5219) );
  NAND2_X1 U4845 ( .A1(n3792), .A2(n3820), .ZN(n6391) );
  INV_X1 U4846 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6393) );
  NOR2_X1 U4847 ( .A1(n3792), .A2(n3791), .ZN(n3810) );
  OR2_X1 U4848 ( .A1(n3810), .A2(n4664), .ZN(n5955) );
  NAND2_X1 U4849 ( .A1(n6393), .A2(n5955), .ZN(n6385) );
  NAND2_X1 U4850 ( .A1(n6391), .A2(n6385), .ZN(n4663) );
  NOR2_X1 U4851 ( .A1(n4664), .A2(n4663), .ZN(n5991) );
  INV_X1 U4852 ( .A(n3810), .ZN(n3793) );
  NAND2_X1 U4853 ( .A1(n6392), .A2(n3793), .ZN(n5995) );
  INV_X1 U4854 ( .A(n5995), .ZN(n3798) );
  NAND2_X1 U4855 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5956) );
  INV_X1 U4856 ( .A(n5956), .ZN(n3794) );
  AND2_X1 U4857 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n3794), .ZN(n5960)
         );
  NAND2_X1 U4858 ( .A1(n5960), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5935) );
  NAND2_X1 U4859 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3815) );
  NOR2_X1 U4860 ( .A1(n5935), .A2(n3815), .ZN(n3799) );
  NOR2_X1 U4861 ( .A1(n6006), .A2(n6365), .ZN(n6005) );
  NAND3_X1 U4862 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n6005), .ZN(n3797) );
  NAND2_X1 U4863 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3796) );
  AOI21_X1 U4864 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4665) );
  NAND2_X1 U4865 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4844) );
  NOR2_X1 U4866 ( .A1(n4665), .A2(n4844), .ZN(n5056) );
  INV_X1 U4867 ( .A(n5888), .ZN(n3795) );
  INV_X1 U4868 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6874) );
  NOR2_X1 U4869 ( .A1(n6874), .A2(n4554), .ZN(n4840) );
  NOR2_X1 U4870 ( .A1(n4844), .A2(n3796), .ZN(n5999) );
  NAND2_X1 U4871 ( .A1(n4840), .A2(n5999), .ZN(n5994) );
  NOR2_X1 U4872 ( .A1(n5994), .A2(n3797), .ZN(n3813) );
  AOI21_X1 U4873 ( .B1(n3813), .B2(n3799), .A(n3798), .ZN(n5890) );
  INV_X1 U4874 ( .A(n5955), .ZN(n3800) );
  NAND2_X1 U4875 ( .A1(n6392), .A2(n6393), .ZN(n4553) );
  INV_X1 U4876 ( .A(n6367), .ZN(n3802) );
  AOI21_X1 U4877 ( .B1(n3802), .B2(n6372), .A(n3801), .ZN(n3803) );
  INV_X1 U4878 ( .A(n5836), .ZN(n3804) );
  NAND2_X1 U4879 ( .A1(n5936), .A2(n3804), .ZN(n3805) );
  NAND2_X1 U4880 ( .A1(n5855), .A2(n3805), .ZN(n5827) );
  INV_X1 U4881 ( .A(n5808), .ZN(n5816) );
  AND2_X1 U4882 ( .A1(n5936), .A2(n5816), .ZN(n3806) );
  OR2_X1 U4883 ( .A1(n5827), .A2(n3806), .ZN(n5813) );
  AND2_X1 U4884 ( .A1(n5936), .A2(n5807), .ZN(n3807) );
  NAND3_X1 U4885 ( .A1(n3810), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n3813), 
        .ZN(n3812) );
  INV_X1 U4886 ( .A(n5931), .ZN(n3811) );
  NAND2_X1 U4887 ( .A1(n3812), .A2(n3811), .ZN(n5958) );
  INV_X1 U4888 ( .A(n3813), .ZN(n5932) );
  NOR2_X1 U4889 ( .A1(n6392), .A2(n5932), .ZN(n3814) );
  INV_X1 U4890 ( .A(n3816), .ZN(n3817) );
  INV_X1 U4891 ( .A(n3818), .ZN(n3819) );
  NAND3_X1 U4892 ( .A1(n5829), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5808), .ZN(n4391) );
  NAND2_X1 U4893 ( .A1(n6368), .A2(REIP_REG_30__SCAN_IN), .ZN(n4427) );
  OAI21_X1 U4894 ( .B1(n4391), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4427), 
        .ZN(n3821) );
  INV_X1 U4895 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4419) );
  NAND2_X1 U4896 ( .A1(n3204), .A2(n4419), .ZN(n4414) );
  NAND2_X1 U4897 ( .A1(n4418), .A2(n3824), .ZN(n3825) );
  OAI22_X1 U4898 ( .A1(n4872), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4410), .ZN(n3826) );
  INV_X1 U4899 ( .A(n3826), .ZN(n3827) );
  INV_X1 U4900 ( .A(n4458), .ZN(n3829) );
  NAND2_X1 U4901 ( .A1(n4449), .A2(n5208), .ZN(n4466) );
  NAND2_X1 U4902 ( .A1(n4369), .A2(n4377), .ZN(n5167) );
  AND2_X1 U4903 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n3830) );
  NAND2_X1 U4904 ( .A1(n4577), .A2(n3830), .ZN(n5206) );
  NAND2_X1 U4905 ( .A1(n5167), .A2(n5206), .ZN(n3831) );
  NAND2_X1 U4906 ( .A1(n6712), .A2(n6435), .ZN(n5230) );
  NAND2_X1 U4907 ( .A1(n5230), .A2(EBX_REG_31__SCAN_IN), .ZN(n3832) );
  NOR2_X1 U4908 ( .A1(n4410), .A2(n3832), .ZN(n3833) );
  NOR2_X1 U4909 ( .A1(n3530), .A2(n5230), .ZN(n3835) );
  AND2_X1 U4910 ( .A1(n3835), .A2(n3834), .ZN(n3836) );
  NAND3_X1 U4911 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n6163) );
  NAND3_X1 U4912 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5483) );
  INV_X1 U4913 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6662) );
  NOR3_X1 U4914 ( .A1(n6163), .A2(n5483), .A3(n6662), .ZN(n5457) );
  NAND2_X1 U4915 ( .A1(n5457), .A2(REIP_REG_8__SCAN_IN), .ZN(n5456) );
  INV_X1 U4916 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6668) );
  NAND3_X1 U4917 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        REIP_REG_11__SCAN_IN), .ZN(n6135) );
  NOR4_X1 U4918 ( .A1(n5456), .A2(n6668), .A3(n6148), .A4(n6135), .ZN(n6121)
         );
  NAND2_X1 U4919 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6121), .ZN(n5424) );
  INV_X1 U4920 ( .A(n5424), .ZN(n5441) );
  AND2_X1 U4921 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n3837) );
  NAND2_X1 U4922 ( .A1(n5441), .A2(n3837), .ZN(n3839) );
  NOR2_X1 U4923 ( .A1(n6206), .A2(n3839), .ZN(n5410) );
  NAND2_X1 U4924 ( .A1(n5410), .A2(REIP_REG_17__SCAN_IN), .ZN(n5395) );
  NAND3_X1 U4925 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n3841) );
  INV_X1 U4926 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6682) );
  INV_X1 U4927 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5691) );
  INV_X1 U4928 ( .A(REIP_REG_23__SCAN_IN), .ZN(n5674) );
  NOR2_X1 U4929 ( .A1(n5319), .A2(n5674), .ZN(n5295) );
  AND2_X1 U4930 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5274) );
  NAND2_X1 U4931 ( .A1(n5274), .A2(REIP_REG_26__SCAN_IN), .ZN(n5265) );
  INV_X1 U4932 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6689) );
  NOR2_X1 U4933 ( .A1(n5265), .A2(n6689), .ZN(n3838) );
  NAND3_X1 U4934 ( .A1(n5254), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .ZN(n5229) );
  INV_X1 U4935 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5228) );
  NOR3_X1 U4936 ( .A1(n5229), .A2(REIP_REG_31__SCAN_IN), .A3(n5228), .ZN(n3854) );
  INV_X1 U4937 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4383) );
  INV_X1 U4938 ( .A(n3839), .ZN(n3840) );
  NAND2_X1 U4939 ( .A1(n6197), .A2(n3840), .ZN(n5377) );
  INV_X1 U4940 ( .A(n3841), .ZN(n3842) );
  NAND2_X1 U4941 ( .A1(REIP_REG_17__SCAN_IN), .A2(n3842), .ZN(n3843) );
  OR2_X1 U4942 ( .A1(n5377), .A2(n3843), .ZN(n3844) );
  NAND2_X1 U4943 ( .A1(n6170), .A2(n3844), .ZN(n5361) );
  NOR2_X1 U4944 ( .A1(n6682), .A2(n5691), .ZN(n5330) );
  NAND2_X1 U4945 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5330), .ZN(n3845) );
  NAND2_X1 U4946 ( .A1(n6170), .A2(n3845), .ZN(n3846) );
  NAND2_X1 U4947 ( .A1(n5361), .A2(n3846), .ZN(n5320) );
  AND2_X1 U4948 ( .A1(n6170), .A2(n5265), .ZN(n3847) );
  OR2_X1 U4949 ( .A1(n5320), .A2(n3847), .ZN(n5275) );
  NAND2_X1 U4950 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n3848) );
  OR2_X1 U4951 ( .A1(n5275), .A2(n3848), .ZN(n3849) );
  NAND2_X1 U4952 ( .A1(n3849), .A2(n6170), .ZN(n5252) );
  OAI211_X1 U4953 ( .C1(REIP_REG_29__SCAN_IN), .C2(n6206), .A(n5252), .B(
        REIP_REG_30__SCAN_IN), .ZN(n5226) );
  NAND3_X1 U4954 ( .A1(n5226), .A2(REIP_REG_31__SCAN_IN), .A3(n6170), .ZN(
        n3852) );
  INV_X1 U4955 ( .A(n6716), .ZN(n6714) );
  INV_X1 U4956 ( .A(n5230), .ZN(n3850) );
  NAND2_X1 U4957 ( .A1(n6714), .A2(n3850), .ZN(n4797) );
  AND2_X1 U4958 ( .A1(n4469), .A2(n4797), .ZN(n5231) );
  NAND3_X1 U4959 ( .A1(n5484), .A2(EBX_REG_31__SCAN_IN), .A3(n5231), .ZN(n3851) );
  OAI211_X1 U4960 ( .C1(n4383), .C2(n6186), .A(n3852), .B(n3851), .ZN(n3853)
         );
  AOI21_X1 U4961 ( .B1(n5504), .B2(n6220), .A(n3855), .ZN(n4376) );
  NAND2_X1 U4962 ( .A1(n3856), .A2(n4018), .ZN(n3861) );
  NOR2_X2 U4963 ( .A1(n4530), .A2(n5165), .ZN(n3913) );
  INV_X1 U4964 ( .A(n3882), .ZN(n4269) );
  AOI22_X1 U4965 ( .A1(n4269), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5165), .ZN(n3859) );
  NAND2_X1 U4966 ( .A1(n3881), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3858) );
  AND2_X1 U4967 ( .A1(n3859), .A2(n3858), .ZN(n3860) );
  NAND2_X1 U4968 ( .A1(n3863), .A2(n4018), .ZN(n3867) );
  AOI22_X1 U4969 ( .A1(n3913), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n5165), .ZN(n3865) );
  NAND2_X1 U4970 ( .A1(n3881), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3864) );
  AND2_X1 U4971 ( .A1(n3865), .A2(n3864), .ZN(n3866) );
  NAND2_X1 U4972 ( .A1(n4515), .A2(n4517), .ZN(n4516) );
  INV_X1 U4973 ( .A(n4517), .ZN(n3868) );
  NAND2_X1 U4974 ( .A1(n3868), .A2(n3908), .ZN(n3869) );
  NAND2_X1 U4975 ( .A1(n3881), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3875) );
  INV_X1 U4976 ( .A(n3891), .ZN(n3870) );
  OAI21_X1 U4977 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3870), .ZN(n6340) );
  NAND2_X1 U4978 ( .A1(n6340), .A2(n3908), .ZN(n3872) );
  NAND2_X1 U4979 ( .A1(n4370), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3871)
         );
  NAND2_X1 U4980 ( .A1(n3872), .A2(n3871), .ZN(n3873) );
  AOI21_X1 U4981 ( .B1(n4269), .B2(EAX_REG_2__SCAN_IN), .A(n3873), .ZN(n3874)
         );
  AND2_X1 U4982 ( .A1(n3875), .A2(n3874), .ZN(n3876) );
  INV_X1 U4983 ( .A(n4370), .ZN(n4225) );
  NAND2_X1 U4984 ( .A1(n4543), .A2(n4546), .ZN(n3880) );
  INV_X1 U4985 ( .A(n4733), .ZN(n3878) );
  INV_X1 U4986 ( .A(n3876), .ZN(n3877) );
  NAND2_X1 U4987 ( .A1(n3878), .A2(n3877), .ZN(n3879) );
  INV_X1 U4988 ( .A(n3881), .ZN(n3890) );
  XNOR2_X1 U4989 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .B(n3891), .ZN(n6201) );
  AOI22_X1 U4990 ( .A1(n4369), .A2(n6201), .B1(n4370), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3884) );
  NAND2_X1 U4991 ( .A1(n3913), .A2(EAX_REG_3__SCAN_IN), .ZN(n3883) );
  OAI211_X1 U4992 ( .C1(n3890), .C2(n4747), .A(n3884), .B(n3883), .ZN(n3885)
         );
  INV_X1 U4993 ( .A(n3885), .ZN(n3886) );
  NAND2_X1 U4994 ( .A1(n3887), .A2(n3886), .ZN(n4549) );
  NAND2_X1 U4995 ( .A1(n4544), .A2(n4549), .ZN(n4547) );
  INV_X1 U4996 ( .A(n4547), .ZN(n3897) );
  NAND2_X1 U4997 ( .A1(n5165), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3889)
         );
  NAND2_X1 U4998 ( .A1(n4269), .A2(EAX_REG_4__SCAN_IN), .ZN(n3888) );
  OAI211_X1 U4999 ( .C1(n3890), .C2(n4784), .A(n3889), .B(n3888), .ZN(n3893)
         );
  OAI21_X1 U5000 ( .B1(n3892), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3899), 
        .ZN(n5482) );
  MUX2_X1 U5001 ( .A(n3893), .B(n5482), .S(n4369), .Z(n3894) );
  AOI21_X1 U5002 ( .B1(n3895), .B2(n4018), .A(n3894), .ZN(n4625) );
  NAND2_X1 U5003 ( .A1(n3897), .A2(n3896), .ZN(n4624) );
  AND2_X1 U5004 ( .A1(n3899), .A2(n6185), .ZN(n3900) );
  OR2_X1 U5005 ( .A1(n3900), .A2(n3906), .ZN(n6196) );
  NAND2_X1 U5006 ( .A1(n6196), .A2(n4369), .ZN(n3901) );
  OAI21_X1 U5007 ( .B1(n6185), .B2(n4225), .A(n3901), .ZN(n3902) );
  AOI21_X1 U5008 ( .B1(n3913), .B2(EAX_REG_5__SCAN_IN), .A(n3902), .ZN(n3903)
         );
  NOR2_X2 U5009 ( .A1(n4624), .A2(n4852), .ZN(n4850) );
  OR2_X1 U5010 ( .A1(n3906), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3907) );
  NAND2_X1 U5011 ( .A1(n3915), .A2(n3907), .ZN(n6184) );
  INV_X1 U5012 ( .A(n6184), .ZN(n3910) );
  AOI22_X1 U5013 ( .A1(n3913), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n5165), .ZN(n3909) );
  MUX2_X1 U5014 ( .A(n3910), .B(n3909), .S(n4339), .Z(n3911) );
  NAND2_X1 U5015 ( .A1(n4850), .A2(n4876), .ZN(n4877) );
  INV_X1 U5016 ( .A(n4877), .ZN(n3922) );
  INV_X1 U5017 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3918) );
  NAND2_X1 U5018 ( .A1(n3915), .A2(n3914), .ZN(n3916) );
  NAND2_X1 U5019 ( .A1(n3923), .A2(n3916), .ZN(n6176) );
  AOI22_X1 U5020 ( .A1(n6176), .A2(n4369), .B1(n4370), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3917) );
  OAI21_X1 U5021 ( .B1(n3882), .B2(n3918), .A(n3917), .ZN(n3919) );
  AOI21_X1 U5022 ( .B1(n3920), .B2(n4018), .A(n3919), .ZN(n5178) );
  INV_X1 U5023 ( .A(n5178), .ZN(n3921) );
  NAND2_X1 U5024 ( .A1(n3922), .A2(n3921), .ZN(n5179) );
  NAND2_X1 U5025 ( .A1(n3913), .A2(EAX_REG_8__SCAN_IN), .ZN(n3939) );
  AOI21_X1 U5026 ( .B1(n6755), .B2(n3923), .A(n3956), .ZN(n6157) );
  INV_X1 U5027 ( .A(n6157), .ZN(n5802) );
  AOI22_X1 U5028 ( .A1(n4370), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n4369), 
        .B2(n5802), .ZN(n3938) );
  AOI22_X1 U5029 ( .A1(n4355), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U5030 ( .A1(n4198), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U5031 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4352), .B1(n4318), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3927) );
  INV_X1 U5032 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3924) );
  INV_X1 U5033 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4739) );
  OAI22_X1 U5034 ( .A1(n3924), .A2(n3467), .B1(n4297), .B2(n4739), .ZN(n3925)
         );
  INV_X1 U5035 ( .A(n3925), .ZN(n3926) );
  NAND4_X1 U5036 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3935)
         );
  AOI22_X1 U5037 ( .A1(n4344), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U5038 ( .A1(n4317), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U5039 ( .A1(n4197), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U5040 ( .A1(n4325), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3930) );
  NAND4_X1 U5041 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3934)
         );
  NOR2_X1 U5042 ( .A1(n3935), .A2(n3934), .ZN(n3936) );
  OR2_X1 U5043 ( .A1(n4052), .A2(n3936), .ZN(n3937) );
  NAND2_X1 U5044 ( .A1(n3913), .A2(EAX_REG_9__SCAN_IN), .ZN(n3955) );
  XNOR2_X1 U5045 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3956), .ZN(n5792) );
  AOI22_X1 U5046 ( .A1(n4369), .A2(n5792), .B1(n4370), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U5047 ( .A1(n4319), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U5048 ( .A1(n4342), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U5049 ( .A1(n4748), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4325), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U5050 ( .A1(n4317), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3942) );
  NAND4_X1 U5051 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3951)
         );
  AOI22_X1 U5052 ( .A1(n4344), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U5053 ( .A1(n4352), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U5054 ( .A1(n4198), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U5055 ( .A1(n4343), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3946) );
  NAND4_X1 U5056 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3950)
         );
  NOR2_X1 U5057 ( .A1(n3951), .A2(n3950), .ZN(n3952) );
  OR2_X1 U5058 ( .A1(n4052), .A2(n3952), .ZN(n3953) );
  XOR2_X1 U5059 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3982), .Z(n6888) );
  AOI22_X1 U5060 ( .A1(n4197), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3962) );
  INV_X1 U5061 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3957) );
  INV_X1 U5062 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4930) );
  OAI22_X1 U5063 ( .A1(n3467), .A2(n3957), .B1(n4296), .B2(n4930), .ZN(n3958)
         );
  INV_X1 U5064 ( .A(n3958), .ZN(n3961) );
  AOI22_X1 U5065 ( .A1(n4343), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U5066 ( .A1(n4352), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3959) );
  NAND4_X1 U5067 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(n3968)
         );
  AOI22_X1 U5068 ( .A1(n4198), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U5069 ( .A1(n4319), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4325), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U5070 ( .A1(n4355), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U5071 ( .A1(n4748), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3963) );
  NAND4_X1 U5072 ( .A1(n3966), .A2(n3965), .A3(n3964), .A4(n3963), .ZN(n3967)
         );
  OR2_X1 U5073 ( .A1(n3968), .A2(n3967), .ZN(n3969) );
  AOI22_X1 U5074 ( .A1(n4018), .A2(n3969), .B1(n4370), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3971) );
  NAND2_X1 U5075 ( .A1(n3913), .A2(EAX_REG_10__SCAN_IN), .ZN(n3970) );
  OAI211_X1 U5076 ( .C1(n6888), .C2(n4339), .A(n3971), .B(n3970), .ZN(n5542)
         );
  AOI22_X1 U5077 ( .A1(n4197), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U5078 ( .A1(n4198), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U5079 ( .A1(n4343), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U5080 ( .A1(n4325), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U5081 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3981)
         );
  AOI22_X1 U5082 ( .A1(n4319), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U5083 ( .A1(n4342), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U5084 ( .A1(n4748), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U5085 ( .A1(n4344), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U5086 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3980)
         );
  NOR2_X1 U5087 ( .A1(n3981), .A2(n3980), .ZN(n3985) );
  XNOR2_X1 U5088 ( .A(n3986), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5772)
         );
  NAND2_X1 U5089 ( .A1(n5772), .A2(n4369), .ZN(n3984) );
  AOI22_X1 U5090 ( .A1(n3913), .A2(EAX_REG_11__SCAN_IN), .B1(n4370), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3983) );
  OAI211_X1 U5091 ( .C1(n3985), .C2(n4052), .A(n3984), .B(n3983), .ZN(n5450)
         );
  XNOR2_X1 U5092 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n4019), .ZN(n6141)
         );
  INV_X1 U5093 ( .A(n6141), .ZN(n5764) );
  AOI22_X1 U5094 ( .A1(n4198), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U5095 ( .A1(n4319), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U5096 ( .A1(n4355), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U5097 ( .A1(n4318), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3987) );
  NAND4_X1 U5098 ( .A1(n3990), .A2(n3989), .A3(n3988), .A4(n3987), .ZN(n3998)
         );
  INV_X1 U5099 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3991) );
  INV_X1 U5100 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4923) );
  OAI22_X1 U5101 ( .A1(n3467), .A2(n3991), .B1(n4296), .B2(n4923), .ZN(n3992)
         );
  INV_X1 U5102 ( .A(n3992), .ZN(n3996) );
  AOI22_X1 U5103 ( .A1(n4197), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U5104 ( .A1(n4352), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4325), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U5105 ( .A1(n4353), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3993) );
  NAND4_X1 U5106 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n3997)
         );
  NOR2_X1 U5107 ( .A1(n3998), .A2(n3997), .ZN(n4001) );
  NAND2_X1 U5108 ( .A1(n3913), .A2(EAX_REG_12__SCAN_IN), .ZN(n4000) );
  NAND2_X1 U5109 ( .A1(n4370), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3999)
         );
  OAI211_X1 U5110 ( .C1(n4001), .C2(n4052), .A(n4000), .B(n3999), .ZN(n4002)
         );
  AOI21_X1 U5111 ( .B1(n5764), .B2(n4369), .A(n4002), .ZN(n5534) );
  AOI22_X1 U5112 ( .A1(n4344), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U5113 ( .A1(n4352), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4009) );
  INV_X1 U5114 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4005) );
  INV_X1 U5115 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4004) );
  OAI22_X1 U5116 ( .A1(n3467), .A2(n4005), .B1(n4297), .B2(n4004), .ZN(n4006)
         );
  INV_X1 U5117 ( .A(n4006), .ZN(n4008) );
  AOI22_X1 U5118 ( .A1(n4325), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4007) );
  NAND4_X1 U5119 ( .A1(n4010), .A2(n4009), .A3(n4008), .A4(n4007), .ZN(n4016)
         );
  AOI22_X1 U5120 ( .A1(n4197), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U5121 ( .A1(n4198), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U5122 ( .A1(n4748), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U5123 ( .A1(n4355), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4011) );
  NAND4_X1 U5124 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(n4015)
         );
  OR2_X1 U5125 ( .A1(n4016), .A2(n4015), .ZN(n4017) );
  AND2_X1 U5126 ( .A1(n4018), .A2(n4017), .ZN(n5436) );
  XNOR2_X1 U5127 ( .A(n4021), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6134)
         );
  AOI22_X1 U5128 ( .A1(n3913), .A2(EAX_REG_13__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4370), .ZN(n4020) );
  OAI21_X1 U5129 ( .B1(n6134), .B2(n4339), .A(n4020), .ZN(n5437) );
  INV_X1 U5130 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4022) );
  XNOR2_X1 U5131 ( .A(n4060), .B(n4022), .ZN(n5738) );
  NAND2_X1 U5132 ( .A1(n5738), .A2(n4369), .ZN(n4039) );
  AOI22_X1 U5133 ( .A1(n4344), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U5134 ( .A1(n4352), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U5135 ( .A1(n4342), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4320), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U5136 ( .A1(n4198), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4325), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U5137 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4033)
         );
  AOI22_X1 U5138 ( .A1(n4319), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5139 ( .A1(n4355), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U5140 ( .A1(n4350), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U5141 ( .A1(n4353), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4028) );
  NAND4_X1 U5142 ( .A1(n4031), .A2(n4030), .A3(n4029), .A4(n4028), .ZN(n4032)
         );
  NOR2_X1 U5143 ( .A1(n4033), .A2(n4032), .ZN(n4036) );
  NAND2_X1 U5144 ( .A1(n3913), .A2(EAX_REG_15__SCAN_IN), .ZN(n4035) );
  NAND2_X1 U5145 ( .A1(n4370), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4034)
         );
  OAI211_X1 U5146 ( .C1(n4036), .C2(n4052), .A(n4035), .B(n4034), .ZN(n4037)
         );
  INV_X1 U5147 ( .A(n4037), .ZN(n4038) );
  NAND2_X1 U5148 ( .A1(n4039), .A2(n4038), .ZN(n5439) );
  XNOR2_X1 U5149 ( .A(n2999), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6124)
         );
  NAND2_X1 U5150 ( .A1(n6124), .A2(n4369), .ZN(n4056) );
  AOI22_X1 U5151 ( .A1(n4198), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5152 ( .A1(n4344), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5153 ( .A1(n4319), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5154 ( .A1(n4352), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4040) );
  NAND4_X1 U5155 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4049)
         );
  AOI22_X1 U5156 ( .A1(n4197), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5157 ( .A1(n4342), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5158 ( .A1(n4343), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4325), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5159 ( .A1(n4748), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4044) );
  NAND4_X1 U5160 ( .A1(n4047), .A2(n4046), .A3(n4045), .A4(n4044), .ZN(n4048)
         );
  NOR2_X1 U5161 ( .A1(n4049), .A2(n4048), .ZN(n4053) );
  NAND2_X1 U5162 ( .A1(n3913), .A2(EAX_REG_14__SCAN_IN), .ZN(n4051) );
  NAND2_X1 U5163 ( .A1(n4370), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4050)
         );
  OAI211_X1 U5164 ( .C1(n4053), .C2(n4052), .A(n4051), .B(n4050), .ZN(n4054)
         );
  INV_X1 U5165 ( .A(n4054), .ZN(n4055) );
  NAND2_X1 U5166 ( .A1(n4056), .A2(n4055), .ZN(n5531) );
  OAI211_X1 U5167 ( .C1(n5436), .C2(n5437), .A(n5439), .B(n5531), .ZN(n4057)
         );
  NAND2_X1 U5168 ( .A1(n4059), .A2(n4058), .ZN(n5416) );
  INV_X1 U5169 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5425) );
  XNOR2_X1 U5170 ( .A(n4089), .B(n5425), .ZN(n5730) );
  AOI22_X1 U5171 ( .A1(n4355), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5172 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4197), .B1(n4198), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4066) );
  INV_X1 U5173 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4062) );
  OAI22_X1 U5174 ( .A1(n4062), .A2(n3467), .B1(n4296), .B2(n5022), .ZN(n4063)
         );
  INV_X1 U5175 ( .A(n4063), .ZN(n4065) );
  AOI22_X1 U5176 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n4352), .B1(n4325), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4064) );
  NAND4_X1 U5177 ( .A1(n4067), .A2(n4066), .A3(n4065), .A4(n4064), .ZN(n4073)
         );
  AOI22_X1 U5178 ( .A1(n4319), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5179 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n4748), .B1(n4353), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U5180 ( .A1(n4199), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5181 ( .A1(n4318), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4068) );
  NAND4_X1 U5182 ( .A1(n4071), .A2(n4070), .A3(n4069), .A4(n4068), .ZN(n4072)
         );
  NOR2_X1 U5183 ( .A1(n4073), .A2(n4072), .ZN(n4075) );
  AOI22_X1 U5184 ( .A1(n3913), .A2(EAX_REG_16__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n4370), .ZN(n4074) );
  OAI21_X1 U5185 ( .B1(n4334), .B2(n4075), .A(n4074), .ZN(n4076) );
  AOI21_X1 U5186 ( .B1(n5730), .B2(n4369), .A(n4076), .ZN(n5417) );
  AOI22_X1 U5187 ( .A1(n4198), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5188 ( .A1(n4319), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U5189 ( .A1(n4342), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5190 ( .A1(n4325), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4077) );
  NAND4_X1 U5191 ( .A1(n4080), .A2(n4079), .A3(n4078), .A4(n4077), .ZN(n4086)
         );
  AOI22_X1 U5192 ( .A1(n4344), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4027), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5193 ( .A1(n4352), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5194 ( .A1(n4350), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5195 ( .A1(n4748), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4081) );
  NAND4_X1 U5196 ( .A1(n4084), .A2(n4083), .A3(n4082), .A4(n4081), .ZN(n4085)
         );
  NOR2_X1 U5197 ( .A1(n4086), .A2(n4085), .ZN(n4088) );
  AOI22_X1 U5198 ( .A1(n3913), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n5165), .ZN(n4087) );
  OAI21_X1 U5199 ( .B1(n4334), .B2(n4088), .A(n4087), .ZN(n4092) );
  NAND2_X1 U5200 ( .A1(n4090), .A2(n6776), .ZN(n4091) );
  NAND2_X1 U5201 ( .A1(n4111), .A2(n4091), .ZN(n5725) );
  MUX2_X1 U5202 ( .A(n4092), .B(n5725), .S(n4369), .Z(n5401) );
  XNOR2_X1 U5203 ( .A(n4111), .B(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5714)
         );
  NAND2_X1 U5204 ( .A1(n5714), .A2(n4369), .ZN(n4110) );
  AOI22_X1 U5205 ( .A1(n4344), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U5206 ( .A1(n4352), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4098) );
  INV_X1 U5207 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4094) );
  INV_X1 U5208 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4093) );
  OAI22_X1 U5209 ( .A1(n3467), .A2(n4094), .B1(n4297), .B2(n4093), .ZN(n4095)
         );
  INV_X1 U5210 ( .A(n4095), .ZN(n4097) );
  AOI22_X1 U5211 ( .A1(n4325), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4096) );
  NAND4_X1 U5212 ( .A1(n4099), .A2(n4098), .A3(n4097), .A4(n4096), .ZN(n4105)
         );
  AOI22_X1 U5213 ( .A1(n4197), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5214 ( .A1(n4198), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5215 ( .A1(n4748), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5216 ( .A1(n4355), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4100) );
  NAND4_X1 U5217 ( .A1(n4103), .A2(n4102), .A3(n4101), .A4(n4100), .ZN(n4104)
         );
  NOR2_X1 U5218 ( .A1(n4105), .A2(n4104), .ZN(n4108) );
  AOI21_X1 U5219 ( .B1(n3073), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4106) );
  AOI21_X1 U5220 ( .B1(n3913), .B2(EAX_REG_18__SCAN_IN), .A(n4106), .ZN(n4107)
         );
  OAI21_X1 U5221 ( .B1(n4334), .B2(n4108), .A(n4107), .ZN(n4109) );
  NAND2_X1 U5222 ( .A1(n4110), .A2(n4109), .ZN(n5389) );
  NAND2_X1 U5223 ( .A1(n4114), .A2(n4113), .ZN(n4115) );
  NAND2_X1 U5224 ( .A1(n4148), .A2(n4115), .ZN(n5706) );
  AOI22_X1 U5225 ( .A1(n4317), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5226 ( .A1(n4342), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5227 ( .A1(n4319), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U5228 ( .A1(n4325), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4116) );
  NAND4_X1 U5229 ( .A1(n4119), .A2(n4118), .A3(n4117), .A4(n4116), .ZN(n4125)
         );
  AOI22_X1 U5230 ( .A1(n4344), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4197), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5231 ( .A1(n4198), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5232 ( .A1(n4748), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5233 ( .A1(n4318), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4120) );
  NAND4_X1 U5234 ( .A1(n4123), .A2(n4122), .A3(n4121), .A4(n4120), .ZN(n4124)
         );
  NOR2_X1 U5235 ( .A1(n4125), .A2(n4124), .ZN(n4127) );
  AOI22_X1 U5236 ( .A1(n3913), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n5165), .ZN(n4126) );
  OAI21_X1 U5237 ( .B1(n4334), .B2(n4127), .A(n4126), .ZN(n4128) );
  MUX2_X1 U5238 ( .A(n5706), .B(n4128), .S(n4339), .Z(n4129) );
  XNOR2_X1 U5239 ( .A(n4148), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5699)
         );
  AOI22_X1 U5240 ( .A1(n4344), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5241 ( .A1(n4352), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4135) );
  INV_X1 U5242 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4131) );
  INV_X1 U5243 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4130) );
  OAI22_X1 U5244 ( .A1(n3467), .A2(n4131), .B1(n4297), .B2(n4130), .ZN(n4132)
         );
  INV_X1 U5245 ( .A(n4132), .ZN(n4134) );
  AOI22_X1 U5246 ( .A1(n4325), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4133) );
  NAND4_X1 U5247 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4142)
         );
  AOI22_X1 U5248 ( .A1(n4197), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5249 ( .A1(n4198), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U5250 ( .A1(n4748), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5251 ( .A1(n4355), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4137) );
  NAND4_X1 U5252 ( .A1(n4140), .A2(n4139), .A3(n4138), .A4(n4137), .ZN(n4141)
         );
  OR2_X1 U5253 ( .A1(n4142), .A2(n4141), .ZN(n4146) );
  INV_X1 U5254 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4144) );
  OAI21_X1 U5255 ( .B1(n6435), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5165), 
        .ZN(n4143) );
  OAI21_X1 U5256 ( .B1(n3882), .B2(n4144), .A(n4143), .ZN(n4145) );
  AOI21_X1 U5257 ( .B1(n4366), .B2(n4146), .A(n4145), .ZN(n4147) );
  AOI21_X1 U5258 ( .B1(n5699), .B2(n4369), .A(n4147), .ZN(n5360) );
  NAND2_X1 U5259 ( .A1(n4149), .A2(n6788), .ZN(n4150) );
  NAND2_X1 U5260 ( .A1(n4182), .A2(n4150), .ZN(n5693) );
  AOI22_X1 U5261 ( .A1(n4197), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5262 ( .A1(n4319), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5263 ( .A1(n4352), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5264 ( .A1(n4748), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4151) );
  NAND4_X1 U5265 ( .A1(n4154), .A2(n4153), .A3(n4152), .A4(n4151), .ZN(n4162)
         );
  INV_X1 U5266 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4155) );
  INV_X1 U5267 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5034) );
  OAI22_X1 U5268 ( .A1(n3408), .A2(n4155), .B1(n4296), .B2(n5034), .ZN(n4156)
         );
  INV_X1 U5269 ( .A(n4156), .ZN(n4160) );
  AOI22_X1 U5270 ( .A1(n4198), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5271 ( .A1(n4353), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5272 ( .A1(n4325), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4157) );
  NAND4_X1 U5273 ( .A1(n4160), .A2(n4159), .A3(n4158), .A4(n4157), .ZN(n4161)
         );
  NOR2_X1 U5274 ( .A1(n4162), .A2(n4161), .ZN(n4164) );
  AOI22_X1 U5275 ( .A1(n4269), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5165), .ZN(n4163) );
  OAI21_X1 U5276 ( .B1(n4334), .B2(n4164), .A(n4163), .ZN(n4165) );
  MUX2_X1 U5277 ( .A(n5693), .B(n4165), .S(n4339), .Z(n4166) );
  XNOR2_X1 U5278 ( .A(n4182), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5686)
         );
  AOI22_X1 U5279 ( .A1(n4355), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5280 ( .A1(n4197), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5281 ( .A1(n4343), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5282 ( .A1(n4342), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4167) );
  NAND4_X1 U5283 ( .A1(n4170), .A2(n4169), .A3(n4168), .A4(n4167), .ZN(n4176)
         );
  AOI22_X1 U5284 ( .A1(n4344), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5285 ( .A1(n4319), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4748), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5286 ( .A1(n4199), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5287 ( .A1(n4325), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4171) );
  NAND4_X1 U5288 ( .A1(n4174), .A2(n4173), .A3(n4172), .A4(n4171), .ZN(n4175)
         );
  OR2_X1 U5289 ( .A1(n4176), .A2(n4175), .ZN(n4179) );
  INV_X1 U5290 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4177) );
  INV_X1 U5291 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5682) );
  OAI22_X1 U5292 ( .A1(n3882), .A2(n4177), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5682), .ZN(n4178) );
  AOI21_X1 U5293 ( .B1(n4366), .B2(n4179), .A(n4178), .ZN(n4180) );
  MUX2_X1 U5294 ( .A(n5686), .B(n4180), .S(n4339), .Z(n5328) );
  NAND2_X1 U5295 ( .A1(n4185), .A2(n4184), .ZN(n4186) );
  NAND2_X1 U5296 ( .A1(n4246), .A2(n4186), .ZN(n5676) );
  AOI22_X1 U5297 ( .A1(n4197), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U5298 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n4343), .B1(n4318), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U5299 ( .A1(n4344), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U5300 ( .A1(n4325), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4187) );
  NAND4_X1 U5301 ( .A1(n4190), .A2(n4189), .A3(n4188), .A4(n4187), .ZN(n4196)
         );
  AOI22_X1 U5302 ( .A1(n4319), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U5303 ( .A1(n4342), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5304 ( .A1(n4320), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U5305 ( .A1(n4355), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4191) );
  NAND4_X1 U5306 ( .A1(n4194), .A2(n4193), .A3(n4192), .A4(n4191), .ZN(n4195)
         );
  NOR2_X1 U5307 ( .A1(n4196), .A2(n4195), .ZN(n4213) );
  AOI22_X1 U5308 ( .A1(n4197), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U5309 ( .A1(n4198), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U5310 ( .A1(n4748), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U5311 ( .A1(n4355), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4200) );
  NAND4_X1 U5312 ( .A1(n4203), .A2(n4202), .A3(n4201), .A4(n4200), .ZN(n4209)
         );
  AOI22_X1 U5313 ( .A1(n4342), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U5314 ( .A1(n4344), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4206) );
  AOI22_X1 U5315 ( .A1(n4352), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U5316 ( .A1(n4325), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4204) );
  NAND4_X1 U5317 ( .A1(n4207), .A2(n4206), .A3(n4205), .A4(n4204), .ZN(n4208)
         );
  NOR2_X1 U5318 ( .A1(n4209), .A2(n4208), .ZN(n4214) );
  XNOR2_X1 U5319 ( .A(n4213), .B(n4214), .ZN(n4211) );
  AOI22_X1 U5320 ( .A1(n3913), .A2(EAX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n5165), .ZN(n4210) );
  OAI21_X1 U5321 ( .B1(n4334), .B2(n4211), .A(n4210), .ZN(n4212) );
  MUX2_X1 U5322 ( .A(n5676), .B(n4212), .S(n4339), .Z(n5315) );
  INV_X1 U5323 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5307) );
  XNOR2_X1 U5324 ( .A(n4246), .B(n5307), .ZN(n5666) );
  NAND2_X1 U5325 ( .A1(n5666), .A2(n4369), .ZN(n4230) );
  OR2_X1 U5326 ( .A1(n4214), .A2(n4213), .ZN(n4233) );
  AOI22_X1 U5327 ( .A1(n4197), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U5328 ( .A1(n4355), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4748), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4217) );
  AOI22_X1 U5329 ( .A1(n4350), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U5330 ( .A1(n4343), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4215) );
  NAND4_X1 U5331 ( .A1(n4218), .A2(n4217), .A3(n4216), .A4(n4215), .ZN(n4224)
         );
  INV_X1 U5332 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n6825) );
  AOI22_X1 U5333 ( .A1(n4319), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U5334 ( .A1(n4342), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U5335 ( .A1(n4344), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4325), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5336 ( .A1(n4352), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4219) );
  NAND4_X1 U5337 ( .A1(n4222), .A2(n4221), .A3(n4220), .A4(n4219), .ZN(n4223)
         );
  XNOR2_X1 U5338 ( .A(n4233), .B(n4231), .ZN(n4228) );
  INV_X1 U5339 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4226) );
  OAI22_X1 U5340 ( .A1(n3882), .A2(n4226), .B1(n5307), .B2(n4225), .ZN(n4227)
         );
  AOI21_X1 U5341 ( .B1(n4366), .B2(n4228), .A(n4227), .ZN(n4229) );
  NAND2_X1 U5342 ( .A1(n4230), .A2(n4229), .ZN(n5302) );
  INV_X1 U5343 ( .A(n4231), .ZN(n4232) );
  AOI22_X1 U5344 ( .A1(n4319), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4198), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4237) );
  AOI22_X1 U5345 ( .A1(n4343), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U5346 ( .A1(n4748), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U5347 ( .A1(n4350), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4234) );
  NAND4_X1 U5348 ( .A1(n4237), .A2(n4236), .A3(n4235), .A4(n4234), .ZN(n4243)
         );
  AOI22_X1 U5349 ( .A1(n4197), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4241) );
  AOI22_X1 U5350 ( .A1(n4344), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4240) );
  AOI22_X1 U5351 ( .A1(n4342), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4239) );
  AOI22_X1 U5352 ( .A1(n4325), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4238) );
  NAND4_X1 U5353 ( .A1(n4241), .A2(n4240), .A3(n4239), .A4(n4238), .ZN(n4242)
         );
  NOR2_X1 U5354 ( .A1(n4243), .A2(n4242), .ZN(n4253) );
  XNOR2_X1 U5355 ( .A(n4252), .B(n4253), .ZN(n4245) );
  AOI22_X1 U5356 ( .A1(n4269), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5165), .ZN(n4244) );
  OAI21_X1 U5357 ( .B1(n4245), .B2(n4334), .A(n4244), .ZN(n4249) );
  NAND2_X1 U5358 ( .A1(n4247), .A2(n5292), .ZN(n4248) );
  NAND2_X1 U5359 ( .A1(n4274), .A2(n4248), .ZN(n5656) );
  MUX2_X1 U5360 ( .A(n4249), .B(n5656), .S(n4369), .Z(n4250) );
  NAND2_X1 U5361 ( .A1(n4251), .A2(n4250), .ZN(n5271) );
  XNOR2_X1 U5362 ( .A(n4274), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5644)
         );
  NAND2_X1 U5363 ( .A1(n5644), .A2(n4369), .ZN(n4273) );
  NOR2_X1 U5364 ( .A1(n4253), .A2(n4252), .ZN(n4290) );
  AOI22_X1 U5365 ( .A1(n4344), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4260) );
  AOI22_X1 U5366 ( .A1(n4352), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4259) );
  INV_X1 U5367 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4255) );
  INV_X1 U5368 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4254) );
  OAI22_X1 U5369 ( .A1(n3467), .A2(n4255), .B1(n4297), .B2(n4254), .ZN(n4256)
         );
  INV_X1 U5370 ( .A(n4256), .ZN(n4258) );
  AOI22_X1 U5371 ( .A1(n4325), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4257) );
  NAND4_X1 U5372 ( .A1(n4260), .A2(n4259), .A3(n4258), .A4(n4257), .ZN(n4266)
         );
  AOI22_X1 U5373 ( .A1(n4197), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4264) );
  AOI22_X1 U5374 ( .A1(n4351), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4263) );
  AOI22_X1 U5375 ( .A1(n4320), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4262) );
  AOI22_X1 U5376 ( .A1(n4355), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4261) );
  NAND4_X1 U5377 ( .A1(n4264), .A2(n4263), .A3(n4262), .A4(n4261), .ZN(n4265)
         );
  XNOR2_X1 U5378 ( .A(n4290), .B(n4289), .ZN(n4271) );
  INV_X1 U5379 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4267) );
  AOI21_X1 U5380 ( .B1(n4267), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4268) );
  AOI21_X1 U5381 ( .B1(n4269), .B2(EAX_REG_26__SCAN_IN), .A(n4268), .ZN(n4270)
         );
  OAI21_X1 U5382 ( .B1(n4271), .B2(n4334), .A(n4270), .ZN(n4272) );
  NAND2_X1 U5383 ( .A1(n4273), .A2(n4272), .ZN(n5273) );
  INV_X1 U5384 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U5385 ( .A1(n4276), .A2(n5264), .ZN(n4277) );
  NAND2_X1 U5386 ( .A1(n4313), .A2(n4277), .ZN(n5637) );
  AOI22_X1 U5387 ( .A1(n4342), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4282) );
  AOI22_X1 U5388 ( .A1(n4355), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4281) );
  AOI22_X1 U5389 ( .A1(n4343), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4280) );
  AOI22_X1 U5390 ( .A1(n4325), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4279) );
  NAND4_X1 U5391 ( .A1(n4282), .A2(n4281), .A3(n4280), .A4(n4279), .ZN(n4288)
         );
  AOI22_X1 U5392 ( .A1(n4351), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4286) );
  AOI22_X1 U5393 ( .A1(n4344), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4285) );
  AOI22_X1 U5394 ( .A1(n4197), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4284) );
  AOI22_X1 U5395 ( .A1(n4320), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4283) );
  NAND4_X1 U5396 ( .A1(n4286), .A2(n4285), .A3(n4284), .A4(n4283), .ZN(n4287)
         );
  NOR2_X1 U5397 ( .A1(n4288), .A2(n4287), .ZN(n4295) );
  NAND2_X1 U5398 ( .A1(n4290), .A2(n4289), .ZN(n4294) );
  XNOR2_X1 U5399 ( .A(n4295), .B(n4294), .ZN(n4292) );
  AOI22_X1 U5400 ( .A1(n3913), .A2(EAX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5165), .ZN(n4291) );
  OAI21_X1 U5401 ( .B1(n4292), .B2(n4334), .A(n4291), .ZN(n4293) );
  MUX2_X1 U5402 ( .A(n5637), .B(n4293), .S(n4339), .Z(n5259) );
  NOR2_X1 U5403 ( .A1(n4295), .A2(n4294), .ZN(n4333) );
  NOR2_X1 U5404 ( .A1(n4296), .A2(n6842), .ZN(n4300) );
  INV_X1 U5405 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4298) );
  OAI22_X1 U5406 ( .A1(n3408), .A2(n4298), .B1(n4297), .B2(n4945), .ZN(n4299)
         );
  AOI211_X1 U5407 ( .C1(INSTQUEUE_REG_6__5__SCAN_IN), .C2(n4343), .A(n4300), 
        .B(n4299), .ZN(n4308) );
  AOI22_X1 U5408 ( .A1(n4197), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4304) );
  AOI22_X1 U5409 ( .A1(n4351), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4303) );
  AOI22_X1 U5410 ( .A1(n4355), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4302) );
  AOI22_X1 U5411 ( .A1(n4320), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4301) );
  AND4_X1 U5412 ( .A1(n4304), .A2(n4303), .A3(n4302), .A4(n4301), .ZN(n4307)
         );
  AOI22_X1 U5413 ( .A1(n4352), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4306) );
  AOI22_X1 U5414 ( .A1(n4325), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4305) );
  NAND4_X1 U5415 ( .A1(n4308), .A2(n4307), .A3(n4306), .A4(n4305), .ZN(n4332)
         );
  XNOR2_X1 U5416 ( .A(n4333), .B(n4332), .ZN(n4310) );
  AOI22_X1 U5417 ( .A1(n3913), .A2(EAX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n5165), .ZN(n4309) );
  OAI21_X1 U5418 ( .B1(n4310), .B2(n4334), .A(n4309), .ZN(n4312) );
  INV_X1 U5419 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4311) );
  XNOR2_X1 U5420 ( .A(n4313), .B(n4311), .ZN(n5628) );
  INV_X1 U5421 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4314) );
  NAND2_X1 U5422 ( .A1(n4315), .A2(n4314), .ZN(n4316) );
  NAND2_X1 U5423 ( .A1(n4374), .A2(n4316), .ZN(n5620) );
  AOI22_X1 U5424 ( .A1(n4351), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4317), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U5425 ( .A1(n4344), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4323) );
  AOI22_X1 U5426 ( .A1(n4319), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U5427 ( .A1(n4320), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4321) );
  NAND4_X1 U5428 ( .A1(n4324), .A2(n4323), .A3(n4322), .A4(n4321), .ZN(n4331)
         );
  AOI22_X1 U5429 ( .A1(n4197), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4355), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4329) );
  AOI22_X1 U5430 ( .A1(n4343), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4352), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4328) );
  AOI22_X1 U5431 ( .A1(n4342), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4327) );
  AOI22_X1 U5432 ( .A1(n4325), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4326) );
  NAND4_X1 U5433 ( .A1(n4329), .A2(n4328), .A3(n4327), .A4(n4326), .ZN(n4330)
         );
  NOR2_X1 U5434 ( .A1(n4331), .A2(n4330), .ZN(n4341) );
  NAND2_X1 U5435 ( .A1(n4333), .A2(n4332), .ZN(n4340) );
  XNOR2_X1 U5436 ( .A(n4341), .B(n4340), .ZN(n4335) );
  NOR2_X1 U5437 ( .A1(n4335), .A2(n4334), .ZN(n4338) );
  INV_X1 U5438 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6807) );
  NOR2_X1 U5439 ( .A1(n6435), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4336)
         );
  OAI22_X1 U5440 ( .A1(n3882), .A2(n6807), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4336), .ZN(n4337) );
  OAI22_X1 U5441 ( .A1(n5620), .A2(n4339), .B1(n4338), .B2(n4337), .ZN(n4402)
         );
  XNOR2_X1 U5442 ( .A(n4374), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5238)
         );
  NOR2_X1 U5443 ( .A1(n4341), .A2(n4340), .ZN(n4363) );
  AOI22_X1 U5444 ( .A1(n4342), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4319), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U5445 ( .A1(n4748), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U5446 ( .A1(n4344), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4343), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4347) );
  AOI22_X1 U5447 ( .A1(n4325), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4345), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4346) );
  NAND4_X1 U5448 ( .A1(n4349), .A2(n4348), .A3(n4347), .A4(n4346), .ZN(n4361)
         );
  AOI22_X1 U5449 ( .A1(n4351), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4350), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4359) );
  AOI22_X1 U5450 ( .A1(n4352), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4318), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4358) );
  AOI22_X1 U5451 ( .A1(n4197), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4353), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4357) );
  AOI22_X1 U5452 ( .A1(n4355), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4354), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4356) );
  NAND4_X1 U5453 ( .A1(n4359), .A2(n4358), .A3(n4357), .A4(n4356), .ZN(n4360)
         );
  NOR2_X1 U5454 ( .A1(n4361), .A2(n4360), .ZN(n4362) );
  XNOR2_X1 U5455 ( .A(n4363), .B(n4362), .ZN(n4367) );
  INV_X1 U5456 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6731) );
  OAI21_X1 U5457 ( .B1(n6435), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5165), 
        .ZN(n4364) );
  OAI21_X1 U5458 ( .B1(n3882), .B2(n6731), .A(n4364), .ZN(n4365) );
  AOI21_X1 U5459 ( .B1(n4367), .B2(n4366), .A(n4365), .ZN(n4368) );
  AOI22_X1 U5460 ( .A1(n4269), .A2(EAX_REG_31__SCAN_IN), .B1(n4370), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4371) );
  INV_X1 U5461 ( .A(n4371), .ZN(n4372) );
  INV_X1 U5462 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U5463 ( .A1(n5215), .A2(n6890), .ZN(n4375) );
  NAND2_X1 U5464 ( .A1(n4376), .A2(n4375), .ZN(U2796) );
  NAND2_X1 U5465 ( .A1(n4377), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6641) );
  NAND2_X1 U5466 ( .A1(n5215), .A2(n5804), .ZN(n4390) );
  NAND2_X1 U5467 ( .A1(n4378), .A2(n6578), .ZN(n4379) );
  NAND2_X1 U5468 ( .A1(n4379), .A2(n6722), .ZN(n4380) );
  NAND2_X1 U5469 ( .A1(n6722), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4382) );
  NAND2_X1 U5470 ( .A1(n6435), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4381) );
  AND2_X1 U5471 ( .A1(n4382), .A2(n4381), .ZN(n4518) );
  INV_X1 U5472 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6699) );
  NOR2_X1 U5473 ( .A1(n3820), .A2(n6699), .ZN(n4392) );
  NOR2_X1 U5474 ( .A1(n5784), .A2(n4383), .ZN(n4384) );
  AOI211_X1 U5475 ( .C1(n5225), .C2(n5787), .A(n4392), .B(n4384), .ZN(n4389)
         );
  NAND2_X1 U5476 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4387) );
  NAND3_X1 U5477 ( .A1(n4385), .A2(n3808), .A3(n5807), .ZN(n4386) );
  OAI22_X1 U5478 ( .A1(n5616), .A2(n4387), .B1(n5651), .B2(n4386), .ZN(n4388)
         );
  NOR3_X1 U5479 ( .A1(n4391), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n3808), 
        .ZN(n4393) );
  AOI21_X1 U5480 ( .B1(n5504), .B2(n6359), .A(n4394), .ZN(n4400) );
  INV_X1 U5481 ( .A(n5936), .ZN(n5996) );
  NOR2_X1 U5482 ( .A1(n5996), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4395)
         );
  OAI21_X1 U5483 ( .B1(n4396), .B2(n4395), .A(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n4399) );
  NAND3_X1 U5484 ( .A1(n4400), .A2(n4399), .A3(n4398), .ZN(U2987) );
  INV_X1 U5485 ( .A(n4425), .ZN(n4404) );
  NAND2_X1 U5486 ( .A1(n4401), .A2(n4402), .ZN(n4403) );
  INV_X1 U5487 ( .A(n5208), .ZN(n4455) );
  NOR2_X1 U5488 ( .A1(n3426), .A2(n4795), .ZN(n4408) );
  NOR2_X1 U5489 ( .A1(n4588), .A2(n4530), .ZN(n4407) );
  NOR2_X1 U5490 ( .A1(n4405), .A2(n3461), .ZN(n4406) );
  NAND4_X1 U5491 ( .A1(n4409), .A2(n4408), .A3(n4407), .A4(n4406), .ZN(n4525)
         );
  INV_X2 U5492 ( .A(n6233), .ZN(n5544) );
  NAND2_X1 U5493 ( .A1(n5622), .A2(n6233), .ZN(n4423) );
  NAND2_X1 U5494 ( .A1(n4413), .A2(n3201), .ZN(n4415) );
  NAND2_X1 U5495 ( .A1(n4415), .A2(n4414), .ZN(n4416) );
  NOR2_X1 U5496 ( .A1(n5250), .A2(n4416), .ZN(n4417) );
  INV_X1 U5497 ( .A(n4530), .ZN(n5558) );
  XNOR2_X2 U5498 ( .A(n4425), .B(n4424), .ZN(n5562) );
  INV_X1 U5499 ( .A(n5562), .ZN(n4426) );
  NAND2_X1 U5500 ( .A1(n5238), .A2(n5787), .ZN(n4428) );
  OAI211_X1 U5501 ( .C1(n5784), .C2(n5235), .A(n4428), .B(n4427), .ZN(n4429)
         );
  INV_X1 U5502 ( .A(HOLD), .ZN(n6750) );
  NAND2_X1 U5503 ( .A1(n4440), .A2(STATE_REG_1__SCAN_IN), .ZN(n4445) );
  NAND2_X1 U5504 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4434) );
  INV_X1 U5505 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6645) );
  INV_X1 U5506 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4436) );
  NOR2_X1 U5507 ( .A1(n6645), .A2(n4436), .ZN(n6648) );
  NAND2_X1 U5508 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6649) );
  INV_X1 U5509 ( .A(n6649), .ZN(n4433) );
  AOI21_X1 U5510 ( .B1(n4434), .B2(n6648), .A(n4433), .ZN(n4435) );
  OAI211_X1 U5511 ( .C1(n6750), .C2(n4445), .A(n6716), .B(n4435), .ZN(U3182)
         );
  INV_X1 U5512 ( .A(NA_N), .ZN(n6647) );
  AOI221_X1 U5513 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6647), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6651) );
  AOI21_X1 U5514 ( .B1(HOLD), .B2(n4437), .A(n4436), .ZN(n4438) );
  OAI22_X1 U5515 ( .A1(n4438), .A2(n6099), .B1(n6712), .B2(n4445), .ZN(n4439)
         );
  OR2_X1 U5516 ( .A1(n6651), .A2(n4439), .ZN(U3181) );
  NAND2_X1 U5517 ( .A1(n6099), .A2(n4440), .ZN(n6698) );
  INV_X1 U5518 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6802) );
  OAI222_X1 U5519 ( .A1(n6694), .A2(n6148), .B1(n6698), .B2(n6668), .C1(n6802), 
        .C2(n6099), .ZN(U3195) );
  INV_X1 U5520 ( .A(REIP_REG_6__SCAN_IN), .ZN(n5059) );
  INV_X1 U5521 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6795) );
  OAI222_X1 U5522 ( .A1(n6698), .A2(n6662), .B1(n6694), .B2(n5059), .C1(n6099), 
        .C2(n6795), .ZN(U3189) );
  INV_X1 U5523 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6786) );
  INV_X1 U5524 ( .A(REIP_REG_20__SCAN_IN), .ZN(n4441) );
  OAI222_X1 U5525 ( .A1(n6698), .A2(n5691), .B1(n6099), .B2(n6786), .C1(n6694), 
        .C2(n4441), .ZN(U3203) );
  INV_X1 U5526 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6672) );
  INV_X1 U5527 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6822) );
  INV_X1 U5528 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6670) );
  OAI222_X1 U5529 ( .A1(n6698), .A2(n6672), .B1(n6099), .B2(n6822), .C1(n6694), 
        .C2(n6670), .ZN(U3198) );
  INV_X1 U5530 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4443) );
  NAND2_X1 U5531 ( .A1(M_IO_N_REG_SCAN_IN), .A2(n6673), .ZN(n4442) );
  OAI21_X1 U5532 ( .B1(n6673), .B2(n4443), .A(n4442), .ZN(U3473) );
  NOR2_X1 U5533 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6100) );
  OAI21_X1 U5534 ( .B1(n6100), .B2(D_C_N_REG_SCAN_IN), .A(n6673), .ZN(n4444)
         );
  OAI21_X1 U5535 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6673), .A(n4444), .ZN(
        U2791) );
  INV_X1 U5536 ( .A(ADS_N_REG_SCAN_IN), .ZN(n4447) );
  NAND2_X1 U5537 ( .A1(n4445), .A2(STATE_REG_0__SCAN_IN), .ZN(n4446) );
  OAI21_X1 U5538 ( .B1(n6099), .B2(n4447), .A(n6644), .ZN(U2789) );
  INV_X1 U5539 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U5540 ( .A1(BE_N_REG_0__SCAN_IN), .A2(n6673), .ZN(n4448) );
  OAI21_X1 U5541 ( .B1(n6673), .B2(n6708), .A(n4448), .ZN(U3448) );
  INV_X1 U5542 ( .A(n4456), .ZN(n4450) );
  OAI22_X1 U5543 ( .A1(n4492), .A2(n5479), .B1(n4450), .B2(n4449), .ZN(n4454)
         );
  OAI21_X1 U5544 ( .B1(n4454), .B2(n4455), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n4452) );
  NAND3_X1 U5545 ( .A1(n5164), .A2(STATE2_REG_0__SCAN_IN), .A3(n5165), .ZN(
        n4451) );
  NAND2_X1 U5546 ( .A1(n4452), .A2(n4451), .ZN(U2790) );
  NAND2_X1 U5547 ( .A1(n6713), .A2(n6711), .ZN(n5220) );
  AOI21_X1 U5548 ( .B1(n5220), .B2(n6716), .A(READY_N), .ZN(n4453) );
  NOR2_X1 U5549 ( .A1(n4454), .A2(n4453), .ZN(n4788) );
  NOR2_X1 U5550 ( .A1(n4788), .A2(n4455), .ZN(n6103) );
  INV_X1 U5551 ( .A(MORE_REG_SCAN_IN), .ZN(n4464) );
  AND3_X1 U5552 ( .A1(n4790), .A2(n4529), .A3(n4456), .ZN(n4457) );
  MUX2_X1 U5553 ( .A(n4457), .B(n4506), .S(n4492), .Z(n4461) );
  NAND2_X1 U5554 ( .A1(n4459), .A2(n4458), .ZN(n4460) );
  AND2_X1 U5555 ( .A1(n4461), .A2(n4460), .ZN(n4791) );
  INV_X1 U5556 ( .A(n4791), .ZN(n4462) );
  NAND2_X1 U5557 ( .A1(n6103), .A2(n4462), .ZN(n4463) );
  OAI21_X1 U5558 ( .B1(n6103), .B2(n4464), .A(n4463), .ZN(U3471) );
  INV_X1 U5559 ( .A(n5219), .ZN(n5375) );
  INV_X1 U5560 ( .A(n4465), .ZN(n4468) );
  AOI211_X1 U5561 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4466), .A(n5375), .B(
        n4468), .ZN(n4467) );
  INV_X1 U5562 ( .A(n4467), .ZN(U2788) );
  OAI21_X1 U5563 ( .B1(n4469), .B2(n6712), .A(n4468), .ZN(n4470) );
  INV_X1 U5564 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n6791) );
  INV_X1 U5565 ( .A(n6324), .ZN(n6285) );
  AOI22_X1 U5566 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6322), .B1(n6285), .B2(
        DATAI_15_), .ZN(n4471) );
  OAI21_X1 U5567 ( .B1(n6273), .B2(n6791), .A(n4471), .ZN(U2954) );
  MUX2_X1 U5568 ( .A(n4506), .B(n4529), .S(n4492), .Z(n4485) );
  NAND2_X1 U5569 ( .A1(n4473), .A2(n6716), .ZN(n4474) );
  NAND2_X1 U5570 ( .A1(n4474), .A2(n6712), .ZN(n4475) );
  AOI21_X1 U5571 ( .B1(n4761), .B2(n3551), .A(n4475), .ZN(n4483) );
  INV_X1 U5572 ( .A(n4476), .ZN(n4477) );
  INV_X1 U5573 ( .A(n4527), .ZN(n4481) );
  INV_X1 U5574 ( .A(n4478), .ZN(n4479) );
  NAND3_X1 U5575 ( .A1(n4481), .A2(n4480), .A3(n4479), .ZN(n4482) );
  AOI21_X1 U5576 ( .B1(n4492), .B2(n4483), .A(n4482), .ZN(n4484) );
  NAND2_X1 U5577 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n6016) );
  NOR2_X1 U5578 ( .A1(n6016), .A2(n6722), .ZN(n6643) );
  AND2_X1 U5579 ( .A1(n6643), .A2(FLUSH_REG_SCAN_IN), .ZN(n4486) );
  AOI21_X1 U5580 ( .B1(n4782), .B2(n5208), .A(n4486), .ZN(n4500) );
  NAND2_X1 U5581 ( .A1(n6722), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4487) );
  INV_X1 U5582 ( .A(n6040), .ZN(n5197) );
  INV_X1 U5583 ( .A(n5498), .ZN(n6515) );
  AND3_X1 U5584 ( .A1(n3784), .A2(n3551), .A3(n3554), .ZN(n4488) );
  NAND2_X1 U5585 ( .A1(n4498), .A2(n4488), .ZN(n4490) );
  OR2_X1 U5586 ( .A1(n4490), .A2(n4489), .ZN(n4763) );
  INV_X1 U5587 ( .A(n4763), .ZN(n4491) );
  OAI22_X1 U5588 ( .A1(n6515), .A2(n4491), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4759), .ZN(n4758) );
  AOI21_X1 U5589 ( .B1(n4758), .B2(n6050), .A(STATE2_REG_1__SCAN_IN), .ZN(
        n4493) );
  AND2_X1 U5590 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        STATE2_REG_1__SCAN_IN), .ZN(n5190) );
  OAI22_X1 U5591 ( .A1(n4493), .A2(n5190), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6036), .ZN(n4494) );
  NOR2_X1 U5592 ( .A1(n4761), .A2(n4472), .ZN(n4757) );
  AOI22_X1 U5593 ( .A1(n5197), .A2(n4494), .B1(n5164), .B2(n4757), .ZN(n4495)
         );
  OAI21_X1 U5594 ( .B1(n4472), .B2(n5197), .A(n4495), .ZN(U3461) );
  INV_X1 U5595 ( .A(n4674), .ZN(n6581) );
  OR2_X1 U5596 ( .A1(n4496), .A2(n6581), .ZN(n4497) );
  XNOR2_X1 U5597 ( .A(n4497), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5491)
         );
  INV_X1 U5598 ( .A(n4498), .ZN(n4780) );
  NAND3_X1 U5599 ( .A1(n5491), .A2(n4780), .A3(n5164), .ZN(n4499) );
  OAI22_X1 U5600 ( .A1(n5197), .A2(n4784), .B1(n4500), .B2(n4499), .ZN(U3455)
         );
  INV_X1 U5601 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4501) );
  AOI22_X1 U5602 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4501), .B2(n4554), .ZN(n5188)
         );
  INV_X1 U5603 ( .A(n4502), .ZN(n4512) );
  NOR3_X1 U5604 ( .A1(n6036), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4512), 
        .ZN(n4511) );
  INV_X1 U5605 ( .A(n4503), .ZN(n6207) );
  XNOR2_X1 U5606 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4505) );
  XNOR2_X1 U5607 ( .A(n4502), .B(n4768), .ZN(n4507) );
  INV_X1 U5608 ( .A(n4507), .ZN(n4504) );
  OAI22_X1 U5609 ( .A1(n4761), .A2(n4505), .B1(n4750), .B2(n4504), .ZN(n4509)
         );
  AND2_X1 U5610 ( .A1(n4506), .A2(n4529), .ZN(n4740) );
  NOR2_X1 U5611 ( .A1(n4740), .A2(n4507), .ZN(n4508) );
  AOI211_X1 U5612 ( .C1(n6207), .C2(n4763), .A(n4509), .B(n4508), .ZN(n4767)
         );
  INV_X1 U5613 ( .A(n5164), .ZN(n6038) );
  NOR2_X1 U5614 ( .A1(n4767), .A2(n6038), .ZN(n4510) );
  AOI211_X1 U5615 ( .C1(n5190), .C2(n5188), .A(n4511), .B(n4510), .ZN(n4514)
         );
  INV_X1 U5616 ( .A(n6036), .ZN(n5193) );
  AOI21_X1 U5617 ( .B1(n5193), .B2(n4512), .A(n6040), .ZN(n4513) );
  OAI22_X1 U5618 ( .A1(n4514), .A2(n6040), .B1(n4513), .B2(n4768), .ZN(U3459)
         );
  OAI21_X1 U5619 ( .B1(n4515), .B2(n4517), .A(n4516), .ZN(n5503) );
  NAND2_X1 U5620 ( .A1(n5784), .A2(n4518), .ZN(n4520) );
  INV_X1 U5621 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4519) );
  NOR2_X1 U5622 ( .A1(n3820), .A2(n4519), .ZN(n6383) );
  AOI21_X1 U5623 ( .B1(n4520), .B2(PHYADDRPOINTER_REG_0__SCAN_IN), .A(n6383), 
        .ZN(n4523) );
  OR2_X1 U5624 ( .A1(n4521), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6382)
         );
  NAND3_X1 U5625 ( .A1(n6382), .A2(n6380), .A3(n6336), .ZN(n4522) );
  OAI211_X1 U5626 ( .C1(n5503), .C2(n5797), .A(n4523), .B(n4522), .ZN(U2986)
         );
  NOR2_X1 U5627 ( .A1(n4525), .A2(n4524), .ZN(n4526) );
  NAND2_X1 U5628 ( .A1(n3431), .A2(n4530), .ZN(n4531) );
  INV_X1 U5629 ( .A(n4531), .ZN(n4532) );
  INV_X1 U5630 ( .A(DATAI_0_), .ZN(n6295) );
  INV_X1 U5631 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6270) );
  OAI222_X1 U5632 ( .A1(n5503), .A2(n5591), .B1(n5180), .B2(n6295), .C1(n5213), 
        .C2(n6270), .ZN(U2891) );
  INV_X1 U5633 ( .A(n6016), .ZN(n4535) );
  NAND2_X1 U5634 ( .A1(n4535), .A2(n6722), .ZN(n6246) );
  INV_X2 U5635 ( .A(n6246), .ZN(n6267) );
  AOI222_X1 U5636 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6239), .B1(n6266), .B2(
        DATAO_REG_30__SCAN_IN), .C1(n6267), .C2(UWORD_REG_14__SCAN_IN), .ZN(
        n4536) );
  INV_X1 U5637 ( .A(n4536), .ZN(U2893) );
  AOI222_X1 U5638 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6239), .B1(n6266), .B2(
        DATAO_REG_27__SCAN_IN), .C1(n6267), .C2(UWORD_REG_11__SCAN_IN), .ZN(
        n4537) );
  INV_X1 U5639 ( .A(n4537), .ZN(U2896) );
  AOI222_X1 U5640 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6239), .B1(n6266), .B2(
        DATAO_REG_24__SCAN_IN), .C1(n6267), .C2(UWORD_REG_8__SCAN_IN), .ZN(
        n4538) );
  INV_X1 U5641 ( .A(n4538), .ZN(U2899) );
  AOI222_X1 U5642 ( .A1(EAX_REG_20__SCAN_IN), .A2(n6239), .B1(n6266), .B2(
        DATAO_REG_20__SCAN_IN), .C1(n6267), .C2(UWORD_REG_4__SCAN_IN), .ZN(
        n4539) );
  INV_X1 U5643 ( .A(n4539), .ZN(U2903) );
  AOI222_X1 U5644 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6239), .B1(n6266), .B2(
        DATAO_REG_25__SCAN_IN), .C1(n6267), .C2(UWORD_REG_9__SCAN_IN), .ZN(
        n4540) );
  INV_X1 U5645 ( .A(n4540), .ZN(U2898) );
  AOI222_X1 U5646 ( .A1(n6266), .A2(DATAO_REG_17__SCAN_IN), .B1(n6239), .B2(
        EAX_REG_17__SCAN_IN), .C1(n6267), .C2(UWORD_REG_1__SCAN_IN), .ZN(n4541) );
  INV_X1 U5647 ( .A(n4541), .ZN(U2906) );
  AOI222_X1 U5648 ( .A1(n6266), .A2(DATAO_REG_29__SCAN_IN), .B1(n6239), .B2(
        EAX_REG_29__SCAN_IN), .C1(n6267), .C2(UWORD_REG_13__SCAN_IN), .ZN(
        n4542) );
  INV_X1 U5649 ( .A(n4542), .ZN(U2894) );
  INV_X1 U5650 ( .A(n4544), .ZN(n4545) );
  OAI21_X1 U5651 ( .B1(n4546), .B2(n4543), .A(n4545), .ZN(n6330) );
  INV_X1 U5652 ( .A(DATAI_2_), .ZN(n6299) );
  INV_X1 U5653 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6810) );
  OAI222_X1 U5654 ( .A1(n6330), .A2(n5591), .B1(n5180), .B2(n6299), .C1(n5213), 
        .C2(n6810), .ZN(U2889) );
  OAI21_X1 U5655 ( .B1(n4544), .B2(n4549), .A(n4548), .ZN(n5069) );
  INV_X1 U5656 ( .A(DATAI_3_), .ZN(n6301) );
  INV_X1 U5657 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6262) );
  OAI222_X1 U5658 ( .A1(n5069), .A2(n5591), .B1(n5180), .B2(n6301), .C1(n5213), 
        .C2(n6262), .ZN(U2888) );
  OAI21_X1 U5659 ( .B1(n4552), .B2(n4551), .A(n4550), .ZN(n5163) );
  INV_X1 U5660 ( .A(n4663), .ZN(n4556) );
  NAND2_X1 U5661 ( .A1(n5936), .A2(n4553), .ZN(n4555) );
  MUX2_X1 U5662 ( .A(n4556), .B(n4555), .S(n4554), .Z(n4561) );
  XNOR2_X1 U5663 ( .A(n4557), .B(n4558), .ZN(n5051) );
  INV_X1 U5664 ( .A(REIP_REG_1__SCAN_IN), .ZN(n4559) );
  NOR2_X1 U5665 ( .A1(n3820), .A2(n4559), .ZN(n5160) );
  AOI21_X1 U5666 ( .B1(n6359), .B2(n5051), .A(n5160), .ZN(n4560) );
  OAI211_X1 U5667 ( .C1(n6015), .C2(n5163), .A(n4561), .B(n4560), .ZN(U3017)
         );
  INV_X1 U5668 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U5669 ( .A1(n6266), .A2(DATAO_REG_28__SCAN_IN), .ZN(n4563) );
  NAND2_X1 U5670 ( .A1(n6267), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4562) );
  OAI211_X1 U5671 ( .C1(n4564), .C2(n4575), .A(n4563), .B(n4562), .ZN(U2895)
         );
  INV_X1 U5672 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U5673 ( .A1(n6266), .A2(DATAO_REG_16__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U5674 ( .A1(n6267), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4565) );
  OAI211_X1 U5675 ( .C1(n4567), .C2(n4575), .A(n4566), .B(n4565), .ZN(U2907)
         );
  INV_X1 U5676 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4570) );
  NAND2_X1 U5677 ( .A1(n6266), .A2(DATAO_REG_18__SCAN_IN), .ZN(n4569) );
  NAND2_X1 U5678 ( .A1(n6267), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4568) );
  OAI211_X1 U5679 ( .C1(n4570), .C2(n4575), .A(n4569), .B(n4568), .ZN(U2905)
         );
  NAND2_X1 U5680 ( .A1(n6266), .A2(DATAO_REG_22__SCAN_IN), .ZN(n4572) );
  NAND2_X1 U5681 ( .A1(n6267), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4571) );
  OAI211_X1 U5682 ( .C1(n4177), .C2(n4575), .A(n4572), .B(n4571), .ZN(U2901)
         );
  INV_X1 U5683 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4576) );
  NAND2_X1 U5684 ( .A1(n6266), .A2(DATAO_REG_21__SCAN_IN), .ZN(n4574) );
  NAND2_X1 U5685 ( .A1(n6267), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4573) );
  OAI211_X1 U5686 ( .C1(n4576), .C2(n4575), .A(n4574), .B(n4573), .ZN(U2902)
         );
  INV_X1 U5687 ( .A(DATAI_6_), .ZN(n6307) );
  INV_X1 U5688 ( .A(n4577), .ZN(n6718) );
  NAND2_X1 U5689 ( .A1(n6718), .A2(n6016), .ZN(n4578) );
  NOR2_X2 U5690 ( .A1(n6307), .A2(n6018), .ZN(n6624) );
  INV_X1 U5691 ( .A(n6624), .ZN(n4893) );
  NOR2_X1 U5692 ( .A1(n4503), .A2(n4583), .ZN(n4806) );
  INV_X1 U5693 ( .A(n4619), .ZN(n4584) );
  AOI21_X1 U5694 ( .B1(n4951), .B2(n4806), .A(n4584), .ZN(n4590) );
  INV_X1 U5695 ( .A(n4590), .ZN(n4585) );
  AOI22_X1 U5696 ( .A1(n4585), .A2(n6437), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4676), .ZN(n4620) );
  NAND2_X1 U5697 ( .A1(n5804), .A2(DATAI_30_), .ZN(n6628) );
  INV_X1 U5698 ( .A(n6628), .ZN(n4976) );
  INV_X1 U5699 ( .A(n4627), .ZN(n4586) );
  INV_X1 U5700 ( .A(n5096), .ZN(n4737) );
  NAND2_X1 U5701 ( .A1(n5804), .A2(DATAI_22_), .ZN(n6558) );
  OR2_X1 U5702 ( .A1(n4618), .A2(n4588), .ZN(n6554) );
  OAI22_X1 U5703 ( .A1(n4941), .A2(n6558), .B1(n4619), .B2(n6554), .ZN(n4589)
         );
  AOI21_X1 U5704 ( .B1(n4976), .B2(n4737), .A(n4589), .ZN(n4594) );
  AOI21_X1 U5705 ( .B1(n4673), .B2(n6021), .A(n5797), .ZN(n4591) );
  OAI21_X1 U5706 ( .B1(n4591), .B2(n6582), .A(n4590), .ZN(n4592) );
  NAND2_X1 U5707 ( .A1(n4616), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4593)
         );
  OAI211_X1 U5708 ( .C1(n4893), .C2(n4620), .A(n4594), .B(n4593), .ZN(U3146)
         );
  NAND2_X1 U5709 ( .A1(n5804), .A2(DATAI_29_), .ZN(n6622) );
  NAND2_X1 U5710 ( .A1(n4616), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4598)
         );
  NAND2_X1 U5711 ( .A1(n5804), .A2(DATAI_21_), .ZN(n6553) );
  INV_X1 U5712 ( .A(DATAI_5_), .ZN(n6305) );
  NOR2_X2 U5713 ( .A1(n6305), .A2(n6018), .ZN(n6618) );
  INV_X1 U5714 ( .A(n6618), .ZN(n4905) );
  OAI22_X1 U5715 ( .A1(n4620), .A2(n4905), .B1(n4619), .B2(n6549), .ZN(n4596)
         );
  AOI21_X1 U5716 ( .B1(n4868), .B2(n6619), .A(n4596), .ZN(n4597) );
  OAI211_X1 U5717 ( .C1(n5096), .C2(n6622), .A(n4598), .B(n4597), .ZN(U3145)
         );
  NAND2_X1 U5718 ( .A1(n5804), .A2(DATAI_28_), .ZN(n6616) );
  NAND2_X1 U5719 ( .A1(n4616), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4602)
         );
  NAND2_X1 U5720 ( .A1(n5804), .A2(DATAI_20_), .ZN(n6545) );
  INV_X1 U5721 ( .A(n6545), .ZN(n6613) );
  INV_X1 U5722 ( .A(DATAI_4_), .ZN(n6303) );
  NOR2_X2 U5723 ( .A1(n6303), .A2(n6018), .ZN(n6612) );
  INV_X1 U5724 ( .A(n6612), .ZN(n4909) );
  OR2_X1 U5725 ( .A1(n4618), .A2(n4599), .ZN(n6544) );
  OAI22_X1 U5726 ( .A1(n4620), .A2(n4909), .B1(n4619), .B2(n6544), .ZN(n4600)
         );
  AOI21_X1 U5727 ( .B1(n4868), .B2(n6613), .A(n4600), .ZN(n4601) );
  OAI211_X1 U5728 ( .C1(n5096), .C2(n6616), .A(n4602), .B(n4601), .ZN(U3144)
         );
  NAND2_X1 U5729 ( .A1(n5804), .A2(DATAI_27_), .ZN(n6610) );
  NAND2_X1 U5730 ( .A1(n4616), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4606)
         );
  NAND2_X1 U5731 ( .A1(n5804), .A2(DATAI_19_), .ZN(n6540) );
  INV_X1 U5732 ( .A(n6540), .ZN(n6607) );
  NOR2_X2 U5733 ( .A1(n6301), .A2(n6018), .ZN(n6606) );
  INV_X1 U5734 ( .A(n6606), .ZN(n4901) );
  OAI22_X1 U5735 ( .A1(n4620), .A2(n4901), .B1(n4619), .B2(n6539), .ZN(n4604)
         );
  AOI21_X1 U5736 ( .B1(n4868), .B2(n6607), .A(n4604), .ZN(n4605) );
  OAI211_X1 U5737 ( .C1(n5096), .C2(n6610), .A(n4606), .B(n4605), .ZN(U3143)
         );
  NAND2_X1 U5738 ( .A1(n5804), .A2(DATAI_24_), .ZN(n6592) );
  NAND2_X1 U5739 ( .A1(n4616), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4609)
         );
  NAND2_X1 U5740 ( .A1(n5804), .A2(DATAI_16_), .ZN(n6528) );
  INV_X1 U5741 ( .A(n6528), .ZN(n6589) );
  INV_X1 U5742 ( .A(n6577), .ZN(n5004) );
  OR2_X1 U5743 ( .A1(n4618), .A2(n3530), .ZN(n6511) );
  OAI22_X1 U5744 ( .A1(n4620), .A2(n5004), .B1(n4619), .B2(n6511), .ZN(n4607)
         );
  AOI21_X1 U5745 ( .B1(n4868), .B2(n6589), .A(n4607), .ZN(n4608) );
  OAI211_X1 U5746 ( .C1(n5096), .C2(n6592), .A(n4609), .B(n4608), .ZN(U3140)
         );
  NAND2_X1 U5747 ( .A1(n5804), .A2(DATAI_25_), .ZN(n6598) );
  NAND2_X1 U5748 ( .A1(n4616), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4612)
         );
  NAND2_X1 U5749 ( .A1(n5804), .A2(DATAI_17_), .ZN(n6530) );
  INV_X1 U5750 ( .A(DATAI_1_), .ZN(n6297) );
  NOR2_X2 U5751 ( .A1(n6297), .A2(n6018), .ZN(n6594) );
  INV_X1 U5752 ( .A(n6594), .ZN(n4917) );
  OR2_X1 U5753 ( .A1(n4618), .A2(n2972), .ZN(n6529) );
  OAI22_X1 U5754 ( .A1(n4620), .A2(n4917), .B1(n4619), .B2(n6529), .ZN(n4610)
         );
  AOI21_X1 U5755 ( .B1(n4868), .B2(n6595), .A(n4610), .ZN(n4611) );
  OAI211_X1 U5756 ( .C1(n5096), .C2(n6598), .A(n4612), .B(n4611), .ZN(U3141)
         );
  NAND2_X1 U5757 ( .A1(n5804), .A2(DATAI_31_), .ZN(n6639) );
  NAND2_X1 U5758 ( .A1(n4616), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4615)
         );
  NAND2_X1 U5759 ( .A1(n5804), .A2(DATAI_23_), .ZN(n6561) );
  INV_X1 U5760 ( .A(DATAI_7_), .ZN(n6837) );
  NOR2_X2 U5761 ( .A1(n6837), .A2(n6018), .ZN(n6631) );
  INV_X1 U5762 ( .A(n6631), .ZN(n4897) );
  OAI22_X1 U5763 ( .A1(n4620), .A2(n4897), .B1(n4619), .B2(n6560), .ZN(n4613)
         );
  AOI21_X1 U5764 ( .B1(n4868), .B2(n6634), .A(n4613), .ZN(n4614) );
  OAI211_X1 U5765 ( .C1(n5096), .C2(n6639), .A(n4615), .B(n4614), .ZN(U3147)
         );
  NAND2_X1 U5766 ( .A1(n5804), .A2(DATAI_26_), .ZN(n6604) );
  NAND2_X1 U5767 ( .A1(n4616), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4623)
         );
  NAND2_X1 U5768 ( .A1(n5804), .A2(DATAI_18_), .ZN(n6535) );
  INV_X1 U5769 ( .A(n6535), .ZN(n6601) );
  NOR2_X2 U5770 ( .A1(n6299), .A2(n6018), .ZN(n6600) );
  INV_X1 U5771 ( .A(n6600), .ZN(n4913) );
  OR2_X1 U5772 ( .A1(n4618), .A2(n4617), .ZN(n6534) );
  OAI22_X1 U5773 ( .A1(n4620), .A2(n4913), .B1(n4619), .B2(n6534), .ZN(n4621)
         );
  AOI21_X1 U5774 ( .B1(n4868), .B2(n6601), .A(n4621), .ZN(n4622) );
  OAI211_X1 U5775 ( .C1(n5096), .C2(n6604), .A(n4623), .B(n4622), .ZN(U3142)
         );
  NAND2_X1 U5776 ( .A1(n4548), .A2(n4625), .ZN(n4626) );
  NAND2_X1 U5777 ( .A1(n4624), .A2(n4626), .ZN(n5497) );
  INV_X1 U5778 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6260) );
  OAI222_X1 U5779 ( .A1(n5497), .A2(n5591), .B1(n5180), .B2(n6303), .C1(n5213), 
        .C2(n6260), .ZN(U2887) );
  NAND2_X1 U5780 ( .A1(n6021), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6513) );
  NOR2_X1 U5781 ( .A1(n4695), .A2(n6513), .ZN(n6027) );
  NOR2_X1 U5782 ( .A1(n6027), .A2(n6578), .ZN(n4633) );
  NAND2_X1 U5783 ( .A1(n4806), .A2(n6581), .ZN(n4804) );
  OR2_X1 U5784 ( .A1(n4804), .A2(n6515), .ZN(n4628) );
  AND2_X1 U5785 ( .A1(n4628), .A2(n4655), .ZN(n4632) );
  INV_X1 U5786 ( .A(n4632), .ZN(n4629) );
  OAI22_X1 U5787 ( .A1(n6474), .A2(n6592), .B1(n4655), .B2(n6511), .ZN(n4631)
         );
  AOI21_X1 U5788 ( .B1(n6589), .B2(n6479), .A(n4631), .ZN(n4636) );
  NAND2_X1 U5789 ( .A1(n4633), .A2(n4632), .ZN(n4634) );
  NAND2_X1 U5790 ( .A1(n4657), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4635) );
  OAI211_X1 U5791 ( .C1(n4660), .C2(n5004), .A(n4636), .B(n4635), .ZN(U3076)
         );
  OAI22_X1 U5792 ( .A1(n6474), .A2(n6622), .B1(n4655), .B2(n6549), .ZN(n4637)
         );
  AOI21_X1 U5793 ( .B1(n6619), .B2(n6479), .A(n4637), .ZN(n4639) );
  NAND2_X1 U5794 ( .A1(n4657), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4638) );
  OAI211_X1 U5795 ( .C1(n4660), .C2(n4905), .A(n4639), .B(n4638), .ZN(U3081)
         );
  OAI22_X1 U5796 ( .A1(n6474), .A2(n6604), .B1(n4655), .B2(n6534), .ZN(n4640)
         );
  AOI21_X1 U5797 ( .B1(n6601), .B2(n6479), .A(n4640), .ZN(n4642) );
  NAND2_X1 U5798 ( .A1(n4657), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4641) );
  OAI211_X1 U5799 ( .C1(n4660), .C2(n4913), .A(n4642), .B(n4641), .ZN(U3078)
         );
  OAI22_X1 U5800 ( .A1(n6474), .A2(n6639), .B1(n4655), .B2(n6560), .ZN(n4643)
         );
  AOI21_X1 U5801 ( .B1(n6634), .B2(n6479), .A(n4643), .ZN(n4645) );
  NAND2_X1 U5802 ( .A1(n4657), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4644) );
  OAI211_X1 U5803 ( .C1(n4660), .C2(n4897), .A(n4645), .B(n4644), .ZN(U3083)
         );
  INV_X1 U5804 ( .A(n6558), .ZN(n6625) );
  OAI22_X1 U5805 ( .A1(n6474), .A2(n6628), .B1(n4655), .B2(n6554), .ZN(n4646)
         );
  AOI21_X1 U5806 ( .B1(n6625), .B2(n6479), .A(n4646), .ZN(n4648) );
  NAND2_X1 U5807 ( .A1(n4657), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4647) );
  OAI211_X1 U5808 ( .C1(n4660), .C2(n4893), .A(n4648), .B(n4647), .ZN(U3082)
         );
  OAI22_X1 U5809 ( .A1(n6474), .A2(n6610), .B1(n4655), .B2(n6539), .ZN(n4649)
         );
  AOI21_X1 U5810 ( .B1(n6607), .B2(n6479), .A(n4649), .ZN(n4651) );
  NAND2_X1 U5811 ( .A1(n4657), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4650) );
  OAI211_X1 U5812 ( .C1(n4660), .C2(n4901), .A(n4651), .B(n4650), .ZN(U3079)
         );
  OAI22_X1 U5813 ( .A1(n6474), .A2(n6616), .B1(n4655), .B2(n6544), .ZN(n4652)
         );
  AOI21_X1 U5814 ( .B1(n6613), .B2(n6479), .A(n4652), .ZN(n4654) );
  NAND2_X1 U5815 ( .A1(n4657), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4653) );
  OAI211_X1 U5816 ( .C1(n4660), .C2(n4909), .A(n4654), .B(n4653), .ZN(U3080)
         );
  OAI22_X1 U5817 ( .A1(n6474), .A2(n6598), .B1(n4655), .B2(n6529), .ZN(n4656)
         );
  AOI21_X1 U5818 ( .B1(n6595), .B2(n6479), .A(n4656), .ZN(n4659) );
  NAND2_X1 U5819 ( .A1(n4657), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4658) );
  OAI211_X1 U5820 ( .C1(n4660), .C2(n4917), .A(n4659), .B(n4658), .ZN(U3077)
         );
  XNOR2_X1 U5821 ( .A(n4662), .B(n4661), .ZN(n5074) );
  INV_X1 U5822 ( .A(n4840), .ZN(n6373) );
  AOI22_X1 U5823 ( .A1(n5995), .A2(n6373), .B1(n6372), .B2(n4663), .ZN(n6378)
         );
  NAND2_X1 U5824 ( .A1(n4664), .A2(n4665), .ZN(n6370) );
  NAND2_X1 U5825 ( .A1(n6378), .A2(n6370), .ZN(n4692) );
  AOI21_X1 U5826 ( .B1(n4840), .B2(n6367), .A(n4664), .ZN(n5058) );
  NOR2_X1 U5827 ( .A1(n4665), .A2(n5058), .ZN(n5998) );
  AOI22_X1 U5828 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4692), .B1(n5998), 
        .B2(n4666), .ZN(n4671) );
  OAI21_X1 U5829 ( .B1(n4667), .B2(n4669), .A(n4668), .ZN(n4875) );
  INV_X1 U5830 ( .A(n4875), .ZN(n6198) );
  INV_X1 U5831 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6792) );
  NOR2_X1 U5832 ( .A1(n3820), .A2(n6792), .ZN(n5070) );
  AOI21_X1 U5833 ( .B1(n6359), .B2(n6198), .A(n5070), .ZN(n4670) );
  OAI211_X1 U5834 ( .C1(n5074), .C2(n6015), .A(n4671), .B(n4670), .ZN(U3015)
         );
  INV_X1 U5835 ( .A(n6021), .ZN(n4672) );
  NAND3_X1 U5836 ( .A1(n5100), .A2(n6437), .A3(n5096), .ZN(n4675) );
  INV_X1 U5837 ( .A(n6582), .ZN(n6033) );
  AOI22_X1 U5838 ( .A1(n4675), .A2(n6033), .B1(n4806), .B2(n4674), .ZN(n4678)
         );
  AND2_X1 U5839 ( .A1(n4676), .A2(n6574), .ZN(n5098) );
  NOR2_X1 U5840 ( .A1(n4679), .A2(n5165), .ZN(n6584) );
  INV_X1 U5841 ( .A(n6584), .ZN(n6055) );
  NAND2_X1 U5842 ( .A1(n6433), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6056) );
  AOI21_X1 U5843 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6056), .A(n6018), .ZN(
        n6049) );
  OAI211_X1 U5844 ( .C1(n5098), .C2(n6050), .A(n6055), .B(n6049), .ZN(n4677)
         );
  INV_X1 U5845 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4686) );
  AND2_X1 U5846 ( .A1(n4581), .A2(n6437), .ZN(n6475) );
  NAND2_X1 U5847 ( .A1(n6475), .A2(n4806), .ZN(n4681) );
  NAND2_X1 U5848 ( .A1(n4679), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6568) );
  OR2_X1 U5849 ( .A1(n6568), .A2(n6056), .ZN(n4680) );
  NAND2_X1 U5850 ( .A1(n4681), .A2(n4680), .ZN(n5097) );
  NOR2_X1 U5851 ( .A1(n5096), .A2(n6558), .ZN(n4684) );
  INV_X1 U5852 ( .A(n5098), .ZN(n4682) );
  OAI22_X1 U5853 ( .A1(n5100), .A2(n6628), .B1(n6554), .B2(n4682), .ZN(n4683)
         );
  AOI211_X1 U5854 ( .C1(n6624), .C2(n5097), .A(n4684), .B(n4683), .ZN(n4685)
         );
  OAI21_X1 U5855 ( .B1(n5075), .B2(n4686), .A(n4685), .ZN(U3138) );
  XNOR2_X1 U5856 ( .A(n4688), .B(n4687), .ZN(n5068) );
  OAI211_X1 U5857 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n5998), .B(n4844), .ZN(n4694) );
  INV_X1 U5858 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6658) );
  NOR2_X1 U5859 ( .A1(n3820), .A2(n6658), .ZN(n4691) );
  OAI21_X1 U5860 ( .B1(n3119), .B2(n3143), .A(n4689), .ZN(n5487) );
  NOR2_X1 U5861 ( .A1(n6387), .A2(n5487), .ZN(n4690) );
  AOI211_X1 U5862 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n4692), .A(n4691), 
        .B(n4690), .ZN(n4693) );
  OAI211_X1 U5863 ( .C1(n6015), .C2(n5068), .A(n4694), .B(n4693), .ZN(U3014)
         );
  AOI21_X1 U5864 ( .B1(n4700), .B2(STATEBS16_REG_SCAN_IN), .A(n6578), .ZN(
        n4703) );
  INV_X1 U5865 ( .A(n4583), .ZN(n6218) );
  NAND2_X1 U5866 ( .A1(n4950), .A2(n6581), .ZN(n6438) );
  INV_X1 U5867 ( .A(n6438), .ZN(n4698) );
  NOR2_X1 U5868 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4696) );
  AND2_X1 U5869 ( .A1(n4696), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6434)
         );
  NAND2_X1 U5870 ( .A1(n6434), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4725) );
  INV_X1 U5871 ( .A(n4725), .ZN(n4697) );
  AOI21_X1 U5872 ( .B1(n4698), .B2(n5498), .A(n4697), .ZN(n4702) );
  INV_X1 U5873 ( .A(n4702), .ZN(n4699) );
  INV_X1 U5874 ( .A(n6592), .ZN(n6470) );
  NAND2_X1 U5875 ( .A1(n4700), .A2(n4587), .ZN(n6436) );
  OAI22_X1 U5876 ( .A1(n6468), .A2(n6528), .B1(n6511), .B2(n4725), .ZN(n4701)
         );
  AOI21_X1 U5877 ( .B1(n6470), .B2(n6460), .A(n4701), .ZN(n4706) );
  NAND2_X1 U5878 ( .A1(n4703), .A2(n4702), .ZN(n4704) );
  NAND2_X1 U5879 ( .A1(n4727), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4705) );
  OAI211_X1 U5880 ( .C1(n4730), .C2(n5004), .A(n4706), .B(n4705), .ZN(U3060)
         );
  INV_X1 U5881 ( .A(n6610), .ZN(n6072) );
  OAI22_X1 U5882 ( .A1(n6468), .A2(n6540), .B1(n6539), .B2(n4725), .ZN(n4707)
         );
  AOI21_X1 U5883 ( .B1(n6072), .B2(n6460), .A(n4707), .ZN(n4709) );
  NAND2_X1 U5884 ( .A1(n4727), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4708) );
  OAI211_X1 U5885 ( .C1(n4730), .C2(n4901), .A(n4709), .B(n4708), .ZN(U3063)
         );
  INV_X1 U5886 ( .A(n6604), .ZN(n6067) );
  OAI22_X1 U5887 ( .A1(n6468), .A2(n6535), .B1(n6534), .B2(n4725), .ZN(n4710)
         );
  AOI21_X1 U5888 ( .B1(n6067), .B2(n6460), .A(n4710), .ZN(n4712) );
  NAND2_X1 U5889 ( .A1(n4727), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4711) );
  OAI211_X1 U5890 ( .C1(n4730), .C2(n4913), .A(n4712), .B(n4711), .ZN(U3062)
         );
  INV_X1 U5891 ( .A(n6639), .ZN(n5140) );
  OAI22_X1 U5892 ( .A1(n6468), .A2(n6561), .B1(n6560), .B2(n4725), .ZN(n4713)
         );
  AOI21_X1 U5893 ( .B1(n5140), .B2(n6460), .A(n4713), .ZN(n4715) );
  NAND2_X1 U5894 ( .A1(n4727), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4714) );
  OAI211_X1 U5895 ( .C1(n4730), .C2(n4897), .A(n4715), .B(n4714), .ZN(U3067)
         );
  INV_X1 U5896 ( .A(n6598), .ZN(n6062) );
  OAI22_X1 U5897 ( .A1(n6468), .A2(n6530), .B1(n6529), .B2(n4725), .ZN(n4716)
         );
  AOI21_X1 U5898 ( .B1(n6062), .B2(n6460), .A(n4716), .ZN(n4718) );
  NAND2_X1 U5899 ( .A1(n4727), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4717) );
  OAI211_X1 U5900 ( .C1(n4730), .C2(n4917), .A(n4718), .B(n4717), .ZN(U3061)
         );
  INV_X1 U5901 ( .A(n6616), .ZN(n6077) );
  OAI22_X1 U5902 ( .A1(n6468), .A2(n6545), .B1(n6544), .B2(n4725), .ZN(n4719)
         );
  AOI21_X1 U5903 ( .B1(n6077), .B2(n6460), .A(n4719), .ZN(n4721) );
  NAND2_X1 U5904 ( .A1(n4727), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4720) );
  OAI211_X1 U5905 ( .C1(n4730), .C2(n4909), .A(n4721), .B(n4720), .ZN(U3064)
         );
  INV_X1 U5906 ( .A(n6622), .ZN(n6082) );
  OAI22_X1 U5907 ( .A1(n6468), .A2(n6553), .B1(n6549), .B2(n4725), .ZN(n4722)
         );
  AOI21_X1 U5908 ( .B1(n6082), .B2(n6460), .A(n4722), .ZN(n4724) );
  NAND2_X1 U5909 ( .A1(n4727), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4723) );
  OAI211_X1 U5910 ( .C1(n4730), .C2(n4905), .A(n4724), .B(n4723), .ZN(U3065)
         );
  OAI22_X1 U5911 ( .A1(n6468), .A2(n6558), .B1(n6554), .B2(n4725), .ZN(n4726)
         );
  AOI21_X1 U5912 ( .B1(n4976), .B2(n6460), .A(n4726), .ZN(n4729) );
  NAND2_X1 U5913 ( .A1(n4727), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4728) );
  OAI211_X1 U5914 ( .C1(n4730), .C2(n4893), .A(n4729), .B(n4728), .ZN(U3066)
         );
  OAI21_X1 U5915 ( .B1(n4731), .B2(n4732), .A(n4734), .ZN(n5157) );
  INV_X1 U5916 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6265) );
  OAI222_X1 U5917 ( .A1(n5157), .A2(n5591), .B1(n5180), .B2(n6297), .C1(n5213), 
        .C2(n6265), .ZN(U2890) );
  AOI22_X1 U5918 ( .A1(n6576), .A2(n5098), .B1(n5097), .B2(n6577), .ZN(n4735)
         );
  OAI21_X1 U5919 ( .B1(n5100), .B2(n6592), .A(n4735), .ZN(n4736) );
  AOI21_X1 U5920 ( .B1(n6589), .B2(n4737), .A(n4736), .ZN(n4738) );
  OAI21_X1 U5921 ( .B1(n5075), .B2(n4739), .A(n4738), .ZN(U3132) );
  NAND2_X1 U5922 ( .A1(n4581), .A2(n4763), .ZN(n4756) );
  INV_X1 U5923 ( .A(n4740), .ZN(n4754) );
  MUX2_X1 U5924 ( .A(n4741), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4502), 
        .Z(n4743) );
  NOR2_X1 U5925 ( .A1(n4743), .A2(n4742), .ZN(n4753) );
  XNOR2_X1 U5926 ( .A(n4744), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4751)
         );
  INV_X1 U5927 ( .A(n4745), .ZN(n4746) );
  OAI21_X1 U5928 ( .B1(n4502), .B2(n4747), .A(n4746), .ZN(n4749) );
  NOR2_X1 U5929 ( .A1(n4749), .A2(n4748), .ZN(n6037) );
  OAI22_X1 U5930 ( .A1(n4761), .A2(n4751), .B1(n6037), .B2(n4750), .ZN(n4752)
         );
  AOI21_X1 U5931 ( .B1(n4754), .B2(n4753), .A(n4752), .ZN(n4755) );
  NAND2_X1 U5932 ( .A1(n4756), .A2(n4755), .ZN(n6035) );
  MUX2_X1 U5933 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6035), .S(n4782), 
        .Z(n4777) );
  INV_X1 U5934 ( .A(n4777), .ZN(n4775) );
  NOR3_X1 U5935 ( .A1(n4758), .A2(n4757), .A3(n6574), .ZN(n4764) );
  OR3_X1 U5936 ( .A1(n4759), .A2(n4502), .A3(n3163), .ZN(n4760) );
  OAI21_X1 U5937 ( .B1(n4761), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4760), 
        .ZN(n4762) );
  AOI21_X1 U5938 ( .B1(n6218), .B2(n4763), .A(n4762), .ZN(n5192) );
  AOI21_X1 U5939 ( .B1(n4764), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n5192), 
        .ZN(n4766) );
  INV_X1 U5940 ( .A(n4764), .ZN(n4765) );
  AOI22_X1 U5941 ( .A1(n4766), .A2(n4782), .B1(n4948), .B2(n4765), .ZN(n4772)
         );
  MUX2_X1 U5942 ( .A(n4768), .B(n4767), .S(n4782), .Z(n4770) );
  INV_X1 U5943 ( .A(n4770), .ZN(n4776) );
  NAND2_X1 U5944 ( .A1(n4776), .A2(n4769), .ZN(n4771) );
  AOI22_X1 U5945 ( .A1(n4772), .A2(n4771), .B1(n4770), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4773) );
  AOI21_X1 U5946 ( .B1(n4777), .B2(n6519), .A(n4773), .ZN(n4774) );
  AOI211_X1 U5947 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n4775), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n4774), .ZN(n4793) );
  INV_X1 U5948 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6102) );
  NAND2_X1 U5949 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6102), .ZN(n4783) );
  INV_X1 U5950 ( .A(n4742), .ZN(n4779) );
  NAND3_X1 U5951 ( .A1(n4777), .A2(n4776), .A3(n4786), .ZN(n4778) );
  OAI21_X1 U5952 ( .B1(n4783), .B2(n4779), .A(n4778), .ZN(n5198) );
  NAND2_X1 U5953 ( .A1(n5491), .A2(n4780), .ZN(n4781) );
  OAI21_X1 U5954 ( .B1(n4782), .B2(n4784), .A(n4781), .ZN(n4787) );
  NOR2_X1 U5955 ( .A1(n4784), .A2(n4783), .ZN(n4785) );
  AOI21_X1 U5956 ( .B1(n4787), .B2(n4786), .A(n4785), .ZN(n5199) );
  OAI21_X1 U5957 ( .B1(MORE_REG_SCAN_IN), .B2(FLUSH_REG_SCAN_IN), .A(n4788), 
        .ZN(n4789) );
  NAND4_X1 U5958 ( .A1(n5199), .A2(n4791), .A3(n4790), .A4(n4789), .ZN(n4792)
         );
  NOR3_X1 U5959 ( .A1(n4793), .A2(n5198), .A3(n4792), .ZN(n5205) );
  AOI21_X1 U5960 ( .B1(n5205), .B2(STATE2_REG_0__SCAN_IN), .A(
        STATE2_REG_1__SCAN_IN), .ZN(n4799) );
  NAND3_X1 U5961 ( .A1(n6722), .A2(STATE2_REG_2__SCAN_IN), .A3(READY_N), .ZN(
        n4794) );
  NAND2_X1 U5962 ( .A1(n4795), .A2(n4794), .ZN(n4796) );
  OAI21_X1 U5963 ( .B1(n4798), .B2(n4797), .A(n4796), .ZN(n5168) );
  OAI21_X1 U5964 ( .B1(n5201), .B2(n6722), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4800) );
  INV_X1 U5965 ( .A(n6643), .ZN(n5212) );
  NAND2_X1 U5966 ( .A1(n4800), .A2(n5212), .ZN(U3453) );
  NAND3_X1 U5967 ( .A1(n6468), .A2(n6437), .A3(n6474), .ZN(n4801) );
  NAND2_X1 U5968 ( .A1(n4801), .A2(n6033), .ZN(n4805) );
  AND2_X1 U5969 ( .A1(n4802), .A2(n6574), .ZN(n6466) );
  NAND2_X1 U5970 ( .A1(n6433), .A2(n6519), .ZN(n5117) );
  AOI21_X1 U5971 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5117), .A(n6018), .ZN(
        n5114) );
  OAI211_X1 U5972 ( .C1(n6466), .C2(n6050), .A(n6055), .B(n5114), .ZN(n4803)
         );
  INV_X1 U5973 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4812) );
  INV_X1 U5974 ( .A(n4581), .ZN(n6482) );
  NAND3_X1 U5975 ( .A1(n6482), .A2(n6437), .A3(n4806), .ZN(n4808) );
  OR2_X1 U5976 ( .A1(n6568), .A2(n5117), .ZN(n4807) );
  NAND2_X1 U5977 ( .A1(n4808), .A2(n4807), .ZN(n6465) );
  AOI22_X1 U5978 ( .A1(n6611), .A2(n6466), .B1(n6465), .B2(n6612), .ZN(n4809)
         );
  OAI21_X1 U5979 ( .B1(n6468), .B2(n6616), .A(n4809), .ZN(n4810) );
  AOI21_X1 U5980 ( .B1(n6613), .B2(n4834), .A(n4810), .ZN(n4811) );
  OAI21_X1 U5981 ( .B1(n6467), .B2(n4812), .A(n4811), .ZN(U3072) );
  INV_X1 U5982 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4817) );
  NOR2_X1 U5983 ( .A1(n6474), .A2(n6558), .ZN(n4815) );
  INV_X1 U5984 ( .A(n6466), .ZN(n4813) );
  OAI22_X1 U5985 ( .A1(n6468), .A2(n6628), .B1(n6554), .B2(n4813), .ZN(n4814)
         );
  AOI211_X1 U5986 ( .C1(n6624), .C2(n6465), .A(n4815), .B(n4814), .ZN(n4816)
         );
  OAI21_X1 U5987 ( .B1(n6467), .B2(n4817), .A(n4816), .ZN(U3074) );
  AOI22_X1 U5988 ( .A1(n6617), .A2(n6466), .B1(n6465), .B2(n6618), .ZN(n4818)
         );
  OAI21_X1 U5989 ( .B1(n6468), .B2(n6622), .A(n4818), .ZN(n4819) );
  AOI21_X1 U5990 ( .B1(n6619), .B2(n4834), .A(n4819), .ZN(n4820) );
  OAI21_X1 U5991 ( .B1(n6467), .B2(n6855), .A(n4820), .ZN(U3073) );
  INV_X1 U5992 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4824) );
  AOI22_X1 U5993 ( .A1(n6593), .A2(n6466), .B1(n6465), .B2(n6594), .ZN(n4821)
         );
  OAI21_X1 U5994 ( .B1(n6468), .B2(n6598), .A(n4821), .ZN(n4822) );
  AOI21_X1 U5995 ( .B1(n6595), .B2(n4834), .A(n4822), .ZN(n4823) );
  OAI21_X1 U5996 ( .B1(n6467), .B2(n4824), .A(n4823), .ZN(U3069) );
  AOI22_X1 U5997 ( .A1(n6599), .A2(n6466), .B1(n6465), .B2(n6600), .ZN(n4825)
         );
  OAI21_X1 U5998 ( .B1(n6468), .B2(n6604), .A(n4825), .ZN(n4826) );
  AOI21_X1 U5999 ( .B1(n6601), .B2(n4834), .A(n4826), .ZN(n4827) );
  OAI21_X1 U6000 ( .B1(n6467), .B2(n6739), .A(n4827), .ZN(U3070) );
  INV_X1 U6001 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4831) );
  AOI22_X1 U6002 ( .A1(n6605), .A2(n6466), .B1(n6465), .B2(n6606), .ZN(n4828)
         );
  OAI21_X1 U6003 ( .B1(n6468), .B2(n6610), .A(n4828), .ZN(n4829) );
  AOI21_X1 U6004 ( .B1(n6607), .B2(n4834), .A(n4829), .ZN(n4830) );
  OAI21_X1 U6005 ( .B1(n6467), .B2(n4831), .A(n4830), .ZN(U3071) );
  INV_X1 U6006 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U6007 ( .A1(n6630), .A2(n6466), .B1(n6465), .B2(n6631), .ZN(n4832)
         );
  OAI21_X1 U6008 ( .B1(n6468), .B2(n6639), .A(n4832), .ZN(n4833) );
  AOI21_X1 U6009 ( .B1(n6634), .B2(n4834), .A(n4833), .ZN(n4835) );
  OAI21_X1 U6010 ( .B1(n6467), .B2(n4836), .A(n4835), .ZN(U3075) );
  XNOR2_X1 U6011 ( .A(n4838), .B(n4837), .ZN(n5110) );
  OAI21_X1 U6012 ( .B1(n4842), .B2(n3024), .A(n5936), .ZN(n4839) );
  NAND2_X1 U6013 ( .A1(n6378), .A2(n4839), .ZN(n5062) );
  NAND2_X1 U6014 ( .A1(n4840), .A2(n6367), .ZN(n4843) );
  OAI211_X1 U6015 ( .C1(n4844), .C2(n4843), .A(n4842), .B(n4841), .ZN(n4845)
         );
  NAND2_X1 U6016 ( .A1(n5062), .A2(n4845), .ZN(n4849) );
  INV_X1 U6017 ( .A(n4996), .ZN(n4846) );
  AOI21_X1 U6018 ( .B1(n4847), .B2(n4689), .A(n4846), .ZN(n6189) );
  INV_X1 U6019 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6660) );
  NOR2_X1 U6020 ( .A1(n3820), .A2(n6660), .ZN(n5106) );
  AOI21_X1 U6021 ( .B1(n6359), .B2(n6189), .A(n5106), .ZN(n4848) );
  OAI211_X1 U6022 ( .C1(n5110), .C2(n6015), .A(n4849), .B(n4848), .ZN(U3013)
         );
  AND2_X1 U6023 ( .A1(n4624), .A2(n4852), .ZN(n4853) );
  OR2_X1 U6024 ( .A1(n4851), .A2(n4853), .ZN(n5105) );
  INV_X1 U6025 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6258) );
  OAI222_X1 U6026 ( .A1(n5105), .A2(n5591), .B1(n5180), .B2(n6305), .C1(n5213), 
        .C2(n6258), .ZN(U2886) );
  INV_X1 U6027 ( .A(n4667), .ZN(n4854) );
  OAI21_X1 U6028 ( .B1(n4856), .B2(n4855), .A(n4854), .ZN(n6371) );
  INV_X1 U6029 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4857) );
  OAI222_X1 U6030 ( .A1(n6371), .A2(n5557), .B1(n4857), .B2(n5552), .C1(n5544), 
        .C2(n6330), .ZN(U2857) );
  INV_X1 U6031 ( .A(EBX_REG_4__SCAN_IN), .ZN(n5488) );
  OAI222_X1 U6032 ( .A1(n5487), .A2(n5557), .B1(n5552), .B2(n5488), .C1(n5544), 
        .C2(n5497), .ZN(U2855) );
  INV_X1 U6033 ( .A(n6024), .ZN(n4859) );
  OAI21_X1 U6034 ( .B1(n5015), .B2(n6578), .A(n6033), .ZN(n5010) );
  NAND2_X1 U6035 ( .A1(n4503), .A2(n4583), .ZN(n6481) );
  OAI211_X1 U6036 ( .C1(n6582), .C2(n4941), .A(n5010), .B(n5006), .ZN(n4862)
         );
  INV_X1 U6037 ( .A(n6433), .ZN(n6569) );
  INV_X1 U6038 ( .A(n6018), .ZN(n4860) );
  OAI21_X1 U6039 ( .B1(n5165), .B2(n6569), .A(n4860), .ZN(n6483) );
  AOI21_X1 U6040 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6476), .A(n6483), .ZN(
        n6441) );
  NOR2_X1 U6041 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U6042 ( .A1(n4881), .A2(n6519), .ZN(n5011) );
  OR2_X1 U6043 ( .A1(n5011), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4919)
         );
  NAND2_X1 U6044 ( .A1(n4919), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4861) );
  NAND4_X1 U6045 ( .A1(n4862), .A2(n6441), .A3(n6568), .A4(n4861), .ZN(n4918)
         );
  NAND2_X1 U6046 ( .A1(n4918), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4865) );
  NAND2_X1 U6047 ( .A1(n6584), .A2(n6569), .ZN(n6477) );
  OAI22_X1 U6048 ( .A1(n5006), .A2(n6578), .B1(n6476), .B2(n6477), .ZN(n4939)
         );
  OAI22_X1 U6049 ( .A1(n4941), .A2(n6628), .B1(n6554), .B2(n4919), .ZN(n4863)
         );
  AOI21_X1 U6050 ( .B1(n6624), .B2(n4939), .A(n4863), .ZN(n4864) );
  OAI211_X1 U6051 ( .C1(n5045), .C2(n6558), .A(n4865), .B(n4864), .ZN(U3026)
         );
  NAND2_X1 U6052 ( .A1(n4918), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4870) );
  INV_X1 U6053 ( .A(n4939), .ZN(n4866) );
  OAI22_X1 U6054 ( .A1(n4866), .A2(n5004), .B1(n6511), .B2(n4919), .ZN(n4867)
         );
  AOI21_X1 U6055 ( .B1(n4868), .B2(n6470), .A(n4867), .ZN(n4869) );
  OAI211_X1 U6056 ( .C1(n5045), .C2(n6528), .A(n4870), .B(n4869), .ZN(U3020)
         );
  OAI21_X1 U6057 ( .B1(n4872), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4871), 
        .ZN(n6386) );
  INV_X1 U6058 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4873) );
  OAI222_X1 U6059 ( .A1(n6386), .A2(n5557), .B1(n5552), .B2(n4873), .C1(n5503), 
        .C2(n5544), .ZN(U2859) );
  INV_X1 U6060 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4874) );
  OAI222_X1 U6061 ( .A1(n4875), .A2(n5557), .B1(n4874), .B2(n5552), .C1(n5069), 
        .C2(n5544), .ZN(U2856) );
  OAI21_X1 U6062 ( .B1(n4851), .B2(n4876), .A(n4878), .ZN(n5173) );
  AOI22_X1 U6063 ( .A1(n5613), .A2(DATAI_6_), .B1(n5612), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n4879) );
  OAI21_X1 U6064 ( .B1(n5173), .B2(n5591), .A(n4879), .ZN(U2885) );
  INV_X1 U6065 ( .A(n4885), .ZN(n4880) );
  OAI21_X1 U6066 ( .B1(n4880), .B2(n6578), .A(n6033), .ZN(n4888) );
  INV_X1 U6067 ( .A(n6481), .ZN(n4883) );
  NAND2_X1 U6068 ( .A1(n4881), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6478) );
  OR2_X1 U6069 ( .A1(n6478), .A2(n6574), .ZN(n4999) );
  INV_X1 U6070 ( .A(n4999), .ZN(n4882) );
  AOI21_X1 U6071 ( .B1(n4951), .B2(n4883), .A(n4882), .ZN(n4887) );
  INV_X1 U6072 ( .A(n4887), .ZN(n4884) );
  INV_X1 U6073 ( .A(n6478), .ZN(n4890) );
  OAI22_X1 U6074 ( .A1(n6091), .A2(n6558), .B1(n6554), .B2(n4999), .ZN(n4886)
         );
  AOI21_X1 U6075 ( .B1(n4976), .B2(n6503), .A(n4886), .ZN(n4892) );
  NAND2_X1 U6076 ( .A1(n4888), .A2(n4887), .ZN(n4889) );
  NAND2_X1 U6077 ( .A1(n5001), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4891) );
  OAI211_X1 U6078 ( .C1(n5005), .C2(n4893), .A(n4892), .B(n4891), .ZN(U3098)
         );
  OAI22_X1 U6079 ( .A1(n6091), .A2(n6561), .B1(n6560), .B2(n4999), .ZN(n4894)
         );
  AOI21_X1 U6080 ( .B1(n5140), .B2(n6503), .A(n4894), .ZN(n4896) );
  NAND2_X1 U6081 ( .A1(n5001), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4895) );
  OAI211_X1 U6082 ( .C1(n5005), .C2(n4897), .A(n4896), .B(n4895), .ZN(U3099)
         );
  OAI22_X1 U6083 ( .A1(n6091), .A2(n6540), .B1(n6539), .B2(n4999), .ZN(n4898)
         );
  AOI21_X1 U6084 ( .B1(n6072), .B2(n6503), .A(n4898), .ZN(n4900) );
  NAND2_X1 U6085 ( .A1(n5001), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4899) );
  OAI211_X1 U6086 ( .C1(n5005), .C2(n4901), .A(n4900), .B(n4899), .ZN(U3095)
         );
  OAI22_X1 U6087 ( .A1(n6091), .A2(n6553), .B1(n6549), .B2(n4999), .ZN(n4902)
         );
  AOI21_X1 U6088 ( .B1(n6082), .B2(n6503), .A(n4902), .ZN(n4904) );
  NAND2_X1 U6089 ( .A1(n5001), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4903) );
  OAI211_X1 U6090 ( .C1(n5005), .C2(n4905), .A(n4904), .B(n4903), .ZN(U3097)
         );
  OAI22_X1 U6091 ( .A1(n6091), .A2(n6545), .B1(n6544), .B2(n4999), .ZN(n4906)
         );
  AOI21_X1 U6092 ( .B1(n6077), .B2(n6503), .A(n4906), .ZN(n4908) );
  NAND2_X1 U6093 ( .A1(n5001), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4907) );
  OAI211_X1 U6094 ( .C1(n5005), .C2(n4909), .A(n4908), .B(n4907), .ZN(U3096)
         );
  OAI22_X1 U6095 ( .A1(n6091), .A2(n6535), .B1(n6534), .B2(n4999), .ZN(n4910)
         );
  AOI21_X1 U6096 ( .B1(n6067), .B2(n6503), .A(n4910), .ZN(n4912) );
  NAND2_X1 U6097 ( .A1(n5001), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4911) );
  OAI211_X1 U6098 ( .C1(n5005), .C2(n4913), .A(n4912), .B(n4911), .ZN(U3094)
         );
  OAI22_X1 U6099 ( .A1(n6091), .A2(n6530), .B1(n6529), .B2(n4999), .ZN(n4914)
         );
  AOI21_X1 U6100 ( .B1(n6062), .B2(n6503), .A(n4914), .ZN(n4916) );
  NAND2_X1 U6101 ( .A1(n5001), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4915) );
  OAI211_X1 U6102 ( .C1(n5005), .C2(n4917), .A(n4916), .B(n4915), .ZN(U3093)
         );
  INV_X1 U6103 ( .A(n4919), .ZN(n4938) );
  AOI22_X1 U6104 ( .A1(n6612), .A2(n4939), .B1(n6611), .B2(n4938), .ZN(n4920)
         );
  OAI21_X1 U6105 ( .B1(n4941), .B2(n6616), .A(n4920), .ZN(n4921) );
  AOI21_X1 U6106 ( .B1(n4943), .B2(n6613), .A(n4921), .ZN(n4922) );
  OAI21_X1 U6107 ( .B1(n4946), .B2(n4923), .A(n4922), .ZN(U3024) );
  AOI22_X1 U6108 ( .A1(n6594), .A2(n4939), .B1(n6593), .B2(n4938), .ZN(n4924)
         );
  OAI21_X1 U6109 ( .B1(n4941), .B2(n6598), .A(n4924), .ZN(n4925) );
  AOI21_X1 U6110 ( .B1(n4943), .B2(n6595), .A(n4925), .ZN(n4926) );
  OAI21_X1 U6111 ( .B1(n4946), .B2(n6825), .A(n4926), .ZN(U3021) );
  AOI22_X1 U6112 ( .A1(n6600), .A2(n4939), .B1(n6599), .B2(n4938), .ZN(n4927)
         );
  OAI21_X1 U6113 ( .B1(n4941), .B2(n6604), .A(n4927), .ZN(n4928) );
  AOI21_X1 U6114 ( .B1(n4943), .B2(n6601), .A(n4928), .ZN(n4929) );
  OAI21_X1 U6115 ( .B1(n4946), .B2(n4930), .A(n4929), .ZN(U3022) );
  AOI22_X1 U6116 ( .A1(n6606), .A2(n4939), .B1(n6605), .B2(n4938), .ZN(n4931)
         );
  OAI21_X1 U6117 ( .B1(n4941), .B2(n6610), .A(n4931), .ZN(n4932) );
  AOI21_X1 U6118 ( .B1(n4943), .B2(n6607), .A(n4932), .ZN(n4933) );
  OAI21_X1 U6119 ( .B1(n4946), .B2(n4254), .A(n4933), .ZN(U3023) );
  AOI22_X1 U6120 ( .A1(n6631), .A2(n4939), .B1(n6630), .B2(n4938), .ZN(n4934)
         );
  OAI21_X1 U6121 ( .B1(n4941), .B2(n6639), .A(n4934), .ZN(n4935) );
  AOI21_X1 U6122 ( .B1(n4943), .B2(n6634), .A(n4935), .ZN(n4936) );
  OAI21_X1 U6123 ( .B1(n4946), .B2(n4937), .A(n4936), .ZN(U3027) );
  AOI22_X1 U6124 ( .A1(n6618), .A2(n4939), .B1(n6617), .B2(n4938), .ZN(n4940)
         );
  OAI21_X1 U6125 ( .B1(n4941), .B2(n6622), .A(n4940), .ZN(n4942) );
  AOI21_X1 U6126 ( .B1(n4943), .B2(n6619), .A(n4942), .ZN(n4944) );
  OAI21_X1 U6127 ( .B1(n4946), .B2(n4945), .A(n4944), .ZN(U3025) );
  INV_X1 U6128 ( .A(n4953), .ZN(n4947) );
  NOR2_X1 U6129 ( .A1(n4947), .A2(n6435), .ZN(n6029) );
  NOR2_X1 U6130 ( .A1(n6029), .A2(n6578), .ZN(n4956) );
  AND2_X1 U6131 ( .A1(n4949), .A2(n4948), .ZN(n6575) );
  AND2_X1 U6132 ( .A1(n6575), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4954)
         );
  AOI21_X1 U6133 ( .B1(n4951), .B2(n4950), .A(n4954), .ZN(n4958) );
  OAI21_X1 U6134 ( .B1(n6575), .B2(n6437), .A(n6400), .ZN(n4952) );
  INV_X1 U6135 ( .A(n4954), .ZN(n4988) );
  OAI22_X1 U6136 ( .A1(n5100), .A2(n6561), .B1(n6560), .B2(n4988), .ZN(n4955)
         );
  AOI21_X1 U6137 ( .B1(n5140), .B2(n6633), .A(n4955), .ZN(n4961) );
  INV_X1 U6138 ( .A(n4956), .ZN(n4959) );
  INV_X1 U6139 ( .A(n6575), .ZN(n4957) );
  NAND2_X1 U6140 ( .A1(n4990), .A2(n6631), .ZN(n4960) );
  OAI211_X1 U6141 ( .C1(n4994), .C2(n4962), .A(n4961), .B(n4960), .ZN(U3131)
         );
  OAI22_X1 U6142 ( .A1(n5100), .A2(n6553), .B1(n6549), .B2(n4988), .ZN(n4963)
         );
  AOI21_X1 U6143 ( .B1(n6082), .B2(n6633), .A(n4963), .ZN(n4965) );
  NAND2_X1 U6144 ( .A1(n4990), .A2(n6618), .ZN(n4964) );
  OAI211_X1 U6145 ( .C1(n4994), .C2(n4966), .A(n4965), .B(n4964), .ZN(U3129)
         );
  OAI22_X1 U6146 ( .A1(n5100), .A2(n6528), .B1(n6511), .B2(n4988), .ZN(n4967)
         );
  AOI21_X1 U6147 ( .B1(n6470), .B2(n6633), .A(n4967), .ZN(n4969) );
  NAND2_X1 U6148 ( .A1(n4990), .A2(n6577), .ZN(n4968) );
  OAI211_X1 U6149 ( .C1(n4994), .C2(n4970), .A(n4969), .B(n4968), .ZN(U3124)
         );
  OAI22_X1 U6150 ( .A1(n5100), .A2(n6535), .B1(n6534), .B2(n4988), .ZN(n4971)
         );
  AOI21_X1 U6151 ( .B1(n6067), .B2(n6633), .A(n4971), .ZN(n4973) );
  NAND2_X1 U6152 ( .A1(n4990), .A2(n6600), .ZN(n4972) );
  OAI211_X1 U6153 ( .C1(n4994), .C2(n4974), .A(n4973), .B(n4972), .ZN(U3126)
         );
  OAI22_X1 U6154 ( .A1(n5100), .A2(n6558), .B1(n6554), .B2(n4988), .ZN(n4975)
         );
  AOI21_X1 U6155 ( .B1(n4976), .B2(n6633), .A(n4975), .ZN(n4978) );
  NAND2_X1 U6156 ( .A1(n4990), .A2(n6624), .ZN(n4977) );
  OAI211_X1 U6157 ( .C1(n4994), .C2(n4979), .A(n4978), .B(n4977), .ZN(U3130)
         );
  OAI22_X1 U6158 ( .A1(n5100), .A2(n6540), .B1(n6539), .B2(n4988), .ZN(n4980)
         );
  AOI21_X1 U6159 ( .B1(n6072), .B2(n6633), .A(n4980), .ZN(n4982) );
  NAND2_X1 U6160 ( .A1(n4990), .A2(n6606), .ZN(n4981) );
  OAI211_X1 U6161 ( .C1(n4994), .C2(n4983), .A(n4982), .B(n4981), .ZN(U3127)
         );
  OAI22_X1 U6162 ( .A1(n5100), .A2(n6545), .B1(n6544), .B2(n4988), .ZN(n4984)
         );
  AOI21_X1 U6163 ( .B1(n6077), .B2(n6633), .A(n4984), .ZN(n4986) );
  NAND2_X1 U6164 ( .A1(n4990), .A2(n6612), .ZN(n4985) );
  OAI211_X1 U6165 ( .C1(n4994), .C2(n4987), .A(n4986), .B(n4985), .ZN(U3128)
         );
  INV_X1 U6166 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4993) );
  OAI22_X1 U6167 ( .A1(n5100), .A2(n6530), .B1(n6529), .B2(n4988), .ZN(n4989)
         );
  AOI21_X1 U6168 ( .B1(n6062), .B2(n6633), .A(n4989), .ZN(n4992) );
  NAND2_X1 U6169 ( .A1(n4990), .A2(n6594), .ZN(n4991) );
  OAI211_X1 U6170 ( .C1(n4994), .C2(n4993), .A(n4992), .B(n4991), .ZN(U3125)
         );
  INV_X1 U6171 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4998) );
  AND2_X1 U6172 ( .A1(n4996), .A2(n4995), .ZN(n4997) );
  OR2_X1 U6173 ( .A1(n4997), .A2(n5554), .ZN(n6179) );
  OAI222_X1 U6174 ( .A1(n5173), .A2(n5544), .B1(n5552), .B2(n4998), .C1(n5557), 
        .C2(n6179), .ZN(U2853) );
  OAI22_X1 U6175 ( .A1(n6091), .A2(n6528), .B1(n6511), .B2(n4999), .ZN(n5000)
         );
  AOI21_X1 U6176 ( .B1(n6470), .B2(n6503), .A(n5000), .ZN(n5003) );
  NAND2_X1 U6177 ( .A1(n5001), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n5002) );
  OAI211_X1 U6178 ( .C1(n5005), .C2(n5004), .A(n5003), .B(n5002), .ZN(U3092)
         );
  INV_X1 U6179 ( .A(n5006), .ZN(n5007) );
  NOR2_X1 U6180 ( .A1(n5011), .A2(n6574), .ZN(n5043) );
  AOI21_X1 U6181 ( .B1(n5007), .B2(n5498), .A(n5043), .ZN(n5012) );
  INV_X1 U6182 ( .A(n5011), .ZN(n5008) );
  OAI21_X1 U6183 ( .B1(n5008), .B2(n6437), .A(n6400), .ZN(n5009) );
  INV_X1 U6184 ( .A(n5010), .ZN(n5013) );
  OAI22_X1 U6185 ( .A1(n5013), .A2(n5012), .B1(n5165), .B2(n5011), .ZN(n5047)
         );
  NAND2_X1 U6186 ( .A1(n5015), .A2(n5014), .ZN(n5120) );
  INV_X1 U6187 ( .A(n6554), .ZN(n6623) );
  AOI22_X1 U6188 ( .A1(n5154), .A2(n6625), .B1(n6623), .B2(n5043), .ZN(n5016)
         );
  OAI21_X1 U6189 ( .B1(n6628), .B2(n5045), .A(n5016), .ZN(n5017) );
  AOI21_X1 U6190 ( .B1(n5047), .B2(n6624), .A(n5017), .ZN(n5018) );
  OAI21_X1 U6191 ( .B1(n5050), .B2(n6869), .A(n5018), .ZN(U3034) );
  AOI22_X1 U6192 ( .A1(n5154), .A2(n6589), .B1(n6576), .B2(n5043), .ZN(n5019)
         );
  OAI21_X1 U6193 ( .B1(n6592), .B2(n5045), .A(n5019), .ZN(n5020) );
  AOI21_X1 U6194 ( .B1(n5047), .B2(n6577), .A(n5020), .ZN(n5021) );
  OAI21_X1 U6195 ( .B1(n5050), .B2(n5022), .A(n5021), .ZN(U3028) );
  INV_X1 U6196 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5026) );
  AOI22_X1 U6197 ( .A1(n5154), .A2(n6613), .B1(n6611), .B2(n5043), .ZN(n5023)
         );
  OAI21_X1 U6198 ( .B1(n6616), .B2(n5045), .A(n5023), .ZN(n5024) );
  AOI21_X1 U6199 ( .B1(n5047), .B2(n6612), .A(n5024), .ZN(n5025) );
  OAI21_X1 U6200 ( .B1(n5050), .B2(n5026), .A(n5025), .ZN(U3032) );
  AOI22_X1 U6201 ( .A1(n5154), .A2(n6601), .B1(n6599), .B2(n5043), .ZN(n5027)
         );
  OAI21_X1 U6202 ( .B1(n6604), .B2(n5045), .A(n5027), .ZN(n5028) );
  AOI21_X1 U6203 ( .B1(n5047), .B2(n6600), .A(n5028), .ZN(n5029) );
  OAI21_X1 U6204 ( .B1(n5050), .B2(n5030), .A(n5029), .ZN(U3030) );
  AOI22_X1 U6205 ( .A1(n5154), .A2(n6619), .B1(n6617), .B2(n5043), .ZN(n5031)
         );
  OAI21_X1 U6206 ( .B1(n6622), .B2(n5045), .A(n5031), .ZN(n5032) );
  AOI21_X1 U6207 ( .B1(n5047), .B2(n6618), .A(n5032), .ZN(n5033) );
  OAI21_X1 U6208 ( .B1(n5050), .B2(n5034), .A(n5033), .ZN(U3033) );
  INV_X1 U6209 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5038) );
  AOI22_X1 U6210 ( .A1(n5154), .A2(n6634), .B1(n6630), .B2(n5043), .ZN(n5035)
         );
  OAI21_X1 U6211 ( .B1(n6639), .B2(n5045), .A(n5035), .ZN(n5036) );
  AOI21_X1 U6212 ( .B1(n5047), .B2(n6631), .A(n5036), .ZN(n5037) );
  OAI21_X1 U6213 ( .B1(n5050), .B2(n5038), .A(n5037), .ZN(U3035) );
  INV_X1 U6214 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n5042) );
  AOI22_X1 U6215 ( .A1(n5154), .A2(n6595), .B1(n6593), .B2(n5043), .ZN(n5039)
         );
  OAI21_X1 U6216 ( .B1(n6598), .B2(n5045), .A(n5039), .ZN(n5040) );
  AOI21_X1 U6217 ( .B1(n5047), .B2(n6594), .A(n5040), .ZN(n5041) );
  OAI21_X1 U6218 ( .B1(n5050), .B2(n5042), .A(n5041), .ZN(U3029) );
  INV_X1 U6219 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5049) );
  AOI22_X1 U6220 ( .A1(n5154), .A2(n6607), .B1(n6605), .B2(n5043), .ZN(n5044)
         );
  OAI21_X1 U6221 ( .B1(n6610), .B2(n5045), .A(n5044), .ZN(n5046) );
  AOI21_X1 U6222 ( .B1(n5047), .B2(n6606), .A(n5046), .ZN(n5048) );
  OAI21_X1 U6223 ( .B1(n5050), .B2(n5049), .A(n5048), .ZN(U3031) );
  AOI22_X1 U6224 ( .A1(n6232), .A2(n5051), .B1(n5518), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n5052) );
  OAI21_X1 U6225 ( .B1(n5157), .B2(n5544), .A(n5052), .ZN(U2858) );
  AOI22_X1 U6226 ( .A1(n6189), .A2(n6232), .B1(n5518), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n5053) );
  OAI21_X1 U6227 ( .B1(n5105), .B2(n5544), .A(n5053), .ZN(U2854) );
  XNOR2_X1 U6228 ( .A(n5055), .B(n5054), .ZN(n5177) );
  NAND2_X1 U6229 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5056), .ZN(n5057)
         );
  NOR3_X1 U6230 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5058), .A3(n5057), 
        .ZN(n5061) );
  OAI22_X1 U6231 ( .A1(n6387), .A2(n6179), .B1(n5059), .B2(n3820), .ZN(n5060)
         );
  AOI211_X1 U6232 ( .C1(n5062), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n5061), 
        .B(n5060), .ZN(n5063) );
  OAI21_X1 U6233 ( .B1(n6015), .B2(n5177), .A(n5063), .ZN(U3012) );
  INV_X1 U6234 ( .A(n5497), .ZN(n5066) );
  AOI22_X1 U6235 ( .A1(n6329), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6368), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n5064) );
  OAI21_X1 U6236 ( .B1(n6341), .B2(n5482), .A(n5064), .ZN(n5065) );
  AOI21_X1 U6237 ( .B1(n5066), .B2(n5804), .A(n5065), .ZN(n5067) );
  OAI21_X1 U6238 ( .B1(n5068), .B2(n6101), .A(n5067), .ZN(U2982) );
  INV_X1 U6239 ( .A(n5069), .ZN(n6203) );
  AOI21_X1 U6240 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5070), 
        .ZN(n5071) );
  OAI21_X1 U6241 ( .B1(n6341), .B2(n6201), .A(n5071), .ZN(n5072) );
  AOI21_X1 U6242 ( .B1(n6203), .B2(n5804), .A(n5072), .ZN(n5073) );
  OAI21_X1 U6243 ( .B1(n5074), .B2(n6101), .A(n5073), .ZN(U2983) );
  NOR2_X1 U6244 ( .A1(n5096), .A2(n6540), .ZN(n5078) );
  AOI22_X1 U6245 ( .A1(n6605), .A2(n5098), .B1(n5097), .B2(n6606), .ZN(n5076)
         );
  OAI21_X1 U6246 ( .B1(n5100), .B2(n6610), .A(n5076), .ZN(n5077) );
  AOI211_X1 U6247 ( .C1(n5103), .C2(INSTQUEUE_REG_14__3__SCAN_IN), .A(n5078), 
        .B(n5077), .ZN(n5079) );
  INV_X1 U6248 ( .A(n5079), .ZN(U3135) );
  NOR2_X1 U6249 ( .A1(n5096), .A2(n6545), .ZN(n5082) );
  AOI22_X1 U6250 ( .A1(n6611), .A2(n5098), .B1(n5097), .B2(n6612), .ZN(n5080)
         );
  OAI21_X1 U6251 ( .B1(n5100), .B2(n6616), .A(n5080), .ZN(n5081) );
  AOI211_X1 U6252 ( .C1(n5103), .C2(INSTQUEUE_REG_14__4__SCAN_IN), .A(n5082), 
        .B(n5081), .ZN(n5083) );
  INV_X1 U6253 ( .A(n5083), .ZN(U3136) );
  NOR2_X1 U6254 ( .A1(n5096), .A2(n6553), .ZN(n5086) );
  AOI22_X1 U6255 ( .A1(n6617), .A2(n5098), .B1(n5097), .B2(n6618), .ZN(n5084)
         );
  OAI21_X1 U6256 ( .B1(n5100), .B2(n6622), .A(n5084), .ZN(n5085) );
  AOI211_X1 U6257 ( .C1(n5103), .C2(INSTQUEUE_REG_14__5__SCAN_IN), .A(n5086), 
        .B(n5085), .ZN(n5087) );
  INV_X1 U6258 ( .A(n5087), .ZN(U3137) );
  NOR2_X1 U6259 ( .A1(n5096), .A2(n6535), .ZN(n5090) );
  AOI22_X1 U6260 ( .A1(n6599), .A2(n5098), .B1(n5097), .B2(n6600), .ZN(n5088)
         );
  OAI21_X1 U6261 ( .B1(n5100), .B2(n6604), .A(n5088), .ZN(n5089) );
  AOI211_X1 U6262 ( .C1(n5103), .C2(INSTQUEUE_REG_14__2__SCAN_IN), .A(n5090), 
        .B(n5089), .ZN(n5091) );
  INV_X1 U6263 ( .A(n5091), .ZN(U3134) );
  NOR2_X1 U6264 ( .A1(n5096), .A2(n6561), .ZN(n5094) );
  AOI22_X1 U6265 ( .A1(n6630), .A2(n5098), .B1(n5097), .B2(n6631), .ZN(n5092)
         );
  OAI21_X1 U6266 ( .B1(n5100), .B2(n6639), .A(n5092), .ZN(n5093) );
  AOI211_X1 U6267 ( .C1(n5103), .C2(INSTQUEUE_REG_14__7__SCAN_IN), .A(n5094), 
        .B(n5093), .ZN(n5095) );
  INV_X1 U6268 ( .A(n5095), .ZN(U3139) );
  NOR2_X1 U6269 ( .A1(n5096), .A2(n6530), .ZN(n5102) );
  AOI22_X1 U6270 ( .A1(n6593), .A2(n5098), .B1(n5097), .B2(n6594), .ZN(n5099)
         );
  OAI21_X1 U6271 ( .B1(n5100), .B2(n6598), .A(n5099), .ZN(n5101) );
  AOI211_X1 U6272 ( .C1(n5103), .C2(INSTQUEUE_REG_14__1__SCAN_IN), .A(n5102), 
        .B(n5101), .ZN(n5104) );
  INV_X1 U6273 ( .A(n5104), .ZN(U3133) );
  INV_X1 U6274 ( .A(n5105), .ZN(n6193) );
  AOI21_X1 U6275 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n5106), 
        .ZN(n5107) );
  OAI21_X1 U6276 ( .B1(n6341), .B2(n6196), .A(n5107), .ZN(n5108) );
  AOI21_X1 U6277 ( .B1(n6193), .B2(n5804), .A(n5108), .ZN(n5109) );
  OAI21_X1 U6278 ( .B1(n6101), .B2(n5110), .A(n5109), .ZN(U2981) );
  AOI21_X1 U6279 ( .B1(n5120), .B2(n6432), .A(n6582), .ZN(n5112) );
  NAND2_X1 U6280 ( .A1(n4503), .A2(n6218), .ZN(n6046) );
  INV_X1 U6281 ( .A(n6399), .ZN(n5111) );
  OAI21_X1 U6282 ( .B1(n5112), .B2(n5111), .A(n6050), .ZN(n5116) );
  NOR2_X1 U6283 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6284 ( .A1(n6522), .A2(n5113), .ZN(n5125) );
  INV_X1 U6285 ( .A(n5114), .ZN(n5115) );
  INV_X1 U6286 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U6287 ( .A1(n6584), .A2(n5118), .ZN(n5119) );
  OAI21_X1 U6288 ( .B1(n6399), .B2(n6578), .A(n5119), .ZN(n5151) );
  OAI22_X1 U6289 ( .A1(n6432), .A2(n6558), .B1(n6554), .B2(n5125), .ZN(n5122)
         );
  NOR2_X1 U6290 ( .A1(n5120), .A2(n6628), .ZN(n5121) );
  AOI211_X1 U6291 ( .C1(n6624), .C2(n5151), .A(n5122), .B(n5121), .ZN(n5123)
         );
  OAI21_X1 U6292 ( .B1(n5156), .B2(n5124), .A(n5123), .ZN(U3042) );
  INV_X1 U6293 ( .A(n5125), .ZN(n5150) );
  AOI22_X1 U6294 ( .A1(n6612), .A2(n5151), .B1(n6611), .B2(n5150), .ZN(n5126)
         );
  OAI21_X1 U6295 ( .B1(n6432), .B2(n6545), .A(n5126), .ZN(n5127) );
  AOI21_X1 U6296 ( .B1(n6077), .B2(n5154), .A(n5127), .ZN(n5128) );
  OAI21_X1 U6297 ( .B1(n5156), .B2(n5129), .A(n5128), .ZN(U3040) );
  INV_X1 U6298 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5133) );
  AOI22_X1 U6299 ( .A1(n6594), .A2(n5151), .B1(n6593), .B2(n5150), .ZN(n5130)
         );
  OAI21_X1 U6300 ( .B1(n6432), .B2(n6530), .A(n5130), .ZN(n5131) );
  AOI21_X1 U6301 ( .B1(n6062), .B2(n5154), .A(n5131), .ZN(n5132) );
  OAI21_X1 U6302 ( .B1(n5156), .B2(n5133), .A(n5132), .ZN(U3037) );
  AOI22_X1 U6303 ( .A1(n6606), .A2(n5151), .B1(n6605), .B2(n5150), .ZN(n5134)
         );
  OAI21_X1 U6304 ( .B1(n6432), .B2(n6540), .A(n5134), .ZN(n5135) );
  AOI21_X1 U6305 ( .B1(n6072), .B2(n5154), .A(n5135), .ZN(n5136) );
  OAI21_X1 U6306 ( .B1(n5156), .B2(n5137), .A(n5136), .ZN(U3039) );
  AOI22_X1 U6307 ( .A1(n6631), .A2(n5151), .B1(n6630), .B2(n5150), .ZN(n5138)
         );
  OAI21_X1 U6308 ( .B1(n6432), .B2(n6561), .A(n5138), .ZN(n5139) );
  AOI21_X1 U6309 ( .B1(n5140), .B2(n5154), .A(n5139), .ZN(n5141) );
  OAI21_X1 U6310 ( .B1(n5156), .B2(n6749), .A(n5141), .ZN(U3043) );
  AOI22_X1 U6311 ( .A1(n6600), .A2(n5151), .B1(n6599), .B2(n5150), .ZN(n5142)
         );
  OAI21_X1 U6312 ( .B1(n6432), .B2(n6535), .A(n5142), .ZN(n5143) );
  AOI21_X1 U6313 ( .B1(n6067), .B2(n5154), .A(n5143), .ZN(n5144) );
  OAI21_X1 U6314 ( .B1(n5156), .B2(n5145), .A(n5144), .ZN(U3038) );
  INV_X1 U6315 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5149) );
  AOI22_X1 U6316 ( .A1(n6577), .A2(n5151), .B1(n6576), .B2(n5150), .ZN(n5146)
         );
  OAI21_X1 U6317 ( .B1(n6432), .B2(n6528), .A(n5146), .ZN(n5147) );
  AOI21_X1 U6318 ( .B1(n6470), .B2(n5154), .A(n5147), .ZN(n5148) );
  OAI21_X1 U6319 ( .B1(n5156), .B2(n5149), .A(n5148), .ZN(U3036) );
  AOI22_X1 U6320 ( .A1(n6618), .A2(n5151), .B1(n6617), .B2(n5150), .ZN(n5152)
         );
  OAI21_X1 U6321 ( .B1(n6432), .B2(n6553), .A(n5152), .ZN(n5153) );
  AOI21_X1 U6322 ( .B1(n6082), .B2(n5154), .A(n5153), .ZN(n5155) );
  OAI21_X1 U6323 ( .B1(n5156), .B2(n6842), .A(n5155), .ZN(U3041) );
  INV_X1 U6324 ( .A(n5157), .ZN(n6226) );
  NAND2_X1 U6325 ( .A1(n6226), .A2(n5804), .ZN(n5162) );
  INV_X1 U6326 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5158) );
  NOR2_X1 U6327 ( .A1(n5784), .A2(n5158), .ZN(n5159) );
  AOI211_X1 U6328 ( .C1(n5787), .C2(n5158), .A(n5160), .B(n5159), .ZN(n5161)
         );
  OAI211_X1 U6329 ( .C1(n5163), .C2(n6101), .A(n5162), .B(n5161), .ZN(U2985)
         );
  NOR2_X1 U6330 ( .A1(READY_N), .A2(n6722), .ZN(n6640) );
  AOI21_X1 U6331 ( .B1(n5164), .B2(n6640), .A(n5208), .ZN(n5172) );
  AOI21_X1 U6332 ( .B1(READY_N), .B2(n5165), .A(n5201), .ZN(n5203) );
  INV_X1 U6333 ( .A(n5203), .ZN(n5166) );
  NAND3_X1 U6334 ( .A1(n5166), .A2(STATE2_REG_1__SCAN_IN), .A3(
        STATE2_REG_0__SCAN_IN), .ZN(n5171) );
  OAI21_X1 U6335 ( .B1(n5168), .B2(n6016), .A(n5167), .ZN(n5169) );
  INV_X1 U6336 ( .A(n5169), .ZN(n5170) );
  OAI211_X1 U6337 ( .C1(n5201), .C2(n5172), .A(n5171), .B(n5170), .ZN(U3149)
         );
  INV_X1 U6338 ( .A(n5173), .ZN(n6181) );
  AOI22_X1 U6339 ( .A1(n6329), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6368), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n5174) );
  OAI21_X1 U6340 ( .B1(n6341), .B2(n6184), .A(n5174), .ZN(n5175) );
  AOI21_X1 U6341 ( .B1(n6181), .B2(n5804), .A(n5175), .ZN(n5176) );
  OAI21_X1 U6342 ( .B1(n5177), .B2(n6101), .A(n5176), .ZN(U2980) );
  AOI21_X1 U6343 ( .B1(n5178), .B2(n4878), .A(n3941), .ZN(n6169) );
  INV_X1 U6344 ( .A(n6169), .ZN(n5556) );
  OAI222_X1 U6345 ( .A1(n5556), .A2(n5591), .B1(n5180), .B2(n6837), .C1(n5213), 
        .C2(n3918), .ZN(U2884) );
  NOR2_X1 U6346 ( .A1(n3820), .A2(n6662), .ZN(n6357) );
  NOR2_X1 U6347 ( .A1(n6341), .A2(n6176), .ZN(n5181) );
  AOI211_X1 U6348 ( .C1(n6329), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6357), 
        .B(n5181), .ZN(n5186) );
  INV_X1 U6349 ( .A(n5183), .ZN(n5184) );
  XNOR2_X1 U6350 ( .A(n5182), .B(n5184), .ZN(n6356) );
  NAND2_X1 U6351 ( .A1(n6356), .A2(n6336), .ZN(n5185) );
  OAI211_X1 U6352 ( .C1(n5556), .C2(n5797), .A(n5186), .B(n5185), .ZN(U2979)
         );
  INV_X1 U6353 ( .A(n5188), .ZN(n5189) );
  AOI22_X1 U6354 ( .A1(n5193), .A2(n5187), .B1(n5190), .B2(n5189), .ZN(n5191)
         );
  OAI21_X1 U6355 ( .B1(n5192), .B2(n6038), .A(n5191), .ZN(n5195) );
  AOI22_X1 U6356 ( .A1(n5197), .A2(n5195), .B1(n5194), .B2(n5193), .ZN(n5196)
         );
  OAI21_X1 U6357 ( .B1(n3146), .B2(n5197), .A(n5196), .ZN(U3460) );
  INV_X1 U6358 ( .A(n5198), .ZN(n5200) );
  OAI21_X1 U6359 ( .B1(n5200), .B2(n3163), .A(n5199), .ZN(n6017) );
  INV_X1 U6360 ( .A(n5201), .ZN(n5202) );
  OAI21_X1 U6361 ( .B1(n6718), .B2(n6036), .A(n5202), .ZN(n5204) );
  MUX2_X1 U6362 ( .A(n5204), .B(n5203), .S(STATE2_REG_0__SCAN_IN), .Z(n5211)
         );
  INV_X1 U6363 ( .A(n5205), .ZN(n5209) );
  INV_X1 U6364 ( .A(n5206), .ZN(n5207) );
  AOI21_X1 U6365 ( .B1(n5209), .B2(n5208), .A(n5207), .ZN(n5210) );
  OAI211_X1 U6366 ( .C1(n5212), .C2(n6017), .A(n5211), .B(n5210), .ZN(U3148)
         );
  AND2_X1 U6367 ( .A1(n5213), .A2(n5558), .ZN(n5214) );
  NAND2_X1 U6368 ( .A1(n5215), .A2(n5214), .ZN(n5218) );
  AOI22_X1 U6369 ( .A1(n5597), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5612), .ZN(n5217) );
  NAND2_X1 U6370 ( .A1(n5218), .A2(n5217), .ZN(U2860) );
  INV_X1 U6371 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6785) );
  NAND2_X1 U6372 ( .A1(n6785), .A2(n5219), .ZN(n5222) );
  INV_X1 U6373 ( .A(n5220), .ZN(n5221) );
  MUX2_X1 U6374 ( .A(n5222), .B(n5221), .S(n6725), .Z(U3474) );
  MUX2_X1 U6375 ( .A(W_R_N_REG_SCAN_IN), .B(n6785), .S(n6099), .Z(U3470) );
  INV_X1 U6376 ( .A(n5223), .ZN(n5224) );
  INV_X1 U6377 ( .A(n5226), .ZN(n5227) );
  AOI21_X1 U6378 ( .B1(n5229), .B2(n5228), .A(n5227), .ZN(n5237) );
  INV_X1 U6379 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6756) );
  NAND2_X1 U6380 ( .A1(n5230), .A2(n6756), .ZN(n5233) );
  INV_X1 U6381 ( .A(n5231), .ZN(n5232) );
  OAI21_X1 U6382 ( .B1(n3530), .B2(n5233), .A(n5232), .ZN(n5234) );
  INV_X1 U6383 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5506) );
  OAI22_X1 U6384 ( .A1(n6229), .A2(n5506), .B1(n5235), .B2(n6186), .ZN(n5236)
         );
  AOI211_X1 U6385 ( .C1(n6889), .C2(n5238), .A(n5237), .B(n5236), .ZN(n5239)
         );
  OAI211_X1 U6386 ( .C1(n5507), .C2(n6899), .A(n5240), .B(n5239), .ZN(U2797)
         );
  INV_X1 U6387 ( .A(n5622), .ZN(n5565) );
  INV_X1 U6388 ( .A(n5811), .ZN(n5245) );
  NOR2_X1 U6389 ( .A1(n6223), .A2(n5620), .ZN(n5244) );
  INV_X1 U6390 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6695) );
  NAND3_X1 U6391 ( .A1(n5254), .A2(REIP_REG_28__SCAN_IN), .A3(n6695), .ZN(
        n5242) );
  AOI22_X1 U6392 ( .A1(n6895), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6894), .ZN(n5241) );
  OAI211_X1 U6393 ( .C1(n5252), .C2(n6695), .A(n5242), .B(n5241), .ZN(n5243)
         );
  AOI211_X1 U6394 ( .C1(n5245), .C2(n6220), .A(n5244), .B(n5243), .ZN(n5246)
         );
  OAI21_X1 U6395 ( .B1(n5565), .B2(n5481), .A(n5246), .ZN(U2798) );
  AND2_X1 U6396 ( .A1(n2982), .A2(n5249), .ZN(n5251) );
  INV_X1 U6397 ( .A(n5508), .ZN(n5820) );
  AOI22_X1 U6398 ( .A1(n6895), .A2(EBX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6894), .ZN(n5256) );
  INV_X1 U6399 ( .A(n5252), .ZN(n5253) );
  OAI21_X1 U6400 ( .B1(n5254), .B2(REIP_REG_28__SCAN_IN), .A(n5253), .ZN(n5255) );
  OAI211_X1 U6401 ( .C1(n6223), .C2(n5628), .A(n5256), .B(n5255), .ZN(n5257)
         );
  AOI21_X1 U6402 ( .B1(n5820), .B2(n6220), .A(n5257), .ZN(n5258) );
  OAI21_X1 U6403 ( .B1(n5626), .B2(n5481), .A(n5258), .ZN(U2799) );
  NAND2_X1 U6404 ( .A1(n5261), .A2(n5262), .ZN(n5263) );
  NAND2_X1 U6405 ( .A1(n2982), .A2(n5263), .ZN(n5510) );
  INV_X1 U6406 ( .A(n5510), .ZN(n5826) );
  INV_X1 U6407 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5511) );
  OAI22_X1 U6408 ( .A1(n6229), .A2(n5511), .B1(n5264), .B2(n6186), .ZN(n5267)
         );
  INV_X1 U6409 ( .A(n5295), .ZN(n5310) );
  NOR3_X1 U6410 ( .A1(n5310), .A2(REIP_REG_27__SCAN_IN), .A3(n5265), .ZN(n5266) );
  AOI211_X1 U6411 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5275), .A(n5267), .B(n5266), .ZN(n5268) );
  OAI21_X1 U6412 ( .B1(n6223), .B2(n5637), .A(n5268), .ZN(n5269) );
  AOI21_X1 U6413 ( .B1(n5826), .B2(n6220), .A(n5269), .ZN(n5270) );
  OAI21_X1 U6414 ( .B1(n5570), .B2(n5481), .A(n5270), .ZN(U2800) );
  AOI21_X1 U6415 ( .B1(n5273), .B2(n5271), .A(n5272), .ZN(n5649) );
  INV_X1 U6416 ( .A(n5649), .ZN(n5573) );
  AOI21_X1 U6417 ( .B1(n5295), .B2(n5274), .A(REIP_REG_26__SCAN_IN), .ZN(n5278) );
  INV_X1 U6418 ( .A(n5275), .ZN(n5277) );
  AOI22_X1 U6419 ( .A1(n6895), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6894), .ZN(n5276) );
  OAI21_X1 U6420 ( .B1(n5278), .B2(n5277), .A(n5276), .ZN(n5282) );
  OAI21_X1 U6421 ( .B1(n5279), .B2(n5280), .A(n5261), .ZN(n5834) );
  NOR2_X1 U6422 ( .A1(n5834), .A2(n6899), .ZN(n5281) );
  AOI211_X1 U6423 ( .C1(n6889), .C2(n5644), .A(n5282), .B(n5281), .ZN(n5283)
         );
  OAI21_X1 U6424 ( .B1(n5573), .B2(n5481), .A(n5283), .ZN(U2801) );
  INV_X1 U6425 ( .A(n5271), .ZN(n5286) );
  AOI21_X1 U6426 ( .B1(n5287), .B2(n5285), .A(n5286), .ZN(n5658) );
  INV_X1 U6427 ( .A(n5658), .ZN(n5576) );
  NOR2_X1 U6428 ( .A1(n5306), .A2(n5289), .ZN(n5290) );
  OR2_X1 U6429 ( .A1(n5279), .A2(n5290), .ZN(n5849) );
  INV_X1 U6430 ( .A(n5849), .ZN(n5299) );
  NAND2_X1 U6431 ( .A1(n6895), .A2(EBX_REG_25__SCAN_IN), .ZN(n5291) );
  OAI21_X1 U6432 ( .B1(n6186), .B2(n5292), .A(n5291), .ZN(n5293) );
  AOI21_X1 U6433 ( .B1(n5320), .B2(REIP_REG_25__SCAN_IN), .A(n5293), .ZN(n5297) );
  INV_X1 U6434 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6684) );
  XNOR2_X1 U6435 ( .A(n6684), .B(REIP_REG_25__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6436 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  OAI211_X1 U6437 ( .C1(n6223), .C2(n5656), .A(n5297), .B(n5296), .ZN(n5298)
         );
  AOI21_X1 U6438 ( .B1(n5299), .B2(n6220), .A(n5298), .ZN(n5300) );
  OAI21_X1 U6439 ( .B1(n5576), .B2(n5481), .A(n5300), .ZN(U2802) );
  OAI21_X1 U6440 ( .B1(n5301), .B2(n5302), .A(n5285), .ZN(n5664) );
  AND2_X1 U6441 ( .A1(n5303), .A2(n5304), .ZN(n5305) );
  NOR2_X1 U6442 ( .A1(n5306), .A2(n5305), .ZN(n5859) );
  NOR2_X1 U6443 ( .A1(n6223), .A2(n5666), .ZN(n5312) );
  INV_X1 U6444 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6805) );
  OAI22_X1 U6445 ( .A1(n6229), .A2(n6805), .B1(n5307), .B2(n6186), .ZN(n5308)
         );
  AOI21_X1 U6446 ( .B1(REIP_REG_24__SCAN_IN), .B2(n5320), .A(n5308), .ZN(n5309) );
  OAI21_X1 U6447 ( .B1(n5310), .B2(REIP_REG_24__SCAN_IN), .A(n5309), .ZN(n5311) );
  AOI211_X1 U6448 ( .C1(n5859), .C2(n6220), .A(n5312), .B(n5311), .ZN(n5313)
         );
  OAI21_X1 U6449 ( .B1(n5664), .B2(n5481), .A(n5313), .ZN(U2803) );
  NOR2_X1 U6450 ( .A1(n5314), .A2(n5315), .ZN(n5316) );
  INV_X1 U6451 ( .A(n5676), .ZN(n5325) );
  NAND2_X1 U6452 ( .A1(n5338), .A2(n5317), .ZN(n5318) );
  AND2_X1 U6453 ( .A1(n5303), .A2(n5318), .ZN(n5863) );
  INV_X1 U6454 ( .A(n5863), .ZN(n5515) );
  AOI22_X1 U6455 ( .A1(n6895), .A2(EBX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6894), .ZN(n5323) );
  INV_X1 U6456 ( .A(n5319), .ZN(n5321) );
  OAI21_X1 U6457 ( .B1(n5321), .B2(REIP_REG_23__SCAN_IN), .A(n5320), .ZN(n5322) );
  OAI211_X1 U6458 ( .C1(n5515), .C2(n6899), .A(n5323), .B(n5322), .ZN(n5324)
         );
  AOI21_X1 U6459 ( .B1(n5325), .B2(n6889), .A(n5324), .ZN(n5326) );
  OAI21_X1 U6460 ( .B1(n5673), .B2(n5481), .A(n5326), .ZN(U2804) );
  AND2_X1 U6461 ( .A1(n5343), .A2(n5328), .ZN(n5329) );
  OR2_X1 U6462 ( .A1(n5329), .A2(n5314), .ZN(n5683) );
  INV_X1 U6463 ( .A(n5352), .ZN(n5332) );
  INV_X1 U6464 ( .A(n5330), .ZN(n5331) );
  OAI211_X1 U6465 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5332), .B(n5331), .ZN(n5335) );
  NOR2_X1 U6466 ( .A1(n6186), .A2(n5682), .ZN(n5333) );
  AOI21_X1 U6467 ( .B1(n6895), .B2(EBX_REG_22__SCAN_IN), .A(n5333), .ZN(n5334)
         );
  OAI211_X1 U6468 ( .C1(n5361), .C2(n6682), .A(n5335), .B(n5334), .ZN(n5340)
         );
  OR2_X1 U6469 ( .A1(n5348), .A2(n5336), .ZN(n5337) );
  NAND2_X1 U6470 ( .A1(n5338), .A2(n5337), .ZN(n5871) );
  NOR2_X1 U6471 ( .A1(n5871), .A2(n6899), .ZN(n5339) );
  AOI211_X1 U6472 ( .C1(n6889), .C2(n5686), .A(n5340), .B(n5339), .ZN(n5341)
         );
  OAI21_X1 U6473 ( .B1(n5683), .B2(n5481), .A(n5341), .ZN(U2805) );
  AOI21_X1 U6474 ( .B1(n5344), .B2(n5342), .A(n5327), .ZN(n5695) );
  INV_X1 U6475 ( .A(n5695), .ZN(n5585) );
  NOR2_X1 U6476 ( .A1(n5346), .A2(n5345), .ZN(n5347) );
  NOR2_X1 U6477 ( .A1(n5348), .A2(n5347), .ZN(n5881) );
  AOI22_X1 U6478 ( .A1(n6895), .A2(EBX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6894), .ZN(n5351) );
  INV_X1 U6479 ( .A(n5361), .ZN(n5349) );
  NAND2_X1 U6480 ( .A1(n5349), .A2(REIP_REG_21__SCAN_IN), .ZN(n5350) );
  OAI211_X1 U6481 ( .C1(n5352), .C2(REIP_REG_21__SCAN_IN), .A(n5351), .B(n5350), .ZN(n5354) );
  NOR2_X1 U6482 ( .A1(n6223), .A2(n5693), .ZN(n5353) );
  AOI211_X1 U6483 ( .C1(n5881), .C2(n6220), .A(n5354), .B(n5353), .ZN(n5355)
         );
  OAI21_X1 U6484 ( .B1(n5585), .B2(n5481), .A(n5355), .ZN(U2806) );
  MUX2_X1 U6485 ( .A(n3190), .B(n5372), .S(n5356), .Z(n5357) );
  XOR2_X1 U6486 ( .A(n5358), .B(n5357), .Z(n5895) );
  XOR2_X1 U6487 ( .A(n5360), .B(n5359), .Z(n5702) );
  NAND2_X1 U6488 ( .A1(n5702), .A2(n6890), .ZN(n5366) );
  INV_X1 U6489 ( .A(n5395), .ZN(n5382) );
  NAND3_X1 U6490 ( .A1(n5382), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .ZN(n5362) );
  AOI21_X1 U6491 ( .B1(n5362), .B2(n4441), .A(n5361), .ZN(n5364) );
  INV_X1 U6492 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5520) );
  OAI22_X1 U6493 ( .A1(n6229), .A2(n5520), .B1(n3074), .B2(n6186), .ZN(n5363)
         );
  AOI211_X1 U6494 ( .C1(n6889), .C2(n5699), .A(n5364), .B(n5363), .ZN(n5365)
         );
  OAI211_X1 U6495 ( .C1(n5895), .C2(n6899), .A(n5366), .B(n5365), .ZN(U2807)
         );
  AND2_X1 U6496 ( .A1(n5367), .A2(n5368), .ZN(n5369) );
  INV_X1 U6497 ( .A(n5706), .ZN(n5385) );
  INV_X1 U6498 ( .A(n5406), .ZN(n5373) );
  MUX2_X1 U6499 ( .A(n5372), .B(n5371), .S(n3190), .Z(n5390) );
  NAND2_X1 U6500 ( .A1(n5373), .A2(n5390), .ZN(n5393) );
  XNOR2_X1 U6501 ( .A(n5393), .B(n5374), .ZN(n5904) );
  XOR2_X1 U6502 ( .A(REIP_REG_18__SCAN_IN), .B(REIP_REG_19__SCAN_IN), .Z(n5381) );
  NAND2_X1 U6503 ( .A1(n6197), .A2(n5375), .ZN(n6896) );
  AOI21_X1 U6504 ( .B1(n6894), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6188), 
        .ZN(n5376) );
  OAI21_X1 U6505 ( .B1(n6229), .B2(n5521), .A(n5376), .ZN(n5380) );
  INV_X1 U6506 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6675) );
  OR2_X1 U6507 ( .A1(n5377), .A2(n6675), .ZN(n5378) );
  NAND2_X1 U6508 ( .A1(n6170), .A2(n5378), .ZN(n5408) );
  INV_X1 U6509 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6679) );
  NOR2_X1 U6510 ( .A1(n5408), .A2(n6679), .ZN(n5379) );
  AOI211_X1 U6511 ( .C1(n5382), .C2(n5381), .A(n5380), .B(n5379), .ZN(n5383)
         );
  OAI21_X1 U6512 ( .B1(n5904), .B2(n6899), .A(n5383), .ZN(n5384) );
  AOI21_X1 U6513 ( .B1(n6889), .B2(n5385), .A(n5384), .ZN(n5386) );
  OAI21_X1 U6514 ( .B1(n5710), .B2(n5481), .A(n5386), .ZN(U2808) );
  INV_X1 U6515 ( .A(n5367), .ZN(n5388) );
  AOI21_X1 U6516 ( .B1(n5389), .B2(n5387), .A(n5388), .ZN(n5718) );
  INV_X1 U6517 ( .A(n5718), .ZN(n5594) );
  INV_X1 U6518 ( .A(n5390), .ZN(n5391) );
  NAND2_X1 U6519 ( .A1(n5406), .A2(n5391), .ZN(n5392) );
  AND2_X1 U6520 ( .A1(n5393), .A2(n5392), .ZN(n5914) );
  INV_X1 U6521 ( .A(n5914), .ZN(n5523) );
  INV_X1 U6522 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6677) );
  AOI21_X1 U6523 ( .B1(n6894), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6188), 
        .ZN(n5394) );
  OAI221_X1 U6524 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5395), .C1(n6677), .C2(
        n5408), .A(n5394), .ZN(n5396) );
  AOI21_X1 U6525 ( .B1(n6895), .B2(EBX_REG_18__SCAN_IN), .A(n5396), .ZN(n5397)
         );
  OAI21_X1 U6526 ( .B1(n5523), .B2(n6899), .A(n5397), .ZN(n5398) );
  AOI21_X1 U6527 ( .B1(n6889), .B2(n5714), .A(n5398), .ZN(n5399) );
  OAI21_X1 U6528 ( .B1(n5594), .B2(n5481), .A(n5399), .ZN(U2809) );
  OR2_X1 U6529 ( .A1(n5400), .A2(n5401), .ZN(n5402) );
  NAND2_X1 U6530 ( .A1(n5387), .A2(n5402), .ZN(n5723) );
  INV_X1 U6531 ( .A(n5725), .ZN(n5414) );
  NAND2_X1 U6532 ( .A1(n5420), .A2(n5404), .ZN(n5405) );
  NAND2_X1 U6533 ( .A1(n5406), .A2(n5405), .ZN(n5925) );
  OAI21_X1 U6534 ( .B1(n6186), .B2(n6776), .A(n6896), .ZN(n5407) );
  AOI21_X1 U6535 ( .B1(n6895), .B2(EBX_REG_17__SCAN_IN), .A(n5407), .ZN(n5412)
         );
  INV_X1 U6536 ( .A(n5408), .ZN(n5409) );
  OAI21_X1 U6537 ( .B1(n5410), .B2(REIP_REG_17__SCAN_IN), .A(n5409), .ZN(n5411) );
  OAI211_X1 U6538 ( .C1(n5925), .C2(n6899), .A(n5412), .B(n5411), .ZN(n5413)
         );
  AOI21_X1 U6539 ( .B1(n6889), .B2(n5414), .A(n5413), .ZN(n5415) );
  OAI21_X1 U6540 ( .B1(n5723), .B2(n5481), .A(n5415), .ZN(U2810) );
  AOI21_X1 U6541 ( .B1(n5417), .B2(n5416), .A(n5400), .ZN(n5418) );
  INV_X1 U6542 ( .A(n5418), .ZN(n5734) );
  INV_X1 U6543 ( .A(n5420), .ZN(n5421) );
  AOI21_X1 U6544 ( .B1(n5422), .B2(n5419), .A(n5421), .ZN(n5941) );
  INV_X1 U6545 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5430) );
  OR2_X1 U6546 ( .A1(n6206), .A2(n5441), .ZN(n6117) );
  NAND2_X1 U6547 ( .A1(n6117), .A2(n6197), .ZN(n6118) );
  NAND2_X1 U6548 ( .A1(n6118), .A2(REIP_REG_16__SCAN_IN), .ZN(n5429) );
  INV_X1 U6549 ( .A(n6206), .ZN(n6217) );
  XNOR2_X1 U6550 ( .A(REIP_REG_16__SCAN_IN), .B(REIP_REG_15__SCAN_IN), .ZN(
        n5423) );
  NOR2_X1 U6551 ( .A1(n5424), .A2(n5423), .ZN(n5427) );
  OAI21_X1 U6552 ( .B1(n6186), .B2(n5425), .A(n6896), .ZN(n5426) );
  AOI21_X1 U6553 ( .B1(n6217), .B2(n5427), .A(n5426), .ZN(n5428) );
  OAI211_X1 U6554 ( .C1(n6229), .C2(n5430), .A(n5429), .B(n5428), .ZN(n5432)
         );
  NOR2_X1 U6555 ( .A1(n6223), .A2(n5730), .ZN(n5431) );
  AOI211_X1 U6556 ( .C1(n5941), .C2(n6220), .A(n5432), .B(n5431), .ZN(n5433)
         );
  OAI21_X1 U6557 ( .B1(n5734), .B2(n5481), .A(n5433), .ZN(U2811) );
  XOR2_X1 U6558 ( .A(n5437), .B(n5435), .Z(n5605) );
  INV_X1 U6559 ( .A(n5436), .ZN(n5604) );
  INV_X1 U6560 ( .A(n5437), .ZN(n5438) );
  OAI22_X1 U6561 ( .A1(n5605), .A2(n5604), .B1(n5438), .B2(n5435), .ZN(n5532)
         );
  NAND2_X1 U6562 ( .A1(n5532), .A2(n5531), .ZN(n5530) );
  INV_X1 U6563 ( .A(n5439), .ZN(n5440) );
  AOI21_X1 U6564 ( .B1(n5530), .B2(n5440), .A(n3128), .ZN(n5740) );
  NAND2_X1 U6565 ( .A1(n5740), .A2(n6890), .ZN(n5448) );
  AOI21_X1 U6566 ( .B1(n6894), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6188), 
        .ZN(n5443) );
  NAND3_X1 U6567 ( .A1(n6217), .A2(n6670), .A3(n5441), .ZN(n5442) );
  OAI211_X1 U6568 ( .C1(n6229), .C2(n5526), .A(n5443), .B(n5442), .ZN(n5446)
         );
  OAI21_X1 U6569 ( .B1(n5528), .B2(n5444), .A(n5419), .ZN(n5946) );
  NOR2_X1 U6570 ( .A1(n5946), .A2(n6899), .ZN(n5445) );
  AOI211_X1 U6571 ( .C1(REIP_REG_15__SCAN_IN), .C2(n6118), .A(n5446), .B(n5445), .ZN(n5447) );
  OAI211_X1 U6572 ( .C1(n6223), .C2(n5738), .A(n5448), .B(n5447), .ZN(U2812)
         );
  OAI21_X1 U6573 ( .B1(n2983), .B2(n5450), .A(n5449), .ZN(n5776) );
  INV_X1 U6574 ( .A(n5772), .ZN(n5464) );
  OR2_X1 U6575 ( .A1(n5452), .A2(n5453), .ZN(n5454) );
  AND2_X1 U6576 ( .A1(n5451), .A2(n5454), .ZN(n6343) );
  AOI22_X1 U6577 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6894), .B1(n6220), 
        .B2(n6343), .ZN(n5455) );
  OAI211_X1 U6578 ( .C1(n6229), .C2(n5537), .A(n5455), .B(n6896), .ZN(n5463)
         );
  INV_X1 U6580 ( .A(n6197), .ZN(n6216) );
  OR2_X1 U6581 ( .A1(n6216), .A2(n5456), .ZN(n5469) );
  OAI21_X1 U6582 ( .B1(n6135), .B2(n5469), .A(n6170), .ZN(n6149) );
  INV_X1 U6583 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6584 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5459) );
  INV_X1 U6585 ( .A(n5457), .ZN(n5458) );
  NOR2_X1 U6586 ( .A1(n6206), .A2(n5458), .ZN(n6154) );
  NAND2_X1 U6587 ( .A1(n6154), .A2(REIP_REG_8__SCAN_IN), .ZN(n6892) );
  OAI33_X1 U6588 ( .A1(1'b0), .A2(n6149), .A3(n5460), .B1(REIP_REG_11__SCAN_IN), .B2(n5459), .B3(n6892), .ZN(n5462) );
  AOI211_X1 U6589 ( .C1(n6889), .C2(n5464), .A(n5463), .B(n5462), .ZN(n5465)
         );
  OAI21_X1 U6590 ( .B1(n5481), .B2(n5776), .A(n5465), .ZN(U2816) );
  AND2_X1 U6591 ( .A1(n5466), .A2(n5467), .ZN(n5468) );
  OR2_X1 U6592 ( .A1(n5468), .A2(n2979), .ZN(n5796) );
  NAND2_X1 U6593 ( .A1(n6170), .A2(n5469), .ZN(n6161) );
  INV_X1 U6594 ( .A(n6161), .ZN(n6902) );
  INV_X1 U6595 ( .A(n6892), .ZN(n5475) );
  INV_X1 U6596 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6893) );
  INV_X1 U6597 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6850) );
  AOI21_X1 U6598 ( .B1(n5472), .B2(n5470), .A(n5471), .ZN(n6350) );
  AOI22_X1 U6599 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6894), .B1(n6220), 
        .B2(n6350), .ZN(n5473) );
  OAI211_X1 U6600 ( .C1(n6229), .C2(n6850), .A(n5473), .B(n6896), .ZN(n5474)
         );
  AOI21_X1 U6601 ( .B1(n5475), .B2(n6893), .A(n5474), .ZN(n5476) );
  OAI21_X1 U6602 ( .B1(n6223), .B2(n5792), .A(n5476), .ZN(n5477) );
  AOI21_X1 U6603 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6902), .A(n5477), .ZN(n5478)
         );
  OAI21_X1 U6604 ( .B1(n5481), .B2(n5796), .A(n5478), .ZN(U2818) );
  NAND2_X1 U6605 ( .A1(n5484), .A2(n5479), .ZN(n5480) );
  NAND2_X1 U6606 ( .A1(n5481), .A2(n5480), .ZN(n6225) );
  INV_X1 U6607 ( .A(n6225), .ZN(n6210) );
  INV_X1 U6608 ( .A(n5482), .ZN(n5495) );
  OAI21_X1 U6609 ( .B1(n6216), .B2(n5483), .A(n6170), .ZN(n6205) );
  NOR2_X1 U6610 ( .A1(n6205), .A2(n6658), .ZN(n5494) );
  OR2_X1 U6611 ( .A1(n6206), .A2(n5483), .ZN(n6190) );
  INV_X1 U6612 ( .A(n5484), .ZN(n5485) );
  NOR2_X1 U6613 ( .A1(n5485), .A2(n6711), .ZN(n6219) );
  INV_X1 U6614 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5486) );
  OAI21_X1 U6615 ( .B1(n6186), .B2(n5486), .A(n6896), .ZN(n5490) );
  OAI22_X1 U6616 ( .A1(n5488), .A2(n6229), .B1(n6899), .B2(n5487), .ZN(n5489)
         );
  AOI211_X1 U6617 ( .C1(n6219), .C2(n5491), .A(n5490), .B(n5489), .ZN(n5492)
         );
  OAI21_X1 U6618 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6190), .A(n5492), .ZN(n5493)
         );
  AOI211_X1 U6619 ( .C1(n6889), .C2(n5495), .A(n5494), .B(n5493), .ZN(n5496)
         );
  OAI21_X1 U6620 ( .B1(n6210), .B2(n5497), .A(n5496), .ZN(U2823) );
  OAI21_X1 U6621 ( .B1(n6889), .B2(n6894), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5502) );
  AOI22_X1 U6622 ( .A1(n6219), .A2(n5498), .B1(n6895), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5499) );
  OAI21_X1 U6623 ( .B1(n6899), .B2(n6386), .A(n5499), .ZN(n5500) );
  AOI21_X1 U6624 ( .B1(REIP_REG_0__SCAN_IN), .B2(n6170), .A(n5500), .ZN(n5501)
         );
  OAI211_X1 U6625 ( .C1(n6210), .C2(n5503), .A(n5502), .B(n5501), .ZN(U2827)
         );
  INV_X1 U6626 ( .A(n5504), .ZN(n5505) );
  OAI22_X1 U6627 ( .A1(n5505), .A2(n5557), .B1(n6756), .B2(n5552), .ZN(U2828)
         );
  OAI222_X1 U6628 ( .A1(n5544), .A2(n5562), .B1(n5557), .B2(n5507), .C1(n5506), 
        .C2(n5552), .ZN(U2829) );
  OAI222_X1 U6629 ( .A1(n5509), .A2(n5552), .B1(n5557), .B2(n5508), .C1(n5626), 
        .C2(n5544), .ZN(U2831) );
  INV_X1 U6630 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5512) );
  OAI222_X1 U6631 ( .A1(n5834), .A2(n5557), .B1(n5512), .B2(n5552), .C1(n5573), 
        .C2(n5544), .ZN(U2833) );
  INV_X1 U6632 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5513) );
  OAI222_X1 U6633 ( .A1(n5849), .A2(n5557), .B1(n5513), .B2(n5552), .C1(n5576), 
        .C2(n5544), .ZN(U2834) );
  INV_X1 U6634 ( .A(n5859), .ZN(n5514) );
  OAI222_X1 U6635 ( .A1(n6805), .A2(n5552), .B1(n5557), .B2(n5514), .C1(n5664), 
        .C2(n5544), .ZN(U2835) );
  OAI222_X1 U6636 ( .A1(n5516), .A2(n5552), .B1(n5557), .B2(n5515), .C1(n5673), 
        .C2(n5544), .ZN(U2836) );
  INV_X1 U6637 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5517) );
  OAI222_X1 U6638 ( .A1(n5517), .A2(n5552), .B1(n5557), .B2(n5871), .C1(n5683), 
        .C2(n5544), .ZN(U2837) );
  AOI22_X1 U6639 ( .A1(n5881), .A2(n6232), .B1(n5518), .B2(EBX_REG_21__SCAN_IN), .ZN(n5519) );
  OAI21_X1 U6640 ( .B1(n5585), .B2(n5544), .A(n5519), .ZN(U2838) );
  INV_X1 U6641 ( .A(n5702), .ZN(n5588) );
  OAI222_X1 U6642 ( .A1(n5588), .A2(n5544), .B1(n5552), .B2(n5520), .C1(n5557), 
        .C2(n5895), .ZN(U2839) );
  OAI222_X1 U6643 ( .A1(n5710), .A2(n5544), .B1(n5557), .B2(n5904), .C1(n5552), 
        .C2(n5521), .ZN(U2840) );
  INV_X1 U6644 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5522) );
  OAI222_X1 U6645 ( .A1(n5523), .A2(n5557), .B1(n5522), .B2(n5552), .C1(n5594), 
        .C2(n5544), .ZN(U2841) );
  OAI222_X1 U6646 ( .A1(n5925), .A2(n5557), .B1(n5524), .B2(n5552), .C1(n5723), 
        .C2(n5544), .ZN(U2842) );
  INV_X1 U6647 ( .A(n5941), .ZN(n5525) );
  OAI222_X1 U6648 ( .A1(n5525), .A2(n5557), .B1(n5552), .B2(n5430), .C1(n5544), 
        .C2(n5734), .ZN(U2843) );
  INV_X1 U6649 ( .A(n5740), .ZN(n5602) );
  OAI222_X1 U6650 ( .A1(n5946), .A2(n5557), .B1(n5526), .B2(n5552), .C1(n5602), 
        .C2(n5544), .ZN(U2844) );
  AND2_X1 U6651 ( .A1(n5973), .A2(n5527), .ZN(n5529) );
  OR2_X1 U6652 ( .A1(n5529), .A2(n5528), .ZN(n6129) );
  INV_X1 U6653 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5533) );
  OAI21_X1 U6654 ( .B1(n5532), .B2(n5531), .A(n5530), .ZN(n6123) );
  OAI222_X1 U6655 ( .A1(n6129), .A2(n5557), .B1(n5552), .B2(n5533), .C1(n5544), 
        .C2(n6123), .ZN(U2845) );
  AOI21_X1 U6656 ( .B1(n5534), .B2(n5449), .A(n4059), .ZN(n6142) );
  INV_X1 U6657 ( .A(n6142), .ZN(n5608) );
  INV_X1 U6658 ( .A(n5535), .ZN(n5972) );
  XNOR2_X1 U6659 ( .A(n5451), .B(n5972), .ZN(n6143) );
  INV_X1 U6660 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5536) );
  OAI222_X1 U6661 ( .A1(n5608), .A2(n5544), .B1(n5557), .B2(n6143), .C1(n5536), 
        .C2(n5552), .ZN(U2847) );
  NOR2_X1 U6662 ( .A1(n5552), .A2(n5537), .ZN(n5538) );
  AOI21_X1 U6663 ( .B1(n6343), .B2(n6232), .A(n5538), .ZN(n5539) );
  OAI21_X1 U6664 ( .B1(n5776), .B2(n5544), .A(n5539), .ZN(U2848) );
  NOR2_X1 U6665 ( .A1(n5471), .A2(n5540), .ZN(n5541) );
  OR2_X1 U6666 ( .A1(n5452), .A2(n5541), .ZN(n6898) );
  INV_X1 U6667 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5545) );
  NOR2_X1 U6668 ( .A1(n2979), .A2(n5542), .ZN(n5543) );
  OR2_X1 U6669 ( .A1(n2983), .A2(n5543), .ZN(n6887) );
  OAI222_X1 U6670 ( .A1(n6898), .A2(n5557), .B1(n5545), .B2(n5552), .C1(n6887), 
        .C2(n5544), .ZN(U2849) );
  INV_X1 U6671 ( .A(n6350), .ZN(n5546) );
  OAI222_X1 U6672 ( .A1(n5546), .A2(n5557), .B1(n5552), .B2(n6850), .C1(n5544), 
        .C2(n5796), .ZN(U2850) );
  NAND2_X1 U6673 ( .A1(n5547), .A2(n5548), .ZN(n5549) );
  NAND2_X1 U6674 ( .A1(n5470), .A2(n5549), .ZN(n6155) );
  INV_X1 U6675 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6794) );
  INV_X1 U6676 ( .A(n5466), .ZN(n5550) );
  AOI21_X1 U6677 ( .B1(n5551), .B2(n5179), .A(n5550), .ZN(n6158) );
  INV_X1 U6678 ( .A(n6158), .ZN(n5615) );
  OAI222_X1 U6679 ( .A1(n6155), .A2(n5557), .B1(n5552), .B2(n6794), .C1(n5544), 
        .C2(n5615), .ZN(U2851) );
  OR2_X1 U6680 ( .A1(n5554), .A2(n5553), .ZN(n5555) );
  AND2_X1 U6681 ( .A1(n5547), .A2(n5555), .ZN(n6358) );
  INV_X1 U6682 ( .A(n6358), .ZN(n6166) );
  INV_X1 U6683 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6808) );
  OAI222_X1 U6684 ( .A1(n6166), .A2(n5557), .B1(n5552), .B2(n6808), .C1(n5544), 
        .C2(n5556), .ZN(U2852) );
  AOI22_X1 U6685 ( .A1(n5597), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5612), .ZN(n5561) );
  NOR3_X1 U6686 ( .A1(n5612), .A2(n5558), .A3(n3426), .ZN(n5559) );
  NAND2_X1 U6687 ( .A1(n5598), .A2(DATAI_14_), .ZN(n5560) );
  OAI211_X1 U6688 ( .C1(n5562), .C2(n5591), .A(n5561), .B(n5560), .ZN(U2861)
         );
  AOI22_X1 U6689 ( .A1(n5597), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n5612), .ZN(n5564) );
  NAND2_X1 U6690 ( .A1(n5598), .A2(DATAI_13_), .ZN(n5563) );
  OAI211_X1 U6691 ( .C1(n5565), .C2(n5591), .A(n5564), .B(n5563), .ZN(U2862)
         );
  AOI22_X1 U6692 ( .A1(n5597), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5612), .ZN(n5567) );
  NAND2_X1 U6693 ( .A1(n5598), .A2(DATAI_12_), .ZN(n5566) );
  OAI211_X1 U6694 ( .C1(n5626), .C2(n5591), .A(n5567), .B(n5566), .ZN(U2863)
         );
  AOI22_X1 U6695 ( .A1(n5597), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5612), .ZN(n5569) );
  NAND2_X1 U6696 ( .A1(n5598), .A2(DATAI_11_), .ZN(n5568) );
  OAI211_X1 U6697 ( .C1(n5570), .C2(n5591), .A(n5569), .B(n5568), .ZN(U2864)
         );
  AOI22_X1 U6698 ( .A1(n5597), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5612), .ZN(n5572) );
  NAND2_X1 U6699 ( .A1(n5598), .A2(DATAI_10_), .ZN(n5571) );
  OAI211_X1 U6700 ( .C1(n5573), .C2(n5591), .A(n5572), .B(n5571), .ZN(U2865)
         );
  AOI22_X1 U6701 ( .A1(n5597), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n5612), .ZN(n5575) );
  NAND2_X1 U6702 ( .A1(n5598), .A2(DATAI_9_), .ZN(n5574) );
  OAI211_X1 U6703 ( .C1(n5576), .C2(n5591), .A(n5575), .B(n5574), .ZN(U2866)
         );
  AOI22_X1 U6704 ( .A1(n5597), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n5612), .ZN(n5578) );
  NAND2_X1 U6705 ( .A1(n5598), .A2(DATAI_8_), .ZN(n5577) );
  OAI211_X1 U6706 ( .C1(n5664), .C2(n5591), .A(n5578), .B(n5577), .ZN(U2867)
         );
  AOI22_X1 U6707 ( .A1(n5597), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n5612), .ZN(n5580) );
  NAND2_X1 U6708 ( .A1(n5598), .A2(DATAI_7_), .ZN(n5579) );
  OAI211_X1 U6709 ( .C1(n5673), .C2(n5591), .A(n5580), .B(n5579), .ZN(U2868)
         );
  AOI22_X1 U6710 ( .A1(n5597), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n5612), .ZN(n5582) );
  NAND2_X1 U6711 ( .A1(n5598), .A2(DATAI_6_), .ZN(n5581) );
  OAI211_X1 U6712 ( .C1(n5683), .C2(n5591), .A(n5582), .B(n5581), .ZN(U2869)
         );
  AOI22_X1 U6713 ( .A1(n5597), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n5612), .ZN(n5584) );
  NAND2_X1 U6714 ( .A1(n5598), .A2(DATAI_5_), .ZN(n5583) );
  OAI211_X1 U6715 ( .C1(n5585), .C2(n5591), .A(n5584), .B(n5583), .ZN(U2870)
         );
  AOI22_X1 U6716 ( .A1(n5597), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n5612), .ZN(n5587) );
  NAND2_X1 U6717 ( .A1(n5598), .A2(DATAI_4_), .ZN(n5586) );
  OAI211_X1 U6718 ( .C1(n5588), .C2(n5591), .A(n5587), .B(n5586), .ZN(U2871)
         );
  AOI22_X1 U6719 ( .A1(n5597), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n5612), .ZN(n5590) );
  NAND2_X1 U6720 ( .A1(n5598), .A2(DATAI_3_), .ZN(n5589) );
  OAI211_X1 U6721 ( .C1(n5710), .C2(n5591), .A(n5590), .B(n5589), .ZN(U2872)
         );
  AOI22_X1 U6722 ( .A1(n5597), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n5612), .ZN(n5593) );
  NAND2_X1 U6723 ( .A1(n5598), .A2(DATAI_2_), .ZN(n5592) );
  OAI211_X1 U6724 ( .C1(n5594), .C2(n5591), .A(n5593), .B(n5592), .ZN(U2873)
         );
  AOI22_X1 U6725 ( .A1(n5597), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n5612), .ZN(n5596) );
  NAND2_X1 U6726 ( .A1(n5598), .A2(DATAI_1_), .ZN(n5595) );
  OAI211_X1 U6727 ( .C1(n5723), .C2(n5591), .A(n5596), .B(n5595), .ZN(U2874)
         );
  AOI22_X1 U6728 ( .A1(n5597), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n5612), .ZN(n5600) );
  NAND2_X1 U6729 ( .A1(n5598), .A2(DATAI_0_), .ZN(n5599) );
  OAI211_X1 U6730 ( .C1(n5734), .C2(n5591), .A(n5600), .B(n5599), .ZN(U2875)
         );
  AOI22_X1 U6731 ( .A1(n5613), .A2(DATAI_15_), .B1(n5612), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5601) );
  OAI21_X1 U6732 ( .B1(n5602), .B2(n5591), .A(n5601), .ZN(U2876) );
  AOI22_X1 U6733 ( .A1(n5613), .A2(DATAI_14_), .B1(n5612), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5603) );
  OAI21_X1 U6734 ( .B1(n6123), .B2(n5591), .A(n5603), .ZN(U2877) );
  XNOR2_X1 U6735 ( .A(n5605), .B(n5604), .ZN(n6133) );
  AOI22_X1 U6736 ( .A1(n5613), .A2(DATAI_13_), .B1(n5612), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5606) );
  OAI21_X1 U6737 ( .B1(n6133), .B2(n5591), .A(n5606), .ZN(U2878) );
  AOI22_X1 U6738 ( .A1(n5613), .A2(DATAI_12_), .B1(n5612), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5607) );
  OAI21_X1 U6739 ( .B1(n5608), .B2(n5591), .A(n5607), .ZN(U2879) );
  AOI22_X1 U6740 ( .A1(n5613), .A2(DATAI_11_), .B1(n5612), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5609) );
  OAI21_X1 U6741 ( .B1(n5776), .B2(n5591), .A(n5609), .ZN(U2880) );
  AOI22_X1 U6742 ( .A1(n5613), .A2(DATAI_10_), .B1(n5612), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5610) );
  OAI21_X1 U6743 ( .B1(n6887), .B2(n5591), .A(n5610), .ZN(U2881) );
  AOI22_X1 U6744 ( .A1(n5613), .A2(DATAI_9_), .B1(n5612), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5611) );
  OAI21_X1 U6745 ( .B1(n5796), .B2(n5591), .A(n5611), .ZN(U2882) );
  AOI22_X1 U6746 ( .A1(n5613), .A2(DATAI_8_), .B1(n5612), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5614) );
  OAI21_X1 U6747 ( .B1(n5615), .B2(n5591), .A(n5614), .ZN(U2883) );
  NAND2_X1 U6748 ( .A1(n5617), .A2(n5616), .ZN(n5618) );
  XNOR2_X1 U6749 ( .A(n5618), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5815)
         );
  NOR2_X1 U6750 ( .A1(n3820), .A2(n6695), .ZN(n5806) );
  AOI21_X1 U6751 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5806), 
        .ZN(n5619) );
  OAI21_X1 U6752 ( .B1(n5620), .B2(n6341), .A(n5619), .ZN(n5621) );
  OAI21_X1 U6753 ( .B1(n5815), .B2(n6101), .A(n5623), .ZN(U2957) );
  INV_X1 U6754 ( .A(n5643), .ZN(n5632) );
  NAND3_X1 U6755 ( .A1(n5632), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5760), .ZN(n5624) );
  NOR2_X1 U6756 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5835) );
  NAND3_X1 U6757 ( .A1(n5653), .A2(n5662), .A3(n5835), .ZN(n5633) );
  AOI22_X1 U6758 ( .A1(n5624), .A2(n5633), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5641), .ZN(n5625) );
  XNOR2_X1 U6759 ( .A(n5625), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5823)
         );
  INV_X1 U6760 ( .A(n5626), .ZN(n5630) );
  INV_X1 U6761 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6873) );
  NOR2_X1 U6762 ( .A1(n3820), .A2(n6873), .ZN(n5819) );
  AOI21_X1 U6763 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5819), 
        .ZN(n5627) );
  OAI21_X1 U6764 ( .B1(n5628), .B2(n6341), .A(n5627), .ZN(n5629) );
  OAI21_X1 U6765 ( .B1(n6101), .B2(n5823), .A(n5631), .ZN(U2958) );
  NAND3_X1 U6766 ( .A1(n5632), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5760), .ZN(n5634) );
  NAND2_X1 U6767 ( .A1(n5634), .A2(n5633), .ZN(n5635) );
  XNOR2_X1 U6768 ( .A(n5635), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5824)
         );
  NOR2_X1 U6769 ( .A1(n3820), .A2(n6689), .ZN(n5825) );
  AOI21_X1 U6770 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5825), 
        .ZN(n5636) );
  OAI21_X1 U6771 ( .B1(n5637), .B2(n6341), .A(n5636), .ZN(n5638) );
  AOI21_X1 U6772 ( .B1(n5639), .B2(n5804), .A(n5638), .ZN(n5640) );
  OAI21_X1 U6773 ( .B1(n5824), .B2(n6101), .A(n5640), .ZN(U2959) );
  XNOR2_X1 U6774 ( .A(n5789), .B(n5641), .ZN(n5642) );
  XNOR2_X1 U6775 ( .A(n5643), .B(n5642), .ZN(n5843) );
  INV_X1 U6776 ( .A(n5644), .ZN(n5647) );
  INV_X1 U6777 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5645) );
  NOR2_X1 U6778 ( .A1(n3820), .A2(n5645), .ZN(n5839) );
  AOI21_X1 U6779 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5839), 
        .ZN(n5646) );
  OAI21_X1 U6780 ( .B1(n5647), .B2(n6341), .A(n5646), .ZN(n5648) );
  AOI21_X1 U6781 ( .B1(n5649), .B2(n5804), .A(n5648), .ZN(n5650) );
  OAI21_X1 U6782 ( .B1(n6101), .B2(n5843), .A(n5650), .ZN(U2960) );
  OAI21_X1 U6783 ( .B1(n5653), .B2(n5652), .A(n5651), .ZN(n5654) );
  INV_X1 U6784 ( .A(n5654), .ZN(n5853) );
  INV_X1 U6785 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6687) );
  NOR2_X1 U6786 ( .A1(n3820), .A2(n6687), .ZN(n5846) );
  AOI21_X1 U6787 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5846), 
        .ZN(n5655) );
  OAI21_X1 U6788 ( .B1(n5656), .B2(n6341), .A(n5655), .ZN(n5657) );
  AOI21_X1 U6789 ( .B1(n5658), .B2(n5804), .A(n5657), .ZN(n5659) );
  OAI21_X1 U6790 ( .B1(n5853), .B2(n6101), .A(n5659), .ZN(U2961) );
  AOI21_X1 U6791 ( .B1(n5662), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5660), 
        .ZN(n5697) );
  XNOR2_X1 U6792 ( .A(n5757), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5698)
         );
  INV_X1 U6793 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5661) );
  AOI22_X2 U6794 ( .A1(n5697), .A2(n5698), .B1(n5760), .B2(n5661), .ZN(n5690)
         );
  XNOR2_X1 U6795 ( .A(n5662), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5689)
         );
  NOR2_X1 U6796 ( .A1(n5757), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5680)
         );
  NAND3_X1 U6797 ( .A1(n5760), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5663) );
  INV_X1 U6798 ( .A(n5664), .ZN(n5668) );
  NOR2_X1 U6799 ( .A1(n3820), .A2(n6684), .ZN(n5858) );
  AOI21_X1 U6800 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5858), 
        .ZN(n5665) );
  OAI21_X1 U6801 ( .B1(n5666), .B2(n6341), .A(n5665), .ZN(n5667) );
  AOI21_X1 U6802 ( .B1(n5668), .B2(n5804), .A(n5667), .ZN(n5669) );
  OAI21_X1 U6803 ( .B1(n5861), .B2(n6101), .A(n5669), .ZN(U2962) );
  NAND2_X1 U6804 ( .A1(n5757), .A2(n5854), .ZN(n5671) );
  OAI21_X1 U6805 ( .B1(n5705), .B2(n5671), .A(n5670), .ZN(n5672) );
  XNOR2_X1 U6806 ( .A(n5672), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5869)
         );
  INV_X1 U6807 ( .A(n5673), .ZN(n5678) );
  NOR2_X1 U6808 ( .A1(n3820), .A2(n5674), .ZN(n5862) );
  AOI21_X1 U6809 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5862), 
        .ZN(n5675) );
  OAI21_X1 U6810 ( .B1(n5676), .B2(n6341), .A(n5675), .ZN(n5677) );
  AOI21_X1 U6811 ( .B1(n5678), .B2(n5804), .A(n5677), .ZN(n5679) );
  OAI21_X1 U6812 ( .B1(n5869), .B2(n6101), .A(n5679), .ZN(U2963) );
  AOI21_X1 U6813 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5757), .A(n5680), 
        .ZN(n5681) );
  XNOR2_X1 U6814 ( .A(n3145), .B(n5681), .ZN(n5879) );
  NAND2_X1 U6815 ( .A1(n6368), .A2(REIP_REG_22__SCAN_IN), .ZN(n5870) );
  OAI21_X1 U6816 ( .B1(n5784), .B2(n5682), .A(n5870), .ZN(n5685) );
  NOR2_X1 U6817 ( .A1(n5683), .A2(n5797), .ZN(n5684) );
  AOI211_X1 U6818 ( .C1(n5787), .C2(n5686), .A(n5685), .B(n5684), .ZN(n5687)
         );
  OAI21_X1 U6819 ( .B1(n5879), .B2(n6101), .A(n5687), .ZN(U2964) );
  AOI21_X1 U6820 ( .B1(n5690), .B2(n5689), .A(n5688), .ZN(n5887) );
  NOR2_X1 U6821 ( .A1(n3820), .A2(n5691), .ZN(n5880) );
  AOI21_X1 U6822 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5880), 
        .ZN(n5692) );
  OAI21_X1 U6823 ( .B1(n5693), .B2(n6341), .A(n5692), .ZN(n5694) );
  AOI21_X1 U6824 ( .B1(n5695), .B2(n5804), .A(n5694), .ZN(n5696) );
  OAI21_X1 U6825 ( .B1(n5887), .B2(n6101), .A(n5696), .ZN(U2965) );
  XOR2_X1 U6826 ( .A(n5698), .B(n5697), .Z(n5902) );
  NAND2_X1 U6827 ( .A1(n5699), .A2(n5787), .ZN(n5700) );
  NAND2_X1 U6828 ( .A1(n6368), .A2(REIP_REG_20__SCAN_IN), .ZN(n5894) );
  OAI211_X1 U6829 ( .C1(n5784), .C2(n3074), .A(n5700), .B(n5894), .ZN(n5701)
         );
  AOI21_X1 U6830 ( .B1(n5702), .B2(n5804), .A(n5701), .ZN(n5703) );
  OAI21_X1 U6831 ( .B1(n5902), .B2(n6101), .A(n5703), .ZN(U2966) );
  XNOR2_X1 U6832 ( .A(n5757), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5704)
         );
  XNOR2_X1 U6833 ( .A(n5705), .B(n5704), .ZN(n5903) );
  NAND2_X1 U6834 ( .A1(n5903), .A2(n6336), .ZN(n5709) );
  NOR2_X1 U6835 ( .A1(n3820), .A2(n6679), .ZN(n5905) );
  NOR2_X1 U6836 ( .A1(n6341), .A2(n5706), .ZN(n5707) );
  AOI211_X1 U6837 ( .C1(n6329), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5905), 
        .B(n5707), .ZN(n5708) );
  OAI211_X1 U6838 ( .C1(n5797), .C2(n5710), .A(n5709), .B(n5708), .ZN(U2967)
         );
  NOR3_X1 U6839 ( .A1(n5711), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5757), 
        .ZN(n5720) );
  NOR3_X1 U6840 ( .A1(n5662), .A2(n5927), .A3(n5944), .ZN(n5712) );
  AOI22_X1 U6841 ( .A1(n5720), .A2(n5927), .B1(n5712), .B2(n5711), .ZN(n5713)
         );
  XNOR2_X1 U6842 ( .A(n5713), .B(n5917), .ZN(n5921) );
  INV_X1 U6843 ( .A(n5714), .ZN(n5716) );
  NOR2_X1 U6844 ( .A1(n3820), .A2(n6677), .ZN(n5913) );
  AOI21_X1 U6845 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5913), 
        .ZN(n5715) );
  OAI21_X1 U6846 ( .B1(n6341), .B2(n5716), .A(n5715), .ZN(n5717) );
  AOI21_X1 U6847 ( .B1(n5718), .B2(n5804), .A(n5717), .ZN(n5719) );
  OAI21_X1 U6848 ( .B1(n5921), .B2(n6101), .A(n5719), .ZN(U2968) );
  NOR2_X1 U6849 ( .A1(n5662), .A2(n5944), .ZN(n5721) );
  AOI21_X1 U6850 ( .B1(n5721), .B2(n5711), .A(n5720), .ZN(n5722) );
  XNOR2_X1 U6851 ( .A(n5722), .B(n5927), .ZN(n5930) );
  INV_X1 U6852 ( .A(n5723), .ZN(n5727) );
  NAND2_X1 U6853 ( .A1(n6368), .A2(REIP_REG_17__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U6854 ( .A1(n6329), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5724)
         );
  OAI211_X1 U6855 ( .C1(n6341), .C2(n5725), .A(n5923), .B(n5724), .ZN(n5726)
         );
  AOI21_X1 U6856 ( .B1(n5727), .B2(n5804), .A(n5726), .ZN(n5728) );
  OAI21_X1 U6857 ( .B1(n5930), .B2(n6101), .A(n5728), .ZN(U2969) );
  XNOR2_X1 U6858 ( .A(n5789), .B(n5944), .ZN(n5729) );
  XNOR2_X1 U6859 ( .A(n5711), .B(n5729), .ZN(n5937) );
  NAND2_X1 U6860 ( .A1(n5937), .A2(n6336), .ZN(n5733) );
  NOR2_X1 U6861 ( .A1(n3820), .A2(n6672), .ZN(n5940) );
  NOR2_X1 U6862 ( .A1(n6341), .A2(n5730), .ZN(n5731) );
  AOI211_X1 U6863 ( .C1(n6329), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5940), 
        .B(n5731), .ZN(n5732) );
  OAI211_X1 U6864 ( .C1(n5797), .C2(n5734), .A(n5733), .B(n5732), .ZN(U2970)
         );
  XNOR2_X1 U6865 ( .A(n5789), .B(n5950), .ZN(n5735) );
  XNOR2_X1 U6866 ( .A(n5736), .B(n5735), .ZN(n5954) );
  NOR2_X1 U6867 ( .A1(n3820), .A2(n6670), .ZN(n5947) );
  AOI21_X1 U6868 ( .B1(n6329), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5947), 
        .ZN(n5737) );
  OAI21_X1 U6869 ( .B1(n6341), .B2(n5738), .A(n5737), .ZN(n5739) );
  AOI21_X1 U6870 ( .B1(n5740), .B2(n5804), .A(n5739), .ZN(n5741) );
  OAI21_X1 U6871 ( .B1(n6101), .B2(n5954), .A(n5741), .ZN(U2971) );
  INV_X1 U6872 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5742) );
  NOR2_X1 U6873 ( .A1(n3820), .A2(n5742), .ZN(n5963) );
  NOR2_X1 U6874 ( .A1(n6341), .A2(n6124), .ZN(n5743) );
  AOI211_X1 U6875 ( .C1(n6329), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5963), 
        .B(n5743), .ZN(n5750) );
  AND2_X1 U6876 ( .A1(n5745), .A2(n5744), .ZN(n5754) );
  XNOR2_X1 U6877 ( .A(n5789), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5753)
         );
  NAND2_X1 U6878 ( .A1(n5754), .A2(n5753), .ZN(n5752) );
  NAND2_X1 U6879 ( .A1(n5752), .A2(n5746), .ZN(n5748) );
  XNOR2_X1 U6880 ( .A(n5789), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5747)
         );
  XNOR2_X1 U6881 ( .A(n5748), .B(n5747), .ZN(n5959) );
  NAND2_X1 U6882 ( .A1(n5959), .A2(n6336), .ZN(n5749) );
  OAI211_X1 U6883 ( .C1(n6123), .C2(n5797), .A(n5750), .B(n5749), .ZN(U2972)
         );
  NAND2_X1 U6884 ( .A1(n6368), .A2(REIP_REG_13__SCAN_IN), .ZN(n5977) );
  OAI21_X1 U6885 ( .B1(n5784), .B2(n6131), .A(n5977), .ZN(n5751) );
  AOI21_X1 U6886 ( .B1(n5787), .B2(n6134), .A(n5751), .ZN(n5756) );
  OAI21_X1 U6887 ( .B1(n5754), .B2(n5753), .A(n5752), .ZN(n5969) );
  NAND2_X1 U6888 ( .A1(n5969), .A2(n6336), .ZN(n5755) );
  OAI211_X1 U6889 ( .C1(n6133), .C2(n5797), .A(n5756), .B(n5755), .ZN(U2973)
         );
  NAND2_X1 U6890 ( .A1(n2991), .A2(n5777), .ZN(n5770) );
  NOR2_X1 U6891 ( .A1(n5757), .A2(n5983), .ZN(n5769) );
  AOI21_X1 U6892 ( .B1(n5770), .B2(n5767), .A(n5769), .ZN(n5762) );
  OAI21_X1 U6893 ( .B1(n5760), .B2(n5759), .A(n5758), .ZN(n5761) );
  XNOR2_X1 U6894 ( .A(n5762), .B(n5761), .ZN(n5990) );
  NAND2_X1 U6895 ( .A1(n6368), .A2(REIP_REG_12__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U6896 ( .A1(n6329), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5763)
         );
  OAI211_X1 U6897 ( .C1(n6341), .C2(n5764), .A(n5986), .B(n5763), .ZN(n5765)
         );
  AOI21_X1 U6898 ( .B1(n6142), .B2(n5804), .A(n5765), .ZN(n5766) );
  OAI21_X1 U6899 ( .B1(n5990), .B2(n6101), .A(n5766), .ZN(U2974) );
  INV_X1 U6900 ( .A(n5767), .ZN(n5768) );
  NOR2_X1 U6901 ( .A1(n5769), .A2(n5768), .ZN(n5771) );
  XOR2_X1 U6902 ( .A(n5771), .B(n5770), .Z(n6345) );
  NAND2_X1 U6903 ( .A1(n6345), .A2(n6336), .ZN(n5775) );
  NOR2_X1 U6904 ( .A1(n3820), .A2(n5460), .ZN(n6342) );
  NOR2_X1 U6905 ( .A1(n6341), .A2(n5772), .ZN(n5773) );
  AOI211_X1 U6906 ( .C1(n6329), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6342), 
        .B(n5773), .ZN(n5774) );
  OAI211_X1 U6907 ( .C1(n5797), .C2(n5776), .A(n5775), .B(n5774), .ZN(U2975)
         );
  INV_X1 U6908 ( .A(n5777), .ZN(n5779) );
  NOR2_X1 U6909 ( .A1(n5779), .A2(n5778), .ZN(n5781) );
  XOR2_X1 U6910 ( .A(n5781), .B(n5780), .Z(n6004) );
  INV_X1 U6911 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5783) );
  INV_X1 U6912 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5782) );
  OAI22_X1 U6913 ( .A1(n5784), .A2(n5783), .B1(n3820), .B2(n5782), .ZN(n5786)
         );
  NOR2_X1 U6914 ( .A1(n6887), .A2(n5797), .ZN(n5785) );
  AOI211_X1 U6915 ( .C1(n5787), .C2(n6888), .A(n5786), .B(n5785), .ZN(n5788)
         );
  OAI21_X1 U6916 ( .B1(n6004), .B2(n6101), .A(n5788), .ZN(U2976) );
  XNOR2_X1 U6917 ( .A(n5789), .B(n6841), .ZN(n5790) );
  XNOR2_X1 U6918 ( .A(n5791), .B(n5790), .ZN(n6351) );
  NAND2_X1 U6919 ( .A1(n6351), .A2(n6336), .ZN(n5795) );
  NOR2_X1 U6920 ( .A1(n3820), .A2(n6893), .ZN(n6349) );
  NOR2_X1 U6921 ( .A1(n6341), .A2(n5792), .ZN(n5793) );
  AOI211_X1 U6922 ( .C1(n6329), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6349), 
        .B(n5793), .ZN(n5794) );
  OAI211_X1 U6923 ( .C1(n5797), .C2(n5796), .A(n5795), .B(n5794), .ZN(U2977)
         );
  XNOR2_X1 U6924 ( .A(n5798), .B(n5799), .ZN(n6014) );
  INV_X1 U6925 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5800) );
  OR2_X1 U6926 ( .A1(n3820), .A2(n5800), .ZN(n6010) );
  NAND2_X1 U6927 ( .A1(n6329), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5801)
         );
  OAI211_X1 U6928 ( .C1(n6341), .C2(n5802), .A(n6010), .B(n5801), .ZN(n5803)
         );
  AOI21_X1 U6929 ( .B1(n6158), .B2(n5804), .A(n5803), .ZN(n5805) );
  OAI21_X1 U6930 ( .B1(n6101), .B2(n6014), .A(n5805), .ZN(U2978) );
  INV_X1 U6931 ( .A(n5806), .ZN(n5810) );
  NAND3_X1 U6932 ( .A1(n5829), .A2(n5808), .A3(n5807), .ZN(n5809) );
  OAI211_X1 U6933 ( .C1(n5811), .C2(n6387), .A(n5810), .B(n5809), .ZN(n5812)
         );
  AOI21_X1 U6934 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5813), .A(n5812), 
        .ZN(n5814) );
  OAI21_X1 U6935 ( .B1(n5815), .B2(n6015), .A(n5814), .ZN(U2989) );
  AND3_X1 U6936 ( .A1(n5829), .A2(n5817), .A3(n5816), .ZN(n5818) );
  AOI211_X1 U6937 ( .C1(n6359), .C2(n5820), .A(n5819), .B(n5818), .ZN(n5822)
         );
  NAND2_X1 U6938 ( .A1(n5827), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5821) );
  OAI211_X1 U6939 ( .C1(n5823), .C2(n6015), .A(n5822), .B(n5821), .ZN(U2990)
         );
  OR2_X1 U6940 ( .A1(n5824), .A2(n6015), .ZN(n5833) );
  AOI21_X1 U6941 ( .B1(n5826), .B2(n6359), .A(n5825), .ZN(n5832) );
  NAND2_X1 U6942 ( .A1(n5827), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U6943 ( .A1(n5829), .A2(n5828), .ZN(n5830) );
  NAND4_X1 U6944 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(U2991)
         );
  INV_X1 U6945 ( .A(n5834), .ZN(n5840) );
  INV_X1 U6946 ( .A(n5845), .ZN(n5837) );
  NOR3_X1 U6947 ( .A1(n5837), .A2(n5836), .A3(n5835), .ZN(n5838) );
  AOI211_X1 U6948 ( .C1(n6359), .C2(n5840), .A(n5839), .B(n5838), .ZN(n5842)
         );
  INV_X1 U6949 ( .A(n5855), .ZN(n5851) );
  NAND2_X1 U6950 ( .A1(n5851), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5841) );
  OAI211_X1 U6951 ( .C1(n5843), .C2(n6015), .A(n5842), .B(n5841), .ZN(U2992)
         );
  INV_X1 U6952 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U6953 ( .A1(n5845), .A2(n5844), .ZN(n5848) );
  INV_X1 U6954 ( .A(n5846), .ZN(n5847) );
  OAI211_X1 U6955 ( .C1(n6387), .C2(n5849), .A(n5848), .B(n5847), .ZN(n5850)
         );
  AOI21_X1 U6956 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5851), .A(n5850), 
        .ZN(n5852) );
  OAI21_X1 U6957 ( .B1(n5853), .B2(n6015), .A(n5852), .ZN(U2993) );
  INV_X1 U6958 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U6959 ( .A1(n5908), .A2(n5854), .ZN(n5865) );
  AOI211_X1 U6960 ( .C1(n6853), .C2(n5865), .A(n5856), .B(n5855), .ZN(n5857)
         );
  AOI211_X1 U6961 ( .C1(n6359), .C2(n5859), .A(n5858), .B(n5857), .ZN(n5860)
         );
  OAI21_X1 U6962 ( .B1(n5861), .B2(n6015), .A(n5860), .ZN(U2994) );
  AOI21_X1 U6963 ( .B1(n5863), .B2(n6359), .A(n5862), .ZN(n5864) );
  OAI21_X1 U6964 ( .B1(n5865), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5864), 
        .ZN(n5866) );
  AOI21_X1 U6965 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5867), .A(n5866), 
        .ZN(n5868) );
  OAI21_X1 U6966 ( .B1(n5869), .B2(n6015), .A(n5868), .ZN(U2995) );
  OAI21_X1 U6967 ( .B1(n5871), .B2(n6387), .A(n5870), .ZN(n5877) );
  INV_X1 U6968 ( .A(n5872), .ZN(n5897) );
  NAND2_X1 U6969 ( .A1(n5908), .A2(n5897), .ZN(n5883) );
  INV_X1 U6970 ( .A(n5873), .ZN(n5875) );
  NOR3_X1 U6971 ( .A1(n5883), .A2(n5875), .A3(n5874), .ZN(n5876) );
  AOI211_X1 U6972 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5885), .A(n5877), .B(n5876), .ZN(n5878) );
  OAI21_X1 U6973 ( .B1(n5879), .B2(n6015), .A(n5878), .ZN(U2996) );
  AOI21_X1 U6974 ( .B1(n5881), .B2(n6359), .A(n5880), .ZN(n5882) );
  OAI21_X1 U6975 ( .B1(n5883), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5882), 
        .ZN(n5884) );
  AOI21_X1 U6976 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5885), .A(n5884), 
        .ZN(n5886) );
  OAI21_X1 U6977 ( .B1(n5887), .B2(n6015), .A(n5886), .ZN(U2997) );
  NOR2_X1 U6978 ( .A1(n5888), .A2(n5927), .ZN(n5889) );
  OR2_X1 U6979 ( .A1(n5991), .A2(n5889), .ZN(n5892) );
  INV_X1 U6980 ( .A(n5890), .ZN(n5891) );
  NAND2_X1 U6981 ( .A1(n5892), .A2(n5891), .ZN(n5922) );
  AND2_X1 U6982 ( .A1(n6367), .A2(n5927), .ZN(n5893) );
  NOR2_X1 U6983 ( .A1(n5922), .A2(n5893), .ZN(n5918) );
  OAI21_X1 U6984 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5996), .A(n5918), 
        .ZN(n5909) );
  OAI21_X1 U6985 ( .B1(n5895), .B2(n6387), .A(n5894), .ZN(n5900) );
  INV_X1 U6986 ( .A(n5908), .ZN(n5898) );
  NOR3_X1 U6987 ( .A1(n5898), .A2(n5897), .A3(n5896), .ZN(n5899) );
  AOI211_X1 U6988 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n5909), .A(n5900), .B(n5899), .ZN(n5901) );
  OAI21_X1 U6989 ( .B1(n5902), .B2(n6015), .A(n5901), .ZN(U2998) );
  INV_X1 U6990 ( .A(n5903), .ZN(n5912) );
  NOR2_X1 U6991 ( .A1(n5904), .A2(n6387), .ZN(n5906) );
  AOI211_X1 U6992 ( .C1(n5908), .C2(n5907), .A(n5906), .B(n5905), .ZN(n5911)
         );
  NAND2_X1 U6993 ( .A1(n5909), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5910) );
  OAI211_X1 U6994 ( .C1(n5912), .C2(n6015), .A(n5911), .B(n5910), .ZN(U2999)
         );
  NAND3_X1 U6995 ( .A1(n5928), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5917), .ZN(n5916) );
  AOI21_X1 U6996 ( .B1(n5914), .B2(n6359), .A(n5913), .ZN(n5915) );
  OAI211_X1 U6997 ( .C1(n5918), .C2(n5917), .A(n5916), .B(n5915), .ZN(n5919)
         );
  INV_X1 U6998 ( .A(n5919), .ZN(n5920) );
  OAI21_X1 U6999 ( .B1(n5921), .B2(n6015), .A(n5920), .ZN(U3000) );
  NAND2_X1 U7000 ( .A1(n5922), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5924) );
  OAI211_X1 U7001 ( .C1(n6387), .C2(n5925), .A(n5924), .B(n5923), .ZN(n5926)
         );
  AOI21_X1 U7002 ( .B1(n5928), .B2(n5927), .A(n5926), .ZN(n5929) );
  OAI21_X1 U7003 ( .B1(n5930), .B2(n6015), .A(n5929), .ZN(U3001) );
  OR2_X1 U7004 ( .A1(n5991), .A2(n5931), .ZN(n5934) );
  NAND2_X1 U7005 ( .A1(n5995), .A2(n5932), .ZN(n5933) );
  NAND2_X1 U7006 ( .A1(n5934), .A2(n5933), .ZN(n6344) );
  AOI21_X1 U7007 ( .B1(n5936), .B2(n5935), .A(n6344), .ZN(n5951) );
  NAND2_X1 U7008 ( .A1(n5937), .A2(n6381), .ZN(n5943) );
  XNOR2_X1 U7009 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5938) );
  NOR2_X1 U7010 ( .A1(n5945), .A2(n5938), .ZN(n5939) );
  AOI211_X1 U7011 ( .C1(n6359), .C2(n5941), .A(n5940), .B(n5939), .ZN(n5942)
         );
  OAI211_X1 U7012 ( .C1(n5951), .C2(n5944), .A(n5943), .B(n5942), .ZN(U3002)
         );
  INV_X1 U7013 ( .A(n5945), .ZN(n5949) );
  NOR2_X1 U7014 ( .A1(n5946), .A2(n6387), .ZN(n5948) );
  AOI211_X1 U7015 ( .C1(n5949), .C2(n5950), .A(n5948), .B(n5947), .ZN(n5953)
         );
  OR2_X1 U7016 ( .A1(n5951), .A2(n5950), .ZN(n5952) );
  OAI211_X1 U7017 ( .C1(n5954), .C2(n6015), .A(n5953), .B(n5952), .ZN(U3003)
         );
  NOR2_X1 U7018 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5956), .ZN(n5980)
         );
  AOI21_X1 U7019 ( .B1(n5956), .B2(n5955), .A(n6344), .ZN(n5957) );
  OAI21_X1 U7020 ( .B1(n6392), .B2(n5960), .A(n5957), .ZN(n5975) );
  AOI21_X1 U7021 ( .B1(n5958), .B2(n5980), .A(n5975), .ZN(n5968) );
  NAND2_X1 U7022 ( .A1(n5959), .A2(n6381), .ZN(n5966) );
  INV_X1 U7023 ( .A(n6129), .ZN(n5964) );
  INV_X1 U7024 ( .A(n5960), .ZN(n5961) );
  NOR3_X1 U7025 ( .A1(n6348), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n5961), 
        .ZN(n5962) );
  AOI211_X1 U7026 ( .C1(n6359), .C2(n5964), .A(n5963), .B(n5962), .ZN(n5965)
         );
  OAI211_X1 U7027 ( .C1(n5968), .C2(n5967), .A(n5966), .B(n5965), .ZN(U3004)
         );
  INV_X1 U7028 ( .A(n5969), .ZN(n5982) );
  INV_X1 U7029 ( .A(n6348), .ZN(n5985) );
  INV_X1 U7030 ( .A(n5970), .ZN(n5971) );
  OAI21_X1 U7031 ( .B1(n5451), .B2(n5972), .A(n5971), .ZN(n5974) );
  AND2_X1 U7032 ( .A1(n5974), .A2(n5973), .ZN(n6231) );
  INV_X1 U7033 ( .A(n6231), .ZN(n5978) );
  NAND2_X1 U7034 ( .A1(n5975), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5976) );
  OAI211_X1 U7035 ( .C1(n5978), .C2(n6387), .A(n5977), .B(n5976), .ZN(n5979)
         );
  AOI21_X1 U7036 ( .B1(n5985), .B2(n5980), .A(n5979), .ZN(n5981) );
  OAI21_X1 U7037 ( .B1(n5982), .B2(n6015), .A(n5981), .ZN(U3005) );
  XNOR2_X1 U7038 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .B(n5983), .ZN(n5984)
         );
  NAND2_X1 U7039 ( .A1(n5985), .A2(n5984), .ZN(n5987) );
  OAI211_X1 U7040 ( .C1(n6143), .C2(n6387), .A(n5987), .B(n5986), .ZN(n5988)
         );
  AOI21_X1 U7041 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6344), .A(n5988), 
        .ZN(n5989) );
  OAI21_X1 U7042 ( .B1(n5990), .B2(n6015), .A(n5989), .ZN(U3006) );
  INV_X1 U7043 ( .A(n5991), .ZN(n5993) );
  AOI22_X1 U7044 ( .A1(n5995), .A2(n5994), .B1(n5993), .B2(n5992), .ZN(n6366)
         );
  OAI21_X1 U7045 ( .B1(n5996), .B2(n6005), .A(n6366), .ZN(n6352) );
  OAI22_X1 U7046 ( .A1(n6898), .A2(n6387), .B1(n5782), .B2(n3820), .ZN(n6002)
         );
  NAND2_X1 U7047 ( .A1(n5999), .A2(n5998), .ZN(n6362) );
  INV_X1 U7048 ( .A(n6362), .ZN(n6007) );
  NAND2_X1 U7049 ( .A1(n6005), .A2(n6007), .ZN(n6355) );
  AOI221_X1 U7050 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n6000), .C2(n6841), .A(n6355), 
        .ZN(n6001) );
  AOI211_X1 U7051 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6352), .A(n6002), .B(n6001), .ZN(n6003) );
  OAI21_X1 U7052 ( .B1(n6015), .B2(n6004), .A(n6003), .ZN(U3008) );
  INV_X1 U7053 ( .A(n6366), .ZN(n6012) );
  AOI21_X1 U7054 ( .B1(n6006), .B2(n6365), .A(n6005), .ZN(n6008) );
  NAND2_X1 U7055 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  OAI211_X1 U7056 ( .C1(n6155), .C2(n6387), .A(n6010), .B(n6009), .ZN(n6011)
         );
  AOI21_X1 U7057 ( .B1(n6012), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6011), 
        .ZN(n6013) );
  OAI21_X1 U7058 ( .B1(n6015), .B2(n6014), .A(n6013), .ZN(U3010) );
  AND2_X1 U7059 ( .A1(n6050), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6030) );
  OAI222_X1 U7060 ( .A1(n6017), .A2(n6016), .B1(n6515), .B2(n6030), .C1(n4587), 
        .C2(n6578), .ZN(n6020) );
  OAI21_X1 U7061 ( .B1(n6017), .B2(FLUSH_REG_SCAN_IN), .A(n6643), .ZN(n6019)
         );
  NAND2_X1 U7062 ( .A1(n6019), .A2(n6018), .ZN(n6394) );
  MUX2_X1 U7063 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n6020), .S(n6394), 
        .Z(U3465) );
  OAI211_X1 U7064 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6021), .A(n6513), .B(
        n6437), .ZN(n6022) );
  OAI21_X1 U7065 ( .B1(n6030), .B2(n4583), .A(n6022), .ZN(n6023) );
  MUX2_X1 U7066 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n6023), .S(n6394), 
        .Z(U3464) );
  XNOR2_X1 U7067 ( .A(n6513), .B(n6024), .ZN(n6025) );
  OAI22_X1 U7068 ( .A1(n6025), .A2(n6578), .B1(n6030), .B2(n4503), .ZN(n6026)
         );
  MUX2_X1 U7069 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n6026), .S(n6394), 
        .Z(U3463) );
  INV_X1 U7070 ( .A(n4858), .ZN(n6032) );
  INV_X1 U7071 ( .A(n6514), .ZN(n6028) );
  NOR3_X1 U7072 ( .A1(n6029), .A2(n6028), .A3(n6027), .ZN(n6031) );
  OAI222_X1 U7073 ( .A1(n6033), .A2(n6032), .B1(n6578), .B2(n6031), .C1(n6030), 
        .C2(n6482), .ZN(n6034) );
  MUX2_X1 U7074 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6034), .S(n6394), 
        .Z(U3462) );
  INV_X1 U7075 ( .A(n6035), .ZN(n6039) );
  OAI22_X1 U7076 ( .A1(n6039), .A2(n6038), .B1(n6037), .B2(n6036), .ZN(n6041)
         );
  MUX2_X1 U7077 ( .A(n6041), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6040), 
        .Z(U3456) );
  INV_X1 U7078 ( .A(n6042), .ZN(n6043) );
  INV_X1 U7079 ( .A(n6567), .ZN(n6044) );
  OAI21_X1 U7080 ( .B1(n6083), .B2(n6044), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6045) );
  NAND2_X1 U7081 ( .A1(n6045), .A2(n6437), .ZN(n6057) );
  INV_X1 U7082 ( .A(n6057), .ZN(n6052) );
  INV_X1 U7083 ( .A(n6046), .ZN(n6047) );
  NAND2_X1 U7084 ( .A1(n6047), .A2(n4581), .ZN(n6516) );
  INV_X1 U7085 ( .A(n6522), .ZN(n6048) );
  NOR3_X1 U7086 ( .A1(n6048), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6519), 
        .ZN(n6053) );
  OAI211_X1 U7087 ( .C1(n6053), .C2(n6050), .A(n6049), .B(n6568), .ZN(n6051)
         );
  INV_X1 U7088 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6060) );
  INV_X1 U7089 ( .A(n6053), .ZN(n6092) );
  OAI22_X1 U7090 ( .A1(n6567), .A2(n6528), .B1(n6092), .B2(n6511), .ZN(n6054)
         );
  AOI21_X1 U7091 ( .B1(n6083), .B2(n6470), .A(n6054), .ZN(n6059) );
  NAND2_X1 U7092 ( .A1(n6095), .A2(n6577), .ZN(n6058) );
  OAI211_X1 U7093 ( .C1(n6098), .C2(n6060), .A(n6059), .B(n6058), .ZN(U3100)
         );
  INV_X1 U7094 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6065) );
  OAI22_X1 U7095 ( .A1(n6567), .A2(n6530), .B1(n6092), .B2(n6529), .ZN(n6061)
         );
  AOI21_X1 U7096 ( .B1(n6083), .B2(n6062), .A(n6061), .ZN(n6064) );
  NAND2_X1 U7097 ( .A1(n6095), .A2(n6594), .ZN(n6063) );
  OAI211_X1 U7098 ( .C1(n6098), .C2(n6065), .A(n6064), .B(n6063), .ZN(U3101)
         );
  INV_X1 U7099 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6070) );
  OAI22_X1 U7100 ( .A1(n6567), .A2(n6535), .B1(n6092), .B2(n6534), .ZN(n6066)
         );
  AOI21_X1 U7101 ( .B1(n6083), .B2(n6067), .A(n6066), .ZN(n6069) );
  NAND2_X1 U7102 ( .A1(n6095), .A2(n6600), .ZN(n6068) );
  OAI211_X1 U7103 ( .C1(n6098), .C2(n6070), .A(n6069), .B(n6068), .ZN(U3102)
         );
  INV_X1 U7104 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6075) );
  OAI22_X1 U7105 ( .A1(n6567), .A2(n6540), .B1(n6092), .B2(n6539), .ZN(n6071)
         );
  AOI21_X1 U7106 ( .B1(n6083), .B2(n6072), .A(n6071), .ZN(n6074) );
  NAND2_X1 U7107 ( .A1(n6095), .A2(n6606), .ZN(n6073) );
  OAI211_X1 U7108 ( .C1(n6098), .C2(n6075), .A(n6074), .B(n6073), .ZN(U3103)
         );
  INV_X1 U7109 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6080) );
  OAI22_X1 U7110 ( .A1(n6567), .A2(n6545), .B1(n6092), .B2(n6544), .ZN(n6076)
         );
  AOI21_X1 U7111 ( .B1(n6083), .B2(n6077), .A(n6076), .ZN(n6079) );
  NAND2_X1 U7112 ( .A1(n6095), .A2(n6612), .ZN(n6078) );
  OAI211_X1 U7113 ( .C1(n6098), .C2(n6080), .A(n6079), .B(n6078), .ZN(U3104)
         );
  INV_X1 U7114 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6086) );
  OAI22_X1 U7115 ( .A1(n6567), .A2(n6553), .B1(n6092), .B2(n6549), .ZN(n6081)
         );
  AOI21_X1 U7116 ( .B1(n6083), .B2(n6082), .A(n6081), .ZN(n6085) );
  NAND2_X1 U7117 ( .A1(n6095), .A2(n6618), .ZN(n6084) );
  OAI211_X1 U7118 ( .C1(n6098), .C2(n6086), .A(n6085), .B(n6084), .ZN(U3105)
         );
  INV_X1 U7119 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6090) );
  NOR2_X1 U7120 ( .A1(n6091), .A2(n6628), .ZN(n6088) );
  OAI22_X1 U7121 ( .A1(n6567), .A2(n6558), .B1(n6092), .B2(n6554), .ZN(n6087)
         );
  AOI211_X1 U7122 ( .C1(n6095), .C2(n6624), .A(n6088), .B(n6087), .ZN(n6089)
         );
  OAI21_X1 U7123 ( .B1(n6098), .B2(n6090), .A(n6089), .ZN(U3106) );
  INV_X1 U7124 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6097) );
  NOR2_X1 U7125 ( .A1(n6091), .A2(n6639), .ZN(n6094) );
  OAI22_X1 U7126 ( .A1(n6567), .A2(n6561), .B1(n6092), .B2(n6560), .ZN(n6093)
         );
  AOI211_X1 U7127 ( .C1(n6095), .C2(n6631), .A(n6094), .B(n6093), .ZN(n6096)
         );
  OAI21_X1 U7128 ( .B1(n6098), .B2(n6097), .A(n6096), .ZN(U3107) );
  MUX2_X1 U7129 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6099), .Z(U3447) );
  MUX2_X1 U7130 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6099), .Z(U3446) );
  MUX2_X1 U7131 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6099), .Z(U3445) );
  INV_X1 U7132 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n6821) );
  NOR2_X1 U7133 ( .A1(n6821), .A2(n6253), .ZN(U2892) );
  OAI21_X1 U7134 ( .B1(n6100), .B2(BS16_N), .A(n6702), .ZN(n6701) );
  OAI21_X1 U7135 ( .B1(n6702), .B2(n6435), .A(n6701), .ZN(U2792) );
  OAI21_X1 U7136 ( .B1(n6103), .B2(n6102), .A(n6101), .ZN(U2793) );
  NOR2_X1 U7137 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6733) );
  AOI211_X1 U7138 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_10__SCAN_IN), .B(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n6104) );
  INV_X1 U7139 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6868) );
  INV_X1 U7140 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6804) );
  AND4_X1 U7141 ( .A1(n6733), .A2(n6104), .A3(n6868), .A4(n6804), .ZN(n6112)
         );
  NOR4_X1 U7142 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n6111) );
  NOR4_X1 U7143 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6110) );
  NOR4_X1 U7144 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n6108) );
  NOR4_X1 U7145 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6107) );
  NOR4_X1 U7146 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6106) );
  NOR4_X1 U7147 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6105) );
  AND4_X1 U7148 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n6109)
         );
  NAND4_X1 U7149 ( .A1(n6112), .A2(n6111), .A3(n6110), .A4(n6109), .ZN(n6709)
         );
  INV_X1 U7150 ( .A(n6709), .ZN(n6705) );
  INV_X1 U7151 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6113) );
  INV_X1 U7152 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6865) );
  NAND2_X1 U7153 ( .A1(n6705), .A2(n6865), .ZN(n6116) );
  NOR2_X1 U7154 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(n6116), .ZN(n6703) );
  NAND2_X1 U7155 ( .A1(n6703), .A2(n4519), .ZN(n6114) );
  OAI221_X1 U7156 ( .B1(n6705), .B2(n6113), .C1(n6709), .C2(n4559), .A(n6114), 
        .ZN(U2794) );
  NAND2_X1 U7157 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(n6709), .ZN(n6115) );
  OAI211_X1 U7158 ( .C1(REIP_REG_1__SCAN_IN), .C2(n6116), .A(n6115), .B(n6114), 
        .ZN(U2795) );
  INV_X1 U7159 ( .A(n6117), .ZN(n6122) );
  AOI22_X1 U7160 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6895), .B1(
        REIP_REG_14__SCAN_IN), .B2(n6118), .ZN(n6119) );
  OAI211_X1 U7161 ( .C1(n6186), .C2(n3069), .A(n6119), .B(n6896), .ZN(n6120)
         );
  AOI21_X1 U7162 ( .B1(n6122), .B2(n6121), .A(n6120), .ZN(n6128) );
  INV_X1 U7163 ( .A(n6123), .ZN(n6126) );
  INV_X1 U7164 ( .A(n6124), .ZN(n6125) );
  AOI22_X1 U7165 ( .A1(n6126), .A2(n6890), .B1(n6125), .B2(n6889), .ZN(n6127)
         );
  OAI211_X1 U7166 ( .C1(n6899), .C2(n6129), .A(n6128), .B(n6127), .ZN(U2813)
         );
  AOI22_X1 U7167 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6895), .B1(n6220), .B2(n6231), .ZN(n6140) );
  OR4_X1 U7168 ( .A1(n6892), .A2(REIP_REG_13__SCAN_IN), .A3(n6135), .A4(n6148), 
        .ZN(n6130) );
  OAI211_X1 U7169 ( .C1(n6186), .C2(n6131), .A(n6130), .B(n6896), .ZN(n6132)
         );
  INV_X1 U7170 ( .A(n6132), .ZN(n6139) );
  INV_X1 U7171 ( .A(n6133), .ZN(n6234) );
  AOI22_X1 U7172 ( .A1(n6234), .A2(n6890), .B1(n6889), .B2(n6134), .ZN(n6138)
         );
  INV_X1 U7173 ( .A(n6149), .ZN(n6136) );
  NOR3_X1 U7174 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6135), .A3(n6892), .ZN(n6151) );
  OAI21_X1 U7175 ( .B1(n6136), .B2(n6151), .A(REIP_REG_13__SCAN_IN), .ZN(n6137) );
  NAND4_X1 U7176 ( .A1(n6140), .A2(n6139), .A3(n6138), .A4(n6137), .ZN(U2814)
         );
  AOI22_X1 U7177 ( .A1(n6142), .A2(n6890), .B1(n6889), .B2(n6141), .ZN(n6153)
         );
  INV_X1 U7178 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6148) );
  INV_X1 U7179 ( .A(n6143), .ZN(n6146) );
  OAI21_X1 U7180 ( .B1(n6186), .B2(n6144), .A(n6896), .ZN(n6145) );
  AOI21_X1 U7181 ( .B1(n6146), .B2(n6220), .A(n6145), .ZN(n6147) );
  OAI21_X1 U7182 ( .B1(n6149), .B2(n6148), .A(n6147), .ZN(n6150) );
  AOI211_X1 U7183 ( .C1(n6895), .C2(EBX_REG_12__SCAN_IN), .A(n6151), .B(n6150), 
        .ZN(n6152) );
  NAND2_X1 U7184 ( .A1(n6153), .A2(n6152), .ZN(U2815) );
  NOR2_X1 U7185 ( .A1(n6154), .A2(REIP_REG_8__SCAN_IN), .ZN(n6162) );
  OAI22_X1 U7186 ( .A1(n6899), .A2(n6155), .B1(n6755), .B2(n6186), .ZN(n6156)
         );
  AOI211_X1 U7187 ( .C1(n6895), .C2(EBX_REG_8__SCAN_IN), .A(n6188), .B(n6156), 
        .ZN(n6160) );
  AOI22_X1 U7188 ( .A1(n6890), .A2(n6158), .B1(n6889), .B2(n6157), .ZN(n6159)
         );
  OAI211_X1 U7189 ( .C1(n6162), .C2(n6161), .A(n6160), .B(n6159), .ZN(U2819)
         );
  NOR3_X1 U7190 ( .A1(n6190), .A2(REIP_REG_7__SCAN_IN), .A3(n6163), .ZN(n6168)
         );
  OAI21_X1 U7191 ( .B1(n6186), .B2(n3914), .A(n6896), .ZN(n6164) );
  AOI21_X1 U7192 ( .B1(n6895), .B2(EBX_REG_7__SCAN_IN), .A(n6164), .ZN(n6165)
         );
  OAI21_X1 U7193 ( .B1(n6899), .B2(n6166), .A(n6165), .ZN(n6167) );
  AOI211_X1 U7194 ( .C1(n6890), .C2(n6169), .A(n6168), .B(n6167), .ZN(n6175)
         );
  NAND2_X1 U7195 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .ZN(
        n6171) );
  NOR3_X1 U7196 ( .A1(n6190), .A2(REIP_REG_6__SCAN_IN), .A3(n6171), .ZN(n6177)
         );
  INV_X1 U7197 ( .A(n6170), .ZN(n6173) );
  INV_X1 U7198 ( .A(n6171), .ZN(n6172) );
  OAI21_X1 U7199 ( .B1(n6173), .B2(n6172), .A(n6205), .ZN(n6192) );
  OAI21_X1 U7200 ( .B1(n6177), .B2(n6192), .A(REIP_REG_7__SCAN_IN), .ZN(n6174)
         );
  OAI211_X1 U7201 ( .C1(n6223), .C2(n6176), .A(n6175), .B(n6174), .ZN(U2820)
         );
  AOI211_X1 U7202 ( .C1(n6894), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6188), 
        .B(n6177), .ZN(n6178) );
  OAI21_X1 U7203 ( .B1(n6899), .B2(n6179), .A(n6178), .ZN(n6180) );
  AOI21_X1 U7204 ( .B1(EBX_REG_6__SCAN_IN), .B2(n6895), .A(n6180), .ZN(n6183)
         );
  AOI22_X1 U7205 ( .A1(n6890), .A2(n6181), .B1(REIP_REG_6__SCAN_IN), .B2(n6192), .ZN(n6182) );
  OAI211_X1 U7206 ( .C1(n6184), .C2(n6223), .A(n6183), .B(n6182), .ZN(U2821)
         );
  OAI22_X1 U7207 ( .A1(n6229), .A2(n6839), .B1(n6186), .B2(n6185), .ZN(n6187)
         );
  AOI211_X1 U7208 ( .C1(n6220), .C2(n6189), .A(n6188), .B(n6187), .ZN(n6195)
         );
  OAI21_X1 U7209 ( .B1(n6190), .B2(n6658), .A(n6660), .ZN(n6191) );
  AOI22_X1 U7210 ( .A1(n6225), .A2(n6193), .B1(n6192), .B2(n6191), .ZN(n6194)
         );
  OAI211_X1 U7211 ( .C1(n6196), .C2(n6223), .A(n6195), .B(n6194), .ZN(U2822)
         );
  OAI211_X1 U7212 ( .C1(n6206), .C2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .B(n6197), .ZN(n6214) );
  AOI22_X1 U7213 ( .A1(n6219), .A2(n4581), .B1(n6894), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6200) );
  AOI22_X1 U7214 ( .A1(n6220), .A2(n6198), .B1(n6895), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n6199) );
  OAI211_X1 U7215 ( .C1(n6223), .C2(n6201), .A(n6200), .B(n6199), .ZN(n6202)
         );
  AOI21_X1 U7216 ( .B1(n6203), .B2(n6225), .A(n6202), .ZN(n6204) );
  OAI221_X1 U7217 ( .B1(n6205), .B2(n6792), .C1(n6205), .C2(n6214), .A(n6204), 
        .ZN(U2824) );
  INV_X1 U7218 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6655) );
  OAI21_X1 U7219 ( .B1(n6206), .B2(n4559), .A(n6655), .ZN(n6213) );
  AOI22_X1 U7220 ( .A1(n6219), .A2(n6207), .B1(n6894), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7221 ( .A1(n6895), .A2(EBX_REG_2__SCAN_IN), .ZN(n6208) );
  OAI211_X1 U7222 ( .C1(n6899), .C2(n6371), .A(n6209), .B(n6208), .ZN(n6212)
         );
  NOR2_X1 U7223 ( .A1(n6210), .A2(n6330), .ZN(n6211) );
  AOI211_X1 U7224 ( .C1(n6214), .C2(n6213), .A(n6212), .B(n6211), .ZN(n6215)
         );
  OAI21_X1 U7225 ( .B1(n6340), .B2(n6223), .A(n6215), .ZN(U2825) );
  AOI22_X1 U7226 ( .A1(n6894), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6216), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6228) );
  AOI22_X1 U7227 ( .A1(n6219), .A2(n6218), .B1(n6217), .B2(n4559), .ZN(n6222)
         );
  NAND2_X1 U7228 ( .A1(n6220), .A2(n4557), .ZN(n6221) );
  OAI211_X1 U7229 ( .C1(n6223), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n6222), 
        .B(n6221), .ZN(n6224) );
  AOI21_X1 U7230 ( .B1(n6226), .B2(n6225), .A(n6224), .ZN(n6227) );
  OAI211_X1 U7231 ( .C1(n6230), .C2(n6229), .A(n6228), .B(n6227), .ZN(U2826)
         );
  AOI22_X1 U7232 ( .A1(n6234), .A2(n6233), .B1(n6232), .B2(n6231), .ZN(n6235)
         );
  OAI21_X1 U7233 ( .B1(n6236), .B2(n5552), .A(n6235), .ZN(U2846) );
  INV_X1 U7234 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n6828) );
  AOI22_X1 U7235 ( .A1(n6239), .A2(EAX_REG_26__SCAN_IN), .B1(n6267), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6237) );
  OAI21_X1 U7236 ( .B1(n6828), .B2(n6253), .A(n6237), .ZN(U2897) );
  INV_X1 U7237 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n6761) );
  AOI22_X1 U7238 ( .A1(n6266), .A2(DATAO_REG_23__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6239), .ZN(n6238) );
  OAI21_X1 U7239 ( .B1(n6761), .B2(n6246), .A(n6238), .ZN(U2900) );
  INV_X1 U7240 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n6858) );
  AOI22_X1 U7241 ( .A1(n6266), .A2(DATAO_REG_19__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6239), .ZN(n6240) );
  OAI21_X1 U7242 ( .B1(n6858), .B2(n6246), .A(n6240), .ZN(U2904) );
  AOI22_X1 U7243 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6251), .B1(n6266), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6241) );
  OAI21_X1 U7244 ( .B1(n6791), .B2(n6246), .A(n6241), .ZN(U2908) );
  INV_X1 U7245 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6328) );
  AOI22_X1 U7246 ( .A1(n6267), .A2(LWORD_REG_14__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6242) );
  OAI21_X1 U7247 ( .B1(n6328), .B2(n6269), .A(n6242), .ZN(U2909) );
  INV_X1 U7248 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6244) );
  AOI22_X1 U7249 ( .A1(n6267), .A2(LWORD_REG_13__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6243) );
  OAI21_X1 U7250 ( .B1(n6244), .B2(n6269), .A(n6243), .ZN(U2910) );
  INV_X1 U7251 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6760) );
  AOI22_X1 U7252 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6251), .B1(n6266), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6245) );
  OAI21_X1 U7253 ( .B1(n6760), .B2(n6246), .A(n6245), .ZN(U2911) );
  INV_X1 U7254 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6319) );
  AOI22_X1 U7255 ( .A1(n6267), .A2(LWORD_REG_11__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6247) );
  OAI21_X1 U7256 ( .B1(n6319), .B2(n6269), .A(n6247), .ZN(U2912) );
  INV_X1 U7257 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6249) );
  AOI22_X1 U7258 ( .A1(n6267), .A2(LWORD_REG_10__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6248) );
  OAI21_X1 U7259 ( .B1(n6249), .B2(n6269), .A(n6248), .ZN(U2913) );
  INV_X1 U7260 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6314) );
  AOI22_X1 U7261 ( .A1(n6267), .A2(LWORD_REG_9__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6250) );
  OAI21_X1 U7262 ( .B1(n6314), .B2(n6269), .A(n6250), .ZN(U2914) );
  INV_X1 U7263 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6777) );
  AOI22_X1 U7264 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6251), .B1(n6267), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6252) );
  OAI21_X1 U7265 ( .B1(n6777), .B2(n6253), .A(n6252), .ZN(U2915) );
  AOI22_X1 U7266 ( .A1(n6267), .A2(LWORD_REG_7__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6254) );
  OAI21_X1 U7267 ( .B1(n3918), .B2(n6269), .A(n6254), .ZN(U2916) );
  INV_X1 U7268 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6256) );
  AOI22_X1 U7269 ( .A1(n6267), .A2(LWORD_REG_6__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6255) );
  OAI21_X1 U7270 ( .B1(n6256), .B2(n6269), .A(n6255), .ZN(U2917) );
  AOI22_X1 U7271 ( .A1(n6267), .A2(LWORD_REG_5__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6257) );
  OAI21_X1 U7272 ( .B1(n6258), .B2(n6269), .A(n6257), .ZN(U2918) );
  AOI22_X1 U7273 ( .A1(n6267), .A2(LWORD_REG_4__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7274 ( .B1(n6260), .B2(n6269), .A(n6259), .ZN(U2919) );
  AOI22_X1 U7275 ( .A1(n6267), .A2(LWORD_REG_3__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6261) );
  OAI21_X1 U7276 ( .B1(n6262), .B2(n6269), .A(n6261), .ZN(U2920) );
  AOI22_X1 U7277 ( .A1(n6267), .A2(LWORD_REG_2__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6263) );
  OAI21_X1 U7278 ( .B1(n6810), .B2(n6269), .A(n6263), .ZN(U2921) );
  AOI22_X1 U7279 ( .A1(n6267), .A2(LWORD_REG_1__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6264) );
  OAI21_X1 U7280 ( .B1(n6265), .B2(n6269), .A(n6264), .ZN(U2922) );
  AOI22_X1 U7281 ( .A1(n6267), .A2(LWORD_REG_0__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6268) );
  OAI21_X1 U7282 ( .B1(n6270), .B2(n6269), .A(n6268), .ZN(U2923) );
  AOI22_X1 U7283 ( .A1(n4470), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6322), .ZN(n6271) );
  OAI21_X1 U7284 ( .B1(n6324), .B2(n6295), .A(n6271), .ZN(U2924) );
  AOI22_X1 U7285 ( .A1(n4470), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6322), .ZN(n6272) );
  OAI21_X1 U7286 ( .B1(n6324), .B2(n6297), .A(n6272), .ZN(U2925) );
  AOI22_X1 U7287 ( .A1(n6320), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6322), .ZN(n6274) );
  OAI21_X1 U7288 ( .B1(n6324), .B2(n6299), .A(n6274), .ZN(U2926) );
  AOI22_X1 U7289 ( .A1(n6320), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6322), .ZN(n6275) );
  OAI21_X1 U7290 ( .B1(n6324), .B2(n6301), .A(n6275), .ZN(U2927) );
  AOI22_X1 U7291 ( .A1(n6320), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6322), .ZN(n6276) );
  OAI21_X1 U7292 ( .B1(n6324), .B2(n6303), .A(n6276), .ZN(U2928) );
  AOI22_X1 U7293 ( .A1(n4470), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6322), .ZN(n6277) );
  OAI21_X1 U7294 ( .B1(n6324), .B2(n6305), .A(n6277), .ZN(U2929) );
  AOI22_X1 U7295 ( .A1(n4470), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6322), .ZN(n6278) );
  OAI21_X1 U7296 ( .B1(n6324), .B2(n6307), .A(n6278), .ZN(U2930) );
  AOI22_X1 U7297 ( .A1(n4470), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6322), .ZN(n6279) );
  OAI21_X1 U7298 ( .B1(n6324), .B2(n6837), .A(n6279), .ZN(U2931) );
  INV_X1 U7299 ( .A(DATAI_8_), .ZN(n6280) );
  NOR2_X1 U7300 ( .A1(n6324), .A2(n6280), .ZN(n6309) );
  AOI21_X1 U7301 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n4470), .A(n6309), .ZN(n6281) );
  OAI21_X1 U7302 ( .B1(n4226), .B2(n6327), .A(n6281), .ZN(U2932) );
  INV_X1 U7303 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6284) );
  INV_X1 U7304 ( .A(DATAI_9_), .ZN(n6282) );
  NOR2_X1 U7305 ( .A1(n6324), .A2(n6282), .ZN(n6312) );
  AOI21_X1 U7306 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n4470), .A(n6312), .ZN(n6283) );
  OAI21_X1 U7307 ( .B1(n6284), .B2(n6327), .A(n6283), .ZN(U2933) );
  AOI22_X1 U7308 ( .A1(n6320), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n6322), .ZN(n6286) );
  NAND2_X1 U7309 ( .A1(n6285), .A2(DATAI_10_), .ZN(n6315) );
  NAND2_X1 U7310 ( .A1(n6286), .A2(n6315), .ZN(U2934) );
  INV_X1 U7311 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6289) );
  INV_X1 U7312 ( .A(DATAI_11_), .ZN(n6287) );
  NOR2_X1 U7313 ( .A1(n6324), .A2(n6287), .ZN(n6317) );
  AOI21_X1 U7314 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n4470), .A(n6317), .ZN(
        n6288) );
  OAI21_X1 U7315 ( .B1(n6289), .B2(n6327), .A(n6288), .ZN(U2935) );
  INV_X1 U7316 ( .A(DATAI_12_), .ZN(n6759) );
  AOI22_X1 U7317 ( .A1(n6320), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n6322), .ZN(n6290) );
  OAI21_X1 U7318 ( .B1(n6324), .B2(n6759), .A(n6290), .ZN(U2936) );
  INV_X1 U7319 ( .A(DATAI_13_), .ZN(n6773) );
  AOI22_X1 U7320 ( .A1(n6320), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6322), .ZN(n6291) );
  OAI21_X1 U7321 ( .B1(n6324), .B2(n6773), .A(n6291), .ZN(U2937) );
  INV_X1 U7322 ( .A(DATAI_14_), .ZN(n6292) );
  NOR2_X1 U7323 ( .A1(n6324), .A2(n6292), .ZN(n6325) );
  AOI21_X1 U7324 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n4470), .A(n6325), .ZN(
        n6293) );
  OAI21_X1 U7325 ( .B1(n6731), .B2(n6327), .A(n6293), .ZN(U2938) );
  AOI22_X1 U7326 ( .A1(n6320), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6322), .ZN(n6294) );
  OAI21_X1 U7327 ( .B1(n6324), .B2(n6295), .A(n6294), .ZN(U2939) );
  AOI22_X1 U7328 ( .A1(n6320), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6322), .ZN(n6296) );
  OAI21_X1 U7329 ( .B1(n6324), .B2(n6297), .A(n6296), .ZN(U2940) );
  AOI22_X1 U7330 ( .A1(n6320), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6322), .ZN(n6298) );
  OAI21_X1 U7331 ( .B1(n6324), .B2(n6299), .A(n6298), .ZN(U2941) );
  AOI22_X1 U7332 ( .A1(n6320), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6322), .ZN(n6300) );
  OAI21_X1 U7333 ( .B1(n6324), .B2(n6301), .A(n6300), .ZN(U2942) );
  AOI22_X1 U7334 ( .A1(n6320), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6322), .ZN(n6302) );
  OAI21_X1 U7335 ( .B1(n6324), .B2(n6303), .A(n6302), .ZN(U2943) );
  AOI22_X1 U7336 ( .A1(n6320), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6322), .ZN(n6304) );
  OAI21_X1 U7337 ( .B1(n6324), .B2(n6305), .A(n6304), .ZN(U2944) );
  AOI22_X1 U7338 ( .A1(n6320), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6322), .ZN(n6306) );
  OAI21_X1 U7339 ( .B1(n6324), .B2(n6307), .A(n6306), .ZN(U2945) );
  AOI22_X1 U7340 ( .A1(n6320), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6322), .ZN(n6308) );
  OAI21_X1 U7341 ( .B1(n6324), .B2(n6837), .A(n6308), .ZN(U2946) );
  INV_X1 U7342 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6311) );
  AOI21_X1 U7343 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6320), .A(n6309), .ZN(n6310) );
  OAI21_X1 U7344 ( .B1(n6311), .B2(n6327), .A(n6310), .ZN(U2947) );
  AOI21_X1 U7345 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6320), .A(n6312), .ZN(n6313) );
  OAI21_X1 U7346 ( .B1(n6314), .B2(n6327), .A(n6313), .ZN(U2948) );
  AOI22_X1 U7347 ( .A1(n6320), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6322), .ZN(n6316) );
  NAND2_X1 U7348 ( .A1(n6316), .A2(n6315), .ZN(U2949) );
  AOI21_X1 U7349 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6320), .A(n6317), .ZN(
        n6318) );
  OAI21_X1 U7350 ( .B1(n6319), .B2(n6327), .A(n6318), .ZN(U2950) );
  AOI22_X1 U7351 ( .A1(n6320), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n6322), .ZN(n6321) );
  OAI21_X1 U7352 ( .B1(n6324), .B2(n6759), .A(n6321), .ZN(U2951) );
  AOI22_X1 U7353 ( .A1(n4470), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6322), .ZN(n6323) );
  OAI21_X1 U7354 ( .B1(n6324), .B2(n6773), .A(n6323), .ZN(U2952) );
  AOI21_X1 U7355 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6320), .A(n6325), .ZN(
        n6326) );
  OAI21_X1 U7356 ( .B1(n6328), .B2(n6327), .A(n6326), .ZN(U2953) );
  AOI22_X1 U7357 ( .A1(n6368), .A2(REIP_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6329), .ZN(n6339) );
  INV_X1 U7358 ( .A(n6330), .ZN(n6337) );
  INV_X1 U7359 ( .A(n6332), .ZN(n6334) );
  NAND2_X1 U7360 ( .A1(n6334), .A2(n6333), .ZN(n6335) );
  XNOR2_X1 U7361 ( .A(n6331), .B(n6335), .ZN(n6376) );
  AOI22_X1 U7362 ( .A1(n6337), .A2(n5804), .B1(n6376), .B2(n6336), .ZN(n6338)
         );
  OAI211_X1 U7363 ( .C1(n6341), .C2(n6340), .A(n6339), .B(n6338), .ZN(U2984)
         );
  AOI21_X1 U7364 ( .B1(n6343), .B2(n6359), .A(n6342), .ZN(n6347) );
  AOI22_X1 U7365 ( .A1(n6345), .A2(n6381), .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6344), .ZN(n6346) );
  OAI211_X1 U7366 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6348), .A(n6347), .B(n6346), .ZN(U3007) );
  AOI21_X1 U7367 ( .B1(n6350), .B2(n6359), .A(n6349), .ZN(n6354) );
  AOI22_X1 U7368 ( .A1(n6352), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n6351), 
        .B2(n6381), .ZN(n6353) );
  OAI211_X1 U7369 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6355), .A(n6354), 
        .B(n6353), .ZN(U3009) );
  NAND2_X1 U7370 ( .A1(n6356), .A2(n6381), .ZN(n6361) );
  AOI21_X1 U7371 ( .B1(n6359), .B2(n6358), .A(n6357), .ZN(n6360) );
  OAI211_X1 U7372 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6362), .A(n6361), 
        .B(n6360), .ZN(n6363) );
  INV_X1 U7373 ( .A(n6363), .ZN(n6364) );
  OAI21_X1 U7374 ( .B1(n6366), .B2(n6365), .A(n6364), .ZN(U3011) );
  NAND2_X1 U7375 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6367), .ZN(n6379)
         );
  NAND2_X1 U7376 ( .A1(n6368), .A2(REIP_REG_2__SCAN_IN), .ZN(n6369) );
  OAI211_X1 U7377 ( .C1(n6371), .C2(n6387), .A(n6370), .B(n6369), .ZN(n6375)
         );
  NOR3_X1 U7378 ( .A1(n6373), .A2(n6372), .A3(n6393), .ZN(n6374) );
  AOI211_X1 U7379 ( .C1(n6381), .C2(n6376), .A(n6375), .B(n6374), .ZN(n6377)
         );
  OAI221_X1 U7380 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6379), .C1(n6874), .C2(n6378), .A(n6377), .ZN(U3016) );
  AND3_X1 U7381 ( .A1(n6382), .A2(n6381), .A3(n6380), .ZN(n6389) );
  INV_X1 U7382 ( .A(n6383), .ZN(n6384) );
  OAI211_X1 U7383 ( .C1(n6387), .C2(n6386), .A(n6385), .B(n6384), .ZN(n6388)
         );
  NOR2_X1 U7384 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  OAI221_X1 U7385 ( .B1(n6393), .B2(n6392), .C1(n6393), .C2(n6391), .A(n6390), 
        .ZN(U3018) );
  NOR2_X1 U7386 ( .A1(n6395), .A2(n6394), .ZN(U3019) );
  OR2_X1 U7387 ( .A1(n6510), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6426)
         );
  OAI22_X1 U7388 ( .A1(n6432), .A2(n6592), .B1(n6511), .B2(n6426), .ZN(n6397)
         );
  INV_X1 U7389 ( .A(n6397), .ZN(n6407) );
  OAI21_X1 U7390 ( .B1(n6398), .B2(n6513), .A(n6437), .ZN(n6405) );
  OAI21_X1 U7391 ( .B1(n6399), .B2(n6515), .A(n6426), .ZN(n6402) );
  OAI21_X1 U7392 ( .B1(n6522), .B2(n6437), .A(n6400), .ZN(n6518) );
  NOR2_X1 U7393 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6518), .ZN(n6401)
         );
  OAI21_X1 U7394 ( .B1(n6405), .B2(n6402), .A(n6401), .ZN(n6429) );
  INV_X1 U7395 ( .A(n6402), .ZN(n6404) );
  NAND3_X1 U7396 ( .A1(n6522), .A2(STATE2_REG_2__SCAN_IN), .A3(n6519), .ZN(
        n6403) );
  AOI22_X1 U7397 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6429), .B1(n6428), 
        .B2(n6577), .ZN(n6406) );
  OAI211_X1 U7398 ( .C1(n6528), .C2(n6464), .A(n6407), .B(n6406), .ZN(U3044)
         );
  OAI22_X1 U7399 ( .A1(n6432), .A2(n6598), .B1(n6529), .B2(n6426), .ZN(n6408)
         );
  INV_X1 U7400 ( .A(n6408), .ZN(n6410) );
  AOI22_X1 U7401 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6429), .B1(n6428), 
        .B2(n6594), .ZN(n6409) );
  OAI211_X1 U7402 ( .C1(n6530), .C2(n6464), .A(n6410), .B(n6409), .ZN(U3045)
         );
  OAI22_X1 U7403 ( .A1(n6464), .A2(n6535), .B1(n6534), .B2(n6426), .ZN(n6411)
         );
  INV_X1 U7404 ( .A(n6411), .ZN(n6413) );
  AOI22_X1 U7405 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6429), .B1(n6428), 
        .B2(n6600), .ZN(n6412) );
  OAI211_X1 U7406 ( .C1(n6432), .C2(n6604), .A(n6413), .B(n6412), .ZN(U3046)
         );
  OAI22_X1 U7407 ( .A1(n6432), .A2(n6610), .B1(n6539), .B2(n6426), .ZN(n6414)
         );
  INV_X1 U7408 ( .A(n6414), .ZN(n6416) );
  AOI22_X1 U7409 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6429), .B1(n6428), 
        .B2(n6606), .ZN(n6415) );
  OAI211_X1 U7410 ( .C1(n6540), .C2(n6464), .A(n6416), .B(n6415), .ZN(U3047)
         );
  OAI22_X1 U7411 ( .A1(n6464), .A2(n6545), .B1(n6544), .B2(n6426), .ZN(n6417)
         );
  INV_X1 U7412 ( .A(n6417), .ZN(n6419) );
  AOI22_X1 U7413 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6429), .B1(n6428), 
        .B2(n6612), .ZN(n6418) );
  OAI211_X1 U7414 ( .C1(n6432), .C2(n6616), .A(n6419), .B(n6418), .ZN(U3048)
         );
  OAI22_X1 U7415 ( .A1(n6432), .A2(n6622), .B1(n6549), .B2(n6426), .ZN(n6420)
         );
  INV_X1 U7416 ( .A(n6420), .ZN(n6422) );
  AOI22_X1 U7417 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6429), .B1(n6428), 
        .B2(n6618), .ZN(n6421) );
  OAI211_X1 U7418 ( .C1(n6553), .C2(n6464), .A(n6422), .B(n6421), .ZN(U3049)
         );
  OAI22_X1 U7419 ( .A1(n6432), .A2(n6628), .B1(n6554), .B2(n6426), .ZN(n6423)
         );
  INV_X1 U7420 ( .A(n6423), .ZN(n6425) );
  AOI22_X1 U7421 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6429), .B1(n6428), 
        .B2(n6624), .ZN(n6424) );
  OAI211_X1 U7422 ( .C1(n6558), .C2(n6464), .A(n6425), .B(n6424), .ZN(U3050)
         );
  OAI22_X1 U7423 ( .A1(n6464), .A2(n6561), .B1(n6560), .B2(n6426), .ZN(n6427)
         );
  INV_X1 U7424 ( .A(n6427), .ZN(n6431) );
  AOI22_X1 U7425 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6429), .B1(n6428), 
        .B2(n6631), .ZN(n6430) );
  OAI211_X1 U7426 ( .C1(n6432), .C2(n6639), .A(n6431), .B(n6430), .ZN(U3051)
         );
  OAI33_X1 U7427 ( .A1(n4581), .A2(n6580), .A3(n6578), .B1(n6433), .B2(n6568), 
        .B3(n6476), .ZN(n6459) );
  NAND2_X1 U7428 ( .A1(n6434), .A2(n6574), .ZN(n6439) );
  INV_X1 U7429 ( .A(n6439), .ZN(n6458) );
  AOI22_X1 U7430 ( .A1(n3007), .A2(n6577), .B1(n6576), .B2(n6458), .ZN(n6445)
         );
  AOI21_X1 U7431 ( .B1(n6464), .B2(n6436), .A(n6435), .ZN(n6443) );
  NAND2_X1 U7432 ( .A1(n6438), .A2(n6437), .ZN(n6442) );
  AOI21_X1 U7433 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6439), .A(n6584), .ZN(
        n6440) );
  AOI22_X1 U7434 ( .A1(n6461), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6589), 
        .B2(n6460), .ZN(n6444) );
  OAI211_X1 U7435 ( .C1(n6592), .C2(n6464), .A(n6445), .B(n6444), .ZN(U3052)
         );
  AOI22_X1 U7436 ( .A1(n3007), .A2(n6594), .B1(n6593), .B2(n6458), .ZN(n6447)
         );
  AOI22_X1 U7437 ( .A1(n6461), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6595), 
        .B2(n6460), .ZN(n6446) );
  OAI211_X1 U7438 ( .C1(n6598), .C2(n6464), .A(n6447), .B(n6446), .ZN(U3053)
         );
  AOI22_X1 U7439 ( .A1(n3007), .A2(n6600), .B1(n6599), .B2(n6458), .ZN(n6449)
         );
  AOI22_X1 U7440 ( .A1(n6461), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6601), 
        .B2(n6460), .ZN(n6448) );
  OAI211_X1 U7441 ( .C1(n6604), .C2(n6464), .A(n6449), .B(n6448), .ZN(U3054)
         );
  AOI22_X1 U7442 ( .A1(n3007), .A2(n6606), .B1(n6605), .B2(n6458), .ZN(n6451)
         );
  AOI22_X1 U7443 ( .A1(n6461), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6607), 
        .B2(n6460), .ZN(n6450) );
  OAI211_X1 U7444 ( .C1(n6610), .C2(n6464), .A(n6451), .B(n6450), .ZN(U3055)
         );
  AOI22_X1 U7445 ( .A1(n3007), .A2(n6612), .B1(n6611), .B2(n6458), .ZN(n6453)
         );
  AOI22_X1 U7446 ( .A1(n6461), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6613), 
        .B2(n6460), .ZN(n6452) );
  OAI211_X1 U7447 ( .C1(n6616), .C2(n6464), .A(n6453), .B(n6452), .ZN(U3056)
         );
  AOI22_X1 U7448 ( .A1(n3007), .A2(n6618), .B1(n6617), .B2(n6458), .ZN(n6455)
         );
  AOI22_X1 U7449 ( .A1(n6461), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6619), 
        .B2(n6460), .ZN(n6454) );
  OAI211_X1 U7450 ( .C1(n6622), .C2(n6464), .A(n6455), .B(n6454), .ZN(U3057)
         );
  AOI22_X1 U7451 ( .A1(n6624), .A2(n3007), .B1(n6623), .B2(n6458), .ZN(n6457)
         );
  AOI22_X1 U7452 ( .A1(n6461), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6625), 
        .B2(n6460), .ZN(n6456) );
  OAI211_X1 U7453 ( .C1(n6628), .C2(n6464), .A(n6457), .B(n6456), .ZN(U3058)
         );
  AOI22_X1 U7454 ( .A1(n3007), .A2(n6631), .B1(n6630), .B2(n6458), .ZN(n6463)
         );
  AOI22_X1 U7455 ( .A1(n6461), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6634), 
        .B2(n6460), .ZN(n6462) );
  OAI211_X1 U7456 ( .C1(n6639), .C2(n6464), .A(n6463), .B(n6462), .ZN(U3059)
         );
  AOI22_X1 U7457 ( .A1(n6576), .A2(n6466), .B1(n6465), .B2(n6577), .ZN(n6473)
         );
  INV_X1 U7458 ( .A(n6467), .ZN(n6471) );
  INV_X1 U7459 ( .A(n6468), .ZN(n6469) );
  AOI22_X1 U7460 ( .A1(n6471), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6470), 
        .B2(n6469), .ZN(n6472) );
  OAI211_X1 U7461 ( .C1(n6528), .C2(n6474), .A(n6473), .B(n6472), .ZN(U3068)
         );
  INV_X1 U7462 ( .A(n6475), .ZN(n6573) );
  INV_X1 U7463 ( .A(n6476), .ZN(n6572) );
  OAI22_X1 U7464 ( .A1(n6573), .A2(n6481), .B1(n6572), .B2(n6477), .ZN(n6502)
         );
  OR2_X1 U7465 ( .A1(n6478), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6484)
         );
  INV_X1 U7466 ( .A(n6484), .ZN(n6501) );
  AOI22_X1 U7467 ( .A1(n6502), .A2(n6577), .B1(n6576), .B2(n6501), .ZN(n6488)
         );
  OAI21_X1 U7468 ( .B1(n6503), .B2(n6479), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6480) );
  OAI211_X1 U7469 ( .C1(n6482), .C2(n6481), .A(n6480), .B(n6437), .ZN(n6486)
         );
  AOI21_X1 U7470 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6572), .A(n6483), .ZN(
        n6587) );
  NAND2_X1 U7471 ( .A1(n6484), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6485) );
  NAND4_X1 U7472 ( .A1(n6486), .A2(n6587), .A3(n6568), .A4(n6485), .ZN(n6504)
         );
  AOI22_X1 U7473 ( .A1(n6504), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6589), 
        .B2(n6503), .ZN(n6487) );
  OAI211_X1 U7474 ( .C1(n6592), .C2(n6507), .A(n6488), .B(n6487), .ZN(U3084)
         );
  AOI22_X1 U7475 ( .A1(n6502), .A2(n6594), .B1(n6593), .B2(n6501), .ZN(n6490)
         );
  AOI22_X1 U7476 ( .A1(n6504), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6595), 
        .B2(n6503), .ZN(n6489) );
  OAI211_X1 U7477 ( .C1(n6598), .C2(n6507), .A(n6490), .B(n6489), .ZN(U3085)
         );
  AOI22_X1 U7478 ( .A1(n6502), .A2(n6600), .B1(n6599), .B2(n6501), .ZN(n6492)
         );
  AOI22_X1 U7479 ( .A1(n6504), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6601), 
        .B2(n6503), .ZN(n6491) );
  OAI211_X1 U7480 ( .C1(n6604), .C2(n6507), .A(n6492), .B(n6491), .ZN(U3086)
         );
  AOI22_X1 U7481 ( .A1(n6502), .A2(n6606), .B1(n6605), .B2(n6501), .ZN(n6494)
         );
  AOI22_X1 U7482 ( .A1(n6504), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6607), 
        .B2(n6503), .ZN(n6493) );
  OAI211_X1 U7483 ( .C1(n6610), .C2(n6507), .A(n6494), .B(n6493), .ZN(U3087)
         );
  AOI22_X1 U7484 ( .A1(n6502), .A2(n6612), .B1(n6611), .B2(n6501), .ZN(n6496)
         );
  AOI22_X1 U7485 ( .A1(n6504), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6613), 
        .B2(n6503), .ZN(n6495) );
  OAI211_X1 U7486 ( .C1(n6616), .C2(n6507), .A(n6496), .B(n6495), .ZN(U3088)
         );
  AOI22_X1 U7487 ( .A1(n6502), .A2(n6618), .B1(n6617), .B2(n6501), .ZN(n6498)
         );
  AOI22_X1 U7488 ( .A1(n6504), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6619), 
        .B2(n6503), .ZN(n6497) );
  OAI211_X1 U7489 ( .C1(n6622), .C2(n6507), .A(n6498), .B(n6497), .ZN(U3089)
         );
  AOI22_X1 U7490 ( .A1(n6624), .A2(n6502), .B1(n6623), .B2(n6501), .ZN(n6500)
         );
  AOI22_X1 U7491 ( .A1(n6504), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6625), 
        .B2(n6503), .ZN(n6499) );
  OAI211_X1 U7492 ( .C1(n6628), .C2(n6507), .A(n6500), .B(n6499), .ZN(U3090)
         );
  AOI22_X1 U7493 ( .A1(n6502), .A2(n6631), .B1(n6630), .B2(n6501), .ZN(n6506)
         );
  AOI22_X1 U7494 ( .A1(n6504), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6634), 
        .B2(n6503), .ZN(n6505) );
  OAI211_X1 U7495 ( .C1(n6639), .C2(n6507), .A(n6506), .B(n6505), .ZN(U3091)
         );
  INV_X1 U7496 ( .A(n6508), .ZN(n6509) );
  OR2_X1 U7497 ( .A1(n6510), .A2(n6519), .ZN(n6559) );
  OAI22_X1 U7498 ( .A1(n6567), .A2(n6592), .B1(n6511), .B2(n6559), .ZN(n6512)
         );
  INV_X1 U7499 ( .A(n6512), .ZN(n6527) );
  OAI21_X1 U7500 ( .B1(n6514), .B2(n6513), .A(n6437), .ZN(n6525) );
  OR2_X1 U7501 ( .A1(n6516), .A2(n6515), .ZN(n6517) );
  NAND2_X1 U7502 ( .A1(n6517), .A2(n6559), .ZN(n6521) );
  NOR2_X1 U7503 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  OAI21_X1 U7504 ( .B1(n6525), .B2(n6521), .A(n6520), .ZN(n6564) );
  INV_X1 U7505 ( .A(n6521), .ZN(n6524) );
  NAND3_X1 U7506 ( .A1(n6522), .A2(STATE2_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6523) );
  AOI22_X1 U7507 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6564), .B1(n6563), 
        .B2(n6577), .ZN(n6526) );
  OAI211_X1 U7508 ( .C1(n6528), .C2(n6638), .A(n6527), .B(n6526), .ZN(U3108)
         );
  OAI22_X1 U7509 ( .A1(n6638), .A2(n6530), .B1(n6529), .B2(n6559), .ZN(n6531)
         );
  INV_X1 U7510 ( .A(n6531), .ZN(n6533) );
  AOI22_X1 U7511 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6564), .B1(n6563), 
        .B2(n6594), .ZN(n6532) );
  OAI211_X1 U7512 ( .C1(n6598), .C2(n6567), .A(n6533), .B(n6532), .ZN(U3109)
         );
  OAI22_X1 U7513 ( .A1(n6638), .A2(n6535), .B1(n6534), .B2(n6559), .ZN(n6536)
         );
  INV_X1 U7514 ( .A(n6536), .ZN(n6538) );
  AOI22_X1 U7515 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6564), .B1(n6563), 
        .B2(n6600), .ZN(n6537) );
  OAI211_X1 U7516 ( .C1(n6604), .C2(n6567), .A(n6538), .B(n6537), .ZN(U3110)
         );
  OAI22_X1 U7517 ( .A1(n6638), .A2(n6540), .B1(n6539), .B2(n6559), .ZN(n6541)
         );
  INV_X1 U7518 ( .A(n6541), .ZN(n6543) );
  AOI22_X1 U7519 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6564), .B1(n6563), 
        .B2(n6606), .ZN(n6542) );
  OAI211_X1 U7520 ( .C1(n6610), .C2(n6567), .A(n6543), .B(n6542), .ZN(U3111)
         );
  OAI22_X1 U7521 ( .A1(n6638), .A2(n6545), .B1(n6544), .B2(n6559), .ZN(n6546)
         );
  INV_X1 U7522 ( .A(n6546), .ZN(n6548) );
  AOI22_X1 U7523 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6564), .B1(n6563), 
        .B2(n6612), .ZN(n6547) );
  OAI211_X1 U7524 ( .C1(n6616), .C2(n6567), .A(n6548), .B(n6547), .ZN(U3112)
         );
  OAI22_X1 U7525 ( .A1(n6567), .A2(n6622), .B1(n6549), .B2(n6559), .ZN(n6550)
         );
  INV_X1 U7526 ( .A(n6550), .ZN(n6552) );
  AOI22_X1 U7527 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6564), .B1(n6563), 
        .B2(n6618), .ZN(n6551) );
  OAI211_X1 U7528 ( .C1(n6553), .C2(n6638), .A(n6552), .B(n6551), .ZN(U3113)
         );
  OAI22_X1 U7529 ( .A1(n6567), .A2(n6628), .B1(n6554), .B2(n6559), .ZN(n6555)
         );
  INV_X1 U7530 ( .A(n6555), .ZN(n6557) );
  AOI22_X1 U7531 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6564), .B1(n6563), 
        .B2(n6624), .ZN(n6556) );
  OAI211_X1 U7532 ( .C1(n6558), .C2(n6638), .A(n6557), .B(n6556), .ZN(U3114)
         );
  OAI22_X1 U7533 ( .A1(n6638), .A2(n6561), .B1(n6560), .B2(n6559), .ZN(n6562)
         );
  INV_X1 U7534 ( .A(n6562), .ZN(n6566) );
  AOI22_X1 U7535 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6564), .B1(n6563), 
        .B2(n6631), .ZN(n6565) );
  OAI211_X1 U7536 ( .C1(n6639), .C2(n6567), .A(n6566), .B(n6565), .ZN(U3115)
         );
  INV_X1 U7537 ( .A(n6568), .ZN(n6570) );
  NAND2_X1 U7538 ( .A1(n6570), .A2(n6569), .ZN(n6571) );
  OAI22_X1 U7539 ( .A1(n6573), .A2(n6580), .B1(n6572), .B2(n6571), .ZN(n6632)
         );
  NAND2_X1 U7540 ( .A1(n6575), .A2(n6574), .ZN(n6585) );
  INV_X1 U7541 ( .A(n6585), .ZN(n6629) );
  AOI22_X1 U7542 ( .A1(n6632), .A2(n6577), .B1(n6576), .B2(n6629), .ZN(n6591)
         );
  INV_X1 U7543 ( .A(n6638), .ZN(n6579) );
  NOR3_X1 U7544 ( .A1(n6633), .A2(n6579), .A3(n6578), .ZN(n6583) );
  OAI22_X1 U7545 ( .A1(n6583), .A2(n6582), .B1(n6581), .B2(n6580), .ZN(n6588)
         );
  AOI21_X1 U7546 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6585), .A(n6584), .ZN(
        n6586) );
  NAND3_X1 U7547 ( .A1(n6588), .A2(n6587), .A3(n6586), .ZN(n6635) );
  AOI22_X1 U7548 ( .A1(n6635), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n6589), 
        .B2(n6633), .ZN(n6590) );
  OAI211_X1 U7549 ( .C1(n6592), .C2(n6638), .A(n6591), .B(n6590), .ZN(U3116)
         );
  AOI22_X1 U7550 ( .A1(n6632), .A2(n6594), .B1(n6593), .B2(n6629), .ZN(n6597)
         );
  AOI22_X1 U7551 ( .A1(n6635), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n6595), 
        .B2(n6633), .ZN(n6596) );
  OAI211_X1 U7552 ( .C1(n6598), .C2(n6638), .A(n6597), .B(n6596), .ZN(U3117)
         );
  AOI22_X1 U7553 ( .A1(n6632), .A2(n6600), .B1(n6599), .B2(n6629), .ZN(n6603)
         );
  AOI22_X1 U7554 ( .A1(n6635), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n6601), 
        .B2(n6633), .ZN(n6602) );
  OAI211_X1 U7555 ( .C1(n6604), .C2(n6638), .A(n6603), .B(n6602), .ZN(U3118)
         );
  AOI22_X1 U7556 ( .A1(n6632), .A2(n6606), .B1(n6605), .B2(n6629), .ZN(n6609)
         );
  AOI22_X1 U7557 ( .A1(n6635), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n6607), 
        .B2(n6633), .ZN(n6608) );
  OAI211_X1 U7558 ( .C1(n6610), .C2(n6638), .A(n6609), .B(n6608), .ZN(U3119)
         );
  AOI22_X1 U7559 ( .A1(n6632), .A2(n6612), .B1(n6611), .B2(n6629), .ZN(n6615)
         );
  AOI22_X1 U7560 ( .A1(n6635), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n6613), 
        .B2(n6633), .ZN(n6614) );
  OAI211_X1 U7561 ( .C1(n6616), .C2(n6638), .A(n6615), .B(n6614), .ZN(U3120)
         );
  AOI22_X1 U7562 ( .A1(n6632), .A2(n6618), .B1(n6617), .B2(n6629), .ZN(n6621)
         );
  AOI22_X1 U7563 ( .A1(n6635), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n6619), 
        .B2(n6633), .ZN(n6620) );
  OAI211_X1 U7564 ( .C1(n6622), .C2(n6638), .A(n6621), .B(n6620), .ZN(U3121)
         );
  AOI22_X1 U7565 ( .A1(n6624), .A2(n6632), .B1(n6623), .B2(n6629), .ZN(n6627)
         );
  AOI22_X1 U7566 ( .A1(n6635), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n6625), 
        .B2(n6633), .ZN(n6626) );
  OAI211_X1 U7567 ( .C1(n6628), .C2(n6638), .A(n6627), .B(n6626), .ZN(U3122)
         );
  AOI22_X1 U7568 ( .A1(n6632), .A2(n6631), .B1(n6630), .B2(n6629), .ZN(n6637)
         );
  AOI22_X1 U7569 ( .A1(n6635), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n6634), 
        .B2(n6633), .ZN(n6636) );
  OAI211_X1 U7570 ( .C1(n6639), .C2(n6638), .A(n6637), .B(n6636), .ZN(U3123)
         );
  AOI21_X1 U7571 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6640), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n6642) );
  OAI21_X1 U7572 ( .B1(n6643), .B2(n6642), .A(n6641), .ZN(U3150) );
  AND2_X1 U7573 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6644), .ZN(U3151) );
  AND2_X1 U7574 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6644), .ZN(U3152) );
  AND2_X1 U7575 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6644), .ZN(U3153) );
  INV_X1 U7576 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6851) );
  NOR2_X1 U7577 ( .A1(n6702), .A2(n6851), .ZN(U3154) );
  NOR2_X1 U7578 ( .A1(n6702), .A2(n6868), .ZN(U3155) );
  INV_X1 U7579 ( .A(DATAWIDTH_REG_26__SCAN_IN), .ZN(n6856) );
  NOR2_X1 U7580 ( .A1(n6702), .A2(n6856), .ZN(U3156) );
  AND2_X1 U7581 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6644), .ZN(U3157) );
  AND2_X1 U7582 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6644), .ZN(U3158) );
  AND2_X1 U7583 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6644), .ZN(U3159) );
  AND2_X1 U7584 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6644), .ZN(U3160) );
  AND2_X1 U7585 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6644), .ZN(U3161) );
  AND2_X1 U7586 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6644), .ZN(U3162) );
  NOR2_X1 U7587 ( .A1(n6702), .A2(n6804), .ZN(U3163) );
  AND2_X1 U7588 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6644), .ZN(U3164) );
  AND2_X1 U7589 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6644), .ZN(U3165) );
  AND2_X1 U7590 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6644), .ZN(U3166) );
  AND2_X1 U7591 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6644), .ZN(U3167) );
  AND2_X1 U7592 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6644), .ZN(U3168) );
  AND2_X1 U7593 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6644), .ZN(U3169) );
  AND2_X1 U7594 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6644), .ZN(U3170) );
  AND2_X1 U7595 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6644), .ZN(U3171) );
  INV_X1 U7596 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6871) );
  NOR2_X1 U7597 ( .A1(n6702), .A2(n6871), .ZN(U3172) );
  AND2_X1 U7598 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6644), .ZN(U3173) );
  AND2_X1 U7599 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6644), .ZN(U3174) );
  AND2_X1 U7600 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6644), .ZN(U3175) );
  AND2_X1 U7601 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6644), .ZN(U3176) );
  AND2_X1 U7602 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6644), .ZN(U3177) );
  AND2_X1 U7603 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6644), .ZN(U3178) );
  AND2_X1 U7604 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6644), .ZN(U3179) );
  AND2_X1 U7605 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6644), .ZN(U3180) );
  AOI221_X1 U7606 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6712), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6646) );
  AOI221_X1 U7607 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6646), .C2(HOLD), .A(n6645), .ZN(n6652) );
  AOI21_X1 U7608 ( .B1(n6648), .B2(n6647), .A(STATE_REG_2__SCAN_IN), .ZN(n6650) );
  OAI22_X1 U7609 ( .A1(n6652), .A2(n6651), .B1(n6650), .B2(n6649), .ZN(U3183)
         );
  AOI22_X1 U7610 ( .A1(n6692), .A2(REIP_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6673), .ZN(n6653) );
  OAI21_X1 U7611 ( .B1(n4559), .B2(n6694), .A(n6653), .ZN(U3184) );
  AOI22_X1 U7612 ( .A1(n6692), .A2(REIP_REG_3__SCAN_IN), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6673), .ZN(n6654) );
  OAI21_X1 U7613 ( .B1(n6655), .B2(n6694), .A(n6654), .ZN(U3185) );
  AOI22_X1 U7614 ( .A1(n6692), .A2(REIP_REG_4__SCAN_IN), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6673), .ZN(n6656) );
  OAI21_X1 U7615 ( .B1(n6792), .B2(n6694), .A(n6656), .ZN(U3186) );
  AOI22_X1 U7616 ( .A1(n6692), .A2(REIP_REG_5__SCAN_IN), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6673), .ZN(n6657) );
  OAI21_X1 U7617 ( .B1(n6658), .B2(n6694), .A(n6657), .ZN(U3187) );
  AOI22_X1 U7618 ( .A1(n6692), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6673), .ZN(n6659) );
  OAI21_X1 U7619 ( .B1(n6660), .B2(n6694), .A(n6659), .ZN(U3188) );
  AOI22_X1 U7620 ( .A1(n6692), .A2(REIP_REG_8__SCAN_IN), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6673), .ZN(n6661) );
  OAI21_X1 U7621 ( .B1(n6662), .B2(n6694), .A(n6661), .ZN(U3190) );
  INV_X1 U7622 ( .A(n6694), .ZN(n6696) );
  AOI22_X1 U7623 ( .A1(n6696), .A2(REIP_REG_8__SCAN_IN), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6673), .ZN(n6663) );
  OAI21_X1 U7624 ( .B1(n6893), .B2(n6698), .A(n6663), .ZN(U3191) );
  AOI22_X1 U7625 ( .A1(n6696), .A2(REIP_REG_9__SCAN_IN), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6673), .ZN(n6664) );
  OAI21_X1 U7626 ( .B1(n5782), .B2(n6698), .A(n6664), .ZN(U3192) );
  AOI22_X1 U7627 ( .A1(n6692), .A2(REIP_REG_11__SCAN_IN), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6673), .ZN(n6665) );
  OAI21_X1 U7628 ( .B1(n5782), .B2(n6694), .A(n6665), .ZN(U3193) );
  AOI22_X1 U7629 ( .A1(n6696), .A2(REIP_REG_11__SCAN_IN), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6673), .ZN(n6666) );
  OAI21_X1 U7630 ( .B1(n6148), .B2(n6698), .A(n6666), .ZN(U3194) );
  AOI22_X1 U7631 ( .A1(n6692), .A2(REIP_REG_14__SCAN_IN), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6673), .ZN(n6667) );
  OAI21_X1 U7632 ( .B1(n6668), .B2(n6694), .A(n6667), .ZN(U3196) );
  AOI22_X1 U7633 ( .A1(n6696), .A2(REIP_REG_14__SCAN_IN), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6673), .ZN(n6669) );
  OAI21_X1 U7634 ( .B1(n6670), .B2(n6698), .A(n6669), .ZN(U3197) );
  AOI22_X1 U7635 ( .A1(n6692), .A2(REIP_REG_17__SCAN_IN), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6673), .ZN(n6671) );
  OAI21_X1 U7636 ( .B1(n6672), .B2(n6694), .A(n6671), .ZN(U3199) );
  AOI22_X1 U7637 ( .A1(n6692), .A2(REIP_REG_18__SCAN_IN), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6673), .ZN(n6674) );
  OAI21_X1 U7638 ( .B1(n6675), .B2(n6694), .A(n6674), .ZN(U3200) );
  AOI22_X1 U7639 ( .A1(n6692), .A2(REIP_REG_19__SCAN_IN), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6673), .ZN(n6676) );
  OAI21_X1 U7640 ( .B1(n6677), .B2(n6694), .A(n6676), .ZN(U3201) );
  AOI22_X1 U7641 ( .A1(n6692), .A2(REIP_REG_20__SCAN_IN), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6673), .ZN(n6678) );
  OAI21_X1 U7642 ( .B1(n6679), .B2(n6694), .A(n6678), .ZN(U3202) );
  AOI22_X1 U7643 ( .A1(n6696), .A2(REIP_REG_21__SCAN_IN), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6673), .ZN(n6680) );
  OAI21_X1 U7644 ( .B1(n6682), .B2(n6698), .A(n6680), .ZN(U3204) );
  AOI22_X1 U7645 ( .A1(n6692), .A2(REIP_REG_23__SCAN_IN), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6673), .ZN(n6681) );
  OAI21_X1 U7646 ( .B1(n6682), .B2(n6694), .A(n6681), .ZN(U3205) );
  AOI22_X1 U7647 ( .A1(n6696), .A2(REIP_REG_23__SCAN_IN), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6673), .ZN(n6683) );
  OAI21_X1 U7648 ( .B1(n6684), .B2(n6698), .A(n6683), .ZN(U3206) );
  AOI22_X1 U7649 ( .A1(n6696), .A2(REIP_REG_24__SCAN_IN), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6673), .ZN(n6685) );
  OAI21_X1 U7650 ( .B1(n6687), .B2(n6698), .A(n6685), .ZN(U3207) );
  AOI22_X1 U7651 ( .A1(n6692), .A2(REIP_REG_26__SCAN_IN), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6673), .ZN(n6686) );
  OAI21_X1 U7652 ( .B1(n6687), .B2(n6694), .A(n6686), .ZN(U3208) );
  AOI22_X1 U7653 ( .A1(n6696), .A2(REIP_REG_26__SCAN_IN), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6673), .ZN(n6688) );
  OAI21_X1 U7654 ( .B1(n6689), .B2(n6698), .A(n6688), .ZN(U3209) );
  AOI22_X1 U7655 ( .A1(n6696), .A2(REIP_REG_27__SCAN_IN), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6673), .ZN(n6690) );
  OAI21_X1 U7656 ( .B1(n6873), .B2(n6698), .A(n6690), .ZN(U3210) );
  AOI22_X1 U7657 ( .A1(n6692), .A2(REIP_REG_29__SCAN_IN), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6673), .ZN(n6691) );
  OAI21_X1 U7658 ( .B1(n6873), .B2(n6694), .A(n6691), .ZN(U3211) );
  AOI22_X1 U7659 ( .A1(n6692), .A2(REIP_REG_30__SCAN_IN), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6673), .ZN(n6693) );
  OAI21_X1 U7660 ( .B1(n6695), .B2(n6694), .A(n6693), .ZN(U3212) );
  AOI22_X1 U7661 ( .A1(n6696), .A2(REIP_REG_30__SCAN_IN), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6673), .ZN(n6697) );
  OAI21_X1 U7662 ( .B1(n6699), .B2(n6698), .A(n6697), .ZN(U3213) );
  OAI21_X1 U7663 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6702), .A(n6701), .ZN(
        n6700) );
  INV_X1 U7664 ( .A(n6700), .ZN(U3451) );
  OAI21_X1 U7665 ( .B1(n6702), .B2(n6865), .A(n6701), .ZN(U3452) );
  NOR2_X1 U7666 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6709), .ZN(n6710) );
  AOI21_X1 U7667 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6710), .A(n6703), .ZN(
        n6707) );
  OAI21_X1 U7668 ( .B1(n4519), .B2(n4559), .A(n6705), .ZN(n6704) );
  OAI21_X1 U7669 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6705), .A(n6704), .ZN(
        n6706) );
  OAI21_X1 U7670 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6707), .A(n6706), .ZN(U3468)
         );
  AOI22_X1 U7671 ( .A1(n6710), .A2(n4559), .B1(n6709), .B2(n6708), .ZN(U3469)
         );
  INV_X1 U7672 ( .A(n6711), .ZN(n6717) );
  NAND2_X1 U7673 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6712), .ZN(n6720) );
  AOI21_X1 U7674 ( .B1(n6714), .B2(STATEBS16_REG_SCAN_IN), .A(n6713), .ZN(
        n6715) );
  AOI211_X1 U7675 ( .C1(n6717), .C2(n6716), .A(n6720), .B(n6715), .ZN(n6719)
         );
  OAI21_X1 U7676 ( .B1(n6719), .B2(n6722), .A(n6718), .ZN(n6727) );
  INV_X1 U7677 ( .A(n6720), .ZN(n6721) );
  AND3_X1 U7678 ( .A1(n6722), .A2(STATE2_REG_1__SCAN_IN), .A3(n6721), .ZN(
        n6723) );
  NOR4_X1 U7679 ( .A1(n6725), .A2(n6724), .A3(n6437), .A4(n6723), .ZN(n6726)
         );
  MUX2_X1 U7680 ( .A(n6727), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6726), .Z(
        U3472) );
  NAND3_X1 U7681 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(DATAI_12_), .A3(
        LWORD_REG_12__SCAN_IN), .ZN(n6728) );
  NOR4_X1 U7682 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n6728), .A3(
        PHYADDRPOINTER_REG_8__SCAN_IN), .A4(DATAI_13_), .ZN(n6729) );
  NAND3_X1 U7683 ( .A1(n6729), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .A3(n6770), 
        .ZN(n6730) );
  NOR3_X1 U7684 ( .A1(n6730), .A2(DATAO_REG_8__SCAN_IN), .A3(n6761), .ZN(n6734) );
  NOR4_X1 U7685 ( .A1(n6731), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .A3(
        EBX_REG_31__SCAN_IN), .A4(UWORD_REG_14__SCAN_IN), .ZN(n6732) );
  AND3_X1 U7686 ( .A1(n6734), .A2(n6733), .A3(n6732), .ZN(n6886) );
  NAND4_X1 U7687 ( .A1(DATAI_25_), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .A3(
        ADDRESS_REG_19__SCAN_IN), .A4(n6785), .ZN(n6738) );
  NAND4_X1 U7688 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        REIP_REG_3__SCAN_IN), .A3(LWORD_REG_15__SCAN_IN), .A4(n6789), .ZN(
        n6737) );
  INV_X1 U7689 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6801) );
  NAND4_X1 U7690 ( .A1(ADDRESS_REG_5__SCAN_IN), .A2(ADDRESS_REG_11__SCAN_IN), 
        .A3(n6801), .A4(n6794), .ZN(n6736) );
  NAND4_X1 U7691 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6805), .A3(n6808), 
        .A4(n6807), .ZN(n6735) );
  NOR4_X1 U7692 ( .A1(n6738), .A2(n6737), .A3(n6736), .A4(n6735), .ZN(n6745)
         );
  NOR4_X1 U7693 ( .A1(EAX_REG_2__SCAN_IN), .A2(DATAI_27_), .A3(n6839), .A4(
        n4255), .ZN(n6744) );
  INV_X1 U7694 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6842) );
  NOR4_X1 U7695 ( .A1(DATAI_23_), .A2(n6825), .A3(n6842), .A4(n6841), .ZN(
        n6743) );
  INV_X1 U7696 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6836) );
  NAND4_X1 U7697 ( .A1(STATE_REG_2__SCAN_IN), .A2(DATAI_7_), .A3(n6836), .A4(
        n6739), .ZN(n6741) );
  NAND2_X1 U7698 ( .A1(DATAO_REG_26__SCAN_IN), .A2(DATAO_REG_31__SCAN_IN), 
        .ZN(n6740) );
  NOR4_X1 U7699 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(
        ADDRESS_REG_14__SCAN_IN), .A3(n6741), .A4(n6740), .ZN(n6742) );
  NAND4_X1 U7700 ( .A1(n6745), .A2(n6744), .A3(n6743), .A4(n6742), .ZN(n6753)
         );
  NOR4_X1 U7701 ( .A1(M_IO_N_REG_SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), .A3(
        n6873), .A4(n6874), .ZN(n6748) );
  NOR4_X1 U7702 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .A3(EAX_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6747) );
  INV_X1 U7703 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6855) );
  NOR3_X1 U7704 ( .A1(EBX_REG_9__SCAN_IN), .A2(BE_N_REG_0__SCAN_IN), .A3(n6855), .ZN(n6746) );
  NAND4_X1 U7705 ( .A1(n6748), .A2(n6747), .A3(UWORD_REG_3__SCAN_IN), .A4(
        n6746), .ZN(n6752) );
  NAND4_X1 U7706 ( .A1(n6750), .A2(n6749), .A3(n6869), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6751) );
  NOR3_X1 U7707 ( .A1(n6753), .A2(n6752), .A3(n6751), .ZN(n6885) );
  AOI22_X1 U7708 ( .A1(n6756), .A2(keyinput59), .B1(n6755), .B2(keyinput32), 
        .ZN(n6754) );
  OAI221_X1 U7709 ( .B1(n6756), .B2(keyinput59), .C1(n6755), .C2(keyinput32), 
        .A(n6754), .ZN(n6768) );
  INV_X1 U7710 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n6758) );
  AOI22_X1 U7711 ( .A1(n6759), .A2(keyinput38), .B1(keyinput56), .B2(n6758), 
        .ZN(n6757) );
  OAI221_X1 U7712 ( .B1(n6759), .B2(keyinput38), .C1(n6758), .C2(keyinput56), 
        .A(n6757), .ZN(n6767) );
  XOR2_X1 U7713 ( .A(n6760), .B(keyinput40), .Z(n6765) );
  XOR2_X1 U7714 ( .A(n6761), .B(keyinput16), .Z(n6764) );
  XNOR2_X1 U7715 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .B(keyinput24), .ZN(n6763) );
  XNOR2_X1 U7716 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .B(keyinput47), .ZN(n6762)
         );
  NAND4_X1 U7717 ( .A1(n6765), .A2(n6764), .A3(n6763), .A4(n6762), .ZN(n6766)
         );
  NOR3_X1 U7718 ( .A1(n6768), .A2(n6767), .A3(n6766), .ZN(n6819) );
  INV_X1 U7719 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6771) );
  AOI22_X1 U7720 ( .A1(n6771), .A2(keyinput45), .B1(n6770), .B2(keyinput54), 
        .ZN(n6769) );
  OAI221_X1 U7721 ( .B1(n6771), .B2(keyinput45), .C1(n6770), .C2(keyinput54), 
        .A(n6769), .ZN(n6783) );
  AOI22_X1 U7722 ( .A1(n6731), .A2(keyinput53), .B1(keyinput12), .B2(n6773), 
        .ZN(n6772) );
  OAI221_X1 U7723 ( .B1(n6731), .B2(keyinput53), .C1(n6773), .C2(keyinput12), 
        .A(n6772), .ZN(n6782) );
  INV_X1 U7724 ( .A(DATAI_25_), .ZN(n6775) );
  AOI22_X1 U7725 ( .A1(n6776), .A2(keyinput26), .B1(keyinput28), .B2(n6775), 
        .ZN(n6774) );
  OAI221_X1 U7726 ( .B1(n6776), .B2(keyinput26), .C1(n6775), .C2(keyinput28), 
        .A(n6774), .ZN(n6781) );
  XOR2_X1 U7727 ( .A(n6777), .B(keyinput22), .Z(n6779) );
  XNOR2_X1 U7728 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .B(keyinput51), .ZN(n6778) );
  NAND2_X1 U7729 ( .A1(n6779), .A2(n6778), .ZN(n6780) );
  NOR4_X1 U7730 ( .A1(n6783), .A2(n6782), .A3(n6781), .A4(n6780), .ZN(n6818)
         );
  AOI22_X1 U7731 ( .A1(n6786), .A2(keyinput7), .B1(keyinput30), .B2(n6785), 
        .ZN(n6784) );
  OAI221_X1 U7732 ( .B1(n6786), .B2(keyinput7), .C1(n6785), .C2(keyinput30), 
        .A(n6784), .ZN(n6799) );
  AOI22_X1 U7733 ( .A1(n6789), .A2(keyinput63), .B1(n6788), .B2(keyinput15), 
        .ZN(n6787) );
  OAI221_X1 U7734 ( .B1(n6789), .B2(keyinput63), .C1(n6788), .C2(keyinput15), 
        .A(n6787), .ZN(n6798) );
  AOI22_X1 U7735 ( .A1(n6792), .A2(keyinput34), .B1(keyinput57), .B2(n6791), 
        .ZN(n6790) );
  OAI221_X1 U7736 ( .B1(n6792), .B2(keyinput34), .C1(n6791), .C2(keyinput57), 
        .A(n6790), .ZN(n6797) );
  AOI22_X1 U7737 ( .A1(n6795), .A2(keyinput11), .B1(n6794), .B2(keyinput10), 
        .ZN(n6793) );
  OAI221_X1 U7738 ( .B1(n6795), .B2(keyinput11), .C1(n6794), .C2(keyinput10), 
        .A(n6793), .ZN(n6796) );
  NOR4_X1 U7739 ( .A1(n6799), .A2(n6798), .A3(n6797), .A4(n6796), .ZN(n6817)
         );
  AOI22_X1 U7740 ( .A1(n6802), .A2(keyinput61), .B1(n6801), .B2(keyinput14), 
        .ZN(n6800) );
  OAI221_X1 U7741 ( .B1(n6802), .B2(keyinput61), .C1(n6801), .C2(keyinput14), 
        .A(n6800), .ZN(n6815) );
  AOI22_X1 U7742 ( .A1(n6805), .A2(keyinput48), .B1(keyinput18), .B2(n6804), 
        .ZN(n6803) );
  OAI221_X1 U7743 ( .B1(n6805), .B2(keyinput48), .C1(n6804), .C2(keyinput18), 
        .A(n6803), .ZN(n6814) );
  AOI22_X1 U7744 ( .A1(n6808), .A2(keyinput0), .B1(keyinput21), .B2(n6807), 
        .ZN(n6806) );
  OAI221_X1 U7745 ( .B1(n6808), .B2(keyinput0), .C1(n6807), .C2(keyinput21), 
        .A(n6806), .ZN(n6813) );
  INV_X1 U7746 ( .A(DATAI_27_), .ZN(n6811) );
  AOI22_X1 U7747 ( .A1(n6811), .A2(keyinput20), .B1(n6810), .B2(keyinput36), 
        .ZN(n6809) );
  OAI221_X1 U7748 ( .B1(n6811), .B2(keyinput20), .C1(n6810), .C2(keyinput36), 
        .A(n6809), .ZN(n6812) );
  NOR4_X1 U7749 ( .A1(n6815), .A2(n6814), .A3(n6813), .A4(n6812), .ZN(n6816)
         );
  NAND4_X1 U7750 ( .A1(n6819), .A2(n6818), .A3(n6817), .A4(n6816), .ZN(n6884)
         );
  AOI22_X1 U7751 ( .A1(n6822), .A2(keyinput62), .B1(keyinput35), .B2(n6821), 
        .ZN(n6820) );
  OAI221_X1 U7752 ( .B1(n6822), .B2(keyinput62), .C1(n6821), .C2(keyinput35), 
        .A(n6820), .ZN(n6834) );
  INV_X1 U7753 ( .A(DATAI_23_), .ZN(n6824) );
  AOI22_X1 U7754 ( .A1(n6825), .A2(keyinput8), .B1(keyinput25), .B2(n6824), 
        .ZN(n6823) );
  OAI221_X1 U7755 ( .B1(n6825), .B2(keyinput8), .C1(n6824), .C2(keyinput25), 
        .A(n6823), .ZN(n6833) );
  INV_X1 U7756 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6827) );
  AOI22_X1 U7757 ( .A1(n6828), .A2(keyinput37), .B1(n6827), .B2(keyinput13), 
        .ZN(n6826) );
  OAI221_X1 U7758 ( .B1(n6828), .B2(keyinput37), .C1(n6827), .C2(keyinput13), 
        .A(n6826), .ZN(n6832) );
  XOR2_X1 U7759 ( .A(n6750), .B(keyinput31), .Z(n6830) );
  XNOR2_X1 U7760 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .B(keyinput43), .ZN(n6829)
         );
  NAND2_X1 U7761 ( .A1(n6830), .A2(n6829), .ZN(n6831) );
  NOR4_X1 U7762 ( .A1(n6834), .A2(n6833), .A3(n6832), .A4(n6831), .ZN(n6882)
         );
  AOI22_X1 U7763 ( .A1(n6837), .A2(keyinput3), .B1(n6836), .B2(keyinput58), 
        .ZN(n6835) );
  OAI221_X1 U7764 ( .B1(n6837), .B2(keyinput3), .C1(n6836), .C2(keyinput58), 
        .A(n6835), .ZN(n6848) );
  AOI22_X1 U7765 ( .A1(n6839), .A2(keyinput27), .B1(n4255), .B2(keyinput2), 
        .ZN(n6838) );
  OAI221_X1 U7766 ( .B1(n6839), .B2(keyinput27), .C1(n4255), .C2(keyinput2), 
        .A(n6838), .ZN(n6847) );
  AOI22_X1 U7767 ( .A1(n6842), .A2(keyinput46), .B1(keyinput49), .B2(n6841), 
        .ZN(n6840) );
  OAI221_X1 U7768 ( .B1(n6842), .B2(keyinput46), .C1(n6841), .C2(keyinput49), 
        .A(n6840), .ZN(n6846) );
  XNOR2_X1 U7769 ( .A(STATE_REG_2__SCAN_IN), .B(keyinput4), .ZN(n6844) );
  XNOR2_X1 U7770 ( .A(keyinput17), .B(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6843)
         );
  NAND2_X1 U7771 ( .A1(n6844), .A2(n6843), .ZN(n6845) );
  NOR4_X1 U7772 ( .A1(n6848), .A2(n6847), .A3(n6846), .A4(n6845), .ZN(n6881)
         );
  AOI22_X1 U7773 ( .A1(n6851), .A2(keyinput60), .B1(n6850), .B2(keyinput33), 
        .ZN(n6849) );
  OAI221_X1 U7774 ( .B1(n6851), .B2(keyinput60), .C1(n6850), .C2(keyinput33), 
        .A(n6849), .ZN(n6863) );
  AOI22_X1 U7775 ( .A1(n6853), .A2(keyinput1), .B1(keyinput23), .B2(n4144), 
        .ZN(n6852) );
  OAI221_X1 U7776 ( .B1(n6853), .B2(keyinput1), .C1(n4144), .C2(keyinput23), 
        .A(n6852), .ZN(n6862) );
  AOI22_X1 U7777 ( .A1(n6856), .A2(keyinput6), .B1(n6855), .B2(keyinput9), 
        .ZN(n6854) );
  OAI221_X1 U7778 ( .B1(n6856), .B2(keyinput6), .C1(n6855), .C2(keyinput9), 
        .A(n6854), .ZN(n6861) );
  INV_X1 U7779 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6859) );
  AOI22_X1 U7780 ( .A1(n6859), .A2(keyinput44), .B1(keyinput42), .B2(n6858), 
        .ZN(n6857) );
  OAI221_X1 U7781 ( .B1(n6859), .B2(keyinput44), .C1(n6858), .C2(keyinput42), 
        .A(n6857), .ZN(n6860) );
  NOR4_X1 U7782 ( .A1(n6863), .A2(n6862), .A3(n6861), .A4(n6860), .ZN(n6880)
         );
  INV_X1 U7783 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6866) );
  AOI22_X1 U7784 ( .A1(n6866), .A2(keyinput39), .B1(keyinput41), .B2(n6865), 
        .ZN(n6864) );
  OAI221_X1 U7785 ( .B1(n6866), .B2(keyinput39), .C1(n6865), .C2(keyinput41), 
        .A(n6864), .ZN(n6878) );
  AOI22_X1 U7786 ( .A1(n6869), .A2(keyinput52), .B1(keyinput29), .B2(n6868), 
        .ZN(n6867) );
  OAI221_X1 U7787 ( .B1(n6869), .B2(keyinput52), .C1(n6868), .C2(keyinput29), 
        .A(n6867), .ZN(n6877) );
  AOI22_X1 U7788 ( .A1(n6871), .A2(keyinput19), .B1(n3991), .B2(keyinput5), 
        .ZN(n6870) );
  OAI221_X1 U7789 ( .B1(n6871), .B2(keyinput19), .C1(n3991), .C2(keyinput5), 
        .A(n6870), .ZN(n6876) );
  AOI22_X1 U7790 ( .A1(n6874), .A2(keyinput55), .B1(keyinput50), .B2(n6873), 
        .ZN(n6872) );
  OAI221_X1 U7791 ( .B1(n6874), .B2(keyinput55), .C1(n6873), .C2(keyinput50), 
        .A(n6872), .ZN(n6875) );
  NOR4_X1 U7792 ( .A1(n6878), .A2(n6877), .A3(n6876), .A4(n6875), .ZN(n6879)
         );
  NAND4_X1 U7793 ( .A1(n6882), .A2(n6881), .A3(n6880), .A4(n6879), .ZN(n6883)
         );
  AOI211_X1 U7794 ( .C1(n6886), .C2(n6885), .A(n6884), .B(n6883), .ZN(n6906)
         );
  INV_X1 U7795 ( .A(n6887), .ZN(n6891) );
  AOI22_X1 U7796 ( .A1(n6891), .A2(n6890), .B1(n6889), .B2(n6888), .ZN(n6904)
         );
  AOI221_X1 U7797 ( .B1(REIP_REG_10__SCAN_IN), .B2(REIP_REG_9__SCAN_IN), .C1(
        n5782), .C2(n6893), .A(n6892), .ZN(n6901) );
  AOI22_X1 U7798 ( .A1(n6895), .A2(EBX_REG_10__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n6894), .ZN(n6897) );
  OAI211_X1 U7799 ( .C1(n6899), .C2(n6898), .A(n6897), .B(n6896), .ZN(n6900)
         );
  AOI211_X1 U7800 ( .C1(n6902), .C2(REIP_REG_10__SCAN_IN), .A(n6901), .B(n6900), .ZN(n6903) );
  NAND2_X1 U7801 ( .A1(n6904), .A2(n6903), .ZN(n6905) );
  XOR2_X1 U7802 ( .A(n6906), .B(n6905), .Z(U2817) );
  AND4_X1 U3442 ( .A1(n3311), .A2(n3310), .A3(n3309), .A4(n3308), .ZN(n3312)
         );
  CLKBUF_X1 U3443 ( .A(n3455), .Z(n3857) );
  NAND2_X2 U3450 ( .A1(n3313), .A2(n3312), .ZN(n3426) );
  CLKBUF_X1 U34600 ( .A(n3400), .Z(n2972) );
  CLKBUF_X1 U34640 ( .A(n3108), .Z(n2970) );
  CLKBUF_X1 U3546 ( .A(n3908), .Z(n4369) );
  CLKBUF_X2 U3700 ( .A(n3421), .Z(n3530) );
  CLKBUF_X1 U4122 ( .A(n5260), .Z(n5272) );
  CLKBUF_X1 U4399 ( .A(n3856), .Z(n6021) );
  INV_X1 U4400 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4472) );
endmodule

