

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, 
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, 
        keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, 
        keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, 
        keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, 
        keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, 
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, 
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, 
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, 
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, 
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, 
        keyinput124, keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183;

  INV_X1 U3561 ( .A(n6463), .ZN(n6449) );
  NAND2_X1 U3562 ( .A1(n3859), .A2(n3858), .ZN(n4951) );
  INV_X1 U3563 ( .A(n5638), .ZN(n5626) );
  OR2_X1 U3564 ( .A1(n4340), .A2(n5456), .ZN(n4442) );
  CLKBUF_X2 U3565 ( .A(n3536), .Z(n3478) );
  CLKBUF_X1 U3566 ( .A(n3421), .Z(n4333) );
  INV_X1 U3567 ( .A(n3434), .ZN(n3590) );
  CLKBUF_X1 U3568 ( .A(n3450), .Z(n3786) );
  INV_X1 U3570 ( .A(n3427), .ZN(n4334) );
  AND2_X1 U3571 ( .A1(n3432), .A2(n3155), .ZN(n3477) );
  OR2_X1 U3572 ( .A1(n4830), .A2(n3603), .ZN(n3609) );
  AND2_X2 U3573 ( .A1(n3307), .A2(n4715), .ZN(n3479) );
  INV_X1 U3574 ( .A(n4360), .ZN(n4800) );
  NAND2_X1 U3575 ( .A1(n3609), .A2(n3608), .ZN(n4774) );
  NAND2_X1 U3576 ( .A1(n5526), .A2(n5525), .ZN(n5528) );
  NOR2_X1 U3577 ( .A1(n7064), .A2(n3848), .ZN(n3863) );
  AND2_X1 U3578 ( .A1(n3612), .A2(n3613), .ZN(n4779) );
  OR2_X1 U3579 ( .A1(n4755), .A2(n5363), .ZN(n6545) );
  INV_X2 U3580 ( .A(n3710), .ZN(n3113) );
  XNOR2_X2 U3581 ( .A(n3522), .B(n3523), .ZN(n3587) );
  NAND2_X2 U3582 ( .A1(n3476), .A2(n3475), .ZN(n3522) );
  OAI22_X2 U3583 ( .A1(n3734), .A2(n3735), .B1(n3732), .B2(n3746), .ZN(n3739)
         );
  OAI21_X1 U3584 ( .B1(n4460), .B2(n5524), .A(n5523), .ZN(n5869) );
  NAND2_X1 U3585 ( .A1(n3857), .A2(n4816), .ZN(n4817) );
  NOR2_X1 U3586 ( .A1(n3441), .A2(n3440), .ZN(n3442) );
  NOR2_X1 U3587 ( .A1(n3431), .A2(n3430), .ZN(n4332) );
  NAND2_X1 U3589 ( .A1(n3355), .A2(n3300), .ZN(n3209) );
  OR2_X1 U3590 ( .A1(n3783), .A2(n3182), .ZN(n3446) );
  NAND3_X1 U3592 ( .A1(n3124), .A2(n3354), .A3(n3353), .ZN(n4340) );
  CLKBUF_X2 U3593 ( .A(n3467), .Z(n4254) );
  BUF_X2 U3594 ( .A(n3537), .Z(n4280) );
  CLKBUF_X2 U3595 ( .A(n3484), .Z(n4253) );
  AND2_X2 U3596 ( .A1(n4720), .A2(n4895), .ZN(n3467) );
  AND2_X2 U3597 ( .A1(n3308), .A2(n3310), .ZN(n3392) );
  NAND2_X1 U3598 ( .A1(n6345), .A2(n4909), .ZN(n6722) );
  XNOR2_X1 U3599 ( .A(n3210), .B(n6184), .ZN(n6177) );
  OR2_X1 U3600 ( .A1(n5918), .A2(n3251), .ZN(n3249) );
  AND2_X1 U3601 ( .A1(n4469), .A2(n4468), .ZN(n5804) );
  OAI21_X1 U3602 ( .B1(n5869), .B2(n6054), .A(n5868), .ZN(n3146) );
  OR2_X1 U3603 ( .A1(n5971), .A2(n5975), .ZN(n3210) );
  CLKBUF_X1 U3604 ( .A(n4466), .Z(n5523) );
  NAND2_X1 U3605 ( .A1(n3151), .A2(n3715), .ZN(n5954) );
  NAND2_X1 U3606 ( .A1(n3239), .A2(n3237), .ZN(n3151) );
  OAI21_X1 U3607 ( .B1(n5993), .B2(n3272), .A(n3274), .ZN(n3720) );
  AOI21_X1 U3608 ( .B1(n5492), .B2(n6439), .A(n3159), .ZN(n3158) );
  NAND2_X1 U3609 ( .A1(n4452), .A2(n5626), .ZN(n4517) );
  OR2_X1 U3610 ( .A1(n3936), .A2(n3935), .ZN(n3951) );
  AND2_X1 U3611 ( .A1(n6134), .A2(n5899), .ZN(n6117) );
  AND3_X1 U3612 ( .A1(n3178), .A2(n3288), .A3(n5761), .ZN(n3173) );
  AND2_X1 U3613 ( .A1(n6140), .A2(n6142), .ZN(n6134) );
  OR2_X1 U3614 ( .A1(n4223), .A2(n4222), .ZN(n4266) );
  NAND2_X1 U3615 ( .A1(n3638), .A2(n3637), .ZN(n3639) );
  XNOR2_X1 U3616 ( .A(n3654), .B(n3662), .ZN(n3787) );
  NAND2_X1 U3617 ( .A1(n3579), .A2(n3578), .ZN(n3620) );
  CLKBUF_X1 U3618 ( .A(n3835), .Z(n6287) );
  NAND2_X1 U3619 ( .A1(n3856), .A2(n3855), .ZN(n4816) );
  NAND2_X1 U3620 ( .A1(n3641), .A2(n3663), .ZN(n3654) );
  NAND2_X1 U3621 ( .A1(n3680), .A2(n3679), .ZN(n3678) );
  XNOR2_X1 U3622 ( .A(n3621), .B(n4913), .ZN(n3835) );
  AND2_X1 U3623 ( .A1(n4782), .A2(n4781), .ZN(n4784) );
  NAND3_X1 U3624 ( .A1(n3552), .A2(n3580), .A3(n4913), .ZN(n3665) );
  CLKBUF_X1 U3625 ( .A(n4828), .Z(n6283) );
  NAND2_X1 U3626 ( .A1(n3575), .A2(n3574), .ZN(n4913) );
  NAND2_X1 U3627 ( .A1(n6218), .A2(n6221), .ZN(n6651) );
  AND2_X1 U3628 ( .A1(n5498), .A2(n4406), .ZN(n5703) );
  CLKBUF_X1 U3629 ( .A(n3839), .Z(n6278) );
  CLKBUF_X1 U3630 ( .A(n4329), .Z(n5839) );
  OR2_X1 U3631 ( .A1(n4537), .A2(n4731), .ZN(n6238) );
  AOI21_X1 U3632 ( .B1(n4728), .B2(n6938), .A(n3548), .ZN(n3551) );
  NAND2_X1 U3633 ( .A1(n3555), .A2(n3554), .ZN(n4692) );
  NAND2_X2 U3634 ( .A1(n6481), .A2(n4853), .ZN(n5802) );
  XNOR2_X1 U3635 ( .A(n3528), .B(n3283), .ZN(n4711) );
  CLKBUF_X2 U3636 ( .A(n3495), .Z(n3498) );
  NAND2_X1 U3637 ( .A1(n3442), .A2(n4332), .ZN(n3496) );
  OAI21_X1 U3638 ( .B1(n3772), .B2(n3764), .A(n3477), .ZN(n3775) );
  NAND2_X1 U3639 ( .A1(n3777), .A2(n4318), .ZN(n3778) );
  NAND2_X1 U3640 ( .A1(n3520), .A2(n3519), .ZN(n3600) );
  AND2_X1 U3641 ( .A1(n4493), .A2(n4698), .ZN(n3430) );
  AND3_X1 U3642 ( .A1(n3494), .A2(n3493), .A3(n3492), .ZN(n3523) );
  AND2_X1 U3643 ( .A1(n4800), .A2(n4371), .ZN(n4378) );
  NAND4_X1 U3644 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3447)
         );
  OR2_X1 U3645 ( .A1(n4321), .A2(n4488), .ZN(n4509) );
  CLKBUF_X1 U3646 ( .A(n4334), .Z(n4843) );
  AND2_X1 U3647 ( .A1(n3416), .A2(n4353), .ZN(n3443) );
  AND2_X1 U3648 ( .A1(n3386), .A2(n4353), .ZN(n3389) );
  OR2_X1 U3649 ( .A1(n4333), .A2(n3433), .ZN(n4347) );
  NOR2_X1 U3650 ( .A1(n4335), .A2(n3591), .ZN(n3782) );
  AND2_X1 U3651 ( .A1(n3182), .A2(n3435), .ZN(n3434) );
  NAND2_X1 U3652 ( .A1(n4334), .A2(n4340), .ZN(n3591) );
  OR2_X1 U3653 ( .A1(n3512), .A2(n3511), .ZN(n3606) );
  OR2_X1 U3654 ( .A1(n3490), .A2(n3489), .ZN(n3699) );
  CLKBUF_X2 U3655 ( .A(n3391), .Z(n5455) );
  NAND2_X1 U3656 ( .A1(n3474), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3562) );
  NAND2_X1 U3657 ( .A1(n5456), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3561) );
  NAND3_X1 U3658 ( .A1(n3316), .A2(n3315), .A3(n3314), .ZN(n3391) );
  AND4_X2 U3659 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3474)
         );
  AND3_X2 U3660 ( .A1(n3365), .A2(n3114), .A3(n3364), .ZN(n3436) );
  OR2_X1 U3661 ( .A1(n3385), .A2(n3384), .ZN(n3427) );
  AND4_X1 U3662 ( .A1(n3306), .A2(n3305), .A3(n3304), .A4(n3303), .ZN(n3316)
         );
  AND4_X1 U3663 ( .A1(n3329), .A2(n3328), .A3(n3327), .A4(n3326), .ZN(n3345)
         );
  AND4_X1 U3664 ( .A1(n3337), .A2(n3336), .A3(n3335), .A4(n3334), .ZN(n3343)
         );
  AND4_X1 U3665 ( .A1(n3333), .A2(n3332), .A3(n3331), .A4(n3330), .ZN(n3344)
         );
  AND4_X1 U3666 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3414)
         );
  AND4_X1 U3667 ( .A1(n3341), .A2(n3340), .A3(n3339), .A4(n3338), .ZN(n3342)
         );
  AND4_X1 U3668 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3413)
         );
  AND4_X1 U3669 ( .A1(n3410), .A2(n3409), .A3(n3408), .A4(n3407), .ZN(n3411)
         );
  BUF_X2 U3670 ( .A(n3392), .Z(n4270) );
  AND4_X1 U3671 ( .A1(n3404), .A2(n3403), .A3(n3402), .A4(n3401), .ZN(n3412)
         );
  AND3_X1 U3672 ( .A1(n3313), .A2(n3312), .A3(n3311), .ZN(n3314) );
  AND4_X1 U3673 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3365)
         );
  AND4_X1 U3674 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3325)
         );
  AOI22_X1 U3675 ( .A1(n3405), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U3676 ( .A1(n3567), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3360) );
  BUF_X2 U3677 ( .A(n3479), .Z(n3500) );
  BUF_X2 U3678 ( .A(n3499), .Z(n4203) );
  BUF_X2 U3679 ( .A(n3567), .Z(n3506) );
  BUF_X2 U3680 ( .A(n3505), .Z(n4269) );
  AND2_X2 U3681 ( .A1(n4881), .A2(n4715), .ZN(n3536) );
  AND2_X2 U3682 ( .A1(n4720), .A2(n4881), .ZN(n3567) );
  NAND2_X2 U3683 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6825), .ZN(n4639) );
  AND2_X2 U3684 ( .A1(n3308), .A2(n3307), .ZN(n3505) );
  AND2_X2 U3685 ( .A1(n4720), .A2(n3307), .ZN(n3499) );
  AND2_X2 U3686 ( .A1(n3308), .A2(n4895), .ZN(n3537) );
  BUF_X2 U3687 ( .A(n3461), .Z(n4251) );
  AND2_X2 U3688 ( .A1(n3302), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3308)
         );
  AND2_X2 U3689 ( .A1(n3309), .A2(n3310), .ZN(n3461) );
  AND2_X2 U3690 ( .A1(n3301), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4881)
         );
  CLKBUF_X1 U3692 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n4749) );
  AND2_X2 U3693 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4715) );
  INV_X2 U3694 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3757) );
  AOI21_X1 U3695 ( .B1(n5550), .B2(n5548), .A(n5549), .ZN(n5883) );
  NAND2_X4 U3696 ( .A1(n3602), .A2(n3601), .ZN(n4830) );
  NAND2_X4 U3697 ( .A1(n3182), .A2(n5455), .ZN(n4360) );
  XNOR2_X2 U3698 ( .A(n3620), .B(n6640), .ZN(n4950) );
  OR2_X1 U3699 ( .A1(n4537), .A2(n4878), .ZN(n6218) );
  NAND2_X1 U3700 ( .A1(n3130), .A2(n3715), .ZN(n3276) );
  INV_X1 U3701 ( .A(n3589), .ZN(n3491) );
  AND2_X1 U3704 ( .A1(n5297), .A2(n3834), .ZN(n3178) );
  NAND2_X1 U3705 ( .A1(n3633), .A2(n3632), .ZN(n3663) );
  CLKBUF_X1 U3706 ( .A(n3405), .Z(n4271) );
  NOR2_X1 U3707 ( .A1(n3716), .A2(n3128), .ZN(n3277) );
  AOI22_X1 U3708 ( .A1(n3477), .A2(n4333), .B1(n3422), .B2(n5455), .ZN(n3423)
         );
  NAND2_X1 U3709 ( .A1(n3495), .A2(n3496), .ZN(n3199) );
  INV_X1 U3710 ( .A(n4175), .ZN(n4289) );
  NAND2_X1 U3711 ( .A1(n3135), .A2(n5496), .ZN(n3287) );
  AND2_X1 U3712 ( .A1(n3985), .A2(n3968), .ZN(n3969) );
  NOR2_X1 U3713 ( .A1(n4347), .A2(n6938), .ZN(n4175) );
  NAND2_X1 U3714 ( .A1(n3710), .A2(n3703), .ZN(n3704) );
  INV_X1 U3715 ( .A(n5925), .ZN(n3252) );
  INV_X1 U3716 ( .A(n3260), .ZN(n3152) );
  NAND2_X1 U3717 ( .A1(n3154), .A2(n3153), .ZN(n3202) );
  NAND2_X1 U3718 ( .A1(n3205), .A2(n3115), .ZN(n3153) );
  NOR2_X1 U3719 ( .A1(n3591), .A2(n4328), .ZN(n3444) );
  AOI21_X1 U3720 ( .B1(n3597), .B2(n3600), .A(n3521), .ZN(n3586) );
  AND3_X1 U3721 ( .A1(n3352), .A2(n3351), .A3(n3350), .ZN(n3354) );
  NAND2_X1 U3722 ( .A1(n6433), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5458) );
  AND2_X1 U3723 ( .A1(n3449), .A2(n4334), .ZN(n4349) );
  NOR2_X1 U3724 ( .A1(n4340), .A2(n3448), .ZN(n3449) );
  NAND2_X1 U3725 ( .A1(n3186), .A2(n5572), .ZN(n3185) );
  INV_X1 U3726 ( .A(n3187), .ZN(n3186) );
  INV_X1 U3727 ( .A(n3720), .ZN(n5864) );
  AND3_X1 U3728 ( .A1(n3197), .A2(n4545), .A3(n6157), .ZN(n6137) );
  NAND2_X1 U3729 ( .A1(n6155), .A2(n6156), .ZN(n3197) );
  INV_X1 U3730 ( .A(n3113), .ZN(n6020) );
  NAND2_X1 U3731 ( .A1(n4506), .A2(n6355), .ZN(n4537) );
  CLKBUF_X1 U3732 ( .A(n4486), .Z(n4487) );
  OR2_X1 U3733 ( .A1(n6287), .A2(n6283), .ZN(n5107) );
  NAND2_X1 U3734 ( .A1(n3161), .A2(n3160), .ZN(n3159) );
  INV_X1 U3735 ( .A(n5489), .ZN(n3160) );
  OR2_X1 U3736 ( .A1(n6080), .A2(n5802), .ZN(n4566) );
  NAND2_X1 U3737 ( .A1(n3182), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3730) );
  INV_X1 U3738 ( .A(n3783), .ZN(n3355) );
  AOI22_X1 U3739 ( .A1(n3567), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3383) );
  OR2_X1 U3740 ( .A1(n4121), .A2(n4120), .ZN(n4140) );
  OR2_X1 U3741 ( .A1(n3473), .A2(n3472), .ZN(n3589) );
  NAND2_X1 U3742 ( .A1(n5510), .A2(n3179), .ZN(n3428) );
  CLKBUF_X1 U3743 ( .A(n3529), .Z(n3530) );
  AOI22_X1 U3744 ( .A1(n3537), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3479), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U3745 ( .A1(n3499), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3322) );
  NAND2_X1 U3746 ( .A1(n3221), .A2(n4369), .ZN(n3220) );
  INV_X1 U3747 ( .A(n5548), .ZN(n3293) );
  OR2_X1 U3748 ( .A1(n4169), .A2(n4168), .ZN(n4182) );
  NAND2_X1 U3749 ( .A1(n3132), .A2(n3188), .ZN(n3187) );
  INV_X1 U3750 ( .A(n5623), .ZN(n3188) );
  INV_X1 U3751 ( .A(n3281), .ZN(n3280) );
  INV_X1 U3752 ( .A(n3815), .ZN(n4197) );
  NOR2_X1 U3753 ( .A1(n4019), .A2(n3967), .ZN(n3985) );
  AND2_X1 U3754 ( .A1(n3289), .A2(n3891), .ZN(n3288) );
  NOR2_X1 U3755 ( .A1(n5472), .A2(n3290), .ZN(n3289) );
  INV_X1 U3756 ( .A(n4294), .ZN(n4154) );
  NOR2_X2 U3757 ( .A1(n3786), .A2(n6345), .ZN(n4030) );
  AND2_X1 U3758 ( .A1(n3299), .A2(n3270), .ZN(n3269) );
  INV_X1 U3759 ( .A(n6089), .ZN(n3270) );
  AND2_X1 U3760 ( .A1(n5563), .A2(n3230), .ZN(n3229) );
  INV_X1 U3761 ( .A(n5551), .ZN(n3230) );
  NAND2_X1 U3762 ( .A1(n3278), .A2(n3273), .ZN(n3272) );
  INV_X1 U3763 ( .A(n3275), .ZN(n3274) );
  INV_X1 U3764 ( .A(n5599), .ZN(n3216) );
  NAND2_X1 U3765 ( .A1(n5944), .A2(n3256), .ZN(n3255) );
  NOR2_X1 U3766 ( .A1(n5995), .A2(n3241), .ZN(n3240) );
  INV_X1 U3767 ( .A(n3711), .ZN(n3241) );
  NOR2_X1 U3768 ( .A1(n5737), .A2(n5719), .ZN(n5498) );
  INV_X1 U3769 ( .A(n4378), .ZN(n4441) );
  OR2_X1 U3770 ( .A1(n5427), .A2(n6247), .ZN(n3233) );
  NAND2_X1 U3771 ( .A1(n3678), .A2(n3700), .ZN(n3710) );
  INV_X1 U3772 ( .A(n3698), .ZN(n3265) );
  AND2_X1 U3773 ( .A1(n5292), .A2(n6428), .ZN(n3221) );
  AND2_X1 U3774 ( .A1(n4976), .A2(n5476), .ZN(n4370) );
  INV_X1 U3775 ( .A(n5477), .ZN(n4369) );
  AND2_X1 U3776 ( .A1(n5455), .A2(n4328), .ZN(n3763) );
  NOR2_X1 U3777 ( .A1(n5456), .A2(n6938), .ZN(n3155) );
  NAND2_X1 U3778 ( .A1(n3699), .A2(n3474), .ZN(n3517) );
  NAND2_X1 U3779 ( .A1(n3526), .A2(n3525), .ZN(n3581) );
  OR2_X1 U3780 ( .A1(n3522), .A2(n3524), .ZN(n3525) );
  XNOR2_X1 U3781 ( .A(n4692), .B(n4691), .ZN(n4831) );
  NAND2_X1 U3782 ( .A1(n3198), .A2(n3527), .ZN(n3553) );
  AND2_X1 U3783 ( .A1(n3556), .A2(n4943), .ZN(n5145) );
  NAND2_X1 U3784 ( .A1(n4394), .A2(n3294), .ZN(n5797) );
  XNOR2_X1 U3785 ( .A(n4298), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5426)
         );
  NOR2_X1 U3786 ( .A1(n4297), .A2(n6918), .ZN(n4298) );
  OR2_X1 U3787 ( .A1(n4266), .A2(n5517), .ZN(n4297) );
  AND2_X1 U3788 ( .A1(n4244), .A2(n4243), .ZN(n5524) );
  OR2_X1 U3789 ( .A1(n4137), .A2(n4153), .ZN(n4177) );
  NAND2_X1 U3790 ( .A1(n4109), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4137)
         );
  INV_X1 U3791 ( .A(n4110), .ZN(n4109) );
  NAND2_X1 U3792 ( .A1(n4055), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4092)
         );
  NOR2_X1 U3793 ( .A1(n3287), .A2(n3286), .ZN(n3285) );
  INV_X1 U3794 ( .A(n5636), .ZN(n3286) );
  NAND2_X1 U3795 ( .A1(n3969), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4053)
         );
  NAND2_X1 U3796 ( .A1(n6557), .A2(n3689), .ZN(n6065) );
  NAND2_X1 U3797 ( .A1(n3794), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3869)
         );
  INV_X1 U3798 ( .A(n4952), .ZN(n3859) );
  OR2_X1 U3799 ( .A1(n4496), .A2(n3783), .ZN(n5351) );
  NAND2_X1 U3800 ( .A1(n4709), .A2(n6355), .ZN(n4755) );
  AND2_X1 U3801 ( .A1(n3269), .A2(n4536), .ZN(n3268) );
  NAND2_X1 U3802 ( .A1(n6078), .A2(n4554), .ZN(n6071) );
  NOR2_X2 U3803 ( .A1(n5587), .A2(n5575), .ZN(n5574) );
  AOI21_X1 U3804 ( .B1(n3250), .B2(n3257), .A(INSTADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n3248) );
  AND2_X1 U3805 ( .A1(n3250), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3245)
         );
  NOR2_X1 U3806 ( .A1(n5919), .A2(n6133), .ZN(n3246) );
  AND2_X1 U3807 ( .A1(n4417), .A2(n4416), .ZN(n5642) );
  INV_X1 U3808 ( .A(n5953), .ZN(n5895) );
  INV_X1 U3809 ( .A(n5954), .ZN(n5896) );
  NAND2_X1 U3810 ( .A1(n3214), .A2(n3213), .ZN(n5674) );
  INV_X1 U3811 ( .A(n5672), .ZN(n3213) );
  INV_X1 U3812 ( .A(n5686), .ZN(n3214) );
  AND2_X1 U3813 ( .A1(n5703), .A2(n5702), .ZN(n5705) );
  XNOR2_X1 U3814 ( .A(n6018), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6011)
         );
  NAND3_X1 U3815 ( .A1(n3261), .A2(n3263), .A3(n3705), .ZN(n3260) );
  INV_X1 U3816 ( .A(n3709), .ZN(n3263) );
  INV_X1 U3817 ( .A(n6063), .ZN(n3262) );
  NAND2_X1 U3818 ( .A1(n3131), .A2(n3259), .ZN(n3258) );
  INV_X2 U3819 ( .A(n3113), .ZN(n6018) );
  AND2_X1 U3820 ( .A1(n6268), .A2(n4532), .ZN(n6220) );
  NAND2_X1 U3821 ( .A1(n3234), .A2(n3640), .ZN(n5053) );
  NOR2_X1 U3822 ( .A1(n6645), .A2(n4538), .ZN(n6216) );
  INV_X1 U3823 ( .A(n5306), .ZN(n5019) );
  CLKBUF_X1 U3824 ( .A(n4711), .Z(n4712) );
  CLKBUF_X1 U3825 ( .A(n4831), .Z(n4832) );
  INV_X1 U3826 ( .A(n5107), .ZN(n5100) );
  AND2_X1 U3827 ( .A1(n5015), .A2(n5216), .ZN(n6660) );
  AND2_X1 U3828 ( .A1(n6283), .A2(n4981), .ZN(n5015) );
  AND2_X1 U3829 ( .A1(n6278), .A2(n6659), .ZN(n5016) );
  AND2_X1 U3830 ( .A1(n4728), .A2(n6280), .ZN(n5149) );
  AND2_X1 U3831 ( .A1(n5022), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6713) );
  AND3_X1 U3832 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n5387) );
  AOI21_X1 U3833 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6718), .A(n5019), .ZN(
        n6668) );
  AND2_X1 U3834 ( .A1(n5357), .A2(n4898), .ZN(n4905) );
  OR2_X1 U3835 ( .A1(n5488), .A2(n5487), .ZN(n3162) );
  NAND2_X1 U3836 ( .A1(n3129), .A2(n3165), .ZN(n5678) );
  INV_X1 U3837 ( .A(n5706), .ZN(n3165) );
  INV_X1 U3838 ( .A(n6424), .ZN(n6411) );
  OR2_X1 U3839 ( .A1(n5458), .A2(n4585), .ZN(n6452) );
  NAND2_X1 U3840 ( .A1(n4455), .A2(n4454), .ZN(n6073) );
  OR3_X1 U3841 ( .A1(n4709), .A2(n6365), .A3(n4731), .ZN(n4352) );
  NOR2_X2 U3842 ( .A1(n5850), .A2(n4488), .ZN(n5838) );
  NAND2_X1 U3843 ( .A1(n4326), .A2(n6516), .ZN(n5856) );
  AOI21_X1 U3844 ( .B1(n4687), .B2(n6355), .A(n4324), .ZN(n4326) );
  INV_X1 U3845 ( .A(n5851), .ZN(n5860) );
  INV_X2 U3846 ( .A(n5856), .ZN(n5850) );
  XNOR2_X1 U3847 ( .A(n4310), .B(n4296), .ZN(n4584) );
  INV_X1 U3848 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6918) );
  INV_X1 U3849 ( .A(n6586), .ZN(n5979) );
  OR2_X1 U3850 ( .A1(n4755), .A2(n5351), .ZN(n6372) );
  INV_X1 U3851 ( .A(n5981), .ZN(n6578) );
  XNOR2_X1 U3852 ( .A(n4520), .B(n4519), .ZN(n5777) );
  OAI21_X1 U3853 ( .B1(n4518), .B2(n4561), .A(n4517), .ZN(n4520) );
  INV_X1 U3854 ( .A(n3194), .ZN(n3193) );
  OAI21_X1 U3855 ( .B1(n6073), .B2(n6252), .A(n6072), .ZN(n3194) );
  NAND2_X1 U3856 ( .A1(n6071), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3195) );
  XNOR2_X1 U3857 ( .A(n4575), .B(n4574), .ZN(n6076) );
  AOI21_X1 U3858 ( .B1(n4573), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4572), 
        .ZN(n4575) );
  NAND2_X1 U3859 ( .A1(n4561), .A2(n3227), .ZN(n6080) );
  OR2_X1 U3860 ( .A1(n4563), .A2(n4562), .ZN(n3227) );
  NAND2_X1 U3861 ( .A1(n3150), .A2(n3149), .ZN(n3148) );
  NAND2_X1 U3862 ( .A1(n5865), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U3863 ( .A1(n5871), .A2(n5866), .ZN(n3150) );
  NAND2_X1 U3864 ( .A1(n6130), .A2(n4549), .ZN(n6124) );
  OR2_X1 U3865 ( .A1(n6178), .A2(n6184), .ZN(n6172) );
  OR2_X1 U3866 ( .A1(n4537), .A2(n4511), .ZN(n6275) );
  NAND2_X1 U3867 ( .A1(n4508), .A2(n3142), .ZN(n4510) );
  INV_X1 U3868 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6718) );
  INV_X1 U3869 ( .A(n6722), .ZN(n6304) );
  OAI21_X1 U3870 ( .B1(n6337), .B2(n6312), .A(n6311), .ZN(n6336) );
  NAND2_X1 U3871 ( .A1(n5015), .A2(n5016), .ZN(n5222) );
  INV_X1 U3872 ( .A(n3180), .ZN(n3179) );
  OAI21_X1 U3873 ( .B1(n3783), .B2(n3182), .A(n3181), .ZN(n3180) );
  NAND2_X1 U3874 ( .A1(n3182), .A2(n4334), .ZN(n3181) );
  INV_X1 U3875 ( .A(n5731), .ZN(n3290) );
  OAI21_X1 U3876 ( .B1(n3277), .B2(n3276), .A(n3719), .ZN(n3275) );
  INV_X1 U3877 ( .A(n3276), .ZN(n3273) );
  OR2_X1 U3878 ( .A1(n3675), .A2(n3674), .ZN(n3692) );
  INV_X1 U3879 ( .A(n3665), .ZN(n3641) );
  OR2_X1 U3880 ( .A1(n3491), .A2(n3562), .ZN(n3475) );
  NAND2_X1 U3881 ( .A1(n3459), .A2(n3297), .ZN(n3200) );
  AND2_X2 U3882 ( .A1(n3757), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3307)
         );
  INV_X1 U3883 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3302) );
  OR2_X1 U3884 ( .A1(n3573), .A2(n3572), .ZN(n3634) );
  NAND2_X1 U3885 ( .A1(n3192), .A2(n3751), .ZN(n3772) );
  OR2_X1 U3886 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  OAI21_X1 U3887 ( .B1(n3741), .B2(n3740), .A(n3748), .ZN(n3192) );
  NAND2_X1 U3888 ( .A1(n3293), .A2(n3291), .ZN(n4466) );
  AND2_X1 U3889 ( .A1(n5524), .A2(n3292), .ZN(n3291) );
  NOR2_X1 U3890 ( .A1(n4459), .A2(n5550), .ZN(n3292) );
  OR2_X1 U3891 ( .A1(n3282), .A2(n5597), .ZN(n3281) );
  INV_X1 U3892 ( .A(n3138), .ZN(n3282) );
  NAND2_X1 U3893 ( .A1(n3912), .A2(n3911), .ZN(n3929) );
  INV_X1 U3894 ( .A(n3910), .ZN(n3912) );
  NOR2_X1 U3895 ( .A1(n3176), .A2(n3175), .ZN(n3892) );
  NAND2_X1 U3896 ( .A1(n3178), .A2(n5761), .ZN(n3175) );
  NAND2_X1 U3897 ( .A1(n3120), .A2(n3174), .ZN(n3176) );
  NOR2_X1 U3898 ( .A1(n3547), .A2(n3546), .ZN(n3582) );
  INV_X1 U3899 ( .A(n3860), .ZN(n3852) );
  CLKBUF_X1 U3900 ( .A(n3815), .Z(n4240) );
  OR3_X1 U3901 ( .A1(n6020), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n6090), 
        .ZN(n4472) );
  AOI21_X1 U3902 ( .B1(n3240), .B2(n3712), .A(n3238), .ZN(n3237) );
  INV_X1 U3903 ( .A(n3277), .ZN(n3238) );
  OR2_X1 U3904 ( .A1(n6018), .A2(n6002), .ZN(n3711) );
  INV_X1 U3905 ( .A(n3712), .ZN(n3203) );
  INV_X1 U3906 ( .A(n3209), .ZN(n4343) );
  NAND2_X1 U3907 ( .A1(n3620), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3236)
         );
  INV_X1 U3908 ( .A(n4442), .ZN(n4430) );
  AND3_X1 U3909 ( .A1(n4493), .A2(n5455), .A3(n4347), .ZN(n3441) );
  NAND2_X1 U3910 ( .A1(n3439), .A2(n3122), .ZN(n3440) );
  INV_X1 U3911 ( .A(n3199), .ZN(n3283) );
  NAND2_X1 U3912 ( .A1(n3527), .A2(n3200), .ZN(n3528) );
  INV_X1 U3913 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3301) );
  NAND2_X2 U3914 ( .A1(n3474), .A2(n3448), .ZN(n3783) );
  OAI21_X1 U3915 ( .B1(n3427), .B2(n3474), .A(n4322), .ZN(n3390) );
  NAND2_X1 U3916 ( .A1(n3560), .A2(n3559), .ZN(n4691) );
  INV_X1 U3917 ( .A(n6278), .ZN(n5216) );
  AND2_X1 U3918 ( .A1(n3768), .A2(n3767), .ZN(n4318) );
  OR2_X1 U3919 ( .A1(n3766), .A2(n3765), .ZN(n3768) );
  AND2_X1 U3920 ( .A1(n7116), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3765)
         );
  NAND2_X1 U3921 ( .A1(n3477), .A2(n3763), .ZN(n3776) );
  AND2_X2 U3922 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4895) );
  AND2_X1 U3923 ( .A1(n5344), .A2(n5343), .ZN(n5347) );
  CLKBUF_X1 U3924 ( .A(n4498), .Z(n4499) );
  NAND2_X1 U3925 ( .A1(n6463), .A2(n5490), .ZN(n3161) );
  OR2_X1 U3926 ( .A1(n5568), .A2(n4634), .ZN(n5542) );
  INV_X1 U3927 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4153) );
  AND2_X1 U3928 ( .A1(n5629), .A2(n4602), .ZN(n5588) );
  NOR2_X1 U3929 ( .A1(n6402), .A2(n6388), .ZN(n5740) );
  INV_X1 U3930 ( .A(n3220), .ZN(n3218) );
  AND3_X1 U3931 ( .A1(n4385), .A2(n4370), .A3(n5750), .ZN(n3217) );
  AND2_X1 U3932 ( .A1(n4438), .A2(n4437), .ZN(n5551) );
  MUX2_X1 U3933 ( .A(n4378), .B(n5638), .S(EBX_REG_3__SCAN_IN), .Z(n4355) );
  AOI21_X1 U3934 ( .B1(n5490), .B2(n4261), .A(n4293), .ZN(n4308) );
  OR2_X1 U3935 ( .A1(n4323), .A2(n4322), .ZN(n4348) );
  NAND2_X1 U3936 ( .A1(n4709), .A2(n3167), .ZN(n4663) );
  AND2_X1 U3937 ( .A1(n3168), .A2(n6355), .ZN(n3167) );
  OAI21_X1 U3938 ( .B1(n5513), .B2(n3814), .A(n4265), .ZN(n4467) );
  NAND2_X1 U3939 ( .A1(n4178), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4180)
         );
  INV_X1 U3940 ( .A(n4177), .ZN(n4178) );
  OR2_X1 U3941 ( .A1(n4180), .A2(n4179), .ZN(n4220) );
  AOI21_X1 U3942 ( .B1(n5893), .B2(n4261), .A(n4176), .ZN(n5561) );
  AND2_X1 U3943 ( .A1(n4136), .A2(n4135), .ZN(n5582) );
  OR2_X1 U3944 ( .A1(n5921), .A2(n3814), .ZN(n4136) );
  OR2_X1 U3945 ( .A1(n4092), .A2(n4091), .ZN(n4110) );
  AND2_X1 U3946 ( .A1(n4054), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4055)
         );
  INV_X1 U3947 ( .A(n4053), .ZN(n4054) );
  OR2_X1 U3948 ( .A1(n5947), .A2(n3814), .ZN(n4074) );
  INV_X1 U3949 ( .A(n5494), .ZN(n3284) );
  NOR2_X1 U3950 ( .A1(n5495), .A2(n5701), .ZN(n5700) );
  NAND2_X1 U3951 ( .A1(n3930), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3931)
         );
  INV_X1 U3952 ( .A(n3929), .ZN(n3930) );
  INV_X1 U3953 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3933) );
  OR2_X1 U3954 ( .A1(n3931), .A2(n3933), .ZN(n4019) );
  AND3_X1 U3955 ( .A1(n3909), .A2(n3908), .A3(n3907), .ZN(n5472) );
  OR2_X1 U3956 ( .A1(n3831), .A2(n7025), .ZN(n3910) );
  OR2_X1 U3957 ( .A1(n3871), .A2(n3829), .ZN(n3831) );
  NAND2_X1 U3958 ( .A1(n3812), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3871)
         );
  INV_X1 U3959 ( .A(n3869), .ZN(n3812) );
  AND2_X1 U3960 ( .A1(n3793), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3794)
         );
  INV_X1 U3961 ( .A(n3862), .ZN(n3793) );
  NAND2_X1 U3962 ( .A1(n3801), .A2(n3800), .ZN(n5297) );
  AND2_X1 U3963 ( .A1(n5298), .A2(n5297), .ZN(n5760) );
  NAND2_X1 U3964 ( .A1(n3617), .A2(n3616), .ZN(n3618) );
  NAND2_X1 U3965 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3848) );
  NAND2_X1 U3966 ( .A1(n3843), .A2(n3842), .ZN(n4782) );
  NOR2_X1 U3967 ( .A1(n4474), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4572)
         );
  NAND2_X1 U3968 ( .A1(n3720), .A2(n3172), .ZN(n4474) );
  INV_X1 U3969 ( .A(n4472), .ZN(n3172) );
  INV_X1 U3970 ( .A(n4572), .ZN(n4475) );
  OR2_X1 U3971 ( .A1(n5528), .A2(n4560), .ZN(n4561) );
  NAND2_X1 U3972 ( .A1(n5864), .A2(n3201), .ZN(n5866) );
  AND2_X1 U3973 ( .A1(n6018), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3201)
         );
  AND2_X1 U3974 ( .A1(n5574), .A2(n3141), .ZN(n5526) );
  INV_X1 U3975 ( .A(n4461), .ZN(n3228) );
  NAND2_X1 U3976 ( .A1(n5574), .A2(n3229), .ZN(n5553) );
  NAND2_X1 U3977 ( .A1(n5574), .A2(n5563), .ZN(n5562) );
  NAND2_X1 U3978 ( .A1(n5624), .A2(n3119), .ZN(n5587) );
  INV_X1 U3979 ( .A(n5585), .ZN(n3215) );
  NOR2_X1 U3980 ( .A1(n5974), .A2(n3137), .ZN(n5971) );
  AOI21_X1 U3981 ( .B1(n3240), .B2(n3712), .A(n3128), .ZN(n3212) );
  NAND2_X1 U3982 ( .A1(n5705), .A2(n5684), .ZN(n5686) );
  AND2_X1 U3983 ( .A1(n4409), .A2(n4408), .ZN(n5702) );
  NAND2_X1 U3984 ( .A1(n3242), .A2(n3240), .ZN(n5963) );
  INV_X1 U3985 ( .A(n5499), .ZN(n4406) );
  INV_X1 U3986 ( .A(n3233), .ZN(n3232) );
  NOR2_X1 U3987 ( .A1(n5797), .A2(n3233), .ZN(n6246) );
  OR2_X1 U3988 ( .A1(n5797), .A2(n5427), .ZN(n6248) );
  NOR2_X1 U3989 ( .A1(n5368), .A2(n6645), .ZN(n6267) );
  NAND2_X1 U3990 ( .A1(n4442), .A2(n4371), .ZN(n4791) );
  OR2_X1 U3991 ( .A1(n6216), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4793)
         );
  NAND2_X1 U3992 ( .A1(n3190), .A2(n3432), .ZN(n3189) );
  INV_X1 U3993 ( .A(n4509), .ZN(n3190) );
  AND3_X1 U3994 ( .A1(n3518), .A2(n3517), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3519) );
  INV_X1 U3995 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n4909) );
  INV_X1 U3996 ( .A(n4749), .ZN(n4744) );
  AND2_X1 U3997 ( .A1(n4487), .A2(n3140), .ZN(n3208) );
  INV_X1 U3998 ( .A(n3553), .ZN(n3555) );
  OR3_X1 U3999 ( .A1(n4688), .A2(n4687), .A3(n4686), .ZN(n5335) );
  OR2_X1 U4000 ( .A1(n5254), .A2(n4832), .ZN(n5180) );
  AND3_X1 U4001 ( .A1(n5345), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6719) );
  NOR2_X1 U4002 ( .A1(n5302), .A2(n6722), .ZN(n5305) );
  AND2_X1 U4003 ( .A1(n5101), .A2(n4832), .ZN(n5308) );
  INV_X1 U4004 ( .A(n4830), .ZN(n6659) );
  NAND2_X1 U4005 ( .A1(n5306), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4866) );
  INV_X1 U4006 ( .A(READY_N), .ZN(n6838) );
  INV_X1 U4007 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4621) );
  NAND2_X1 U4008 ( .A1(n4663), .A2(n4664), .ZN(n6842) );
  NOR2_X1 U4009 ( .A1(n3164), .A2(n3163), .ZN(n5589) );
  INV_X1 U4010 ( .A(n4593), .ZN(n3163) );
  OR2_X1 U4011 ( .A1(n5709), .A2(n4601), .ZN(n5667) );
  OR2_X1 U4012 ( .A1(n5504), .A2(n5503), .ZN(n5709) );
  NAND2_X1 U4013 ( .A1(n3166), .A2(n3127), .ZN(n5706) );
  INV_X1 U4014 ( .A(n6394), .ZN(n3166) );
  OR2_X1 U4015 ( .A1(n5458), .A2(n5436), .ZN(n6443) );
  AND2_X1 U4016 ( .A1(n6433), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U4017 ( .A1(n3184), .A2(n3183), .ZN(n5812) );
  NAND2_X1 U4018 ( .A1(n4458), .A2(n4459), .ZN(n3183) );
  INV_X1 U4019 ( .A(n4460), .ZN(n3184) );
  AND2_X1 U4020 ( .A1(n5856), .A2(n4806), .ZN(n5851) );
  NAND2_X2 U4021 ( .A1(n5856), .A2(n4805), .ZN(n5859) );
  INV_X1 U4022 ( .A(n6497), .ZN(n6492) );
  OR3_X1 U4023 ( .A1(n4755), .A2(n4754), .A3(n4753), .ZN(n6500) );
  AND2_X1 U4024 ( .A1(n4878), .A2(n5363), .ZN(n4754) );
  AND2_X1 U4025 ( .A1(n6500), .A2(n4770), .ZN(n6497) );
  OR3_X1 U4026 ( .A1(n4663), .A2(n3435), .A3(READY_N), .ZN(n6516) );
  INV_X1 U4027 ( .A(n6545), .ZN(n6552) );
  INV_X1 U4028 ( .A(n5812), .ZN(n5877) );
  OAI21_X1 U4029 ( .B1(n5560), .B2(n5561), .A(n5548), .ZN(n5890) );
  OR2_X1 U4030 ( .A1(n5560), .A2(n5573), .ZN(n5915) );
  AND2_X1 U4031 ( .A1(n3987), .A2(n3986), .ZN(n5978) );
  CLKBUF_X1 U4032 ( .A(n5715), .Z(n5716) );
  NAND2_X1 U4033 ( .A1(n6063), .A2(n3698), .ZN(n6057) );
  INV_X1 U4034 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n7064) );
  XNOR2_X1 U4035 ( .A(n3271), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4559)
         );
  NAND2_X1 U4036 ( .A1(n3267), .A2(n3266), .ZN(n3271) );
  NAND2_X1 U4037 ( .A1(n5885), .A2(n3126), .ZN(n3267) );
  INV_X1 U4038 ( .A(n6079), .ZN(n3226) );
  NAND2_X1 U4039 ( .A1(n6083), .A2(n6082), .ZN(n3224) );
  OR2_X1 U4040 ( .A1(n6124), .A2(n4551), .ZN(n6100) );
  NAND2_X1 U4041 ( .A1(n5864), .A2(n3299), .ZN(n5870) );
  XNOR2_X1 U4042 ( .A(n5864), .B(n5879), .ZN(n6111) );
  AND2_X1 U4043 ( .A1(n5885), .A2(n3724), .ZN(n5886) );
  NAND2_X1 U4044 ( .A1(n5902), .A2(n5901), .ZN(n5911) );
  AND2_X1 U4045 ( .A1(n6137), .A2(n4547), .ZN(n6130) );
  NAND2_X1 U4046 ( .A1(n5918), .A2(n3246), .ZN(n3243) );
  NAND2_X1 U4047 ( .A1(n3253), .A2(n3245), .ZN(n3244) );
  OAI211_X1 U4048 ( .C1(n5945), .C2(n5919), .A(n3249), .B(n3248), .ZN(n3247)
         );
  XNOR2_X1 U4049 ( .A(n5929), .B(n5928), .ZN(n6146) );
  INV_X1 U4050 ( .A(n5927), .ZN(n5928) );
  AND2_X1 U4051 ( .A1(n5624), .A2(n4423), .ZN(n5611) );
  NAND2_X1 U4052 ( .A1(n3254), .A2(n3256), .ZN(n5937) );
  AND2_X1 U4053 ( .A1(n5661), .A2(n5660), .ZN(n6181) );
  OR2_X1 U4054 ( .A1(n6239), .A2(n4543), .ZN(n4534) );
  AND2_X1 U4055 ( .A1(n3258), .A2(n3708), .ZN(n3207) );
  OR2_X1 U4056 ( .A1(n3262), .A2(n3260), .ZN(n3206) );
  NOR2_X1 U4057 ( .A1(n6220), .A2(n6195), .ZN(n6253) );
  NAND2_X1 U4058 ( .A1(n5051), .A2(n3661), .ZN(n6559) );
  OR2_X1 U4059 ( .A1(n4537), .A2(n4524), .ZN(n6252) );
  NAND2_X1 U4060 ( .A1(n4521), .A2(n3474), .ZN(n4522) );
  NAND2_X1 U4061 ( .A1(n4793), .A2(n4794), .ZN(n5368) );
  INV_X1 U4062 ( .A(n6566), .ZN(n6577) );
  AND2_X1 U4063 ( .A1(n6278), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6282) );
  OR2_X1 U4064 ( .A1(n6722), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6307) );
  AND2_X1 U4065 ( .A1(n4956), .A2(n6287), .ZN(n6289) );
  INV_X1 U4066 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7116) );
  OAI21_X1 U4067 ( .B1(n4904), .B2(n5365), .A(n5019), .ZN(n6656) );
  INV_X1 U4068 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4696) );
  INV_X1 U4069 ( .A(n6308), .ZN(n6344) );
  NOR2_X2 U4070 ( .A1(n5107), .A2(n5106), .ZN(n6341) );
  NAND2_X1 U4071 ( .A1(n5021), .A2(n5020), .ZN(n5044) );
  INV_X1 U4072 ( .A(n6716), .ZN(n6762) );
  OAI21_X1 U4073 ( .B1(n5221), .B2(n5220), .A(n5219), .ZN(n5246) );
  INV_X1 U4074 ( .A(n5301), .ZN(n6856) );
  AOI22_X1 U4075 ( .A1(n5305), .A2(n5308), .B1(n6303), .B2(n5392), .ZN(n6861)
         );
  AND2_X1 U4076 ( .A1(n6571), .A2(DATAI_28_), .ZN(n6855) );
  NAND2_X1 U4077 ( .A1(n6289), .A2(n5105), .ZN(n6853) );
  NOR2_X1 U4078 ( .A1(n4836), .A2(n6659), .ZN(n5175) );
  OAI211_X1 U4079 ( .C1(n6304), .C2(n5143), .A(n4835), .B(n6668), .ZN(n4865)
         );
  AND2_X1 U4080 ( .A1(n5394), .A2(n5393), .ZN(n5418) );
  NAND2_X1 U4081 ( .A1(n5306), .A2(DATAI_0_), .ZN(n6717) );
  OR2_X1 U4082 ( .A1(n4866), .A2(n3435), .ZN(n6770) );
  INV_X1 U4083 ( .A(n6773), .ZN(n6678) );
  OR2_X1 U4084 ( .A1(n4866), .A2(n4843), .ZN(n6777) );
  INV_X1 U4085 ( .A(n6780), .ZN(n6683) );
  INV_X1 U4086 ( .A(n6794), .ZN(n6697) );
  INV_X1 U4087 ( .A(n6804), .ZN(n6702) );
  OR2_X1 U4088 ( .A1(n4919), .A2(n6659), .ZN(n5382) );
  OR2_X1 U4089 ( .A1(n4866), .A2(n4853), .ZN(n6704) );
  INV_X1 U4090 ( .A(n5063), .ZN(n5096) );
  OAI211_X1 U4091 ( .C1(n4918), .C2(n4920), .A(n6668), .B(n4917), .ZN(n4942)
         );
  NAND2_X1 U4092 ( .A1(n4709), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6349) );
  INV_X1 U4093 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6359) );
  NOR2_X1 U4094 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6357) );
  AND2_X1 U4095 ( .A1(n3780), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6355) );
  INV_X2 U4096 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6345) );
  AND3_X1 U4097 ( .A1(n6938), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n4617) );
  NOR2_X1 U4098 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6844) );
  AND2_X1 U4099 ( .A1(n6815), .A2(STATE_REG_1__SCAN_IN), .ZN(n6825) );
  OAI21_X1 U4100 ( .B1(n5777), .B2(n6452), .A(n4609), .ZN(n4610) );
  NOR2_X1 U4101 ( .A1(n3157), .A2(n3156), .ZN(n5493) );
  NOR2_X1 U4102 ( .A1(n5491), .A2(REIP_REG_30__SCAN_IN), .ZN(n3156) );
  NAND2_X1 U4103 ( .A1(n3162), .A2(n3158), .ZN(n3157) );
  OAI22_X1 U4104 ( .A1(n6073), .A2(n5802), .B1(n6481), .B2(n5486), .ZN(n4456)
         );
  AND2_X1 U4105 ( .A1(n4566), .A2(n4565), .ZN(n4567) );
  NAND2_X1 U4106 ( .A1(n4465), .A2(n4464), .ZN(U2832) );
  INV_X1 U4107 ( .A(n4463), .ZN(n4464) );
  NAND2_X1 U4108 ( .A1(n5877), .A2(n6479), .ZN(n4465) );
  OAI22_X1 U4109 ( .A1(n6096), .A2(n5802), .B1(n6945), .B2(n6481), .ZN(n4463)
         );
  NOR2_X1 U4110 ( .A1(n4330), .A2(n3296), .ZN(n4331) );
  INV_X1 U4111 ( .A(n4327), .ZN(n4330) );
  AOI21_X1 U4112 ( .B1(n5490), .B2(n5979), .A(n4576), .ZN(n4580) );
  NAND2_X1 U4113 ( .A1(n3147), .A2(n3145), .ZN(U2958) );
  INV_X1 U4114 ( .A(n3146), .ZN(n3145) );
  NAND2_X1 U4115 ( .A1(n6085), .A2(n3784), .ZN(n3147) );
  NAND2_X1 U4116 ( .A1(n6177), .A2(n3784), .ZN(n5969) );
  OAI211_X1 U4117 ( .C1(n6077), .C2(n3196), .A(n3195), .B(n3193), .ZN(n6074)
         );
  NAND2_X1 U4118 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n4574), .ZN(n3196) );
  OAI21_X1 U4119 ( .B1(n6084), .B2(n6275), .A(n3222), .ZN(U2989) );
  INV_X1 U4120 ( .A(n3223), .ZN(n3222) );
  OAI211_X1 U4121 ( .C1(n6080), .C2(n6252), .A(n3225), .B(n3224), .ZN(n3223)
         );
  NOR2_X1 U4122 ( .A1(n6081), .A2(n3226), .ZN(n3225) );
  OR2_X1 U4123 ( .A1(n5609), .A2(n3282), .ZN(n5596) );
  NOR2_X1 U4124 ( .A1(n3284), .A2(n3287), .ZN(n5635) );
  INV_X2 U4125 ( .A(n5456), .ZN(n3182) );
  AND3_X1 U4126 ( .A1(n3363), .A2(n3362), .A3(n3361), .ZN(n3114) );
  NAND2_X1 U4127 ( .A1(n6018), .A2(n7166), .ZN(n3115) );
  XNOR2_X1 U4128 ( .A(n3704), .B(n4386), .ZN(n6056) );
  NOR2_X1 U4129 ( .A1(n5621), .A2(n3187), .ZN(n3116) );
  INV_X1 U4130 ( .A(n3279), .ZN(n5583) );
  AND2_X1 U4131 ( .A1(n3715), .A2(n3143), .ZN(n3117) );
  NAND2_X1 U4132 ( .A1(n5624), .A2(n3134), .ZN(n5598) );
  AND2_X1 U4133 ( .A1(n3134), .A2(n3216), .ZN(n3118) );
  AND2_X1 U4134 ( .A1(n3118), .A2(n3215), .ZN(n3119) );
  AND2_X1 U4135 ( .A1(n4340), .A2(n3391), .ZN(n3300) );
  INV_X1 U4136 ( .A(n3300), .ZN(n4371) );
  AND2_X1 U4137 ( .A1(n3177), .A2(n5054), .ZN(n3120) );
  NOR2_X1 U4138 ( .A1(n5377), .A2(n5472), .ZN(n5473) );
  INV_X1 U4139 ( .A(n3164), .ZN(n5617) );
  OR2_X1 U4140 ( .A1(n5678), .A2(n4592), .ZN(n3164) );
  NAND2_X1 U4141 ( .A1(n5624), .A2(n3118), .ZN(n3121) );
  AND2_X1 U4142 ( .A1(n3209), .A2(n3438), .ZN(n3122) );
  AND2_X1 U4143 ( .A1(n5936), .A2(n3255), .ZN(n3123) );
  AND4_X1 U4144 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3124)
         );
  NAND2_X1 U4145 ( .A1(n3892), .A2(n3891), .ZN(n5377) );
  INV_X1 U4146 ( .A(n3705), .ZN(n3264) );
  NAND2_X1 U4147 ( .A1(n3202), .A2(n3204), .ZN(n6001) );
  AND2_X1 U4148 ( .A1(n3261), .A2(n3705), .ZN(n3125) );
  INV_X1 U4149 ( .A(n5550), .ZN(n4200) );
  NAND2_X1 U4150 ( .A1(n3242), .A2(n3711), .ZN(n5993) );
  NAND2_X1 U4151 ( .A1(n6057), .A2(n6056), .ZN(n6055) );
  AND2_X1 U4152 ( .A1(n3726), .A2(n3724), .ZN(n3126) );
  OR2_X1 U4153 ( .A1(n6402), .A2(n4590), .ZN(n3127) );
  OR2_X1 U4154 ( .A1(n5609), .A2(n3281), .ZN(n3279) );
  AND2_X1 U4155 ( .A1(n6018), .A2(n7117), .ZN(n3128) );
  NOR2_X1 U4156 ( .A1(n4951), .A2(n5178), .ZN(n5055) );
  NAND2_X1 U4157 ( .A1(n6435), .A2(n4601), .ZN(n3129) );
  OR2_X1 U4158 ( .A1(n6020), .A2(n3717), .ZN(n3130) );
  NOR2_X1 U4159 ( .A1(n3709), .A2(n3264), .ZN(n3131) );
  AND2_X1 U4160 ( .A1(n3280), .A2(n5582), .ZN(n3132) );
  AND2_X1 U4161 ( .A1(n3232), .A2(n5736), .ZN(n3133) );
  INV_X1 U4162 ( .A(n3251), .ZN(n3250) );
  NAND2_X1 U4163 ( .A1(n3123), .A2(n3252), .ZN(n3251) );
  INV_X1 U4164 ( .A(n3191), .ZN(n6850) );
  NOR2_X1 U4165 ( .A1(n4866), .A2(n3474), .ZN(n3191) );
  AND2_X1 U4166 ( .A1(n4423), .A2(n5610), .ZN(n3134) );
  AND4_X1 U4167 ( .A1(n5657), .A2(n5655), .A3(n5696), .A4(n5654), .ZN(n3135)
         );
  NAND2_X1 U4168 ( .A1(n5053), .A2(n5052), .ZN(n5051) );
  INV_X1 U4169 ( .A(n3257), .ZN(n3256) );
  NOR2_X1 U4170 ( .A1(n6018), .A2(n6107), .ZN(n3136) );
  OR2_X1 U4171 ( .A1(n3113), .A2(n6937), .ZN(n3137) );
  INV_X1 U4172 ( .A(n4325), .ZN(n3168) );
  AND2_X1 U4173 ( .A1(n4090), .A2(n4089), .ZN(n3138) );
  INV_X1 U4174 ( .A(n4817), .ZN(n3858) );
  AND2_X1 U4175 ( .A1(n4312), .A2(n3208), .ZN(n3139) );
  AND2_X1 U4176 ( .A1(n4321), .A2(n3209), .ZN(n3140) );
  AND2_X1 U4177 ( .A1(n3229), .A2(n3228), .ZN(n3141) );
  AND3_X1 U4178 ( .A1(n3221), .A2(n4369), .A3(n4370), .ZN(n5294) );
  INV_X1 U4179 ( .A(n3474), .ZN(n3432) );
  AND2_X1 U4180 ( .A1(n4312), .A2(n3189), .ZN(n3142) );
  NAND2_X1 U4181 ( .A1(n3450), .A2(n3474), .ZN(n4322) );
  NAND2_X1 U4182 ( .A1(n4617), .A2(n6304), .ZN(n6054) );
  INV_X2 U4183 ( .A(n6054), .ZN(n6571) );
  AND3_X1 U4184 ( .A1(n6141), .A2(n6163), .A3(n6122), .ZN(n3143) );
  AND3_X1 U4185 ( .A1(n6142), .A2(n5899), .A3(n6164), .ZN(n3144) );
  AND2_X2 U4186 ( .A1(n4710), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4720)
         );
  NOR4_X2 U4187 ( .A1(n6997), .A2(n6383), .A3(n6382), .A4(n6381), .ZN(n6833)
         );
  XNOR2_X2 U4188 ( .A(n3148), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6085)
         );
  NAND2_X1 U4189 ( .A1(n3151), .A2(n3117), .ZN(n3722) );
  NAND3_X1 U4190 ( .A1(n3152), .A2(n6063), .A3(n6011), .ZN(n3204) );
  NAND2_X2 U4191 ( .A1(n6065), .A2(n6064), .ZN(n6063) );
  NAND3_X1 U4192 ( .A1(n3258), .A2(n3708), .A3(n3115), .ZN(n3154) );
  NOR2_X2 U4193 ( .A1(n3665), .A2(n3664), .ZN(n3680) );
  NAND2_X2 U4194 ( .A1(n3779), .A2(n3778), .ZN(n4709) );
  NAND2_X1 U4195 ( .A1(n3169), .A2(n3661), .ZN(n3170) );
  INV_X1 U4196 ( .A(n5052), .ZN(n3169) );
  NAND3_X1 U4197 ( .A1(n3171), .A2(n6558), .A3(n3170), .ZN(n6557) );
  NAND3_X1 U4198 ( .A1(n3661), .A2(n3640), .A3(n3234), .ZN(n3171) );
  NAND3_X1 U4199 ( .A1(n3204), .A2(n3202), .A3(n3203), .ZN(n3242) );
  NAND3_X1 U4200 ( .A1(n3173), .A2(n3120), .A3(n3174), .ZN(n3936) );
  INV_X1 U4201 ( .A(n4951), .ZN(n3174) );
  INV_X1 U4202 ( .A(n5178), .ZN(n3177) );
  INV_X1 U4203 ( .A(n3892), .ZN(n5378) );
  OR2_X1 U4204 ( .A1(n5621), .A2(n5623), .ZN(n5609) );
  NOR2_X2 U4205 ( .A1(n5621), .A2(n3185), .ZN(n5560) );
  NAND2_X1 U4206 ( .A1(n3426), .A2(n3425), .ZN(n3495) );
  NAND3_X1 U4207 ( .A1(n3455), .A2(n3457), .A3(n3456), .ZN(n3527) );
  NAND3_X1 U4208 ( .A1(n3199), .A2(n3200), .A3(n3527), .ZN(n3198) );
  XNOR2_X2 U4209 ( .A(n3551), .B(n3550), .ZN(n3580) );
  INV_X1 U4210 ( .A(n6011), .ZN(n3205) );
  NAND2_X1 U4211 ( .A1(n3206), .A2(n3207), .ZN(n6010) );
  OAI21_X1 U4212 ( .B1(n3451), .B2(n4328), .A(n3209), .ZN(n3356) );
  NAND2_X1 U4213 ( .A1(n3240), .A2(n6001), .ZN(n3211) );
  NAND2_X1 U4214 ( .A1(n3211), .A2(n3212), .ZN(n5961) );
  NAND2_X1 U4215 ( .A1(n3421), .A2(n4340), .ZN(n3388) );
  NAND2_X1 U4216 ( .A1(n3218), .A2(n3217), .ZN(n5748) );
  NOR2_X1 U4217 ( .A1(n3220), .A2(n3219), .ZN(n5749) );
  NAND2_X1 U4218 ( .A1(n4385), .A2(n4370), .ZN(n3219) );
  NAND2_X1 U4219 ( .A1(n4369), .A2(n4370), .ZN(n6429) );
  INV_X1 U4220 ( .A(n5797), .ZN(n3231) );
  NAND2_X1 U4221 ( .A1(n3231), .A2(n3133), .ZN(n5737) );
  NAND2_X1 U4222 ( .A1(n3235), .A2(n6567), .ZN(n3234) );
  NAND2_X1 U4223 ( .A1(n4948), .A2(n3236), .ZN(n3235) );
  NAND2_X1 U4224 ( .A1(n6569), .A2(n6567), .ZN(n6568) );
  NAND2_X1 U4225 ( .A1(n4948), .A2(n3236), .ZN(n6569) );
  NAND2_X2 U4226 ( .A1(n4950), .A2(n4949), .ZN(n4948) );
  NAND2_X1 U4227 ( .A1(n6001), .A2(n3240), .ZN(n3239) );
  NAND3_X1 U4228 ( .A1(n3247), .A2(n3244), .A3(n3243), .ZN(n6136) );
  NAND2_X2 U4229 ( .A1(n5918), .A2(n3256), .ZN(n3253) );
  OR2_X1 U4230 ( .A1(n5918), .A2(n5944), .ZN(n3254) );
  NAND2_X2 U4231 ( .A1(n3253), .A2(n3123), .ZN(n5935) );
  NOR2_X1 U4232 ( .A1(n3113), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3257)
         );
  INV_X1 U4233 ( .A(n6056), .ZN(n3259) );
  NAND2_X1 U4234 ( .A1(n6056), .A2(n3265), .ZN(n3261) );
  OAI21_X1 U4235 ( .B1(n6063), .B2(n3259), .A(n3125), .ZN(n6019) );
  NAND2_X1 U4236 ( .A1(n5864), .A2(n3268), .ZN(n3266) );
  AND2_X1 U4237 ( .A1(n5864), .A2(n3269), .ZN(n4573) );
  NAND2_X2 U4238 ( .A1(n3723), .A2(n3722), .ZN(n5885) );
  INV_X1 U4239 ( .A(n5995), .ZN(n3278) );
  NAND3_X1 U4240 ( .A1(n4305), .A2(n4306), .A3(n4304), .ZN(U2955) );
  NAND2_X1 U4241 ( .A1(n5494), .A2(n3285), .ZN(n5621) );
  NAND2_X1 U4242 ( .A1(n5494), .A2(n5496), .ZN(n5495) );
  NAND2_X1 U4243 ( .A1(n3936), .A2(n3935), .ZN(n3937) );
  AND2_X1 U4244 ( .A1(n3293), .A2(n3292), .ZN(n4460) );
  NAND2_X1 U4245 ( .A1(n3293), .A2(n4200), .ZN(n4458) );
  NAND2_X1 U4246 ( .A1(n3552), .A2(n3580), .ZN(n3621) );
  NAND2_X1 U4247 ( .A1(n5935), .A2(n3295), .ZN(n5929) );
  NAND2_X1 U4248 ( .A1(n5935), .A2(n5904), .ZN(n5910) );
  AOI21_X1 U4249 ( .B1(n4830), .B2(n3844), .A(n6345), .ZN(n4773) );
  NAND2_X1 U4250 ( .A1(n5523), .A2(n4467), .ZN(n4469) );
  INV_X1 U4251 ( .A(n5804), .ZN(n5807) );
  NAND2_X1 U4252 ( .A1(n5804), .A2(n6479), .ZN(n4568) );
  AOI21_X2 U4253 ( .B1(n4780), .B2(n4779), .A(n3614), .ZN(n6579) );
  AOI22_X1 U4254 ( .A1(n4279), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4255 ( .A1(n3406), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3505), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3370) );
  NAND2_X1 U4256 ( .A1(n4307), .A2(n4308), .ZN(n4310) );
  XNOR2_X1 U4257 ( .A(n3587), .B(n3586), .ZN(n3839) );
  AND2_X1 U4258 ( .A1(n6481), .A2(n4353), .ZN(n6479) );
  AND2_X1 U4259 ( .A1(n4393), .A2(n4392), .ZN(n3294) );
  NAND2_X2 U4260 ( .A1(n4352), .A2(n4351), .ZN(n6481) );
  INV_X1 U4261 ( .A(n6481), .ZN(n4564) );
  INV_X1 U4262 ( .A(n4832), .ZN(n6453) );
  OR2_X1 U4263 ( .A1(n3113), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3295)
         );
  INV_X1 U4264 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6815) );
  AND2_X1 U4265 ( .A1(n5839), .A2(DATAI_14_), .ZN(n3296) );
  OR2_X1 U4266 ( .A1(n3458), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3297)
         );
  AND3_X1 U4267 ( .A1(n3323), .A2(n3322), .A3(n3321), .ZN(n3298) );
  AND2_X1 U4268 ( .A1(n6018), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3299)
         );
  AND2_X1 U4269 ( .A1(n6357), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3438) );
  AND2_X1 U4270 ( .A1(n4315), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3735) );
  AND2_X1 U4271 ( .A1(n6718), .A2(n4749), .ZN(n3742) );
  AND2_X1 U4272 ( .A1(n3454), .A2(n3453), .ZN(n3457) );
  AOI22_X1 U4273 ( .A1(n3536), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3362) );
  OR2_X1 U4274 ( .A1(n4131), .A2(n4130), .ZN(n4139) );
  OR2_X1 U4275 ( .A1(n3631), .A2(n3630), .ZN(n3682) );
  AOI22_X1 U4276 ( .A1(n3467), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3357) );
  AND3_X1 U4277 ( .A1(n4338), .A2(n4337), .A3(n4336), .ZN(n4339) );
  INV_X1 U4278 ( .A(n5718), .ZN(n3949) );
  OR2_X1 U4279 ( .A1(n4213), .A2(n4212), .ZN(n4236) );
  AND2_X1 U4280 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3911) );
  AND2_X1 U4281 ( .A1(n5795), .A2(n5745), .ZN(n3834) );
  OR2_X1 U4282 ( .A1(n3651), .A2(n3650), .ZN(n3681) );
  AOI22_X1 U4283 ( .A1(n3499), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3479), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3303) );
  INV_X1 U4284 ( .A(n3496), .ZN(n3497) );
  OR3_X1 U4285 ( .A1(n3766), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n7116), 
        .ZN(n4316) );
  INV_X1 U4286 ( .A(n4791), .ZN(n4446) );
  INV_X1 U4287 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4179) );
  AND2_X1 U4288 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3968) );
  INV_X1 U4289 ( .A(n5379), .ZN(n3891) );
  INV_X1 U4290 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3829) );
  AND2_X1 U4291 ( .A1(n3763), .A2(n3699), .ZN(n3700) );
  NAND2_X1 U4292 ( .A1(n4349), .A2(n4666), .ZN(n4321) );
  INV_X1 U4293 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5333) );
  AND2_X1 U4294 ( .A1(n4418), .A2(n5637), .ZN(n5640) );
  NOR2_X1 U4295 ( .A1(n4713), .A2(n4346), .ZN(n4530) );
  NOR2_X1 U4296 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3849) );
  AND2_X1 U4297 ( .A1(n6345), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4294) );
  AND2_X1 U4298 ( .A1(n4521), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3860) );
  AND2_X1 U4299 ( .A1(n4728), .A2(n4712), .ZN(n6714) );
  INV_X1 U4300 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5337) );
  OR2_X1 U4301 ( .A1(n3600), .A2(n3599), .ZN(n3601) );
  INV_X1 U4302 ( .A(n6307), .ZN(n6725) );
  AND2_X2 U4303 ( .A1(n3435), .A2(n5456), .ZN(n4666) );
  INV_X1 U4304 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n7025) );
  INV_X1 U4305 ( .A(n6419), .ZN(n6455) );
  INV_X1 U4306 ( .A(n3814), .ZN(n4261) );
  NAND2_X1 U4307 ( .A1(n4320), .A2(n4319), .ZN(n4687) );
  OR2_X1 U4308 ( .A1(n5862), .A2(n3814), .ZN(n4244) );
  AND4_X1 U4309 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n5379)
         );
  AND2_X1 U4310 ( .A1(n6218), .A2(n4539), .ZN(n6266) );
  AND2_X1 U4311 ( .A1(n5070), .A2(n5069), .ZN(n5094) );
  NAND2_X1 U4312 ( .A1(n5100), .A2(n5216), .ZN(n5183) );
  NAND2_X1 U4313 ( .A1(n5100), .A2(n5016), .ZN(n5134) );
  INV_X1 U4314 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U4315 ( .A1(n6349), .A2(n4833), .ZN(n4834) );
  OR3_X1 U4316 ( .A1(n6288), .A2(n6722), .A3(n4839), .ZN(n4835) );
  OR2_X1 U4317 ( .A1(n4866), .A2(n4861), .ZN(n6791) );
  AND2_X1 U4318 ( .A1(n6359), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3780) );
  OR2_X1 U4319 ( .A1(n4667), .A2(n6365), .ZN(n4664) );
  OR2_X1 U4320 ( .A1(n6366), .A2(n6843), .ZN(n5353) );
  INV_X1 U4321 ( .A(n6443), .ZN(n6458) );
  INV_X1 U4322 ( .A(n6452), .ZN(n6439) );
  INV_X1 U4323 ( .A(n5802), .ZN(n6478) );
  OR2_X1 U4324 ( .A1(n4487), .A2(n3590), .ZN(n5363) );
  INV_X1 U4325 ( .A(n6503), .ZN(n6553) );
  NAND2_X1 U4326 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3863), .ZN(n3862)
         );
  NAND2_X1 U4327 ( .A1(n6372), .A2(n4300), .ZN(n5981) );
  INV_X1 U4328 ( .A(n5918), .ZN(n5945) );
  INV_X1 U4329 ( .A(n6275), .ZN(n6649) );
  INV_X1 U4330 ( .A(n6252), .ZN(n6644) );
  NAND2_X1 U4331 ( .A1(n5066), .A2(n5065), .ZN(n5092) );
  OAI211_X1 U4332 ( .C1(n5188), .C2(n5187), .A(n6668), .B(n5186), .ZN(n5212)
         );
  NOR2_X1 U4333 ( .A1(n5183), .A2(n4830), .ZN(n6308) );
  OAI211_X1 U4334 ( .C1(n5112), .C2(n5111), .A(n6668), .B(n5110), .ZN(n5136)
         );
  INV_X1 U4335 ( .A(n5134), .ZN(n5048) );
  INV_X1 U4336 ( .A(n6671), .ZN(n6707) );
  AND2_X1 U4337 ( .A1(n6660), .A2(n6659), .ZN(n6763) );
  OAI211_X1 U4338 ( .C1(n4988), .C2(n4987), .A(n6668), .B(n4986), .ZN(n5011)
         );
  INV_X1 U4339 ( .A(n6768), .ZN(n6723) );
  INV_X1 U4340 ( .A(n5222), .ZN(n5250) );
  AND2_X1 U4341 ( .A1(n6289), .A2(n5216), .ZN(n5263) );
  OAI211_X1 U4342 ( .C1(n5262), .C2(n5261), .A(n6668), .B(n5260), .ZN(n5285)
         );
  INV_X1 U4343 ( .A(n6790), .ZN(n6744) );
  OAI211_X1 U4344 ( .C1(n5309), .C2(n5308), .A(n6311), .B(n5307), .ZN(n6857)
         );
  AND2_X1 U4345 ( .A1(n6278), .A2(n4830), .ZN(n5105) );
  AND2_X1 U4346 ( .A1(n4834), .A2(n6938), .ZN(n5306) );
  NAND2_X1 U4347 ( .A1(n5147), .A2(n5146), .ZN(n5171) );
  INV_X1 U4348 ( .A(n5423), .ZN(n5383) );
  INV_X1 U4349 ( .A(n5382), .ZN(n5420) );
  INV_X1 U4350 ( .A(n6785), .ZN(n6685) );
  INV_X1 U4351 ( .A(n6800), .ZN(n6699) );
  OR4_X1 U4352 ( .A1(n5357), .A2(n5356), .A3(n5355), .A4(n5354), .ZN(n5358) );
  INV_X1 U4353 ( .A(n6825), .ZN(n4660) );
  INV_X1 U4354 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6371) );
  INV_X1 U4355 ( .A(n4610), .ZN(n4611) );
  OR2_X4 U4356 ( .A1(n5426), .A2(n5424), .ZN(n6424) );
  INV_X1 U4357 ( .A(n6446), .ZN(n6460) );
  OR2_X1 U4358 ( .A1(n5760), .A2(n5299), .ZN(n6561) );
  OR2_X1 U4359 ( .A1(n4784), .A2(n4783), .ZN(n5465) );
  OR2_X1 U4360 ( .A1(n4906), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4770) );
  INV_X1 U4361 ( .A(n6549), .ZN(n6503) );
  NAND2_X1 U4362 ( .A1(n5981), .A2(n4775), .ZN(n6586) );
  NAND2_X1 U4363 ( .A1(n5062), .A2(n4830), .ZN(n5210) );
  AOI22_X1 U4364 ( .A1(n5182), .A2(n5187), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5181), .ZN(n5215) );
  AOI22_X1 U4365 ( .A1(n5109), .A2(n5111), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5104), .ZN(n5139) );
  NAND2_X1 U4366 ( .A1(n6660), .A2(n4830), .ZN(n6671) );
  AOI22_X1 U4367 ( .A1(n6664), .A2(n6669), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6665), .ZN(n6711) );
  NAND2_X1 U4368 ( .A1(n5015), .A2(n5105), .ZN(n6768) );
  AOI22_X1 U4369 ( .A1(n4984), .A2(n4987), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6719), .ZN(n5014) );
  NAND2_X1 U4370 ( .A1(n5263), .A2(n4830), .ZN(n5287) );
  AOI22_X1 U4371 ( .A1(n5258), .A2(n5261), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5257), .ZN(n5291) );
  INV_X1 U4372 ( .A(n6787), .ZN(n6688) );
  NAND2_X1 U4373 ( .A1(n5306), .A2(DATAI_4_), .ZN(n6860) );
  NAND2_X1 U4374 ( .A1(n5306), .A2(DATAI_7_), .ZN(n6758) );
  NAND2_X1 U4375 ( .A1(n6289), .A2(n5016), .ZN(n6801) );
  INV_X1 U4376 ( .A(n5175), .ZN(n4872) );
  OR2_X1 U4377 ( .A1(n4836), .A2(n4830), .ZN(n5423) );
  INV_X1 U4378 ( .A(n6855), .ZN(n6329) );
  INV_X1 U4379 ( .A(n6764), .ZN(n6343) );
  INV_X1 U4380 ( .A(n6829), .ZN(n6809) );
  AND2_X1 U4381 ( .A1(n4623), .A2(n6849), .ZN(n6829) );
  INV_X1 U4382 ( .A(n6825), .ZN(n6849) );
  NAND2_X1 U4383 ( .A1(n4568), .A2(n4567), .ZN(U2830) );
  NOR2_X4 U4384 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3309) );
  AND2_X2 U4385 ( .A1(n4881), .A2(n3309), .ZN(n3405) );
  INV_X1 U4386 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4710) );
  AOI22_X1 U4387 ( .A1(n3405), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3306) );
  NOR2_X4 U4388 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4389 ( .A1(n3537), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3305) );
  AND2_X4 U4390 ( .A1(n3309), .A2(n4895), .ZN(n3484) );
  AOI22_X1 U4391 ( .A1(n3505), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3304) );
  AND2_X4 U4392 ( .A1(n3307), .A2(n3309), .ZN(n3535) );
  AND2_X4 U4393 ( .A1(n3308), .A2(n4881), .ZN(n4279) );
  AOI22_X1 U4394 ( .A1(n3535), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3315) );
  AND2_X4 U4395 ( .A1(n4720), .A2(n3310), .ZN(n3460) );
  AOI22_X1 U4396 ( .A1(n3567), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3313) );
  AND2_X4 U4397 ( .A1(n4895), .A2(n4715), .ZN(n3406) );
  AOI22_X1 U4398 ( .A1(n3461), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3312) );
  AND2_X4 U4399 ( .A1(n4715), .A2(n3310), .ZN(n3462) );
  AOI22_X1 U4400 ( .A1(n3536), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3311) );
  XNOR2_X1 U4401 ( .A(n4621), .B(STATE_REG_1__SCAN_IN), .ZN(n4482) );
  NOR2_X1 U4402 ( .A1(n5455), .A2(n4482), .ZN(n3451) );
  AOI22_X1 U4403 ( .A1(n3567), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4404 ( .A1(n3536), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4405 ( .A1(n3505), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4406 ( .A1(n3461), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3321) );
  NAND3_X2 U4407 ( .A1(n3325), .A2(n3298), .A3(n3324), .ZN(n3448) );
  NAND2_X1 U4408 ( .A1(n4279), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3329)
         );
  NAND2_X1 U4409 ( .A1(n3536), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3328)
         );
  NAND2_X1 U4410 ( .A1(n3535), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3327) );
  NAND2_X1 U4411 ( .A1(n3392), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3326) );
  NAND2_X1 U4412 ( .A1(n3460), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3333) );
  NAND2_X1 U4413 ( .A1(n3567), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4414 ( .A1(n3505), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3331) );
  NAND2_X1 U4415 ( .A1(n3484), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3330)
         );
  NAND2_X1 U4416 ( .A1(n3537), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3337)
         );
  NAND2_X1 U4417 ( .A1(n3499), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3336) );
  NAND2_X1 U4418 ( .A1(n3479), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3335) );
  NAND2_X1 U4419 ( .A1(n3462), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U4420 ( .A1(n3467), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3341)
         );
  NAND2_X1 U4421 ( .A1(n3405), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3340) );
  NAND2_X1 U4422 ( .A1(n3406), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3339)
         );
  NAND2_X1 U4423 ( .A1(n3461), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4424 ( .A1(n3537), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4425 ( .A1(n3405), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4426 ( .A1(n3505), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4427 ( .A1(n3567), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4428 ( .A1(n3467), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4429 ( .A1(n3499), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3479), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4430 ( .A1(n3536), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4431 ( .A1(n4279), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3353) );
  INV_X1 U4432 ( .A(n3356), .ZN(n3419) );
  AOI22_X1 U4433 ( .A1(n3405), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4434 ( .A1(n3460), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4435 ( .A1(n3499), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3479), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4436 ( .A1(n3537), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4437 ( .A1(n4279), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3364) );
  NAND2_X1 U4438 ( .A1(n3436), .A2(n3448), .ZN(n3421) );
  AOI22_X1 U4439 ( .A1(n3392), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3479), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4440 ( .A1(n3405), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4441 ( .A1(n4279), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3536), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4442 ( .A1(n3567), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3366) );
  NAND4_X1 U4443 ( .A1(n3369), .A2(n3368), .A3(n3367), .A4(n3366), .ZN(n3375)
         );
  AOI22_X1 U4444 ( .A1(n3499), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3537), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4445 ( .A1(n3535), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4446 ( .A1(n3484), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3371) );
  NAND4_X1 U4447 ( .A1(n3373), .A2(n3372), .A3(n3371), .A4(n3370), .ZN(n3374)
         );
  OR2_X2 U4448 ( .A1(n3375), .A2(n3374), .ZN(n4353) );
  OAI21_X1 U4449 ( .B1(n3421), .B2(n3432), .A(n4353), .ZN(n4335) );
  AOI22_X1 U4450 ( .A1(n4279), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4451 ( .A1(n3536), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3392), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4452 ( .A1(n3499), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3479), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4453 ( .A1(n3537), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3376) );
  NAND4_X1 U4454 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n3385)
         );
  AOI22_X1 U4455 ( .A1(n3405), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3461), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4456 ( .A1(n3460), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4457 ( .A1(n3467), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3380) );
  NAND4_X1 U4458 ( .A1(n3383), .A2(n3382), .A3(n3381), .A4(n3380), .ZN(n3384)
         );
  INV_X2 U4459 ( .A(n3436), .ZN(n3450) );
  INV_X1 U4460 ( .A(n3448), .ZN(n4861) );
  NAND2_X1 U4461 ( .A1(n4861), .A2(n3427), .ZN(n3386) );
  NAND3_X1 U4462 ( .A1(n4334), .A2(n3448), .A3(n3450), .ZN(n3387) );
  INV_X2 U4463 ( .A(n3391), .ZN(n3435) );
  NAND2_X1 U4464 ( .A1(n4279), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3396)
         );
  NAND2_X1 U4465 ( .A1(n3536), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3395)
         );
  NAND2_X1 U4466 ( .A1(n3535), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3394) );
  NAND2_X1 U4467 ( .A1(n3392), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3393) );
  NAND2_X1 U4468 ( .A1(n3460), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3400) );
  NAND2_X1 U4469 ( .A1(n3567), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3399) );
  NAND2_X1 U4470 ( .A1(n3505), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3398) );
  NAND2_X1 U4471 ( .A1(n3484), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3397)
         );
  NAND2_X1 U4472 ( .A1(n3537), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3404)
         );
  NAND2_X1 U4473 ( .A1(n3499), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3403) );
  NAND2_X1 U4474 ( .A1(n3479), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3402) );
  NAND2_X1 U4475 ( .A1(n3462), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3401) );
  NAND2_X1 U4476 ( .A1(n3467), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3410)
         );
  NAND2_X1 U4477 ( .A1(n3405), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3409) );
  NAND2_X1 U4478 ( .A1(n3406), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3408)
         );
  NAND2_X1 U4479 ( .A1(n3461), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3407) );
  AND4_X4 U4480 ( .A1(n3414), .A2(n3413), .A3(n3412), .A4(n3411), .ZN(n5456)
         );
  NAND2_X1 U4481 ( .A1(n3447), .A2(n4666), .ZN(n3429) );
  NAND2_X1 U4482 ( .A1(n3436), .A2(n3474), .ZN(n3415) );
  NAND2_X1 U4483 ( .A1(n3783), .A2(n3415), .ZN(n3416) );
  INV_X1 U4484 ( .A(n3443), .ZN(n3417) );
  NAND2_X1 U4485 ( .A1(n3417), .A2(n3434), .ZN(n3418) );
  NAND4_X1 U4486 ( .A1(n3419), .A2(n3782), .A3(n3429), .A4(n3418), .ZN(n3420)
         );
  NAND2_X1 U4487 ( .A1(n3420), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3424) );
  INV_X1 U4488 ( .A(n3561), .ZN(n3422) );
  NAND2_X1 U4489 ( .A1(n3424), .A2(n3423), .ZN(n3529) );
  NAND2_X1 U4490 ( .A1(n3529), .A2(n4749), .ZN(n3426) );
  NAND2_X1 U4491 ( .A1(n6357), .A2(n6938), .ZN(n4299) );
  MUX2_X1 U4492 ( .A(n3780), .B(n4299), .S(n6718), .Z(n3425) );
  INV_X2 U4493 ( .A(n4666), .ZN(n5510) );
  NAND2_X1 U4494 ( .A1(n3429), .A2(n3428), .ZN(n3431) );
  NAND2_X1 U4495 ( .A1(n4333), .A2(n3443), .ZN(n4493) );
  NAND2_X1 U4496 ( .A1(n3432), .A2(n4353), .ZN(n3433) );
  NAND2_X1 U4497 ( .A1(n3436), .A2(n4353), .ZN(n4345) );
  NAND3_X1 U4498 ( .A1(n3590), .A2(n3435), .A3(n4345), .ZN(n3437) );
  INV_X1 U4499 ( .A(n4340), .ZN(n4857) );
  NAND2_X1 U4500 ( .A1(n3437), .A2(n4857), .ZN(n3439) );
  NAND2_X1 U4501 ( .A1(n3529), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3455) );
  NAND2_X1 U4502 ( .A1(n3444), .A2(n3443), .ZN(n4486) );
  INV_X1 U4503 ( .A(n4486), .ZN(n3445) );
  NAND2_X1 U4504 ( .A1(n3445), .A2(n3182), .ZN(n4325) );
  NOR2_X2 U4505 ( .A1(n3447), .A2(n3446), .ZN(n4498) );
  NAND2_X1 U4506 ( .A1(n4498), .A2(n3435), .ZN(n4312) );
  NAND2_X1 U4507 ( .A1(n4353), .A2(n3786), .ZN(n4488) );
  OAI211_X1 U4508 ( .C1(n4325), .C2(n3451), .A(n4312), .B(n4509), .ZN(n3452)
         );
  NAND2_X1 U4509 ( .A1(n3452), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3456) );
  INV_X1 U4510 ( .A(n4299), .ZN(n3558) );
  XNOR2_X1 U4511 ( .A(n5337), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6301)
         );
  NAND2_X1 U4512 ( .A1(n3558), .A2(n6301), .ZN(n3454) );
  INV_X1 U4513 ( .A(n3780), .ZN(n3532) );
  NAND2_X1 U4514 ( .A1(n3532), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3453) );
  INV_X1 U4515 ( .A(n3456), .ZN(n3459) );
  INV_X1 U4516 ( .A(n3457), .ZN(n3458) );
  NAND2_X1 U4517 ( .A1(n4711), .A2(n6938), .ZN(n3476) );
  BUF_X1 U4518 ( .A(n3460), .Z(n4273) );
  AOI22_X1 U4519 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n3506), .B1(n4273), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4520 ( .A1(n4279), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4521 ( .A1(n4271), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4522 ( .A1(n4203), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3463) );
  NAND4_X1 U4523 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3473)
         );
  BUF_X1 U4524 ( .A(n3535), .Z(n4278) );
  AOI22_X1 U4525 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n3478), .B1(n4278), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4526 ( .A1(n4280), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4527 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n4269), .B1(n4253), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4529 ( .A1(n4254), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3468) );
  NAND4_X1 U4530 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3472)
         );
  NAND2_X1 U4531 ( .A1(n3477), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4532 ( .A1(n3478), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4533 ( .A1(n4203), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4534 ( .A1(n4273), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4535 ( .A1(n4269), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3480) );
  NAND4_X1 U4536 ( .A1(n3483), .A2(n3482), .A3(n3481), .A4(n3480), .ZN(n3490)
         );
  AOI22_X1 U4537 ( .A1(n3506), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3467), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U4538 ( .A1(n4279), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4539 ( .A1(n4271), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U4540 ( .A1(n3484), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3485) );
  NAND4_X1 U4541 ( .A1(n3488), .A2(n3487), .A3(n3486), .A4(n3485), .ZN(n3489)
         );
  OR2_X1 U4542 ( .A1(n3562), .A2(n3699), .ZN(n3493) );
  OR2_X1 U4543 ( .A1(n3491), .A2(n3561), .ZN(n3492) );
  XNOR2_X2 U4544 ( .A(n3498), .B(n3497), .ZN(n3845) );
  NAND2_X1 U4545 ( .A1(n3845), .A2(n6938), .ZN(n3516) );
  INV_X1 U4546 ( .A(n3562), .ZN(n3515) );
  AOI22_X1 U4547 ( .A1(n4254), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4548 ( .A1(n4203), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4549 ( .A1(n4271), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3502) );
  BUF_X1 U4550 ( .A(n3462), .Z(n4272) );
  AOI22_X1 U4551 ( .A1(n3478), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3501) );
  NAND4_X1 U4552 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(n3512)
         );
  AOI22_X1 U4553 ( .A1(n4225), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4554 ( .A1(n4280), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4555 ( .A1(n4269), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4556 ( .A1(n3506), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3507) );
  NAND4_X1 U4557 ( .A1(n3510), .A2(n3509), .A3(n3508), .A4(n3507), .ZN(n3511)
         );
  INV_X1 U4558 ( .A(n3606), .ZN(n3513) );
  XNOR2_X1 U4559 ( .A(n3513), .B(n3699), .ZN(n3514) );
  NAND2_X1 U4560 ( .A1(n3515), .A2(n3514), .ZN(n3598) );
  NAND2_X1 U4561 ( .A1(n3516), .A2(n3598), .ZN(n3597) );
  NAND2_X1 U4562 ( .A1(n3477), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3520) );
  NAND2_X1 U4563 ( .A1(n5456), .A2(n3606), .ZN(n3518) );
  INV_X1 U4564 ( .A(n3699), .ZN(n3701) );
  NOR2_X1 U4565 ( .A1(n3562), .A2(n3701), .ZN(n3521) );
  NAND2_X1 U4566 ( .A1(n3587), .A2(n3586), .ZN(n3526) );
  INV_X1 U4567 ( .A(n3523), .ZN(n3524) );
  INV_X1 U4568 ( .A(n3581), .ZN(n3552) );
  NAND2_X1 U4569 ( .A1(n3530), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3534) );
  NAND2_X1 U4570 ( .A1(n5333), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5102) );
  MUX2_X1 U4571 ( .A(n5102), .B(n5333), .S(n6718), .Z(n3531) );
  NAND2_X1 U4572 ( .A1(n5337), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U4573 ( .A1(n3531), .A2(n5018), .ZN(n5022) );
  AOI22_X1 U4574 ( .A1(n5022), .A2(n3558), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3532), .ZN(n3533) );
  NAND2_X1 U4575 ( .A1(n3534), .A2(n3533), .ZN(n3554) );
  XNOR2_X2 U4576 ( .A(n3553), .B(n3554), .ZN(n4728) );
  AOI22_X1 U4577 ( .A1(n4279), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4578 ( .A1(n3478), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4579 ( .A1(n4203), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4580 ( .A1(n4280), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3538) );
  NAND4_X1 U4581 ( .A1(n3541), .A2(n3540), .A3(n3539), .A4(n3538), .ZN(n3547)
         );
  AOI22_X1 U4582 ( .A1(n3506), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3545) );
  AOI22_X1 U4583 ( .A1(n4271), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4584 ( .A1(n4273), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4585 ( .A1(n4254), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3542) );
  NAND4_X1 U4586 ( .A1(n3545), .A2(n3544), .A3(n3543), .A4(n3542), .ZN(n3546)
         );
  NOR2_X1 U4587 ( .A1(n3562), .A2(n3582), .ZN(n3548) );
  NAND2_X1 U4588 ( .A1(n3477), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3549) );
  OAI21_X1 U4589 ( .B1(n3582), .B2(n3561), .A(n3549), .ZN(n3550) );
  NAND2_X1 U4590 ( .A1(n3530), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3560) );
  NAND2_X1 U4591 ( .A1(n6719), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U4592 ( .A1(n5009), .A2(n5345), .ZN(n3556) );
  NAND2_X1 U4593 ( .A1(n5387), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4943) );
  NOR2_X1 U4594 ( .A1(n3780), .A2(n5345), .ZN(n3557) );
  AOI21_X1 U4595 ( .B1(n5145), .B2(n3558), .A(n3557), .ZN(n3559) );
  NAND2_X1 U4596 ( .A1(n4831), .A2(n6938), .ZN(n3575) );
  NAND2_X2 U4597 ( .A1(n3562), .A2(n3561), .ZN(n3769) );
  INV_X1 U4598 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6985) );
  AOI22_X1 U4599 ( .A1(n4225), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4600 ( .A1(n3478), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4601 ( .A1(n4203), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4602 ( .A1(n4280), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4603 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3573)
         );
  AOI22_X1 U4604 ( .A1(n3506), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4605 ( .A1(n4271), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4606 ( .A1(n4273), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4607 ( .A1(n4254), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3568) );
  NAND4_X1 U4608 ( .A1(n3571), .A2(n3570), .A3(n3569), .A4(n3568), .ZN(n3572)
         );
  AOI22_X1 U4609 ( .A1(n3769), .A2(n3634), .B1(n3477), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3574) );
  NAND2_X1 U4610 ( .A1(n3835), .A2(n3763), .ZN(n3579) );
  NAND2_X1 U4611 ( .A1(n3589), .A2(n3606), .ZN(n3588) );
  NAND2_X1 U4612 ( .A1(n3588), .A2(n3582), .ZN(n3635) );
  INV_X1 U4613 ( .A(n3634), .ZN(n3576) );
  XNOR2_X1 U4614 ( .A(n3635), .B(n3576), .ZN(n3577) );
  NAND2_X1 U4615 ( .A1(n3577), .A2(n4698), .ZN(n3578) );
  INV_X1 U4616 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6640) );
  XNOR2_X1 U4617 ( .A(n3581), .B(n3580), .ZN(n4828) );
  NAND2_X1 U4618 ( .A1(n4828), .A2(n3763), .ZN(n3585) );
  XNOR2_X1 U4619 ( .A(n3588), .B(n3582), .ZN(n3583) );
  AND2_X1 U4620 ( .A1(n5456), .A2(n4340), .ZN(n3604) );
  AOI21_X1 U4621 ( .B1(n3583), .B2(n4698), .A(n3604), .ZN(n3584) );
  NAND2_X1 U4622 ( .A1(n3585), .A2(n3584), .ZN(n6580) );
  NAND2_X1 U4623 ( .A1(n6580), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3615)
         );
  NAND2_X1 U4624 ( .A1(n3839), .A2(n3763), .ZN(n3596) );
  OAI21_X1 U4625 ( .B1(n3606), .B2(n3589), .A(n3588), .ZN(n3593) );
  INV_X1 U4626 ( .A(n3591), .ZN(n3592) );
  OAI211_X1 U4627 ( .C1(n3593), .C2(n3590), .A(n3592), .B(n4328), .ZN(n3594)
         );
  INV_X1 U4628 ( .A(n3594), .ZN(n3595) );
  NAND2_X1 U4629 ( .A1(n3596), .A2(n3595), .ZN(n4780) );
  NAND2_X1 U4630 ( .A1(n3597), .A2(n3600), .ZN(n3602) );
  INV_X1 U4631 ( .A(n3598), .ZN(n3599) );
  INV_X1 U4632 ( .A(n3763), .ZN(n3603) );
  INV_X1 U4633 ( .A(n3604), .ZN(n3605) );
  OAI21_X1 U4634 ( .B1(n3590), .B2(n3606), .A(n3605), .ZN(n3607) );
  INV_X1 U4635 ( .A(n3607), .ZN(n3608) );
  NAND2_X1 U4636 ( .A1(n4774), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3610)
         );
  INV_X1 U4637 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n7101) );
  NAND2_X1 U4638 ( .A1(n3610), .A2(n7101), .ZN(n3612) );
  AND2_X1 U4639 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3611) );
  NAND2_X1 U4640 ( .A1(n4774), .A2(n3611), .ZN(n3613) );
  INV_X1 U4641 ( .A(n3613), .ZN(n3614) );
  NAND2_X1 U4642 ( .A1(n3615), .A2(n6579), .ZN(n3619) );
  INV_X1 U4643 ( .A(n6580), .ZN(n3617) );
  INV_X1 U4644 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3616) );
  AND2_X2 U4645 ( .A1(n3619), .A2(n3618), .ZN(n4949) );
  AOI22_X1 U4646 ( .A1(n3478), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4647 ( .A1(n3506), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4254), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4648 ( .A1(n4203), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4649 ( .A1(n3500), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3622) );
  NAND4_X1 U4650 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(n3631)
         );
  AOI22_X1 U4651 ( .A1(n4225), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4652 ( .A1(n4271), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4653 ( .A1(n4273), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4654 ( .A1(n4269), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3626) );
  NAND4_X1 U4655 ( .A1(n3629), .A2(n3628), .A3(n3627), .A4(n3626), .ZN(n3630)
         );
  NAND2_X1 U4656 ( .A1(n3769), .A2(n3682), .ZN(n3633) );
  NAND2_X1 U4657 ( .A1(n3477), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3632) );
  XNOR2_X1 U4658 ( .A(n3665), .B(n3663), .ZN(n3868) );
  NAND2_X1 U4659 ( .A1(n3868), .A2(n3763), .ZN(n3638) );
  NAND2_X1 U4660 ( .A1(n3635), .A2(n3634), .ZN(n3684) );
  XNOR2_X1 U4661 ( .A(n3684), .B(n3682), .ZN(n3636) );
  NAND2_X1 U4662 ( .A1(n3636), .A2(n4698), .ZN(n3637) );
  INV_X1 U4663 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6629) );
  XNOR2_X1 U4664 ( .A(n3639), .B(n6629), .ZN(n6567) );
  NAND2_X1 U4665 ( .A1(n3639), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3640)
         );
  AOI22_X1 U4666 ( .A1(n4225), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4667 ( .A1(n3478), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4668 ( .A1(n4203), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4669 ( .A1(n4280), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3642) );
  NAND4_X1 U4670 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(n3651)
         );
  AOI22_X1 U4671 ( .A1(n3506), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4672 ( .A1(n4252), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4673 ( .A1(n4273), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3647) );
  INV_X1 U4674 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n6987) );
  AOI22_X1 U4675 ( .A1(n4254), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3646) );
  NAND4_X1 U4676 ( .A1(n3649), .A2(n3648), .A3(n3647), .A4(n3646), .ZN(n3650)
         );
  NAND2_X1 U4677 ( .A1(n3769), .A2(n3681), .ZN(n3653) );
  NAND2_X1 U4678 ( .A1(n3477), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3652) );
  NAND2_X1 U4679 ( .A1(n3653), .A2(n3652), .ZN(n3662) );
  NAND2_X1 U4680 ( .A1(n3787), .A2(n3763), .ZN(n3659) );
  INV_X1 U4681 ( .A(n3682), .ZN(n3655) );
  OR2_X1 U4682 ( .A1(n3684), .A2(n3655), .ZN(n3656) );
  XNOR2_X1 U4683 ( .A(n3656), .B(n3681), .ZN(n3657) );
  NAND2_X1 U4684 ( .A1(n3657), .A2(n4698), .ZN(n3658) );
  NAND2_X1 U4685 ( .A1(n3659), .A2(n3658), .ZN(n3660) );
  INV_X1 U4686 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n7150) );
  XNOR2_X1 U4687 ( .A(n3660), .B(n7150), .ZN(n5052) );
  NAND2_X1 U4688 ( .A1(n3660), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3661)
         );
  NAND2_X1 U4689 ( .A1(n3663), .A2(n3662), .ZN(n3664) );
  AOI22_X1 U4690 ( .A1(n4225), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4691 ( .A1(n3478), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4692 ( .A1(n4203), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4693 ( .A1(n4280), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3666) );
  NAND4_X1 U4694 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3675)
         );
  AOI22_X1 U4695 ( .A1(n3506), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4696 ( .A1(n4252), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4697 ( .A1(n4273), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4698 ( .A1(n4254), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3670) );
  NAND4_X1 U4699 ( .A1(n3673), .A2(n3672), .A3(n3671), .A4(n3670), .ZN(n3674)
         );
  NAND2_X1 U4700 ( .A1(n3769), .A2(n3692), .ZN(n3677) );
  NAND2_X1 U4701 ( .A1(n3477), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3676) );
  NAND2_X1 U4702 ( .A1(n3677), .A2(n3676), .ZN(n3679) );
  OR2_X1 U4703 ( .A1(n3680), .A2(n3679), .ZN(n3792) );
  NAND3_X1 U4704 ( .A1(n3678), .A2(n3763), .A3(n3792), .ZN(n3687) );
  NAND2_X1 U4705 ( .A1(n3682), .A2(n3681), .ZN(n3683) );
  OR2_X1 U4706 ( .A1(n3684), .A2(n3683), .ZN(n3691) );
  XNOR2_X1 U4707 ( .A(n3691), .B(n3692), .ZN(n3685) );
  NAND2_X1 U4708 ( .A1(n3685), .A2(n4698), .ZN(n3686) );
  NAND2_X1 U4709 ( .A1(n3687), .A2(n3686), .ZN(n3688) );
  INV_X1 U4710 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6620) );
  XNOR2_X1 U4711 ( .A(n3688), .B(n6620), .ZN(n6558) );
  NAND2_X1 U4712 ( .A1(n3688), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3689)
         );
  AOI22_X1 U4713 ( .A1(n3769), .A2(n3699), .B1(n3477), .B2(
        INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3690) );
  XNOR2_X2 U4714 ( .A(n3678), .B(n3690), .ZN(n3876) );
  OR2_X1 U4715 ( .A1(n3876), .A2(n3603), .ZN(n3696) );
  INV_X1 U4716 ( .A(n3691), .ZN(n3693) );
  NAND2_X1 U4717 ( .A1(n3693), .A2(n3692), .ZN(n3702) );
  XNOR2_X1 U4718 ( .A(n3702), .B(n3699), .ZN(n3694) );
  NAND2_X1 U4719 ( .A1(n3694), .A2(n4698), .ZN(n3695) );
  NAND2_X1 U4720 ( .A1(n3696), .A2(n3695), .ZN(n3697) );
  INV_X1 U4721 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4380) );
  XNOR2_X1 U4722 ( .A(n3697), .B(n4380), .ZN(n6064) );
  NAND2_X1 U4723 ( .A1(n3697), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3698)
         );
  OR3_X1 U4724 ( .A1(n3702), .A2(n3590), .A3(n3701), .ZN(n3703) );
  INV_X1 U4725 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4386) );
  NAND2_X1 U4726 ( .A1(n3704), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3705)
         );
  INV_X1 U4727 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6593) );
  INV_X1 U4728 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6240) );
  INV_X1 U4729 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6021) );
  INV_X1 U4730 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n7018) );
  AND4_X1 U4731 ( .A1(n6593), .A2(n6240), .A3(n6021), .A4(n7018), .ZN(n3706)
         );
  NOR2_X1 U4732 ( .A1(n6020), .A2(n3706), .ZN(n3709) );
  NAND2_X1 U4733 ( .A1(n6020), .A2(n6593), .ZN(n6047) );
  NAND2_X1 U4734 ( .A1(n6018), .A2(n7018), .ZN(n6017) );
  NAND2_X1 U4735 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U4736 ( .A1(n6018), .A2(n6023), .ZN(n3707) );
  AND3_X1 U4737 ( .A1(n6047), .A2(n6017), .A3(n3707), .ZN(n3708) );
  INV_X1 U4738 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n7166) );
  INV_X1 U4739 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6002) );
  AND2_X1 U4740 ( .A1(n6018), .A2(n6002), .ZN(n3712) );
  INV_X1 U4741 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n7117) );
  XNOR2_X1 U4742 ( .A(n6018), .B(n7117), .ZN(n5995) );
  NAND3_X1 U4743 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n3713) );
  AND2_X1 U4744 ( .A1(n6018), .A2(n3713), .ZN(n3716) );
  INV_X1 U4745 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n7144) );
  INV_X1 U4746 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6937) );
  INV_X1 U4747 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6184) );
  NAND3_X1 U4748 ( .A1(n7144), .A2(n6937), .A3(n6184), .ZN(n3714) );
  NAND2_X1 U4749 ( .A1(n3113), .A2(n3714), .ZN(n3715) );
  NOR2_X1 U4750 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6163) );
  NOR2_X1 U4751 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6141) );
  NOR2_X1 U4752 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6122) );
  INV_X1 U4753 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6116) );
  AND4_X1 U4754 ( .A1(n6163), .A2(n6141), .A3(n6122), .A4(n6116), .ZN(n3717)
         );
  AND2_X1 U4755 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6142) );
  AND2_X1 U4756 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6164) );
  AND2_X1 U4757 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5899) );
  NAND4_X1 U4758 ( .A1(n6142), .A2(n6164), .A3(n5899), .A4(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3718) );
  NAND2_X1 U4759 ( .A1(n6018), .A2(n3718), .ZN(n3719) );
  NAND2_X1 U4760 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6089) );
  AND2_X1 U4761 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4536) );
  NAND2_X1 U4762 ( .A1(n5954), .A2(n3144), .ZN(n3721) );
  NAND2_X1 U4763 ( .A1(n3721), .A2(n6020), .ZN(n3723) );
  XOR2_X1 U4764 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n6020), .Z(n5887) );
  INV_X1 U4765 ( .A(n5887), .ZN(n3724) );
  INV_X1 U4766 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5867) );
  INV_X1 U4767 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3725) );
  NAND2_X1 U4768 ( .A1(n5867), .A2(n3725), .ZN(n6090) );
  NOR3_X1 U4769 ( .A1(n4472), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3726) );
  INV_X1 U4770 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4721) );
  INV_X1 U4771 ( .A(n4559), .ZN(n3785) );
  NAND2_X1 U4772 ( .A1(n3769), .A2(n5455), .ZN(n3727) );
  NAND2_X1 U4773 ( .A1(n3727), .A2(n4328), .ZN(n3734) );
  INV_X1 U4774 ( .A(n3742), .ZN(n3728) );
  XNOR2_X1 U4775 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3743) );
  XNOR2_X1 U4776 ( .A(n3728), .B(n3743), .ZN(n4315) );
  AND2_X1 U4777 ( .A1(n4744), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3729)
         );
  NOR2_X1 U4778 ( .A1(n3742), .A2(n3729), .ZN(n3733) );
  AOI21_X1 U4779 ( .B1(n3783), .B2(n3733), .A(n3730), .ZN(n3732) );
  NAND2_X1 U4780 ( .A1(n3435), .A2(n4328), .ZN(n3731) );
  NAND2_X1 U4781 ( .A1(n5510), .A2(n3731), .ZN(n3746) );
  NAND2_X1 U4782 ( .A1(n3769), .A2(n3733), .ZN(n3738) );
  INV_X1 U4783 ( .A(n3734), .ZN(n3737) );
  INV_X1 U4784 ( .A(n3735), .ZN(n3736) );
  OAI22_X1 U4785 ( .A1(n3739), .A2(n3738), .B1(n3737), .B2(n3736), .ZN(n3741)
         );
  AOI21_X1 U4786 ( .B1(n3739), .B2(n4315), .A(n3776), .ZN(n3740) );
  NAND2_X1 U4787 ( .A1(n3743), .A2(n3742), .ZN(n3745) );
  NAND2_X1 U4788 ( .A1(n5337), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3744) );
  NAND2_X1 U4789 ( .A1(n3745), .A2(n3744), .ZN(n3754) );
  XNOR2_X1 U4790 ( .A(n5333), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3752)
         );
  XNOR2_X1 U4791 ( .A(n3754), .B(n3752), .ZN(n4314) );
  INV_X1 U4792 ( .A(n3477), .ZN(n3747) );
  NAND2_X1 U4793 ( .A1(n3769), .A2(n4314), .ZN(n3749) );
  INV_X1 U4794 ( .A(n3746), .ZN(n3750) );
  OAI211_X1 U4795 ( .C1(n4314), .C2(n3747), .A(n3749), .B(n3750), .ZN(n3748)
         );
  INV_X1 U4796 ( .A(n3752), .ZN(n3753) );
  NAND2_X1 U4797 ( .A1(n3754), .A2(n3753), .ZN(n3756) );
  NAND2_X1 U4798 ( .A1(n5333), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U4799 ( .A1(n3756), .A2(n3755), .ZN(n3762) );
  XNOR2_X1 U4800 ( .A(n3757), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3761)
         );
  INV_X1 U4801 ( .A(n3761), .ZN(n3758) );
  NAND2_X1 U4802 ( .A1(n3762), .A2(n3758), .ZN(n3760) );
  NAND2_X1 U4803 ( .A1(n5345), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3759) );
  NAND2_X1 U4804 ( .A1(n3760), .A2(n3759), .ZN(n3766) );
  XNOR2_X1 U4805 ( .A(n3762), .B(n3761), .ZN(n4313) );
  NAND2_X1 U4806 ( .A1(n4316), .A2(n4313), .ZN(n3770) );
  AND2_X1 U4807 ( .A1(n3763), .A2(n3770), .ZN(n3764) );
  NAND2_X1 U4808 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4696), .ZN(n3767) );
  AOI22_X1 U4809 ( .A1(n3769), .A2(n4318), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6938), .ZN(n3774) );
  INV_X1 U4810 ( .A(n3770), .ZN(n3771) );
  NAND2_X1 U4811 ( .A1(n3772), .A2(n3771), .ZN(n3773) );
  NAND3_X1 U4812 ( .A1(n3775), .A2(n3774), .A3(n3773), .ZN(n3779) );
  INV_X1 U4813 ( .A(n3776), .ZN(n3777) );
  NAND2_X1 U4814 ( .A1(n4347), .A2(n5456), .ZN(n3781) );
  NAND2_X1 U4815 ( .A1(n3782), .A2(n3781), .ZN(n4496) );
  INV_X1 U4816 ( .A(n6372), .ZN(n3784) );
  NAND2_X1 U4817 ( .A1(n3785), .A2(n3784), .ZN(n4306) );
  NAND2_X1 U4818 ( .A1(n3787), .A2(n4030), .ZN(n3791) );
  NOR2_X2 U4819 ( .A1(n4353), .A2(n6345), .ZN(n3815) );
  XNOR2_X1 U4820 ( .A(n3862), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5058) );
  INV_X1 U4821 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3788) );
  OAI22_X1 U4822 ( .A1(n5058), .A2(n3814), .B1(n3788), .B2(n4154), .ZN(n3789)
         );
  AOI21_X1 U4823 ( .B1(n4240), .B2(EAX_REG_5__SCAN_IN), .A(n3789), .ZN(n3790)
         );
  NAND2_X1 U4824 ( .A1(n3791), .A2(n3790), .ZN(n5054) );
  NAND2_X1 U4825 ( .A1(n3792), .A2(n4030), .ZN(n3801) );
  INV_X1 U4826 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6494) );
  INV_X1 U4827 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3795) );
  OAI22_X1 U4828 ( .A1(n4197), .A2(n6494), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3795), .ZN(n3799) );
  INV_X1 U4829 ( .A(n3794), .ZN(n3796) );
  NAND2_X1 U4830 ( .A1(n3796), .A2(n3795), .ZN(n3797) );
  NAND2_X1 U4831 ( .A1(n3869), .A2(n3797), .ZN(n6565) );
  AND2_X1 U4832 ( .A1(n6565), .A2(n3849), .ZN(n3798) );
  AOI21_X1 U4833 ( .B1(n3799), .B2(n3814), .A(n3798), .ZN(n3800) );
  INV_X1 U4834 ( .A(n4030), .ZN(n3875) );
  AOI22_X1 U4835 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n3478), .B1(n4278), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4836 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n4203), .B1(n4270), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4837 ( .A1(n4269), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4838 ( .A1(n3500), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3802) );
  NAND4_X1 U4839 ( .A1(n3805), .A2(n3804), .A3(n3803), .A4(n3802), .ZN(n3811)
         );
  AOI22_X1 U4840 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3506), .B1(n4254), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4841 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n4273), .B1(n4280), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4842 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n4279), .B1(n4272), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4843 ( .A1(n4252), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3806) );
  NAND4_X1 U4844 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(n3810)
         );
  NOR2_X1 U4845 ( .A1(n3811), .A2(n3810), .ZN(n3818) );
  NAND2_X1 U4846 ( .A1(n3831), .A2(n7025), .ZN(n3813) );
  NAND2_X1 U4847 ( .A1(n3910), .A2(n3813), .ZN(n6409) );
  INV_X1 U4848 ( .A(n3849), .ZN(n3814) );
  AOI22_X1 U4849 ( .A1(n6409), .A2(n4261), .B1(PHYADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n4294), .ZN(n3817) );
  NAND2_X1 U4850 ( .A1(n3815), .A2(EAX_REG_9__SCAN_IN), .ZN(n3816) );
  OAI211_X1 U4851 ( .C1(n3875), .C2(n3818), .A(n3817), .B(n3816), .ZN(n5795)
         );
  INV_X1 U4852 ( .A(EAX_REG_8__SCAN_IN), .ZN(n5854) );
  AOI22_X1 U4853 ( .A1(n3478), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4854 ( .A1(n4254), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4855 ( .A1(n4203), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4856 ( .A1(n4280), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4857 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3828)
         );
  AOI22_X1 U4858 ( .A1(n4225), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4859 ( .A1(n4252), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4860 ( .A1(n4273), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4861 ( .A1(n3506), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4862 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3827)
         );
  OAI21_X1 U4863 ( .B1(n3828), .B2(n3827), .A(n4030), .ZN(n3833) );
  NAND2_X1 U4864 ( .A1(n3871), .A2(n3829), .ZN(n3830) );
  NAND2_X1 U4865 ( .A1(n3831), .A2(n3830), .ZN(n6059) );
  AOI22_X1 U4866 ( .A1(n6059), .A2(n4261), .B1(PHYADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n4294), .ZN(n3832) );
  OAI211_X1 U4867 ( .C1(n4197), .C2(n5854), .A(n3833), .B(n3832), .ZN(n5745)
         );
  INV_X1 U4868 ( .A(n4488), .ZN(n4521) );
  AOI21_X1 U4869 ( .B1(n7064), .B2(n3848), .A(n3863), .ZN(n6464) );
  OAI22_X1 U4870 ( .A1(n6464), .A2(n3814), .B1(n4154), .B2(n7064), .ZN(n3836)
         );
  AOI21_X1 U4871 ( .B1(n3815), .B2(EAX_REG_3__SCAN_IN), .A(n3836), .ZN(n3837)
         );
  OAI21_X1 U4872 ( .B1(n3757), .B2(n3852), .A(n3837), .ZN(n3838) );
  AOI21_X1 U4873 ( .B1(n3835), .B2(n4030), .A(n3838), .ZN(n4952) );
  AOI21_X1 U4874 ( .B1(n4828), .B2(n4030), .A(n4294), .ZN(n4818) );
  NAND2_X1 U4875 ( .A1(n3839), .A2(n4030), .ZN(n3843) );
  AOI22_X1 U4876 ( .A1(n3815), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6345), .ZN(n3841) );
  NAND2_X1 U4877 ( .A1(n3860), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3840) );
  AND2_X1 U4878 ( .A1(n3841), .A2(n3840), .ZN(n3842) );
  INV_X1 U4879 ( .A(n4345), .ZN(n3844) );
  NAND2_X1 U4880 ( .A1(n3845), .A2(n4030), .ZN(n3847) );
  AOI22_X1 U4881 ( .A1(n4240), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6345), .ZN(n3846) );
  OAI211_X1 U4882 ( .C1(n3852), .C2(n4744), .A(n3847), .B(n3846), .ZN(n4772)
         );
  MUX2_X1 U4883 ( .A(n3849), .B(n4773), .S(n4772), .Z(n4781) );
  INV_X1 U4884 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4742) );
  OAI21_X1 U4885 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3848), .ZN(n6585) );
  AOI22_X1 U4886 ( .A1(n4294), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n3849), 
        .B2(n6585), .ZN(n3851) );
  NAND2_X1 U4887 ( .A1(n4240), .A2(EAX_REG_2__SCAN_IN), .ZN(n3850) );
  OAI211_X1 U4888 ( .C1(n3852), .C2(n4742), .A(n3851), .B(n3850), .ZN(n3854)
         );
  NAND2_X1 U4889 ( .A1(n4784), .A2(n3854), .ZN(n3853) );
  NAND2_X1 U4890 ( .A1(n4818), .A2(n3853), .ZN(n3857) );
  INV_X1 U4891 ( .A(n4784), .ZN(n3856) );
  INV_X1 U4892 ( .A(n3854), .ZN(n3855) );
  NAND2_X1 U4893 ( .A1(n3860), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3866) );
  INV_X1 U4894 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6431) );
  AOI21_X1 U4895 ( .B1(n6431), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3861) );
  AOI21_X1 U4896 ( .B1(n3815), .B2(EAX_REG_4__SCAN_IN), .A(n3861), .ZN(n3865)
         );
  OAI21_X1 U4897 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3863), .A(n3862), 
        .ZN(n6575) );
  NOR2_X1 U4898 ( .A1(n6575), .A2(n3814), .ZN(n3864) );
  AOI21_X1 U4899 ( .B1(n3866), .B2(n3865), .A(n3864), .ZN(n3867) );
  AOI21_X1 U4900 ( .B1(n3868), .B2(n4030), .A(n3867), .ZN(n5178) );
  INV_X1 U4901 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n7159) );
  NAND2_X1 U4902 ( .A1(n3869), .A2(n7159), .ZN(n3870) );
  NAND2_X1 U4903 ( .A1(n3871), .A2(n3870), .ZN(n6067) );
  NAND2_X1 U4904 ( .A1(n6067), .A2(n4261), .ZN(n3872) );
  OAI21_X1 U4905 ( .B1(n4154), .B2(n7159), .A(n3872), .ZN(n3873) );
  AOI21_X1 U4906 ( .B1(n4240), .B2(EAX_REG_7__SCAN_IN), .A(n3873), .ZN(n3874)
         );
  OAI21_X4 U4907 ( .B1(n3876), .B2(n3875), .A(n3874), .ZN(n5761) );
  AOI22_X1 U4908 ( .A1(n3506), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4909 ( .A1(n4225), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4910 ( .A1(n4254), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4911 ( .A1(n3500), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3877) );
  NAND4_X1 U4912 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3886)
         );
  AOI22_X1 U4913 ( .A1(n4203), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4914 ( .A1(n3478), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4915 ( .A1(n4280), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4916 ( .A1(n4252), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3881) );
  NAND4_X1 U4917 ( .A1(n3884), .A2(n3883), .A3(n3882), .A4(n3881), .ZN(n3885)
         );
  OAI21_X1 U4918 ( .B1(n3886), .B2(n3885), .A(n4030), .ZN(n3890) );
  NAND2_X1 U4919 ( .A1(n3815), .A2(EAX_REG_10__SCAN_IN), .ZN(n3889) );
  INV_X1 U4920 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3893) );
  XNOR2_X1 U4921 ( .A(n3910), .B(n3893), .ZN(n6042) );
  NAND2_X1 U4922 ( .A1(n6042), .A2(n4261), .ZN(n3888) );
  NAND2_X1 U4923 ( .A1(n4294), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3887)
         );
  NOR2_X1 U4924 ( .A1(n3910), .A2(n3893), .ZN(n3894) );
  XNOR2_X1 U4925 ( .A(n3894), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6395)
         );
  NAND2_X1 U4926 ( .A1(n6395), .A2(n4261), .ZN(n3909) );
  AOI22_X1 U4927 ( .A1(n4225), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4928 ( .A1(n3506), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4929 ( .A1(n4203), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4930 ( .A1(n3478), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3895) );
  NAND4_X1 U4931 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3895), .ZN(n3904)
         );
  AOI22_X1 U4932 ( .A1(n4270), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4933 ( .A1(n4252), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4934 ( .A1(n4273), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4935 ( .A1(n4254), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3899) );
  NAND4_X1 U4936 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n3903)
         );
  OR2_X1 U4937 ( .A1(n3904), .A2(n3903), .ZN(n3906) );
  INV_X1 U4938 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6392) );
  NOR2_X1 U4939 ( .A1(n4154), .A2(n6392), .ZN(n3905) );
  AOI21_X1 U4940 ( .B1(n4030), .B2(n3906), .A(n3905), .ZN(n3908) );
  NAND2_X1 U4941 ( .A1(n3815), .A2(EAX_REG_11__SCAN_IN), .ZN(n3907) );
  XNOR2_X1 U4942 ( .A(n3929), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5732)
         );
  NAND2_X1 U4943 ( .A1(n5732), .A2(n4261), .ZN(n3916) );
  INV_X1 U4944 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5847) );
  INV_X1 U4945 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5734) );
  AOI21_X1 U4946 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5734), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3913) );
  INV_X1 U4947 ( .A(n3913), .ZN(n3914) );
  OAI21_X1 U4948 ( .B1(n4197), .B2(n5847), .A(n3914), .ZN(n3915) );
  NAND2_X1 U4949 ( .A1(n3916), .A2(n3915), .ZN(n3928) );
  AOI22_X1 U4950 ( .A1(n4225), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4951 ( .A1(n4203), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4952 ( .A1(n3460), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4953 ( .A1(n4269), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3917) );
  NAND4_X1 U4954 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3926)
         );
  AOI22_X1 U4955 ( .A1(n3506), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4254), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4956 ( .A1(n3478), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4957 ( .A1(n4252), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4958 ( .A1(n4253), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3921) );
  NAND4_X1 U4959 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3925)
         );
  OAI21_X1 U4960 ( .B1(n3926), .B2(n3925), .A(n4030), .ZN(n3927) );
  NAND2_X1 U4961 ( .A1(n3928), .A2(n3927), .ZN(n5731) );
  NAND2_X1 U4962 ( .A1(n3931), .A2(n3933), .ZN(n3932) );
  NAND2_X1 U4963 ( .A1(n4019), .A2(n3932), .ZN(n6013) );
  INV_X1 U4964 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5845) );
  OAI22_X1 U4965 ( .A1(n4197), .A2(n5845), .B1(n3933), .B2(n4154), .ZN(n3934)
         );
  AOI21_X1 U4966 ( .B1(n6013), .B2(n3849), .A(n3934), .ZN(n3935) );
  NAND2_X1 U4967 ( .A1(n3951), .A2(n3937), .ZN(n5714) );
  INV_X1 U4968 ( .A(n5714), .ZN(n3950) );
  AOI22_X1 U4969 ( .A1(n4279), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3478), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4970 ( .A1(n4203), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4971 ( .A1(n4280), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4972 ( .A1(n4254), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3938) );
  NAND4_X1 U4973 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(n3947)
         );
  AOI22_X1 U4974 ( .A1(n3506), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4975 ( .A1(n4270), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4976 ( .A1(n3500), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4977 ( .A1(n4252), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3942) );
  NAND4_X1 U4978 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3946)
         );
  OR2_X1 U4979 ( .A1(n3947), .A2(n3946), .ZN(n3948) );
  NAND2_X1 U4980 ( .A1(n4030), .A2(n3948), .ZN(n5718) );
  NAND2_X1 U4981 ( .A1(n3950), .A2(n3949), .ZN(n5715) );
  NAND2_X1 U4982 ( .A1(n5715), .A2(n3951), .ZN(n5494) );
  INV_X1 U4983 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4018) );
  XNOR2_X1 U4984 ( .A(n4019), .B(n4018), .ZN(n6006) );
  NAND2_X1 U4985 ( .A1(n6006), .A2(n3849), .ZN(n3966) );
  AOI22_X1 U4986 ( .A1(n4270), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4987 ( .A1(n3506), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4252), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4988 ( .A1(n4273), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4989 ( .A1(n4280), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3952) );
  NAND4_X1 U4990 ( .A1(n3955), .A2(n3954), .A3(n3953), .A4(n3952), .ZN(n3961)
         );
  AOI22_X1 U4991 ( .A1(n4279), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3478), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4992 ( .A1(n4254), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4993 ( .A1(n4203), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4994 ( .A1(n4251), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3956) );
  NAND4_X1 U4995 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3960)
         );
  OAI21_X1 U4996 ( .B1(n3961), .B2(n3960), .A(n4030), .ZN(n3964) );
  NAND2_X1 U4997 ( .A1(n3815), .A2(EAX_REG_14__SCAN_IN), .ZN(n3963) );
  NAND2_X1 U4998 ( .A1(n4294), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3962)
         );
  AND3_X1 U4999 ( .A1(n3964), .A2(n3963), .A3(n3962), .ZN(n3965) );
  NAND2_X1 U5000 ( .A1(n3966), .A2(n3965), .ZN(n5496) );
  NAND2_X1 U5001 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3967) );
  INV_X1 U5002 ( .A(n3969), .ZN(n3986) );
  INV_X1 U5003 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U5004 ( .A1(n3986), .A2(n5965), .ZN(n3970) );
  AND2_X1 U5005 ( .A1(n4053), .A2(n3970), .ZN(n5967) );
  AOI22_X1 U5006 ( .A1(n4203), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3460), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U5007 ( .A1(n4254), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U5008 ( .A1(n4225), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U5009 ( .A1(n3478), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3971) );
  NAND4_X1 U5010 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n3980)
         );
  AOI22_X1 U5011 ( .A1(n4280), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U5012 ( .A1(n4252), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U5013 ( .A1(n3500), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U5014 ( .A1(n3506), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U5015 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3979)
         );
  OR2_X1 U5016 ( .A1(n3980), .A2(n3979), .ZN(n3983) );
  INV_X1 U5017 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6509) );
  OAI21_X1 U5018 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6371), .A(n6345), 
        .ZN(n3981) );
  OAI21_X1 U5019 ( .B1(n4197), .B2(n6509), .A(n3981), .ZN(n3982) );
  AOI21_X1 U5020 ( .B1(n4175), .B2(n3983), .A(n3982), .ZN(n3984) );
  AOI21_X1 U5021 ( .B1(n5967), .B2(n3849), .A(n3984), .ZN(n5657) );
  INV_X1 U5022 ( .A(n3985), .ZN(n4021) );
  INV_X1 U5023 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4012) );
  INV_X1 U5024 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n7046) );
  OAI21_X1 U5025 ( .B1(n4021), .B2(n4012), .A(n7046), .ZN(n3987) );
  AOI22_X1 U5026 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n3478), .B1(n4279), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U5027 ( .A1(n4252), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4254), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U5028 ( .A1(n4203), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U5029 ( .A1(n4270), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3988) );
  NAND4_X1 U5030 ( .A1(n3991), .A2(n3990), .A3(n3989), .A4(n3988), .ZN(n3997)
         );
  AOI22_X1 U5031 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n3506), .B1(n4273), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U5032 ( .A1(n4280), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U5033 ( .A1(n3500), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U5034 ( .A1(n4251), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3992) );
  NAND4_X1 U5035 ( .A1(n3995), .A2(n3994), .A3(n3993), .A4(n3992), .ZN(n3996)
         );
  OR2_X1 U5036 ( .A1(n3997), .A2(n3996), .ZN(n4000) );
  NAND2_X1 U5037 ( .A1(n4240), .A2(EAX_REG_17__SCAN_IN), .ZN(n3998) );
  OAI211_X1 U5038 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n7046), .A(n3998), .B(
        n3814), .ZN(n3999) );
  AOI21_X1 U5039 ( .B1(n4175), .B2(n4000), .A(n3999), .ZN(n4001) );
  AOI21_X1 U5040 ( .B1(n5978), .B2(n3849), .A(n4001), .ZN(n5655) );
  XNOR2_X1 U5041 ( .A(n4021), .B(n4012), .ZN(n5988) );
  NAND2_X1 U5042 ( .A1(n5988), .A2(n3849), .ZN(n4017) );
  AOI22_X1 U5043 ( .A1(n4279), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U5044 ( .A1(n3460), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U5045 ( .A1(n4203), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U5046 ( .A1(n4254), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4002) );
  NAND4_X1 U5047 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4011)
         );
  AOI22_X1 U5048 ( .A1(n4280), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U5049 ( .A1(n3478), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U5050 ( .A1(n3506), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U5051 ( .A1(n4252), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4006) );
  NAND4_X1 U5052 ( .A1(n4009), .A2(n4008), .A3(n4007), .A4(n4006), .ZN(n4010)
         );
  OR2_X1 U5053 ( .A1(n4011), .A2(n4010), .ZN(n4015) );
  INV_X1 U5054 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4013) );
  OAI22_X1 U5055 ( .A1(n4197), .A2(n4013), .B1(n4012), .B2(n4154), .ZN(n4014)
         );
  AOI21_X1 U5056 ( .B1(n4175), .B2(n4015), .A(n4014), .ZN(n4016) );
  NAND2_X1 U5057 ( .A1(n4017), .A2(n4016), .ZN(n5696) );
  INV_X1 U5058 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6955) );
  OAI21_X1 U5059 ( .B1(n4019), .B2(n4018), .A(n6955), .ZN(n4020) );
  NAND2_X1 U5060 ( .A1(n4021), .A2(n4020), .ZN(n5997) );
  NAND2_X1 U5061 ( .A1(n5997), .A2(n4261), .ZN(n4037) );
  AOI22_X1 U5062 ( .A1(n3478), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U5063 ( .A1(n4203), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U5064 ( .A1(n4254), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U5065 ( .A1(n4251), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4022) );
  NAND4_X1 U5066 ( .A1(n4025), .A2(n4024), .A3(n4023), .A4(n4022), .ZN(n4032)
         );
  AOI22_X1 U5067 ( .A1(n4273), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U5068 ( .A1(n3506), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4252), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U5069 ( .A1(n4279), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U5070 ( .A1(n4270), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4026) );
  NAND4_X1 U5071 ( .A1(n4029), .A2(n4028), .A3(n4027), .A4(n4026), .ZN(n4031)
         );
  OAI21_X1 U5072 ( .B1(n4032), .B2(n4031), .A(n4030), .ZN(n4035) );
  NAND2_X1 U5073 ( .A1(n3815), .A2(EAX_REG_15__SCAN_IN), .ZN(n4034) );
  NAND2_X1 U5074 ( .A1(n4294), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4033)
         );
  AND3_X1 U5075 ( .A1(n4035), .A2(n4034), .A3(n4033), .ZN(n4036) );
  NAND2_X1 U5076 ( .A1(n4037), .A2(n4036), .ZN(n5654) );
  XNOR2_X1 U5077 ( .A(n4053), .B(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5959)
         );
  AOI22_X1 U5078 ( .A1(n4225), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5079 ( .A1(n3478), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5080 ( .A1(n4203), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U5081 ( .A1(n4280), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4038) );
  NAND4_X1 U5082 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4038), .ZN(n4047)
         );
  AOI22_X1 U5083 ( .A1(n3506), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5084 ( .A1(n4252), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5085 ( .A1(n3460), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5086 ( .A1(n4254), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U5087 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4046)
         );
  OR2_X1 U5088 ( .A1(n4047), .A2(n4046), .ZN(n4051) );
  INV_X1 U5089 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4049) );
  OAI21_X1 U5090 ( .B1(n6371), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6345), 
        .ZN(n4048) );
  OAI21_X1 U5091 ( .B1(n4197), .B2(n4049), .A(n4048), .ZN(n4050) );
  AOI21_X1 U5092 ( .B1(n4175), .B2(n4051), .A(n4050), .ZN(n4052) );
  AOI21_X1 U5093 ( .B1(n5959), .B2(n3849), .A(n4052), .ZN(n5636) );
  INV_X1 U5094 ( .A(n4055), .ZN(n4057) );
  INV_X1 U5095 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4056) );
  NAND2_X1 U5096 ( .A1(n4057), .A2(n4056), .ZN(n4058) );
  NAND2_X1 U5097 ( .A1(n4092), .A2(n4058), .ZN(n5947) );
  AOI22_X1 U5098 ( .A1(n3478), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5099 ( .A1(n3506), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4254), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5100 ( .A1(n4203), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5101 ( .A1(n4252), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4059) );
  NAND4_X1 U5102 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4068)
         );
  AOI22_X1 U5103 ( .A1(n4225), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5104 ( .A1(n4280), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5105 ( .A1(n3460), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5106 ( .A1(n4269), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4063) );
  NAND4_X1 U5107 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4067)
         );
  NOR2_X1 U5108 ( .A1(n4068), .A2(n4067), .ZN(n4072) );
  NAND2_X1 U5109 ( .A1(n6345), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4069)
         );
  NAND2_X1 U5110 ( .A1(n3814), .A2(n4069), .ZN(n4070) );
  AOI21_X1 U5111 ( .B1(n3815), .B2(EAX_REG_20__SCAN_IN), .A(n4070), .ZN(n4071)
         );
  OAI21_X1 U5112 ( .B1(n4289), .B2(n4072), .A(n4071), .ZN(n4073) );
  NAND2_X1 U5113 ( .A1(n4074), .A2(n4073), .ZN(n5623) );
  XNOR2_X1 U5114 ( .A(n4092), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5940)
         );
  NAND2_X1 U5115 ( .A1(n5940), .A2(n4261), .ZN(n4090) );
  AOI22_X1 U5116 ( .A1(n4225), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5117 ( .A1(n3506), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4254), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5118 ( .A1(n4270), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5119 ( .A1(n4252), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4075) );
  NAND4_X1 U5120 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4084)
         );
  AOI22_X1 U5121 ( .A1(n4203), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5122 ( .A1(n3478), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5123 ( .A1(n4273), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5124 ( .A1(n4269), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4079) );
  NAND4_X1 U5125 ( .A1(n4082), .A2(n4081), .A3(n4080), .A4(n4079), .ZN(n4083)
         );
  NOR2_X1 U5126 ( .A1(n4084), .A2(n4083), .ZN(n4088) );
  NAND2_X1 U5127 ( .A1(n6345), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4085)
         );
  NAND2_X1 U5128 ( .A1(n3814), .A2(n4085), .ZN(n4086) );
  AOI21_X1 U5129 ( .B1(n3815), .B2(EAX_REG_21__SCAN_IN), .A(n4086), .ZN(n4087)
         );
  OAI21_X1 U5130 ( .B1(n4289), .B2(n4088), .A(n4087), .ZN(n4089) );
  INV_X1 U5131 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5938) );
  INV_X1 U5132 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6980) );
  OAI21_X1 U5133 ( .B1(n4092), .B2(n5938), .A(n6980), .ZN(n4093) );
  NAND2_X1 U5134 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4091) );
  AND2_X1 U5135 ( .A1(n4093), .A2(n4110), .ZN(n5930) );
  NAND2_X1 U5136 ( .A1(n5930), .A2(n4261), .ZN(n4108) );
  AOI22_X1 U5137 ( .A1(n4225), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5138 ( .A1(n3506), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4252), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5139 ( .A1(n3460), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U5140 ( .A1(n4203), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4094) );
  NAND4_X1 U5141 ( .A1(n4097), .A2(n4096), .A3(n4095), .A4(n4094), .ZN(n4103)
         );
  AOI22_X1 U5142 ( .A1(n3478), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5143 ( .A1(n4280), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5144 ( .A1(n4254), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U5145 ( .A1(n4251), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4098) );
  NAND4_X1 U5146 ( .A1(n4101), .A2(n4100), .A3(n4099), .A4(n4098), .ZN(n4102)
         );
  NOR2_X1 U5147 ( .A1(n4103), .A2(n4102), .ZN(n4106) );
  OAI21_X1 U5148 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6980), .A(n3814), .ZN(
        n4104) );
  AOI21_X1 U5149 ( .B1(n3815), .B2(EAX_REG_22__SCAN_IN), .A(n4104), .ZN(n4105)
         );
  OAI21_X1 U5150 ( .B1(n4289), .B2(n4106), .A(n4105), .ZN(n4107) );
  NAND2_X1 U5151 ( .A1(n4108), .A2(n4107), .ZN(n5597) );
  INV_X1 U5152 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6901) );
  NAND2_X1 U5153 ( .A1(n4110), .A2(n6901), .ZN(n4111) );
  NAND2_X1 U5154 ( .A1(n4137), .A2(n4111), .ZN(n5921) );
  AOI22_X1 U5155 ( .A1(n4279), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5156 ( .A1(n3478), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5157 ( .A1(n4203), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U5158 ( .A1(n4280), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4112) );
  NAND4_X1 U5159 ( .A1(n4115), .A2(n4114), .A3(n4113), .A4(n4112), .ZN(n4121)
         );
  AOI22_X1 U5160 ( .A1(n3506), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5161 ( .A1(n4252), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5162 ( .A1(n4273), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U5163 ( .A1(n4254), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4116) );
  NAND4_X1 U5164 ( .A1(n4119), .A2(n4118), .A3(n4117), .A4(n4116), .ZN(n4120)
         );
  AOI22_X1 U5165 ( .A1(n4279), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5166 ( .A1(n3478), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5167 ( .A1(n4203), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5168 ( .A1(n4280), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4122) );
  NAND4_X1 U5169 ( .A1(n4125), .A2(n4124), .A3(n4123), .A4(n4122), .ZN(n4131)
         );
  AOI22_X1 U5170 ( .A1(n3506), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5171 ( .A1(n4252), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5172 ( .A1(n3460), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4127) );
  INV_X1 U5173 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n7009) );
  AOI22_X1 U5174 ( .A1(n4254), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4126) );
  NAND4_X1 U5175 ( .A1(n4129), .A2(n4128), .A3(n4127), .A4(n4126), .ZN(n4130)
         );
  XNOR2_X1 U5176 ( .A(n4140), .B(n4139), .ZN(n4134) );
  OAI21_X1 U5177 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6901), .A(n3814), .ZN(
        n4132) );
  AOI21_X1 U5178 ( .B1(n3815), .B2(EAX_REG_23__SCAN_IN), .A(n4132), .ZN(n4133)
         );
  OAI21_X1 U5179 ( .B1(n4289), .B2(n4134), .A(n4133), .ZN(n4135) );
  NAND2_X1 U5180 ( .A1(n4137), .A2(n4153), .ZN(n4138) );
  NAND2_X1 U5181 ( .A1(n4177), .A2(n4138), .ZN(n5912) );
  NAND2_X1 U5182 ( .A1(n5912), .A2(n4261), .ZN(n4159) );
  NAND2_X1 U5183 ( .A1(n4140), .A2(n4139), .ZN(n4152) );
  AOI22_X1 U5184 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n4225), .B1(n4278), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5185 ( .A1(n3478), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U5186 ( .A1(n4203), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5187 ( .A1(n4280), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4141) );
  NAND4_X1 U5188 ( .A1(n4144), .A2(n4143), .A3(n4142), .A4(n4141), .ZN(n4150)
         );
  AOI22_X1 U5189 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n3506), .B1(n4269), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5190 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n4252), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5191 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n4273), .B1(n4253), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5192 ( .A1(n4254), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4145) );
  NAND4_X1 U5193 ( .A1(n4148), .A2(n4147), .A3(n4146), .A4(n4145), .ZN(n4149)
         );
  NOR2_X1 U5194 ( .A1(n4150), .A2(n4149), .ZN(n4151) );
  NOR2_X1 U5195 ( .A1(n4151), .A2(n4152), .ZN(n4183) );
  AOI21_X1 U5196 ( .B1(n4152), .B2(n4151), .A(n4183), .ZN(n4157) );
  INV_X1 U5197 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4155) );
  OAI22_X1 U5198 ( .A1(n4197), .A2(n4155), .B1(n4154), .B2(n4153), .ZN(n4156)
         );
  AOI21_X1 U5199 ( .B1(n4175), .B2(n4157), .A(n4156), .ZN(n4158) );
  NAND2_X1 U5200 ( .A1(n4159), .A2(n4158), .ZN(n5572) );
  XNOR2_X1 U5201 ( .A(n4177), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5893)
         );
  AOI22_X1 U5202 ( .A1(n4225), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U5203 ( .A1(n3478), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U5204 ( .A1(n4203), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U5205 ( .A1(n4280), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4160) );
  NAND4_X1 U5206 ( .A1(n4163), .A2(n4162), .A3(n4161), .A4(n4160), .ZN(n4169)
         );
  AOI22_X1 U5207 ( .A1(n3506), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U5208 ( .A1(n4252), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U5209 ( .A1(n4273), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U5210 ( .A1(n4254), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4164) );
  NAND4_X1 U5211 ( .A1(n4167), .A2(n4166), .A3(n4165), .A4(n4164), .ZN(n4168)
         );
  INV_X1 U5212 ( .A(n4183), .ZN(n4170) );
  XNOR2_X1 U5213 ( .A(n4182), .B(n4170), .ZN(n4174) );
  INV_X1 U5214 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4172) );
  NAND2_X1 U5215 ( .A1(n6345), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4171)
         );
  OAI211_X1 U5216 ( .C1(n4197), .C2(n4172), .A(n3814), .B(n4171), .ZN(n4173)
         );
  AOI21_X1 U5217 ( .B1(n4175), .B2(n4174), .A(n4173), .ZN(n4176) );
  NAND2_X1 U5218 ( .A1(n5560), .A2(n5561), .ZN(n5548) );
  NAND2_X1 U5219 ( .A1(n4180), .A2(n4179), .ZN(n4181) );
  NAND2_X1 U5220 ( .A1(n4220), .A2(n4181), .ZN(n5881) );
  NAND2_X1 U5221 ( .A1(n4183), .A2(n4182), .ZN(n4201) );
  AOI22_X1 U5222 ( .A1(n3478), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U5223 ( .A1(n3506), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4254), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U5224 ( .A1(n4280), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U5225 ( .A1(n4271), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4184) );
  NAND4_X1 U5226 ( .A1(n4187), .A2(n4186), .A3(n4185), .A4(n4184), .ZN(n4194)
         );
  AOI22_X1 U5227 ( .A1(n4279), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U5228 ( .A1(n4203), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U5229 ( .A1(n4273), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U5230 ( .A1(n4269), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4189) );
  NAND4_X1 U5231 ( .A1(n4192), .A2(n4191), .A3(n4190), .A4(n4189), .ZN(n4193)
         );
  NOR2_X1 U5232 ( .A1(n4194), .A2(n4193), .ZN(n4202) );
  XNOR2_X1 U5233 ( .A(n4201), .B(n4202), .ZN(n4195) );
  NOR2_X1 U5234 ( .A1(n4195), .A2(n4289), .ZN(n4199) );
  INV_X1 U5235 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6526) );
  OAI21_X1 U5236 ( .B1(n6371), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6345), 
        .ZN(n4196) );
  OAI21_X1 U5237 ( .B1(n4197), .B2(n6526), .A(n4196), .ZN(n4198) );
  OAI22_X1 U5238 ( .A1(n5881), .A2(n3814), .B1(n4199), .B2(n4198), .ZN(n5550)
         );
  XNOR2_X1 U5239 ( .A(n4220), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5873)
         );
  NAND2_X1 U5240 ( .A1(n5873), .A2(n4261), .ZN(n4219) );
  NOR2_X1 U5241 ( .A1(n4202), .A2(n4201), .ZN(n4237) );
  AOI22_X1 U5242 ( .A1(n4279), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U5243 ( .A1(n3478), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4206) );
  AOI22_X1 U5244 ( .A1(n4203), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U5245 ( .A1(n4280), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4204) );
  NAND4_X1 U5246 ( .A1(n4207), .A2(n4206), .A3(n4205), .A4(n4204), .ZN(n4213)
         );
  AOI22_X1 U5247 ( .A1(n3506), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4211) );
  AOI22_X1 U5248 ( .A1(n4252), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4210) );
  AOI22_X1 U5249 ( .A1(n4273), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U5250 ( .A1(n4254), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4208) );
  NAND4_X1 U5251 ( .A1(n4211), .A2(n4210), .A3(n4209), .A4(n4208), .ZN(n4212)
         );
  XNOR2_X1 U5252 ( .A(n4237), .B(n4236), .ZN(n4217) );
  NAND2_X1 U5253 ( .A1(n6345), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4214)
         );
  NAND2_X1 U5254 ( .A1(n3814), .A2(n4214), .ZN(n4215) );
  AOI21_X1 U5255 ( .B1(n3815), .B2(EAX_REG_27__SCAN_IN), .A(n4215), .ZN(n4216)
         );
  OAI21_X1 U5256 ( .B1(n4217), .B2(n4289), .A(n4216), .ZN(n4218) );
  NAND2_X1 U5257 ( .A1(n4219), .A2(n4218), .ZN(n4459) );
  INV_X1 U5258 ( .A(n4220), .ZN(n4221) );
  NAND2_X1 U5259 ( .A1(n4221), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4223)
         );
  INV_X1 U5260 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4222) );
  NAND2_X1 U5261 ( .A1(n4223), .A2(n4222), .ZN(n4224) );
  NAND2_X1 U5262 ( .A1(n4266), .A2(n4224), .ZN(n5862) );
  AOI22_X1 U5263 ( .A1(n4225), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3478), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4229) );
  AOI22_X1 U5264 ( .A1(n3506), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4254), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U5265 ( .A1(n3460), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4227) );
  AOI22_X1 U5266 ( .A1(n4203), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4226) );
  NAND4_X1 U5267 ( .A1(n4229), .A2(n4228), .A3(n4227), .A4(n4226), .ZN(n4235)
         );
  AOI22_X1 U5268 ( .A1(n4270), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U5269 ( .A1(n4271), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4232) );
  AOI22_X1 U5270 ( .A1(n4280), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4231) );
  AOI22_X1 U5271 ( .A1(n4253), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4230) );
  NAND4_X1 U5272 ( .A1(n4233), .A2(n4232), .A3(n4231), .A4(n4230), .ZN(n4234)
         );
  NOR2_X1 U5273 ( .A1(n4235), .A2(n4234), .ZN(n4246) );
  NAND2_X1 U5274 ( .A1(n4237), .A2(n4236), .ZN(n4245) );
  XNOR2_X1 U5275 ( .A(n4246), .B(n4245), .ZN(n4242) );
  NAND2_X1 U5276 ( .A1(n6345), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4238)
         );
  NAND2_X1 U5277 ( .A1(n3814), .A2(n4238), .ZN(n4239) );
  AOI21_X1 U5278 ( .B1(n4240), .B2(EAX_REG_28__SCAN_IN), .A(n4239), .ZN(n4241)
         );
  OAI21_X1 U5279 ( .B1(n4242), .B2(n4289), .A(n4241), .ZN(n4243) );
  INV_X1 U5280 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5517) );
  XNOR2_X1 U5281 ( .A(n4266), .B(n5517), .ZN(n5513) );
  NOR2_X1 U5282 ( .A1(n4246), .A2(n4245), .ZN(n4268) );
  AOI22_X1 U5283 ( .A1(n4279), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3535), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U5284 ( .A1(n3478), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4249) );
  AOI22_X1 U5285 ( .A1(n4203), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3500), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4248) );
  AOI22_X1 U5286 ( .A1(n4280), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3462), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4247) );
  NAND4_X1 U5287 ( .A1(n4250), .A2(n4249), .A3(n4248), .A4(n4247), .ZN(n4260)
         );
  AOI22_X1 U5288 ( .A1(n3506), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4258) );
  AOI22_X1 U5289 ( .A1(n4252), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4257) );
  AOI22_X1 U5290 ( .A1(n4273), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4253), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4256) );
  AOI22_X1 U5291 ( .A1(n4254), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4255) );
  NAND4_X1 U5292 ( .A1(n4258), .A2(n4257), .A3(n4256), .A4(n4255), .ZN(n4259)
         );
  OR2_X1 U5293 ( .A1(n4260), .A2(n4259), .ZN(n4267) );
  XNOR2_X1 U5294 ( .A(n4268), .B(n4267), .ZN(n4264) );
  AOI21_X1 U5295 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6345), .A(n4261), 
        .ZN(n4263) );
  NAND2_X1 U5296 ( .A1(n3815), .A2(EAX_REG_29__SCAN_IN), .ZN(n4262) );
  OAI211_X1 U5297 ( .C1(n4264), .C2(n4289), .A(n4263), .B(n4262), .ZN(n4265)
         );
  NOR2_X2 U5298 ( .A1(n4466), .A2(n4467), .ZN(n4307) );
  XNOR2_X1 U5299 ( .A(n4297), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5490)
         );
  OAI21_X1 U5300 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6918), .A(n3814), .ZN(
        n4292) );
  NAND2_X1 U5301 ( .A1(n4268), .A2(n4267), .ZN(n4288) );
  AOI22_X1 U5302 ( .A1(n3467), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4269), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U5303 ( .A1(n3478), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U5304 ( .A1(n4271), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U5305 ( .A1(n4273), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4274) );
  NAND4_X1 U5306 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4286)
         );
  AOI22_X1 U5307 ( .A1(n4279), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4278), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4284) );
  AOI22_X1 U5308 ( .A1(n4203), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4283) );
  AOI22_X1 U5309 ( .A1(n3500), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3484), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4282) );
  AOI22_X1 U5310 ( .A1(n3506), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3406), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4281) );
  NAND4_X1 U5311 ( .A1(n4284), .A2(n4283), .A3(n4282), .A4(n4281), .ZN(n4285)
         );
  NOR2_X1 U5312 ( .A1(n4286), .A2(n4285), .ZN(n4287) );
  XNOR2_X1 U5313 ( .A(n4288), .B(n4287), .ZN(n4290) );
  NOR2_X1 U5314 ( .A1(n4290), .A2(n4289), .ZN(n4291) );
  AOI211_X1 U5315 ( .C1(n3815), .C2(EAX_REG_30__SCAN_IN), .A(n4292), .B(n4291), 
        .ZN(n4293) );
  AOI22_X1 U5316 ( .A1(n3815), .A2(EAX_REG_31__SCAN_IN), .B1(n4294), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4295) );
  INV_X1 U5317 ( .A(n4295), .ZN(n4296) );
  NAND2_X1 U5318 ( .A1(n4584), .A2(n6571), .ZN(n4305) );
  NAND2_X1 U5319 ( .A1(n4299), .A2(n6722), .ZN(n6840) );
  NAND2_X1 U5320 ( .A1(n6840), .A2(n6938), .ZN(n4300) );
  NAND2_X1 U5321 ( .A1(n6371), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4581) );
  NAND2_X1 U5322 ( .A1(n6938), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4301) );
  NAND2_X1 U5323 ( .A1(n4581), .A2(n4301), .ZN(n4775) );
  NOR2_X1 U5324 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6360) );
  AND2_X2 U5325 ( .A1(n6357), .A2(n6360), .ZN(n6566) );
  NAND2_X1 U5326 ( .A1(n6566), .A2(REIP_REG_31__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U5327 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4302)
         );
  OAI211_X1 U5328 ( .C1(n5426), .C2(n6586), .A(n4525), .B(n4302), .ZN(n4303)
         );
  INV_X1 U5329 ( .A(n4303), .ZN(n4304) );
  INV_X1 U5330 ( .A(n4307), .ZN(n4468) );
  INV_X1 U5331 ( .A(n4308), .ZN(n4309) );
  NAND2_X1 U5332 ( .A1(n4468), .A2(n4309), .ZN(n4311) );
  NAND2_X1 U5333 ( .A1(n4311), .A2(n4310), .ZN(n4577) );
  NOR2_X1 U5334 ( .A1(n4496), .A2(n5510), .ZN(n4729) );
  NAND2_X1 U5335 ( .A1(n4709), .A2(n4729), .ZN(n4320) );
  AND3_X1 U5336 ( .A1(n4315), .A2(n4314), .A3(n4313), .ZN(n4317) );
  OAI21_X1 U5337 ( .B1(n4318), .B2(n4317), .A(n4316), .ZN(n4673) );
  NAND2_X1 U5338 ( .A1(n4673), .A2(n6838), .ZN(n4483) );
  OR2_X1 U5339 ( .A1(n4312), .A2(n4483), .ZN(n4319) );
  INV_X1 U5340 ( .A(n4353), .ZN(n4853) );
  NAND2_X1 U5341 ( .A1(n4853), .A2(n6355), .ZN(n4323) );
  NOR2_X1 U5342 ( .A1(n4321), .A2(n4348), .ZN(n4324) );
  NAND2_X1 U5343 ( .A1(n4333), .A2(n4353), .ZN(n4805) );
  AOI22_X1 U5344 ( .A1(n5838), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n5850), .ZN(n4327) );
  NOR3_X1 U5345 ( .A1(n5850), .A2(n4853), .A3(n4328), .ZN(n4329) );
  OAI21_X1 U5346 ( .B1(n4577), .B2(n5859), .A(n4331), .ZN(U2861) );
  INV_X1 U5347 ( .A(n6355), .ZN(n6365) );
  AND2_X1 U5348 ( .A1(n4333), .A2(n3182), .ZN(n4494) );
  NAND2_X1 U5349 ( .A1(n4493), .A2(n4494), .ZN(n4338) );
  NAND2_X1 U5350 ( .A1(n4843), .A2(n5456), .ZN(n4341) );
  NOR2_X1 U5351 ( .A1(n4341), .A2(n3435), .ZN(n4683) );
  OAI21_X1 U5352 ( .B1(n4683), .B2(n4791), .A(n3591), .ZN(n4337) );
  INV_X1 U5353 ( .A(n4335), .ZN(n4336) );
  NAND2_X1 U5354 ( .A1(n4332), .A2(n4339), .ZN(n4713) );
  INV_X1 U5355 ( .A(n4347), .ZN(n4745) );
  NOR2_X1 U5356 ( .A1(n4341), .A2(n4340), .ZN(n4342) );
  NAND2_X1 U5357 ( .A1(n4745), .A2(n4342), .ZN(n4887) );
  NAND2_X1 U5358 ( .A1(n4343), .A2(n5456), .ZN(n4344) );
  OAI211_X1 U5359 ( .C1(n4345), .C2(n4321), .A(n4887), .B(n4344), .ZN(n4346)
         );
  NOR2_X1 U5360 ( .A1(n4347), .A2(n3435), .ZN(n4502) );
  NAND2_X1 U5361 ( .A1(n4530), .A2(n4502), .ZN(n4731) );
  INV_X1 U5362 ( .A(n4348), .ZN(n4350) );
  NAND3_X1 U5363 ( .A1(n4350), .A2(n4800), .A3(n4349), .ZN(n4351) );
  INV_X2 U5364 ( .A(n6479), .ZN(n6474) );
  NOR2_X1 U5365 ( .A1(n4791), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4354)
         );
  NOR2_X2 U5366 ( .A1(n4355), .A2(n4354), .ZN(n4976) );
  NAND2_X1 U5367 ( .A1(n4442), .A2(n3616), .ZN(n4356) );
  OAI211_X1 U5368 ( .C1(n4360), .C2(EBX_REG_2__SCAN_IN), .A(n4371), .B(n4356), 
        .ZN(n4358) );
  INV_X1 U5369 ( .A(EBX_REG_2__SCAN_IN), .ZN(n7066) );
  NAND2_X1 U5370 ( .A1(n3300), .A2(n7066), .ZN(n4357) );
  NAND2_X1 U5371 ( .A1(n4358), .A2(n4357), .ZN(n5476) );
  NAND2_X1 U5372 ( .A1(n4442), .A2(n7101), .ZN(n4359) );
  OAI211_X1 U5373 ( .C1(n4360), .C2(EBX_REG_1__SCAN_IN), .A(n4371), .B(n4359), 
        .ZN(n4363) );
  INV_X1 U5374 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4361) );
  NAND2_X1 U5375 ( .A1(n5638), .A2(n4361), .ZN(n4362) );
  NAND2_X1 U5376 ( .A1(n4363), .A2(n4362), .ZN(n4366) );
  NAND2_X1 U5377 ( .A1(n4442), .A2(EBX_REG_0__SCAN_IN), .ZN(n4365) );
  INV_X1 U5378 ( .A(EBX_REG_0__SCAN_IN), .ZN(n7050) );
  NAND2_X1 U5379 ( .A1(n4371), .A2(n7050), .ZN(n4364) );
  NAND2_X1 U5380 ( .A1(n4365), .A2(n4364), .ZN(n4790) );
  XNOR2_X1 U5381 ( .A(n4366), .B(n4790), .ZN(n4801) );
  NAND2_X1 U5382 ( .A1(n4801), .A2(n4800), .ZN(n4802) );
  INV_X1 U5383 ( .A(n4366), .ZN(n4367) );
  NAND2_X1 U5384 ( .A1(n4367), .A2(n4790), .ZN(n4368) );
  NAND2_X1 U5385 ( .A1(n4802), .A2(n4368), .ZN(n5477) );
  INV_X2 U5386 ( .A(n4371), .ZN(n5638) );
  INV_X1 U5387 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4372) );
  MUX2_X1 U5388 ( .A(n5638), .B(n4378), .S(n4372), .Z(n4374) );
  NOR2_X1 U5389 ( .A1(n4791), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4373)
         );
  NOR2_X1 U5390 ( .A1(n4374), .A2(n4373), .ZN(n5292) );
  MUX2_X1 U5391 ( .A(n5638), .B(n4430), .S(EBX_REG_4__SCAN_IN), .Z(n4375) );
  INV_X1 U5392 ( .A(n4375), .ZN(n4377) );
  NAND2_X1 U5393 ( .A1(n4360), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4376)
         );
  NAND2_X1 U5394 ( .A1(n4377), .A2(n4376), .ZN(n6428) );
  MUX2_X1 U5395 ( .A(n4378), .B(n5638), .S(EBX_REG_7__SCAN_IN), .Z(n4379) );
  INV_X1 U5396 ( .A(n4379), .ZN(n4382) );
  NAND2_X1 U5397 ( .A1(n4446), .A2(n4380), .ZN(n4381) );
  NAND2_X1 U5398 ( .A1(n4382), .A2(n4381), .ZN(n5764) );
  MUX2_X1 U5399 ( .A(n5638), .B(n4430), .S(EBX_REG_6__SCAN_IN), .Z(n4384) );
  AND2_X1 U5400 ( .A1(n4360), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4383)
         );
  NOR2_X1 U5401 ( .A1(n4384), .A2(n4383), .ZN(n5763) );
  NOR2_X1 U5402 ( .A1(n5764), .A2(n5763), .ZN(n4385) );
  NAND2_X1 U5403 ( .A1(n4442), .A2(n4386), .ZN(n4387) );
  OAI211_X1 U5404 ( .C1(n4360), .C2(EBX_REG_8__SCAN_IN), .A(n5626), .B(n4387), 
        .ZN(n4390) );
  INV_X1 U5405 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U5406 ( .A1(n5638), .A2(n4388), .ZN(n4389) );
  NAND2_X1 U5407 ( .A1(n4390), .A2(n4389), .ZN(n5750) );
  INV_X1 U5408 ( .A(n5748), .ZN(n4394) );
  MUX2_X1 U5409 ( .A(n4378), .B(n5638), .S(EBX_REG_9__SCAN_IN), .Z(n4391) );
  INV_X1 U5410 ( .A(n4391), .ZN(n4393) );
  NAND2_X1 U5411 ( .A1(n4446), .A2(n6593), .ZN(n4392) );
  MUX2_X1 U5412 ( .A(n5638), .B(n4430), .S(EBX_REG_10__SCAN_IN), .Z(n4396) );
  AND2_X1 U5413 ( .A1(n4360), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4395)
         );
  NOR2_X1 U5414 ( .A1(n4396), .A2(n4395), .ZN(n5427) );
  NAND2_X1 U5415 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4397) );
  OAI211_X1 U5416 ( .C1(n4360), .C2(EBX_REG_11__SCAN_IN), .A(n4442), .B(n4397), 
        .ZN(n4398) );
  OAI21_X1 U5417 ( .B1(n4441), .B2(EBX_REG_11__SCAN_IN), .A(n4398), .ZN(n6247)
         );
  MUX2_X1 U5418 ( .A(n5638), .B(n4430), .S(EBX_REG_12__SCAN_IN), .Z(n4399) );
  INV_X1 U5419 ( .A(n4399), .ZN(n4401) );
  NAND2_X1 U5420 ( .A1(n4360), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4400) );
  NAND2_X1 U5421 ( .A1(n4401), .A2(n4400), .ZN(n5736) );
  NAND2_X1 U5422 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4402) );
  OAI211_X1 U5423 ( .C1(n4360), .C2(EBX_REG_13__SCAN_IN), .A(n4442), .B(n4402), 
        .ZN(n4403) );
  OAI21_X1 U5424 ( .B1(n4441), .B2(EBX_REG_13__SCAN_IN), .A(n4403), .ZN(n5719)
         );
  MUX2_X1 U5425 ( .A(n5638), .B(n4430), .S(EBX_REG_14__SCAN_IN), .Z(n4405) );
  AND2_X1 U5426 ( .A1(n4360), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4404)
         );
  NOR2_X1 U5427 ( .A1(n4405), .A2(n4404), .ZN(n5499) );
  INV_X1 U5428 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U5429 ( .A1(n4378), .A2(n5789), .ZN(n4409) );
  NAND2_X1 U5430 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4407) );
  OAI211_X1 U5431 ( .C1(n4360), .C2(EBX_REG_15__SCAN_IN), .A(n4442), .B(n4407), 
        .ZN(n4408) );
  MUX2_X1 U5432 ( .A(n5638), .B(n4430), .S(EBX_REG_16__SCAN_IN), .Z(n4410) );
  INV_X1 U5433 ( .A(n4410), .ZN(n4412) );
  NAND2_X1 U5434 ( .A1(n4360), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4411) );
  NAND2_X1 U5435 ( .A1(n4412), .A2(n4411), .ZN(n5684) );
  NAND2_X1 U5436 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4413) );
  OAI211_X1 U5437 ( .C1(n4360), .C2(EBX_REG_17__SCAN_IN), .A(n4442), .B(n4413), 
        .ZN(n4414) );
  OAI21_X1 U5438 ( .B1(n4441), .B2(EBX_REG_17__SCAN_IN), .A(n4414), .ZN(n5672)
         );
  INV_X1 U5439 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U5440 ( .A1(n4442), .A2(n5897), .ZN(n4415) );
  OAI211_X1 U5441 ( .C1(n4360), .C2(EBX_REG_19__SCAN_IN), .A(n5626), .B(n4415), 
        .ZN(n4417) );
  INV_X1 U5442 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U5443 ( .A1(n5638), .A2(n5644), .ZN(n4416) );
  NOR2_X2 U5444 ( .A1(n5674), .A2(n5642), .ZN(n5624) );
  INV_X1 U5445 ( .A(EBX_REG_20__SCAN_IN), .ZN(n7141) );
  NAND2_X1 U5446 ( .A1(n4446), .A2(n6184), .ZN(n4418) );
  OR2_X1 U5447 ( .A1(n4360), .A2(EBX_REG_18__SCAN_IN), .ZN(n5637) );
  OR2_X1 U5448 ( .A1(n4360), .A2(EBX_REG_20__SCAN_IN), .ZN(n4419) );
  OAI21_X1 U5449 ( .B1(n4791), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n4419), 
        .ZN(n5627) );
  NAND2_X1 U5450 ( .A1(n5640), .A2(n5627), .ZN(n4421) );
  INV_X1 U5451 ( .A(n5640), .ZN(n5625) );
  NAND2_X1 U5452 ( .A1(n5625), .A2(n5626), .ZN(n4420) );
  OAI211_X1 U5453 ( .C1(n5626), .C2(n7141), .A(n4421), .B(n4420), .ZN(n4422)
         );
  INV_X1 U5454 ( .A(n4422), .ZN(n4423) );
  MUX2_X1 U5455 ( .A(n4378), .B(n5638), .S(EBX_REG_21__SCAN_IN), .Z(n4425) );
  NOR2_X1 U5456 ( .A1(n4791), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4424)
         );
  NOR2_X1 U5457 ( .A1(n4425), .A2(n4424), .ZN(n5610) );
  MUX2_X1 U5458 ( .A(n5638), .B(n4430), .S(EBX_REG_22__SCAN_IN), .Z(n4427) );
  AND2_X1 U5459 ( .A1(n4360), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4426)
         );
  NOR2_X1 U5460 ( .A1(n4427), .A2(n4426), .ZN(n5599) );
  NAND2_X1 U5461 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4428) );
  OAI211_X1 U5462 ( .C1(n4360), .C2(EBX_REG_23__SCAN_IN), .A(n4442), .B(n4428), 
        .ZN(n4429) );
  OAI21_X1 U5463 ( .B1(n4441), .B2(EBX_REG_23__SCAN_IN), .A(n4429), .ZN(n5585)
         );
  MUX2_X1 U5464 ( .A(n5638), .B(n4430), .S(EBX_REG_24__SCAN_IN), .Z(n4432) );
  AND2_X1 U5465 ( .A1(n4360), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4431)
         );
  NOR2_X1 U5466 ( .A1(n4432), .A2(n4431), .ZN(n5575) );
  MUX2_X1 U5467 ( .A(n4378), .B(n5638), .S(EBX_REG_25__SCAN_IN), .Z(n4434) );
  NOR2_X1 U5468 ( .A1(n4791), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4433)
         );
  NOR2_X1 U5469 ( .A1(n4434), .A2(n4433), .ZN(n5563) );
  INV_X1 U5470 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U5471 ( .A1(n4442), .A2(n5865), .ZN(n4435) );
  OAI211_X1 U5472 ( .C1(n4360), .C2(EBX_REG_26__SCAN_IN), .A(n5626), .B(n4435), 
        .ZN(n4438) );
  INV_X1 U5473 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U5474 ( .A1(n5638), .A2(n4436), .ZN(n4437) );
  NAND2_X1 U5475 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4439) );
  OAI211_X1 U5476 ( .C1(n4360), .C2(EBX_REG_27__SCAN_IN), .A(n4442), .B(n4439), 
        .ZN(n4440) );
  OAI21_X1 U5477 ( .B1(n4441), .B2(EBX_REG_27__SCAN_IN), .A(n4440), .ZN(n4461)
         );
  NAND2_X1 U5478 ( .A1(n4442), .A2(n5867), .ZN(n4443) );
  OAI211_X1 U5479 ( .C1(n4360), .C2(EBX_REG_28__SCAN_IN), .A(n5626), .B(n4443), 
        .ZN(n4445) );
  INV_X1 U5480 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U5481 ( .A1(n5638), .A2(n5778), .ZN(n4444) );
  NAND2_X1 U5482 ( .A1(n4445), .A2(n4444), .ZN(n5525) );
  INV_X1 U5483 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U5484 ( .A1(n4446), .A2(n6082), .ZN(n4512) );
  INV_X1 U5485 ( .A(EBX_REG_29__SCAN_IN), .ZN(n7140) );
  NAND2_X1 U5486 ( .A1(n4800), .A2(n7140), .ZN(n4447) );
  NAND2_X1 U5487 ( .A1(n4512), .A2(n4447), .ZN(n4448) );
  OR2_X2 U5488 ( .A1(n5528), .A2(n4448), .ZN(n4452) );
  INV_X1 U5489 ( .A(n4452), .ZN(n4451) );
  NAND2_X1 U5490 ( .A1(n4791), .A2(EBX_REG_30__SCAN_IN), .ZN(n4450) );
  NAND2_X1 U5491 ( .A1(n4360), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U5492 ( .A1(n4450), .A2(n4449), .ZN(n4518) );
  OAI211_X1 U5493 ( .C1(n4451), .C2(n5528), .A(n4517), .B(n4518), .ZN(n4455)
         );
  INV_X1 U5494 ( .A(n5528), .ZN(n4563) );
  INV_X1 U5495 ( .A(n4518), .ZN(n4453) );
  OAI211_X1 U5496 ( .C1(n4563), .C2(n5626), .A(n4453), .B(n4452), .ZN(n4454)
         );
  INV_X1 U5497 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5486) );
  INV_X1 U5498 ( .A(n4456), .ZN(n4457) );
  OAI21_X1 U5499 ( .B1(n4577), .B2(n6474), .A(n4457), .ZN(U2829) );
  AND2_X1 U5500 ( .A1(n5553), .A2(n4461), .ZN(n4462) );
  OR2_X1 U5501 ( .A1(n4462), .A2(n5526), .ZN(n6096) );
  INV_X1 U5502 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6945) );
  NAND2_X1 U5503 ( .A1(n6566), .A2(REIP_REG_29__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U5504 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4470)
         );
  OAI211_X1 U5505 ( .C1(n5513), .C2(n6586), .A(n6079), .B(n4470), .ZN(n4471)
         );
  AOI21_X1 U5506 ( .B1(n5804), .B2(n6571), .A(n4471), .ZN(n4481) );
  INV_X1 U5507 ( .A(n4474), .ZN(n4473) );
  NOR3_X1 U5508 ( .A1(n4573), .A2(n4473), .A3(n6082), .ZN(n4478) );
  NAND2_X1 U5509 ( .A1(n4573), .A2(n6082), .ZN(n4476) );
  NAND2_X1 U5510 ( .A1(n4476), .A2(n4475), .ZN(n4477) );
  NOR2_X1 U5511 ( .A1(n4478), .A2(n4477), .ZN(n6084) );
  INV_X1 U5512 ( .A(n6084), .ZN(n4479) );
  NAND2_X1 U5513 ( .A1(n4479), .A2(n3784), .ZN(n4480) );
  NAND2_X1 U5514 ( .A1(n4481), .A2(n4480), .ZN(U2957) );
  NAND2_X1 U5515 ( .A1(n4482), .A2(n6815), .ZN(n4753) );
  NAND2_X1 U5516 ( .A1(n5455), .A2(n4753), .ZN(n4485) );
  INV_X1 U5517 ( .A(n4483), .ZN(n4484) );
  NAND2_X1 U5518 ( .A1(n4485), .A2(n4484), .ZN(n4492) );
  NAND2_X1 U5519 ( .A1(n3435), .A2(n4753), .ZN(n4587) );
  NAND2_X1 U5520 ( .A1(n4587), .A2(n6838), .ZN(n4489) );
  OAI211_X1 U5521 ( .C1(n4487), .C2(n4489), .A(n3182), .B(n4488), .ZN(n4490)
         );
  NAND2_X1 U5522 ( .A1(n4709), .A2(n4490), .ZN(n4491) );
  MUX2_X1 U5523 ( .A(n4492), .B(n4491), .S(n4843), .Z(n4505) );
  OAI21_X1 U5524 ( .B1(n4698), .B2(n4494), .A(n4493), .ZN(n4495) );
  INV_X1 U5525 ( .A(n4495), .ZN(n4497) );
  OR2_X1 U5526 ( .A1(n4497), .A2(n4496), .ZN(n4501) );
  INV_X1 U5527 ( .A(n4499), .ZN(n4500) );
  NAND2_X1 U5528 ( .A1(n4501), .A2(n4500), .ZN(n4685) );
  INV_X1 U5529 ( .A(n4502), .ZN(n4503) );
  OR2_X1 U5530 ( .A1(n4709), .A2(n4503), .ZN(n4504) );
  NAND3_X1 U5531 ( .A1(n4505), .A2(n4685), .A3(n4504), .ZN(n4506) );
  INV_X1 U5532 ( .A(n5351), .ZN(n4507) );
  OR2_X1 U5533 ( .A1(n4507), .A2(n4729), .ZN(n4671) );
  OR2_X1 U5534 ( .A1(n4487), .A2(n4360), .ZN(n4508) );
  NOR2_X1 U5535 ( .A1(n4671), .A2(n4510), .ZN(n4511) );
  INV_X1 U5536 ( .A(n4512), .ZN(n4513) );
  MUX2_X1 U5537 ( .A(n4513), .B(EBX_REG_29__SCAN_IN), .S(n5638), .Z(n4514) );
  INV_X1 U5538 ( .A(n4514), .ZN(n4516) );
  NAND2_X1 U5539 ( .A1(n4378), .A2(n7140), .ZN(n4515) );
  NAND2_X1 U5540 ( .A1(n4516), .A2(n4515), .ZN(n4560) );
  OAI22_X1 U5541 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n4791), .B1(n4360), .B2(EBX_REG_31__SCAN_IN), .ZN(n4519) );
  OR2_X1 U5542 ( .A1(n4321), .A2(n4522), .ZN(n4523) );
  AND2_X1 U5543 ( .A1(n5363), .A2(n4523), .ZN(n4524) );
  OAI21_X1 U5544 ( .B1(n5777), .B2(n6252), .A(n4525), .ZN(n4526) );
  INV_X1 U5545 ( .A(n4526), .ZN(n4558) );
  INV_X2 U5546 ( .A(n6238), .ZN(n6645) );
  AOI21_X1 U5547 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6647) );
  NAND2_X1 U5548 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6625) );
  NOR2_X1 U5549 ( .A1(n6647), .A2(n6625), .ZN(n5367) );
  NAND2_X1 U5550 ( .A1(n6645), .A2(n5367), .ZN(n5370) );
  NAND2_X1 U5551 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4527) );
  NOR2_X1 U5552 ( .A1(n5370), .A2(n4527), .ZN(n6268) );
  NAND2_X1 U5553 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U5554 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4528) );
  NOR2_X1 U5555 ( .A1(n6595), .A2(n4528), .ZN(n4532) );
  AND2_X1 U5556 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6237) );
  AND2_X1 U5557 ( .A1(n6237), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6217)
         );
  NAND2_X1 U5558 ( .A1(n6217), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U5559 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4529) );
  NOR2_X1 U5560 ( .A1(n6200), .A2(n4529), .ZN(n4533) );
  NAND2_X1 U5561 ( .A1(n6220), .A2(n4533), .ZN(n6156) );
  NAND2_X1 U5562 ( .A1(n4499), .A2(n5455), .ZN(n4878) );
  NOR2_X1 U5563 ( .A1(n4530), .A2(n4537), .ZN(n4538) );
  NAND2_X1 U5564 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4538), .ZN(n6221)
         );
  NOR2_X1 U5565 ( .A1(n7101), .A2(n3616), .ZN(n6646) );
  INV_X1 U5566 ( .A(n6646), .ZN(n4531) );
  NOR2_X1 U5567 ( .A1(n6625), .A2(n4531), .ZN(n5371) );
  AND3_X1 U5568 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n5371), .ZN(n6265) );
  AND2_X1 U5569 ( .A1(n4532), .A2(n6265), .ZN(n6199) );
  NAND2_X1 U5570 ( .A1(n6651), .A2(n6199), .ZN(n6239) );
  INV_X1 U5571 ( .A(n4533), .ZN(n4543) );
  NAND2_X1 U5572 ( .A1(n6156), .A2(n4534), .ZN(n6186) );
  NAND2_X1 U5573 ( .A1(n6186), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6178) );
  INV_X1 U5574 ( .A(n6164), .ZN(n4535) );
  NOR2_X1 U5575 ( .A1(n6172), .A2(n4535), .ZN(n6140) );
  AND2_X1 U5576 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U5577 ( .A1(n6117), .A2(n4550), .ZN(n6097) );
  OR2_X1 U5578 ( .A1(n6097), .A2(n6089), .ZN(n6077) );
  INV_X1 U5579 ( .A(n4536), .ZN(n4553) );
  NOR2_X1 U5580 ( .A1(n6077), .A2(n4553), .ZN(n4555) );
  NAND2_X1 U5581 ( .A1(n4537), .A2(n6577), .ZN(n4794) );
  INV_X1 U5582 ( .A(n6267), .ZN(n6155) );
  INV_X1 U5583 ( .A(n4538), .ZN(n4539) );
  NAND2_X1 U5584 ( .A1(n6266), .A2(n6267), .ZN(n4541) );
  NAND3_X1 U5585 ( .A1(n6164), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4540) );
  NAND2_X1 U5586 ( .A1(n4541), .A2(n4540), .ZN(n4545) );
  INV_X1 U5587 ( .A(n6199), .ZN(n4542) );
  NOR2_X1 U5588 ( .A1(n4543), .A2(n4542), .ZN(n4544) );
  OR2_X1 U5589 ( .A1(n6266), .A2(n4544), .ZN(n6157) );
  NAND2_X1 U5590 ( .A1(n6218), .A2(n6216), .ZN(n6269) );
  INV_X1 U5591 ( .A(n6142), .ZN(n4546) );
  NAND2_X1 U5592 ( .A1(n6269), .A2(n4546), .ZN(n4547) );
  INV_X1 U5593 ( .A(n5899), .ZN(n4548) );
  OAI21_X1 U5594 ( .B1(n6651), .B2(n6645), .A(n4548), .ZN(n4549) );
  INV_X1 U5595 ( .A(n4550), .ZN(n6108) );
  AND2_X1 U5596 ( .A1(n6269), .A2(n6108), .ZN(n4551) );
  AND2_X1 U5597 ( .A1(n6269), .A2(n6089), .ZN(n4552) );
  NOR2_X1 U5598 ( .A1(n6100), .A2(n4552), .ZN(n6078) );
  NAND2_X1 U5599 ( .A1(n6269), .A2(n4553), .ZN(n4554) );
  MUX2_X1 U5600 ( .A(n4555), .B(n6071), .S(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .Z(n4556) );
  INV_X1 U5601 ( .A(n4556), .ZN(n4557) );
  OAI211_X1 U5602 ( .C1(n4559), .C2(n6275), .A(n4558), .B(n4557), .ZN(U2987)
         );
  INV_X1 U5603 ( .A(n4560), .ZN(n4562) );
  NAND2_X1 U5604 ( .A1(n4564), .A2(EBX_REG_29__SCAN_IN), .ZN(n4565) );
  AND2_X1 U5605 ( .A1(n5856), .A2(n4853), .ZN(n4569) );
  NAND2_X1 U5606 ( .A1(n4584), .A2(n4569), .ZN(n4571) );
  AOI22_X1 U5607 ( .A1(n5838), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5850), .ZN(n4570) );
  NAND2_X1 U5608 ( .A1(n4571), .A2(n4570), .ZN(U2860) );
  INV_X1 U5609 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4574) );
  NAND2_X1 U5610 ( .A1(n6566), .A2(REIP_REG_30__SCAN_IN), .ZN(n6072) );
  OAI21_X1 U5611 ( .B1(n5981), .B2(n6918), .A(n6072), .ZN(n4576) );
  INV_X1 U5612 ( .A(n4577), .ZN(n4578) );
  NAND2_X1 U5613 ( .A1(n4578), .A2(n6571), .ZN(n4579) );
  OAI211_X1 U5614 ( .C1(n6076), .C2(n6372), .A(n4580), .B(n4579), .ZN(U2956)
         );
  NAND2_X1 U5615 ( .A1(n4499), .A2(n4673), .ZN(n4667) );
  INV_X1 U5616 ( .A(n4581), .ZN(n4582) );
  NAND2_X1 U5617 ( .A1(n4582), .A2(n6360), .ZN(n6362) );
  NAND3_X1 U5618 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_0__SCAN_IN), 
        .A3(n6844), .ZN(n6352) );
  NAND2_X1 U5619 ( .A1(n6362), .A2(n6352), .ZN(n4583) );
  OR3_X4 U5620 ( .A1(n6842), .A2(n6566), .A3(n4583), .ZN(n6433) );
  NAND2_X1 U5621 ( .A1(n6433), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U5622 ( .A1(n4584), .A2(n6411), .ZN(n4612) );
  NOR2_X1 U5623 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4586) );
  INV_X1 U5624 ( .A(n4586), .ZN(n5432) );
  NAND3_X1 U5625 ( .A1(n4800), .A2(EBX_REG_31__SCAN_IN), .A3(n5432), .ZN(n4585) );
  NAND3_X1 U5626 ( .A1(n4587), .A2(n3182), .A3(n4586), .ZN(n4588) );
  OR2_X2 U5627 ( .A1(n5458), .A2(n4588), .ZN(n6402) );
  INV_X1 U5628 ( .A(n6402), .ZN(n6389) );
  INV_X1 U5629 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5518) );
  INV_X1 U5630 ( .A(REIP_REG_7__SCAN_IN), .ZN(n4646) );
  INV_X1 U5631 ( .A(REIP_REG_5__SCAN_IN), .ZN(n5444) );
  NAND4_X1 U5632 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .A4(REIP_REG_2__SCAN_IN), .ZN(n5445) );
  NOR2_X1 U5633 ( .A1(n5444), .A2(n5445), .ZN(n5771) );
  NAND2_X1 U5634 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5771), .ZN(n5762) );
  NOR2_X1 U5635 ( .A1(n4646), .A2(n5762), .ZN(n5752) );
  NAND2_X1 U5636 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5752), .ZN(n6401) );
  NAND2_X1 U5637 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5430) );
  NOR2_X1 U5638 ( .A1(n6401), .A2(n5430), .ZN(n6387) );
  NAND2_X1 U5639 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6387), .ZN(n6388) );
  INV_X1 U5640 ( .A(n6388), .ZN(n4589) );
  OAI21_X1 U5641 ( .B1(n6402), .B2(n4589), .A(n6433), .ZN(n6394) );
  NAND2_X1 U5642 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5723) );
  AND2_X1 U5643 ( .A1(REIP_REG_14__SCAN_IN), .A2(n4600), .ZN(n4590) );
  NAND2_X1 U5644 ( .A1(n6402), .A2(n6433), .ZN(n6435) );
  NAND3_X1 U5645 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_17__SCAN_IN), .ZN(n4601) );
  NAND2_X1 U5646 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5646) );
  INV_X1 U5647 ( .A(n5646), .ZN(n4591) );
  NAND2_X1 U5648 ( .A1(n4591), .A2(REIP_REG_20__SCAN_IN), .ZN(n5602) );
  AND2_X1 U5649 ( .A1(n6435), .A2(n5602), .ZN(n4592) );
  NAND2_X1 U5650 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .ZN(
        n5564) );
  INV_X1 U5651 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5616) );
  OAI21_X1 U5652 ( .B1(n5564), .B2(n5616), .A(n6435), .ZN(n4593) );
  NAND3_X1 U5653 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4594) );
  NAND2_X1 U5654 ( .A1(n6389), .A2(n4594), .ZN(n4595) );
  AND2_X1 U5655 ( .A1(n5589), .A2(n4595), .ZN(n5538) );
  AND2_X1 U5656 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4597) );
  INV_X1 U5657 ( .A(n6435), .ZN(n4596) );
  AOI21_X1 U5658 ( .B1(n5538), .B2(n4597), .A(n4596), .ZN(n5532) );
  AOI21_X1 U5659 ( .B1(n6389), .B2(n5518), .A(n5532), .ZN(n5488) );
  OAI21_X1 U5660 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6402), .A(n5488), .ZN(n4608) );
  INV_X1 U5661 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4599) );
  OR2_X1 U5662 ( .A1(n4753), .A2(n5432), .ZN(n5362) );
  AND2_X1 U5663 ( .A1(n4698), .A2(n5362), .ZN(n5435) );
  NAND2_X1 U5664 ( .A1(n5435), .A2(EBX_REG_31__SCAN_IN), .ZN(n4598) );
  OAI22_X1 U5665 ( .A1(n6455), .A2(n4599), .B1(n5458), .B2(n4598), .ZN(n4607)
         );
  AND2_X1 U5666 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n4600) );
  NAND2_X1 U5667 ( .A1(n5740), .A2(n4600), .ZN(n5504) );
  INV_X1 U5668 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5503) );
  NOR2_X1 U5669 ( .A1(n5667), .A2(n5646), .ZN(n5629) );
  AND2_X1 U5670 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n4602) );
  INV_X1 U5671 ( .A(n5564), .ZN(n4603) );
  AND2_X1 U5672 ( .A1(REIP_REG_24__SCAN_IN), .A2(n4603), .ZN(n4604) );
  NAND2_X1 U5673 ( .A1(n5588), .A2(n4604), .ZN(n5568) );
  INV_X1 U5674 ( .A(REIP_REG_25__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U5675 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .ZN(
        n4605) );
  NOR2_X1 U5676 ( .A1(n5542), .A2(n4605), .ZN(n5533) );
  NAND3_X1 U5677 ( .A1(n5533), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .ZN(n5491) );
  INV_X1 U5678 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5487) );
  NOR3_X1 U5679 ( .A1(n5491), .A2(REIP_REG_31__SCAN_IN), .A3(n5487), .ZN(n4606) );
  AOI211_X1 U5680 ( .C1(REIP_REG_31__SCAN_IN), .C2(n4608), .A(n4607), .B(n4606), .ZN(n4609) );
  NAND2_X1 U5681 ( .A1(n4612), .A2(n4611), .ZN(U2796) );
  NAND2_X1 U5682 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6814) );
  INV_X1 U5683 ( .A(n6814), .ZN(n4613) );
  AOI21_X1 U5684 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n4613), .ZN(n4615) );
  NAND2_X1 U5685 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6810) );
  INV_X1 U5686 ( .A(n6810), .ZN(n4614) );
  NAND2_X1 U5687 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6817) );
  OAI211_X1 U5688 ( .C1(n4615), .C2(n4614), .A(n6817), .B(n4753), .ZN(U3182)
         );
  AOI211_X1 U5689 ( .C1(READY_N), .C2(n6345), .A(n6844), .B(n6360), .ZN(n4618)
         );
  NAND2_X1 U5690 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n4906) );
  INV_X1 U5691 ( .A(n4906), .ZN(n4616) );
  NAND2_X1 U5692 ( .A1(n4616), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5365) );
  AOI21_X1 U5693 ( .B1(n4618), .B2(n5365), .A(n4617), .ZN(n4619) );
  INV_X1 U5694 ( .A(n4619), .ZN(U3150) );
  INV_X1 U5695 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6041) );
  INV_X1 U5696 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7100) );
  NAND2_X1 U5697 ( .A1(n4621), .A2(n6825), .ZN(n4625) );
  INV_X1 U5698 ( .A(REIP_REG_11__SCAN_IN), .ZN(n4650) );
  OAI222_X1 U5699 ( .A1(n4639), .A2(n6041), .B1(n6825), .B2(n7100), .C1(n4625), 
        .C2(n4650), .ZN(U3193) );
  INV_X1 U5700 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6958) );
  INV_X1 U5701 ( .A(REIP_REG_31__SCAN_IN), .ZN(n4620) );
  OAI222_X1 U5702 ( .A1(n4639), .A2(n5487), .B1(n6825), .B2(n6958), .C1(n4620), 
        .C2(n4625), .ZN(U3213) );
  INV_X1 U5703 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n7075) );
  INV_X1 U5704 ( .A(REIP_REG_22__SCAN_IN), .ZN(n4627) );
  OAI222_X1 U5705 ( .A1(n4639), .A2(n5616), .B1(n6825), .B2(n7075), .C1(n4627), 
        .C2(n4625), .ZN(U3204) );
  INV_X1 U5706 ( .A(ADS_N_REG_SCAN_IN), .ZN(n4624) );
  NAND2_X1 U5707 ( .A1(n4621), .A2(STATE_REG_1__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U5708 ( .A1(n4622), .A2(STATE_REG_0__SCAN_IN), .ZN(n4623) );
  OAI21_X1 U5709 ( .B1(n6825), .B2(n4624), .A(n6809), .ZN(U2789) );
  INV_X1 U5710 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6436) );
  INV_X1 U5711 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n7113) );
  OAI222_X1 U5712 ( .A1(n4625), .A2(n5444), .B1(n4639), .B2(n6436), .C1(n6825), 
        .C2(n7113), .ZN(U3187) );
  INV_X1 U5713 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6910) );
  INV_X1 U5714 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6875) );
  OAI222_X1 U5715 ( .A1(n4625), .A2(n5503), .B1(n6825), .B2(n6910), .C1(n4639), 
        .C2(n6875), .ZN(U3196) );
  INV_X1 U5716 ( .A(n4625), .ZN(n4661) );
  AOI22_X1 U5717 ( .A1(n4661), .A2(REIP_REG_23__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_21__SCAN_IN), .ZN(n4626) );
  OAI21_X1 U5718 ( .B1(n4627), .B2(n4639), .A(n4626), .ZN(U3205) );
  INV_X1 U5719 ( .A(REIP_REG_23__SCAN_IN), .ZN(n4629) );
  AOI22_X1 U5720 ( .A1(n4661), .A2(REIP_REG_24__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_22__SCAN_IN), .ZN(n4628) );
  OAI21_X1 U5721 ( .B1(n4629), .B2(n4639), .A(n4628), .ZN(U3206) );
  INV_X1 U5722 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6467) );
  AOI22_X1 U5723 ( .A1(n4661), .A2(REIP_REG_4__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_2__SCAN_IN), .ZN(n4630) );
  OAI21_X1 U5724 ( .B1(n6467), .B2(n4639), .A(n4630), .ZN(U3186) );
  INV_X1 U5725 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5650) );
  AOI22_X1 U5726 ( .A1(n4661), .A2(REIP_REG_20__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_18__SCAN_IN), .ZN(n4631) );
  OAI21_X1 U5727 ( .B1(n5650), .B2(n4639), .A(n4631), .ZN(U3202) );
  INV_X1 U5728 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5964) );
  AOI22_X1 U5729 ( .A1(n4661), .A2(REIP_REG_19__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_17__SCAN_IN), .ZN(n4632) );
  OAI21_X1 U5730 ( .B1(n5964), .B2(n4639), .A(n4632), .ZN(U3201) );
  AOI22_X1 U5731 ( .A1(n4661), .A2(REIP_REG_26__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_24__SCAN_IN), .ZN(n4633) );
  OAI21_X1 U5732 ( .B1(n4634), .B2(n4639), .A(n4633), .ZN(U3208) );
  INV_X1 U5733 ( .A(REIP_REG_26__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5734 ( .A1(n4661), .A2(REIP_REG_27__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_25__SCAN_IN), .ZN(n4635) );
  OAI21_X1 U5735 ( .B1(n4636), .B2(n4639), .A(n4635), .ZN(U3209) );
  INV_X1 U5736 ( .A(REIP_REG_20__SCAN_IN), .ZN(n4638) );
  AOI22_X1 U5737 ( .A1(n4661), .A2(REIP_REG_21__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_19__SCAN_IN), .ZN(n4637) );
  OAI21_X1 U5738 ( .B1(n4638), .B2(n4639), .A(n4637), .ZN(U3203) );
  AOI22_X1 U5739 ( .A1(n4661), .A2(REIP_REG_30__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_28__SCAN_IN), .ZN(n4640) );
  OAI21_X1 U5740 ( .B1(n5518), .B2(n4639), .A(n4640), .ZN(U3212) );
  INV_X1 U5741 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6926) );
  AOI22_X1 U5742 ( .A1(n4661), .A2(REIP_REG_2__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_0__SCAN_IN), .ZN(n4641) );
  OAI21_X1 U5743 ( .B1(n6926), .B2(n4639), .A(n4641), .ZN(U3184) );
  INV_X1 U5744 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6576) );
  AOI22_X1 U5745 ( .A1(n4661), .A2(REIP_REG_3__SCAN_IN), .B1(n6849), .B2(
        ADDRESS_REG_1__SCAN_IN), .ZN(n4642) );
  OAI21_X1 U5746 ( .B1(n6576), .B2(n4639), .A(n4642), .ZN(U3185) );
  AOI22_X1 U5747 ( .A1(n4661), .A2(REIP_REG_6__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_4__SCAN_IN), .ZN(n4643) );
  OAI21_X1 U5748 ( .B1(n5444), .B2(n4639), .A(n4643), .ZN(U3188) );
  INV_X1 U5749 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6556) );
  AOI22_X1 U5750 ( .A1(n4661), .A2(REIP_REG_7__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_5__SCAN_IN), .ZN(n4644) );
  OAI21_X1 U5751 ( .B1(n6556), .B2(n4639), .A(n4644), .ZN(U3189) );
  AOI22_X1 U5752 ( .A1(n4661), .A2(REIP_REG_8__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_6__SCAN_IN), .ZN(n4645) );
  OAI21_X1 U5753 ( .B1(n4646), .B2(n4639), .A(n4645), .ZN(U3190) );
  INV_X1 U5754 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5755) );
  AOI22_X1 U5755 ( .A1(n4661), .A2(REIP_REG_9__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_7__SCAN_IN), .ZN(n4647) );
  OAI21_X1 U5756 ( .B1(n5755), .B2(n4639), .A(n4647), .ZN(U3191) );
  INV_X1 U5757 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6404) );
  AOI22_X1 U5758 ( .A1(n4661), .A2(REIP_REG_10__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_8__SCAN_IN), .ZN(n4648) );
  OAI21_X1 U5759 ( .B1(n6404), .B2(n4639), .A(n4648), .ZN(U3192) );
  AOI22_X1 U5760 ( .A1(n4661), .A2(REIP_REG_12__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_10__SCAN_IN), .ZN(n4649) );
  OAI21_X1 U5761 ( .B1(n4650), .B2(n4639), .A(n4649), .ZN(U3194) );
  INV_X1 U5762 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5739) );
  AOI22_X1 U5763 ( .A1(n4661), .A2(REIP_REG_13__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_11__SCAN_IN), .ZN(n4651) );
  OAI21_X1 U5764 ( .B1(n5739), .B2(n4639), .A(n4651), .ZN(U3195) );
  AOI22_X1 U5765 ( .A1(n4661), .A2(REIP_REG_15__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_13__SCAN_IN), .ZN(n4652) );
  OAI21_X1 U5766 ( .B1(n5503), .B2(n4639), .A(n4652), .ZN(U3197) );
  INV_X1 U5767 ( .A(REIP_REG_15__SCAN_IN), .ZN(n4654) );
  AOI22_X1 U5768 ( .A1(n4661), .A2(REIP_REG_16__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_14__SCAN_IN), .ZN(n4653) );
  OAI21_X1 U5769 ( .B1(n4654), .B2(n4639), .A(n4653), .ZN(U3198) );
  INV_X1 U5770 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5987) );
  AOI22_X1 U5771 ( .A1(n4661), .A2(REIP_REG_17__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_15__SCAN_IN), .ZN(n4655) );
  OAI21_X1 U5772 ( .B1(n5987), .B2(n4639), .A(n4655), .ZN(U3199) );
  INV_X1 U5773 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5677) );
  AOI22_X1 U5774 ( .A1(n4661), .A2(REIP_REG_18__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_16__SCAN_IN), .ZN(n4656) );
  OAI21_X1 U5775 ( .B1(n5677), .B2(n4639), .A(n4656), .ZN(U3200) );
  INV_X1 U5776 ( .A(REIP_REG_24__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U5777 ( .A1(n4661), .A2(REIP_REG_25__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_23__SCAN_IN), .ZN(n4657) );
  OAI21_X1 U5778 ( .B1(n4658), .B2(n4639), .A(n4657), .ZN(U3207) );
  INV_X1 U5779 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5861) );
  AOI22_X1 U5780 ( .A1(n4661), .A2(REIP_REG_29__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_27__SCAN_IN), .ZN(n4659) );
  OAI21_X1 U5781 ( .B1(n5861), .B2(n4639), .A(n4659), .ZN(U3211) );
  INV_X1 U5782 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5543) );
  AOI22_X1 U5783 ( .A1(n4661), .A2(REIP_REG_28__SCAN_IN), .B1(n4660), .B2(
        ADDRESS_REG_26__SCAN_IN), .ZN(n4662) );
  OAI21_X1 U5784 ( .B1(n5543), .B2(n4639), .A(n4662), .ZN(U3210) );
  NOR2_X1 U5785 ( .A1(n6722), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5509) );
  INV_X1 U5786 ( .A(n4663), .ZN(n4697) );
  AOI211_X1 U5787 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4664), .A(n5509), .B(
        n4697), .ZN(n4665) );
  INV_X1 U5788 ( .A(n4665), .ZN(U2788) );
  OR2_X1 U5789 ( .A1(n4709), .A2(n4666), .ZN(n4669) );
  NAND2_X1 U5790 ( .A1(n4667), .A2(n4325), .ZN(n4668) );
  NAND2_X1 U5791 ( .A1(n4669), .A2(n4668), .ZN(n6366) );
  NAND3_X1 U5792 ( .A1(n4360), .A2(n4753), .A3(n5510), .ZN(n4670) );
  AND2_X1 U5793 ( .A1(n4670), .A2(n6838), .ZN(n6843) );
  AND2_X1 U5794 ( .A1(n5353), .A2(n6355), .ZN(n6374) );
  INV_X1 U5795 ( .A(MORE_REG_SCAN_IN), .ZN(n4678) );
  NOR2_X1 U5796 ( .A1(n4671), .A2(n3168), .ZN(n4672) );
  MUX2_X1 U5797 ( .A(n4672), .B(n4731), .S(n4709), .Z(n4676) );
  INV_X1 U5798 ( .A(n4673), .ZN(n4674) );
  NAND2_X1 U5799 ( .A1(n4499), .A2(n4674), .ZN(n4675) );
  NAND2_X1 U5800 ( .A1(n4676), .A2(n4675), .ZN(n5355) );
  NAND2_X1 U5801 ( .A1(n6374), .A2(n5355), .ZN(n4677) );
  OAI21_X1 U5802 ( .B1(n6374), .B2(n4678), .A(n4677), .ZN(U3471) );
  INV_X1 U5803 ( .A(n4731), .ZN(n4682) );
  AND2_X1 U5804 ( .A1(n4360), .A2(n4753), .ZN(n4679) );
  OAI22_X1 U5805 ( .A1(n4878), .A2(n4753), .B1(n4679), .B2(n4487), .ZN(n4680)
         );
  AND2_X1 U5806 ( .A1(n4680), .A2(n6838), .ZN(n4681) );
  MUX2_X1 U5807 ( .A(n4682), .B(n4681), .S(n4709), .Z(n4688) );
  INV_X1 U5808 ( .A(n4683), .ZN(n4684) );
  NAND2_X1 U5809 ( .A1(n4685), .A2(n4684), .ZN(n4686) );
  INV_X1 U5810 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6373) );
  NOR2_X1 U5811 ( .A1(n5365), .A2(n6373), .ZN(n4689) );
  AOI21_X1 U5812 ( .B1(n5335), .B2(n6355), .A(n4689), .ZN(n4694) );
  NAND2_X1 U5813 ( .A1(n6938), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4690) );
  NAND2_X1 U5814 ( .A1(n4694), .A2(n4690), .ZN(n6299) );
  INV_X1 U5815 ( .A(n4691), .ZN(n5017) );
  OR2_X1 U5816 ( .A1(n4692), .A2(n5017), .ZN(n4693) );
  XNOR2_X1 U5817 ( .A(n4693), .B(n4696), .ZN(n6442) );
  INV_X1 U5818 ( .A(n6357), .ZN(n6297) );
  OR4_X1 U5819 ( .A1(n4694), .A2(n6442), .A3(n6297), .A4(n4312), .ZN(n4695) );
  OAI21_X1 U5820 ( .B1(n6299), .B2(n4696), .A(n4695), .ZN(U3455) );
  INV_X1 U5821 ( .A(DATAI_14_), .ZN(n7059) );
  OAI21_X1 U5822 ( .B1(n4698), .B2(n6838), .A(n4697), .ZN(n6549) );
  AOI22_X1 U5823 ( .A1(n6549), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6552), .ZN(n4699) );
  OAI21_X1 U5824 ( .B1(n7059), .B2(n6516), .A(n4699), .ZN(U2953) );
  INV_X1 U5825 ( .A(DATAI_11_), .ZN(n7157) );
  AOI22_X1 U5826 ( .A1(n6549), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n6552), .ZN(n4700) );
  OAI21_X1 U5827 ( .B1(n7157), .B2(n6516), .A(n4700), .ZN(U2950) );
  INV_X1 U5828 ( .A(DATAI_15_), .ZN(n7024) );
  AOI22_X1 U5829 ( .A1(n6549), .A2(LWORD_REG_15__SCAN_IN), .B1(
        EAX_REG_15__SCAN_IN), .B2(n6552), .ZN(n4701) );
  OAI21_X1 U5830 ( .B1(n7024), .B2(n6516), .A(n4701), .ZN(U2954) );
  INV_X1 U5831 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n7081) );
  INV_X1 U5832 ( .A(DATAI_2_), .ZN(n4702) );
  NOR2_X1 U5833 ( .A1(n6516), .A2(n4702), .ZN(n6507) );
  INV_X1 U5834 ( .A(n6507), .ZN(n4704) );
  NAND2_X1 U5835 ( .A1(n6552), .A2(EAX_REG_2__SCAN_IN), .ZN(n4703) );
  OAI211_X1 U5836 ( .C1(n6503), .C2(n7081), .A(n4704), .B(n4703), .ZN(U2941)
         );
  INV_X1 U5837 ( .A(EAX_REG_7__SCAN_IN), .ZN(n5857) );
  INV_X1 U5838 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n4706) );
  INV_X1 U5839 ( .A(DATAI_7_), .ZN(n4705) );
  OAI222_X1 U5840 ( .A1(n6545), .A2(n5857), .B1(n4706), .B2(n6503), .C1(n6516), 
        .C2(n4705), .ZN(U2946) );
  INV_X1 U5841 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n7043) );
  INV_X1 U5842 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4707) );
  OAI222_X1 U5843 ( .A1(n7059), .A2(n6516), .B1(n7043), .B2(n6503), .C1(n4707), 
        .C2(n6545), .ZN(U2938) );
  INV_X1 U5844 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n4708) );
  OAI222_X1 U5845 ( .A1(n6545), .A2(n6494), .B1(n4708), .B2(n6503), .C1(n6516), 
        .C2(n5300), .ZN(U2945) );
  OAI21_X1 U5846 ( .B1(n4749), .B2(n6349), .A(n6299), .ZN(n4751) );
  INV_X1 U5847 ( .A(n4751), .ZN(n4726) );
  INV_X1 U5848 ( .A(n6299), .ZN(n4741) );
  INV_X1 U5849 ( .A(n4713), .ZN(n4714) );
  NAND2_X1 U5850 ( .A1(n4714), .A2(n3139), .ZN(n4873) );
  NAND2_X1 U5851 ( .A1(n4712), .A2(n4873), .ZN(n4719) );
  INV_X1 U5852 ( .A(n4715), .ZN(n4885) );
  INV_X1 U5853 ( .A(n3309), .ZN(n4898) );
  NAND3_X1 U5854 ( .A1(n4745), .A2(n4885), .A3(n4898), .ZN(n4716) );
  OAI21_X1 U5855 ( .B1(n4878), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4716), 
        .ZN(n4717) );
  INV_X1 U5856 ( .A(n4717), .ZN(n4718) );
  NAND2_X1 U5857 ( .A1(n4719), .A2(n4718), .ZN(n5334) );
  INV_X1 U5858 ( .A(n4720), .ZN(n4723) );
  AOI22_X1 U5859 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4721), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n7101), .ZN(n4737) );
  NAND3_X1 U5860 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n4737), .A3(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4722) );
  OAI21_X1 U5861 ( .B1(n6349), .B2(n4723), .A(n4722), .ZN(n4724) );
  AOI21_X1 U5862 ( .B1(n6357), .B2(n5334), .A(n4724), .ZN(n4725) );
  OAI22_X1 U5863 ( .A1(n4726), .A2(n4710), .B1(n4741), .B2(n4725), .ZN(U3460)
         );
  INV_X1 U5864 ( .A(n6349), .ZN(n4727) );
  AOI21_X1 U5865 ( .B1(n4727), .B2(n4885), .A(n4741), .ZN(n4743) );
  NAND2_X1 U5866 ( .A1(n4728), .A2(n4873), .ZN(n4736) );
  INV_X1 U5867 ( .A(n4729), .ZN(n4730) );
  NAND2_X1 U5868 ( .A1(n4731), .A2(n4730), .ZN(n4875) );
  XNOR2_X1 U5869 ( .A(n4715), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4734)
         );
  XNOR2_X1 U5870 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4732) );
  OAI22_X1 U5871 ( .A1(n4878), .A2(n4732), .B1(n4887), .B2(n4734), .ZN(n4733)
         );
  AOI21_X1 U5872 ( .B1(n4875), .B2(n4734), .A(n4733), .ZN(n4735) );
  NAND2_X1 U5873 ( .A1(n4736), .A2(n4735), .ZN(n4892) );
  INV_X1 U5874 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4821) );
  NOR3_X1 U5875 ( .A1(n6359), .A2(n4821), .A3(n4737), .ZN(n4739) );
  NOR3_X1 U5876 ( .A1(n6349), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4885), 
        .ZN(n4738) );
  AOI211_X1 U5877 ( .C1(n6357), .C2(n4892), .A(n4739), .B(n4738), .ZN(n4740)
         );
  OAI22_X1 U5878 ( .A1(n4743), .A2(n4742), .B1(n4741), .B2(n4740), .ZN(U3459)
         );
  OR2_X1 U5879 ( .A1(n4878), .A2(n4744), .ZN(n5330) );
  NAND2_X1 U5880 ( .A1(n3845), .A2(n4873), .ZN(n4747) );
  NAND2_X1 U5881 ( .A1(n4745), .A2(n4744), .ZN(n4746) );
  NAND2_X1 U5882 ( .A1(n4747), .A2(n4746), .ZN(n5332) );
  INV_X1 U5883 ( .A(n5332), .ZN(n4748) );
  OAI22_X1 U5884 ( .A1(n4748), .A2(n6297), .B1(n6359), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4750) );
  OAI22_X1 U5885 ( .A1(n4751), .A2(n4750), .B1(n4749), .B2(n6299), .ZN(n4752)
         );
  OAI21_X1 U5886 ( .B1(n5330), .B2(n6297), .A(n4752), .ZN(U3461) );
  NOR2_X2 U5887 ( .A1(n6500), .A2(n5456), .ZN(n6482) );
  INV_X2 U5888 ( .A(n4770), .ZN(n6839) );
  AOI222_X1 U5889 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6482), .B1(n6497), .B2(
        DATAO_REG_26__SCAN_IN), .C1(n6839), .C2(UWORD_REG_10__SCAN_IN), .ZN(
        n4756) );
  INV_X1 U5890 ( .A(n4756), .ZN(U2897) );
  INV_X1 U5891 ( .A(n6500), .ZN(n6490) );
  AOI222_X1 U5892 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6839), .B1(n6497), .B2(
        DATAO_REG_11__SCAN_IN), .C1(EAX_REG_11__SCAN_IN), .C2(n6490), .ZN(
        n4757) );
  INV_X1 U5893 ( .A(n4757), .ZN(U2912) );
  AOI222_X1 U5894 ( .A1(EAX_REG_23__SCAN_IN), .A2(n6482), .B1(n6497), .B2(
        DATAO_REG_23__SCAN_IN), .C1(n6839), .C2(UWORD_REG_7__SCAN_IN), .ZN(
        n4758) );
  INV_X1 U5895 ( .A(n4758), .ZN(U2900) );
  AOI222_X1 U5896 ( .A1(EAX_REG_21__SCAN_IN), .A2(n6482), .B1(n6497), .B2(
        DATAO_REG_21__SCAN_IN), .C1(n6839), .C2(UWORD_REG_5__SCAN_IN), .ZN(
        n4759) );
  INV_X1 U5897 ( .A(n4759), .ZN(U2902) );
  AOI222_X1 U5898 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6482), .B1(n6497), .B2(
        DATAO_REG_25__SCAN_IN), .C1(n6839), .C2(UWORD_REG_9__SCAN_IN), .ZN(
        n4760) );
  INV_X1 U5899 ( .A(n4760), .ZN(U2898) );
  AOI222_X1 U5900 ( .A1(EAX_REG_16__SCAN_IN), .A2(n6482), .B1(n6497), .B2(
        DATAO_REG_16__SCAN_IN), .C1(n6839), .C2(UWORD_REG_0__SCAN_IN), .ZN(
        n4761) );
  INV_X1 U5901 ( .A(n4761), .ZN(U2907) );
  AOI222_X1 U5902 ( .A1(EAX_REG_22__SCAN_IN), .A2(n6482), .B1(n6497), .B2(
        DATAO_REG_22__SCAN_IN), .C1(n6839), .C2(UWORD_REG_6__SCAN_IN), .ZN(
        n4762) );
  INV_X1 U5903 ( .A(n4762), .ZN(U2901) );
  INV_X1 U5904 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n7026) );
  OAI22_X1 U5905 ( .A1(n6503), .A2(n7026), .B1(n5854), .B2(n6545), .ZN(n4763)
         );
  INV_X1 U5906 ( .A(DATAI_8_), .ZN(n5853) );
  NOR2_X1 U5907 ( .A1(n6516), .A2(n5853), .ZN(n6520) );
  OR2_X1 U5908 ( .A1(n4763), .A2(n6520), .ZN(U2947) );
  INV_X1 U5909 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6947) );
  OAI22_X1 U5910 ( .A1(n6503), .A2(n6947), .B1(n5847), .B2(n6545), .ZN(n4764)
         );
  INV_X1 U5911 ( .A(DATAI_12_), .ZN(n5849) );
  NOR2_X1 U5912 ( .A1(n6516), .A2(n5849), .ZN(n6528) );
  OR2_X1 U5913 ( .A1(n4764), .A2(n6528), .ZN(U2951) );
  INV_X1 U5914 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n7023) );
  INV_X1 U5915 ( .A(n6482), .ZN(n4769) );
  INV_X1 U5916 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6513) );
  INV_X1 U5917 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6944) );
  OAI222_X1 U5918 ( .A1(n6492), .A2(n7023), .B1(n4769), .B2(n6513), .C1(n4770), 
        .C2(n6944), .ZN(U2903) );
  INV_X1 U5919 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4765) );
  OAI222_X1 U5920 ( .A1(n4765), .A2(n6492), .B1(n4770), .B2(n7026), .C1(n5854), 
        .C2(n6500), .ZN(U2915) );
  INV_X1 U5921 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4766) );
  OAI222_X1 U5922 ( .A1(n4766), .A2(n6492), .B1(n4770), .B2(n6947), .C1(n5847), 
        .C2(n6500), .ZN(U2911) );
  INV_X1 U5923 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4768) );
  INV_X1 U5924 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6878) );
  INV_X1 U5925 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4767) );
  OAI222_X1 U5926 ( .A1(n4768), .A2(n6492), .B1(n4770), .B2(n6878), .C1(n4767), 
        .C2(n6500), .ZN(U2909) );
  INV_X1 U5927 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6939) );
  INV_X1 U5928 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n7134) );
  OAI222_X1 U5929 ( .A1(n4769), .A2(n6509), .B1(n6492), .B2(n6939), .C1(n4770), 
        .C2(n7134), .ZN(U2905) );
  INV_X1 U5930 ( .A(EAX_REG_2__SCAN_IN), .ZN(n4771) );
  INV_X1 U5931 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n6881) );
  OAI222_X1 U5932 ( .A1(n6500), .A2(n4771), .B1(n6492), .B2(n6881), .C1(n4770), 
        .C2(n7081), .ZN(U2921) );
  XNOR2_X1 U5933 ( .A(n4773), .B(n4772), .ZN(n5471) );
  XOR2_X1 U5934 ( .A(n4774), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n4792) );
  NAND2_X1 U5935 ( .A1(n4792), .A2(n3784), .ZN(n4778) );
  OR2_X1 U5936 ( .A1(n6578), .A2(n4775), .ZN(n4776) );
  AOI22_X1 U5937 ( .A1(n4776), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6566), 
        .B2(REIP_REG_0__SCAN_IN), .ZN(n4777) );
  OAI211_X1 U5938 ( .C1(n5471), .C2(n6054), .A(n4778), .B(n4777), .ZN(U2986)
         );
  XNOR2_X1 U5939 ( .A(n4780), .B(n4779), .ZN(n4827) );
  NOR2_X1 U5940 ( .A1(n4782), .A2(n4781), .ZN(n4783) );
  INV_X1 U5941 ( .A(n5465), .ZN(n4788) );
  INV_X1 U5942 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5943 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6566), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4786) );
  OAI21_X1 U5944 ( .B1(n6586), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4786), 
        .ZN(n4787) );
  AOI21_X1 U5945 ( .B1(n4788), .B2(n6571), .A(n4787), .ZN(n4789) );
  OAI21_X1 U5946 ( .B1(n4827), .B2(n6372), .A(n4789), .ZN(U2985) );
  OAI21_X1 U5947 ( .B1(n4791), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4790), 
        .ZN(n5466) );
  OAI222_X1 U5948 ( .A1(n5466), .A2(n5802), .B1(n6474), .B2(n5471), .C1(n7050), 
        .C2(n6481), .ZN(U2859) );
  INV_X1 U5949 ( .A(n4792), .ZN(n4799) );
  INV_X1 U5950 ( .A(n5466), .ZN(n4797) );
  INV_X1 U5951 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6928) );
  OAI21_X1 U5952 ( .B1(n6577), .B2(n6928), .A(n4793), .ZN(n4796) );
  AOI21_X1 U5953 ( .B1(n6218), .B2(n4794), .A(n4821), .ZN(n4795) );
  AOI211_X1 U5954 ( .C1(n4797), .C2(n6644), .A(n4796), .B(n4795), .ZN(n4798)
         );
  OAI21_X1 U5955 ( .B1(n4799), .B2(n6275), .A(n4798), .ZN(U3018) );
  OR2_X1 U5956 ( .A1(n4801), .A2(n4800), .ZN(n4803) );
  AND2_X1 U5957 ( .A1(n4803), .A2(n4802), .ZN(n5454) );
  INV_X1 U5958 ( .A(n5454), .ZN(n4825) );
  AOI22_X1 U5959 ( .A1(n6478), .A2(n4825), .B1(n4564), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4804) );
  OAI21_X1 U5960 ( .B1(n5465), .B2(n6474), .A(n4804), .ZN(U2858) );
  INV_X1 U5961 ( .A(n4805), .ZN(n4806) );
  AOI22_X1 U5962 ( .A1(n5851), .A2(DATAI_1_), .B1(n5850), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n4807) );
  OAI21_X1 U5963 ( .B1(n5465), .B2(n5859), .A(n4807), .ZN(U2890) );
  AOI22_X1 U5964 ( .A1(n5851), .A2(DATAI_0_), .B1(n5850), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n4808) );
  OAI21_X1 U5965 ( .B1(n5471), .B2(n5859), .A(n4808), .ZN(U2891) );
  AOI222_X1 U5966 ( .A1(n6497), .A2(DATAO_REG_1__SCAN_IN), .B1(n6490), .B2(
        EAX_REG_1__SCAN_IN), .C1(n6839), .C2(LWORD_REG_1__SCAN_IN), .ZN(n4809)
         );
  INV_X1 U5967 ( .A(n4809), .ZN(U2922) );
  AOI222_X1 U5968 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6839), .B1(n6497), .B2(
        DATAO_REG_30__SCAN_IN), .C1(EAX_REG_30__SCAN_IN), .C2(n6482), .ZN(
        n4810) );
  INV_X1 U5969 ( .A(n4810), .ZN(U2893) );
  AOI222_X1 U5970 ( .A1(EAX_REG_17__SCAN_IN), .A2(n6482), .B1(n6497), .B2(
        DATAO_REG_17__SCAN_IN), .C1(n6839), .C2(UWORD_REG_1__SCAN_IN), .ZN(
        n4811) );
  INV_X1 U5971 ( .A(n4811), .ZN(U2906) );
  AOI222_X1 U5972 ( .A1(EAX_REG_19__SCAN_IN), .A2(n6482), .B1(n6497), .B2(
        DATAO_REG_19__SCAN_IN), .C1(n6839), .C2(UWORD_REG_3__SCAN_IN), .ZN(
        n4812) );
  INV_X1 U5973 ( .A(n4812), .ZN(U2904) );
  AOI222_X1 U5974 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6482), .B1(n6497), .B2(
        DATAO_REG_24__SCAN_IN), .C1(n6839), .C2(UWORD_REG_8__SCAN_IN), .ZN(
        n4813) );
  INV_X1 U5975 ( .A(n4813), .ZN(U2899) );
  AOI222_X1 U5976 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6482), .B1(n6497), .B2(
        DATAO_REG_27__SCAN_IN), .C1(n6839), .C2(UWORD_REG_11__SCAN_IN), .ZN(
        n4814) );
  INV_X1 U5977 ( .A(n4814), .ZN(U2896) );
  AOI222_X1 U5978 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6482), .B1(n6497), .B2(
        DATAO_REG_28__SCAN_IN), .C1(n6839), .C2(UWORD_REG_12__SCAN_IN), .ZN(
        n4815) );
  INV_X1 U5979 ( .A(n4815), .ZN(U2895) );
  INV_X1 U5980 ( .A(n4816), .ZN(n4819) );
  AOI21_X1 U5981 ( .B1(n4819), .B2(n4818), .A(n3858), .ZN(n6582) );
  INV_X1 U5982 ( .A(n6582), .ZN(n5485) );
  AOI22_X1 U5983 ( .A1(n5851), .A2(DATAI_2_), .B1(n5850), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4820) );
  OAI21_X1 U5984 ( .B1(n5485), .B2(n5859), .A(n4820), .ZN(U2889) );
  NOR2_X1 U5985 ( .A1(n6577), .A2(n6926), .ZN(n4824) );
  OAI21_X1 U5986 ( .B1(n6216), .B2(n4821), .A(n6218), .ZN(n4822) );
  MUX2_X1 U5987 ( .A(n4822), .B(n5368), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4823) );
  AOI211_X1 U5988 ( .C1(n6644), .C2(n4825), .A(n4824), .B(n4823), .ZN(n4826)
         );
  OAI21_X1 U5989 ( .B1(n4827), .B2(n6275), .A(n4826), .ZN(U3017) );
  INV_X1 U5990 ( .A(n4913), .ZN(n4981) );
  NOR2_X1 U5991 ( .A1(n6278), .A2(n4981), .ZN(n4829) );
  NAND2_X1 U5992 ( .A1(n6283), .A2(n4829), .ZN(n4836) );
  NAND2_X1 U5993 ( .A1(n6571), .A2(DATAI_25_), .ZN(n6776) );
  NOR2_X1 U5994 ( .A1(n5018), .A2(n5345), .ZN(n5143) );
  NOR2_X1 U5995 ( .A1(n4836), .A2(n6371), .ZN(n6288) );
  NAND2_X1 U5996 ( .A1(n4832), .A2(n3845), .ZN(n5255) );
  INV_X1 U5997 ( .A(n4712), .ZN(n6280) );
  INV_X1 U5998 ( .A(n5149), .ZN(n5141) );
  NAND2_X1 U5999 ( .A1(n5143), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4867) );
  OAI21_X1 U6000 ( .B1(n5255), .B2(n5141), .A(n4867), .ZN(n4839) );
  INV_X1 U6001 ( .A(n6844), .ZN(n6348) );
  NAND2_X1 U6002 ( .A1(n4906), .A2(n6348), .ZN(n4833) );
  NAND2_X1 U6003 ( .A1(n4865), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4842)
         );
  NAND2_X1 U6004 ( .A1(n6571), .A2(DATAI_17_), .ZN(n6771) );
  INV_X1 U6005 ( .A(n6771), .ZN(n6675) );
  NAND2_X1 U6006 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4837) );
  NOR2_X1 U6007 ( .A1(n5018), .A2(n4837), .ZN(n4838) );
  AOI21_X1 U6008 ( .B1(n4839), .B2(n6304), .A(n4838), .ZN(n4868) );
  AND2_X1 U6009 ( .A1(n5306), .A2(DATAI_1_), .ZN(n6773) );
  OAI22_X1 U6010 ( .A1(n4868), .A2(n6678), .B1(n6770), .B2(n4867), .ZN(n4840)
         );
  AOI21_X1 U6011 ( .B1(n5383), .B2(n6675), .A(n4840), .ZN(n4841) );
  OAI211_X1 U6012 ( .C1(n4872), .C2(n6776), .A(n4842), .B(n4841), .ZN(U3125)
         );
  NAND2_X1 U6013 ( .A1(n6571), .A2(DATAI_26_), .ZN(n6783) );
  NAND2_X1 U6014 ( .A1(n4865), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4846)
         );
  NAND2_X1 U6015 ( .A1(n6571), .A2(DATAI_18_), .ZN(n6778) );
  INV_X1 U6016 ( .A(n6778), .ZN(n6680) );
  AND2_X1 U6017 ( .A1(n5306), .A2(DATAI_2_), .ZN(n6780) );
  OAI22_X1 U6018 ( .A1(n4868), .A2(n6683), .B1(n6777), .B2(n4867), .ZN(n4844)
         );
  AOI21_X1 U6019 ( .B1(n5383), .B2(n6680), .A(n4844), .ZN(n4845) );
  OAI211_X1 U6020 ( .C1(n4872), .C2(n6783), .A(n4846), .B(n4845), .ZN(U3126)
         );
  NAND2_X1 U6021 ( .A1(n4865), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4849)
         );
  NAND2_X1 U6022 ( .A1(n6571), .A2(DATAI_20_), .ZN(n6852) );
  INV_X1 U6023 ( .A(n6852), .ZN(n6690) );
  OAI22_X1 U6024 ( .A1(n4868), .A2(n6860), .B1(n6850), .B2(n4867), .ZN(n4847)
         );
  AOI21_X1 U6025 ( .B1(n5383), .B2(n6690), .A(n4847), .ZN(n4848) );
  OAI211_X1 U6026 ( .C1(n4872), .C2(n6329), .A(n4849), .B(n4848), .ZN(U3128)
         );
  AND2_X1 U6027 ( .A1(n6571), .A2(DATAI_24_), .ZN(n6731) );
  INV_X1 U6028 ( .A(n6731), .ZN(n6316) );
  NAND2_X1 U6029 ( .A1(n4865), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4852)
         );
  NAND2_X1 U6030 ( .A1(n6571), .A2(DATAI_16_), .ZN(n6734) );
  INV_X1 U6031 ( .A(n6734), .ZN(n6663) );
  OR2_X1 U6032 ( .A1(n4866), .A2(n5456), .ZN(n6661) );
  OAI22_X1 U6033 ( .A1(n4868), .A2(n6717), .B1(n6661), .B2(n4867), .ZN(n4850)
         );
  AOI21_X1 U6034 ( .B1(n5383), .B2(n6663), .A(n4850), .ZN(n4851) );
  OAI211_X1 U6035 ( .C1(n4872), .C2(n6316), .A(n4852), .B(n4851), .ZN(U3124)
         );
  AND2_X1 U6036 ( .A1(n6571), .A2(DATAI_31_), .ZN(n6764) );
  NAND2_X1 U6037 ( .A1(n4865), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4856)
         );
  NAND2_X1 U6038 ( .A1(n6571), .A2(DATAI_23_), .ZN(n6769) );
  INV_X1 U6039 ( .A(n6769), .ZN(n6706) );
  OAI22_X1 U6040 ( .A1(n4868), .A2(n6758), .B1(n6704), .B2(n4867), .ZN(n4854)
         );
  AOI21_X1 U6041 ( .B1(n5383), .B2(n6706), .A(n4854), .ZN(n4855) );
  OAI211_X1 U6042 ( .C1(n4872), .C2(n6343), .A(n4856), .B(n4855), .ZN(U3131)
         );
  NAND2_X1 U6043 ( .A1(n6571), .A2(DATAI_27_), .ZN(n6790) );
  NAND2_X1 U6044 ( .A1(n4865), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4860)
         );
  NAND2_X1 U6045 ( .A1(n6571), .A2(DATAI_19_), .ZN(n6785) );
  AND2_X1 U6046 ( .A1(n5306), .A2(DATAI_3_), .ZN(n6787) );
  OR2_X1 U6047 ( .A1(n4866), .A2(n4857), .ZN(n6784) );
  OAI22_X1 U6048 ( .A1(n4868), .A2(n6688), .B1(n6784), .B2(n4867), .ZN(n4858)
         );
  AOI21_X1 U6049 ( .B1(n5383), .B2(n6685), .A(n4858), .ZN(n4859) );
  OAI211_X1 U6050 ( .C1(n4872), .C2(n6790), .A(n4860), .B(n4859), .ZN(U3127)
         );
  NAND2_X1 U6051 ( .A1(n6571), .A2(DATAI_29_), .ZN(n6797) );
  NAND2_X1 U6052 ( .A1(n4865), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4864)
         );
  NAND2_X1 U6053 ( .A1(n6571), .A2(DATAI_21_), .ZN(n6792) );
  INV_X1 U6054 ( .A(n6792), .ZN(n6694) );
  AND2_X1 U6055 ( .A1(n5306), .A2(DATAI_5_), .ZN(n6794) );
  OAI22_X1 U6056 ( .A1(n4868), .A2(n6697), .B1(n6791), .B2(n4867), .ZN(n4862)
         );
  AOI21_X1 U6057 ( .B1(n5383), .B2(n6694), .A(n4862), .ZN(n4863) );
  OAI211_X1 U6058 ( .C1(n4872), .C2(n6797), .A(n4864), .B(n4863), .ZN(U3129)
         );
  NAND2_X1 U6059 ( .A1(n6571), .A2(DATAI_30_), .ZN(n6808) );
  NAND2_X1 U6060 ( .A1(n4865), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4871)
         );
  NAND2_X1 U6061 ( .A1(n6571), .A2(DATAI_22_), .ZN(n6800) );
  AND2_X1 U6062 ( .A1(n5306), .A2(DATAI_6_), .ZN(n6804) );
  OR2_X1 U6063 ( .A1(n4866), .A2(n3436), .ZN(n6799) );
  OAI22_X1 U6064 ( .A1(n4868), .A2(n6702), .B1(n6799), .B2(n4867), .ZN(n4869)
         );
  AOI21_X1 U6065 ( .B1(n5383), .B2(n6699), .A(n4869), .ZN(n4870) );
  OAI211_X1 U6066 ( .C1(n4872), .C2(n6808), .A(n4871), .B(n4870), .ZN(U3130)
         );
  NAND2_X1 U6067 ( .A1(n4832), .A2(n4873), .ZN(n4891) );
  AND2_X1 U6068 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4874) );
  NOR2_X1 U6069 ( .A1(n4878), .A2(n4874), .ZN(n4880) );
  INV_X1 U6070 ( .A(n4874), .ZN(n4877) );
  OAI21_X1 U6071 ( .B1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n4715), .A(n4875), 
        .ZN(n4876) );
  OAI21_X1 U6072 ( .B1(n4878), .B2(n4877), .A(n4876), .ZN(n4879) );
  MUX2_X1 U6073 ( .A(n4880), .B(n4879), .S(n3757), .Z(n4889) );
  INV_X1 U6074 ( .A(n4881), .ZN(n4883) );
  NAND2_X1 U6075 ( .A1(n4885), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4882) );
  NAND2_X1 U6076 ( .A1(n4883), .A2(n4882), .ZN(n4884) );
  NOR2_X1 U6077 ( .A1(n4884), .A2(n3500), .ZN(n6296) );
  NAND2_X1 U6078 ( .A1(n4885), .A2(n4881), .ZN(n4886) );
  OAI21_X1 U6079 ( .B1(n6296), .B2(n4887), .A(n4886), .ZN(n4888) );
  NOR2_X1 U6080 ( .A1(n4889), .A2(n4888), .ZN(n4890) );
  NAND2_X1 U6081 ( .A1(n4891), .A2(n4890), .ZN(n6295) );
  MUX2_X1 U6082 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6295), .S(n5335), 
        .Z(n5346) );
  MUX2_X1 U6083 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n4892), .S(n5335), 
        .Z(n5341) );
  NAND3_X1 U6084 ( .A1(n5346), .A2(n6359), .A3(n5341), .ZN(n4897) );
  NAND2_X1 U6085 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6373), .ZN(n4899) );
  INV_X1 U6086 ( .A(n4899), .ZN(n4894) );
  NAND2_X1 U6087 ( .A1(n4895), .A2(n4894), .ZN(n4896) );
  NAND2_X1 U6088 ( .A1(n4897), .A2(n4896), .ZN(n5357) );
  OAI21_X1 U6089 ( .B1(n5335), .B2(STATE2_REG_1__SCAN_IN), .A(n4899), .ZN(
        n4900) );
  NAND2_X1 U6090 ( .A1(n4900), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4903) );
  OR2_X1 U6091 ( .A1(n4312), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4901) );
  OR2_X1 U6092 ( .A1(n6442), .A2(n4901), .ZN(n4902) );
  NAND2_X1 U6093 ( .A1(n4903), .A2(n4902), .ZN(n5356) );
  NOR3_X1 U6094 ( .A1(n4905), .A2(n5356), .A3(FLUSH_REG_SCAN_IN), .ZN(n4904)
         );
  INV_X1 U6095 ( .A(n4905), .ZN(n4908) );
  NOR2_X1 U6096 ( .A1(n5356), .A2(n4906), .ZN(n4907) );
  NAND2_X1 U6097 ( .A1(n4908), .A2(n4907), .ZN(n6346) );
  INV_X1 U6098 ( .A(n6346), .ZN(n4911) );
  AND2_X1 U6099 ( .A1(n4909), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6291) );
  INV_X1 U6100 ( .A(n3845), .ZN(n6657) );
  OAI22_X1 U6101 ( .A1(n4830), .A2(n6722), .B1(n6291), .B2(n6657), .ZN(n4910)
         );
  OAI21_X1 U6102 ( .B1(n4911), .B2(n4910), .A(n6656), .ZN(n4912) );
  OAI21_X1 U6103 ( .B1(n6656), .B2(n6718), .A(n4912), .ZN(U3465) );
  AND2_X1 U6104 ( .A1(n4913), .A2(n6278), .ZN(n4914) );
  NAND2_X1 U6105 ( .A1(n6283), .A2(n4914), .ZN(n4919) );
  AOI21_X1 U6106 ( .B1(n4919), .B2(n6571), .A(n6725), .ZN(n4918) );
  INV_X1 U6107 ( .A(n6714), .ZN(n5384) );
  OR2_X1 U6108 ( .A1(n5384), .A2(n5255), .ZN(n4915) );
  NAND2_X1 U6109 ( .A1(n4915), .A2(n4943), .ZN(n4920) );
  INV_X1 U6110 ( .A(n5387), .ZN(n4916) );
  NAND2_X1 U6111 ( .A1(n4916), .A2(n6722), .ZN(n4917) );
  NAND2_X1 U6112 ( .A1(n4942), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4923)
         );
  OR2_X1 U6113 ( .A1(n4919), .A2(n4830), .ZN(n5063) );
  AOI22_X1 U6114 ( .A1(n4920), .A2(n6304), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5387), .ZN(n4944) );
  OAI22_X1 U6115 ( .A1(n4944), .A2(n6697), .B1(n4943), .B2(n6791), .ZN(n4921)
         );
  AOI21_X1 U6116 ( .B1(n5096), .B2(n6694), .A(n4921), .ZN(n4922) );
  OAI211_X1 U6117 ( .C1(n5382), .C2(n6797), .A(n4923), .B(n4922), .ZN(U3145)
         );
  NAND2_X1 U6118 ( .A1(n4942), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4926)
         );
  OAI22_X1 U6119 ( .A1(n4944), .A2(n6688), .B1(n4943), .B2(n6784), .ZN(n4924)
         );
  AOI21_X1 U6120 ( .B1(n5096), .B2(n6685), .A(n4924), .ZN(n4925) );
  OAI211_X1 U6121 ( .C1(n5382), .C2(n6790), .A(n4926), .B(n4925), .ZN(U3143)
         );
  NAND2_X1 U6122 ( .A1(n4942), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4929)
         );
  OAI22_X1 U6123 ( .A1(n4944), .A2(n6683), .B1(n4943), .B2(n6777), .ZN(n4927)
         );
  AOI21_X1 U6124 ( .B1(n5096), .B2(n6680), .A(n4927), .ZN(n4928) );
  OAI211_X1 U6125 ( .C1(n5382), .C2(n6783), .A(n4929), .B(n4928), .ZN(U3142)
         );
  NAND2_X1 U6126 ( .A1(n4942), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4932)
         );
  OAI22_X1 U6127 ( .A1(n4944), .A2(n6758), .B1(n4943), .B2(n6704), .ZN(n4930)
         );
  AOI21_X1 U6128 ( .B1(n5096), .B2(n6706), .A(n4930), .ZN(n4931) );
  OAI211_X1 U6129 ( .C1(n5382), .C2(n6343), .A(n4932), .B(n4931), .ZN(U3147)
         );
  NAND2_X1 U6130 ( .A1(n4942), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4935)
         );
  OAI22_X1 U6131 ( .A1(n4944), .A2(n6717), .B1(n4943), .B2(n6661), .ZN(n4933)
         );
  AOI21_X1 U6132 ( .B1(n5096), .B2(n6663), .A(n4933), .ZN(n4934) );
  OAI211_X1 U6133 ( .C1(n5382), .C2(n6316), .A(n4935), .B(n4934), .ZN(U3140)
         );
  NAND2_X1 U6134 ( .A1(n4942), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4938)
         );
  OAI22_X1 U6135 ( .A1(n4944), .A2(n6702), .B1(n4943), .B2(n6799), .ZN(n4936)
         );
  AOI21_X1 U6136 ( .B1(n5096), .B2(n6699), .A(n4936), .ZN(n4937) );
  OAI211_X1 U6137 ( .C1(n5382), .C2(n6808), .A(n4938), .B(n4937), .ZN(U3146)
         );
  NAND2_X1 U6138 ( .A1(n4942), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4941)
         );
  OAI22_X1 U6139 ( .A1(n4944), .A2(n6860), .B1(n4943), .B2(n6850), .ZN(n4939)
         );
  AOI21_X1 U6140 ( .B1(n5096), .B2(n6690), .A(n4939), .ZN(n4940) );
  OAI211_X1 U6141 ( .C1(n5382), .C2(n6329), .A(n4941), .B(n4940), .ZN(U3144)
         );
  NAND2_X1 U6142 ( .A1(n4942), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4947)
         );
  OAI22_X1 U6143 ( .A1(n4944), .A2(n6678), .B1(n4943), .B2(n6770), .ZN(n4945)
         );
  AOI21_X1 U6144 ( .B1(n5096), .B2(n6675), .A(n4945), .ZN(n4946) );
  OAI211_X1 U6145 ( .C1(n5382), .C2(n6776), .A(n4947), .B(n4946), .ZN(U3141)
         );
  OAI21_X1 U6146 ( .B1(n4950), .B2(n4949), .A(n4948), .ZN(n6635) );
  AOI21_X1 U6147 ( .B1(n4952), .B2(n4817), .A(n3174), .ZN(n4974) );
  NAND2_X1 U6148 ( .A1(n5979), .A2(n6464), .ZN(n4953) );
  NAND2_X1 U6149 ( .A1(n6566), .A2(REIP_REG_3__SCAN_IN), .ZN(n6631) );
  OAI211_X1 U6150 ( .C1(n5981), .C2(n7064), .A(n4953), .B(n6631), .ZN(n4954)
         );
  AOI21_X1 U6151 ( .B1(n4974), .B2(n6571), .A(n4954), .ZN(n4955) );
  OAI21_X1 U6152 ( .B1(n6372), .B2(n6635), .A(n4955), .ZN(U2983) );
  INV_X1 U6153 ( .A(n6283), .ZN(n4956) );
  AOI21_X1 U6154 ( .B1(n6289), .B2(n6282), .A(n6722), .ZN(n4962) );
  INV_X1 U6155 ( .A(n4962), .ZN(n4958) );
  NOR2_X1 U6156 ( .A1(n4728), .A2(n6280), .ZN(n5101) );
  NOR2_X1 U6157 ( .A1(n5102), .A2(n5345), .ZN(n5303) );
  AND2_X1 U6158 ( .A1(n5303), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4959)
         );
  AOI21_X1 U6159 ( .B1(n5308), .B2(n3845), .A(n4959), .ZN(n4961) );
  INV_X1 U6160 ( .A(n5303), .ZN(n4957) );
  OAI22_X1 U6161 ( .A1(n4958), .A2(n4961), .B1(n6345), .B2(n4957), .ZN(n6803)
         );
  INV_X1 U6162 ( .A(n6803), .ZN(n4973) );
  INV_X1 U6163 ( .A(n6853), .ZN(n4970) );
  INV_X1 U6164 ( .A(n4959), .ZN(n6798) );
  OAI22_X1 U6165 ( .A1(n6801), .A2(n6734), .B1(n6661), .B2(n6798), .ZN(n4960)
         );
  AOI21_X1 U6166 ( .B1(n4970), .B2(n6731), .A(n4960), .ZN(n4965) );
  NAND2_X1 U6167 ( .A1(n4962), .A2(n4961), .ZN(n4963) );
  OAI211_X1 U6168 ( .C1(n6304), .C2(n5303), .A(n4963), .B(n6668), .ZN(n6805)
         );
  NAND2_X1 U6169 ( .A1(n6805), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4964)
         );
  OAI211_X1 U6170 ( .C1(n4973), .C2(n6717), .A(n4965), .B(n4964), .ZN(U3108)
         );
  OAI22_X1 U6171 ( .A1(n6801), .A2(n6769), .B1(n6704), .B2(n6798), .ZN(n4966)
         );
  AOI21_X1 U6172 ( .B1(n4970), .B2(n6764), .A(n4966), .ZN(n4968) );
  NAND2_X1 U6173 ( .A1(n6805), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4967)
         );
  OAI211_X1 U6174 ( .C1(n4973), .C2(n6758), .A(n4968), .B(n4967), .ZN(U3115)
         );
  OAI22_X1 U6175 ( .A1(n6801), .A2(n6852), .B1(n6850), .B2(n6798), .ZN(n4969)
         );
  AOI21_X1 U6176 ( .B1(n4970), .B2(n6855), .A(n4969), .ZN(n4972) );
  NAND2_X1 U6177 ( .A1(n6805), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4971)
         );
  OAI211_X1 U6178 ( .C1(n4973), .C2(n6860), .A(n4972), .B(n4971), .ZN(U3112)
         );
  INV_X1 U6179 ( .A(n4974), .ZN(n6461) );
  INV_X1 U6180 ( .A(DATAI_3_), .ZN(n4975) );
  INV_X1 U6181 ( .A(EAX_REG_3__SCAN_IN), .ZN(n7160) );
  OAI222_X1 U6182 ( .A1(n6461), .A2(n5859), .B1(n5860), .B2(n4975), .C1(n7160), 
        .C2(n5856), .ZN(U2888) );
  INV_X1 U6183 ( .A(n5476), .ZN(n4978) );
  INV_X1 U6184 ( .A(n4976), .ZN(n4977) );
  OAI21_X1 U6185 ( .B1(n5477), .B2(n4978), .A(n4977), .ZN(n4979) );
  NAND2_X1 U6186 ( .A1(n4979), .A2(n6429), .ZN(n6630) );
  INV_X1 U6187 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4980) );
  OAI222_X1 U6188 ( .A1(n6630), .A2(n5802), .B1(n4980), .B2(n6481), .C1(n6474), 
        .C2(n6461), .ZN(U2856) );
  INV_X1 U6189 ( .A(n5015), .ZN(n4982) );
  INV_X1 U6190 ( .A(n6282), .ZN(n6277) );
  NOR2_X1 U6191 ( .A1(n4982), .A2(n6277), .ZN(n6290) );
  NOR2_X1 U6192 ( .A1(n6290), .A2(n6722), .ZN(n4984) );
  NAND2_X1 U6193 ( .A1(n6714), .A2(n5017), .ZN(n6724) );
  OAI21_X1 U6194 ( .B1(n6724), .B2(n6657), .A(n5009), .ZN(n4987) );
  OAI22_X1 U6195 ( .A1(n5222), .A2(n6785), .B1(n5009), .B2(n6784), .ZN(n4983)
         );
  AOI21_X1 U6196 ( .B1(n6744), .B2(n6723), .A(n4983), .ZN(n4990) );
  INV_X1 U6197 ( .A(n4984), .ZN(n4988) );
  INV_X1 U6198 ( .A(n6719), .ZN(n4985) );
  NAND2_X1 U6199 ( .A1(n4985), .A2(n6722), .ZN(n4986) );
  NAND2_X1 U6200 ( .A1(n5011), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4989) );
  OAI211_X1 U6201 ( .C1(n5014), .C2(n6688), .A(n4990), .B(n4989), .ZN(U3079)
         );
  OAI22_X1 U6202 ( .A1(n5222), .A2(n6734), .B1(n5009), .B2(n6661), .ZN(n4991)
         );
  AOI21_X1 U6203 ( .B1(n6731), .B2(n6723), .A(n4991), .ZN(n4993) );
  NAND2_X1 U6204 ( .A1(n5011), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4992) );
  OAI211_X1 U6205 ( .C1(n5014), .C2(n6717), .A(n4993), .B(n4992), .ZN(U3076)
         );
  INV_X1 U6206 ( .A(n6783), .ZN(n6740) );
  OAI22_X1 U6207 ( .A1(n5222), .A2(n6778), .B1(n5009), .B2(n6777), .ZN(n4994)
         );
  AOI21_X1 U6208 ( .B1(n6740), .B2(n6723), .A(n4994), .ZN(n4996) );
  NAND2_X1 U6209 ( .A1(n5011), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4995) );
  OAI211_X1 U6210 ( .C1(n5014), .C2(n6683), .A(n4996), .B(n4995), .ZN(U3078)
         );
  INV_X1 U6211 ( .A(n6776), .ZN(n6736) );
  OAI22_X1 U6212 ( .A1(n5222), .A2(n6771), .B1(n5009), .B2(n6770), .ZN(n4997)
         );
  AOI21_X1 U6213 ( .B1(n6736), .B2(n6723), .A(n4997), .ZN(n4999) );
  NAND2_X1 U6214 ( .A1(n5011), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4998) );
  OAI211_X1 U6215 ( .C1(n5014), .C2(n6678), .A(n4999), .B(n4998), .ZN(U3077)
         );
  INV_X1 U6216 ( .A(n6797), .ZN(n6751) );
  OAI22_X1 U6217 ( .A1(n5222), .A2(n6792), .B1(n5009), .B2(n6791), .ZN(n5000)
         );
  AOI21_X1 U6218 ( .B1(n6751), .B2(n6723), .A(n5000), .ZN(n5002) );
  NAND2_X1 U6219 ( .A1(n5011), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5001) );
  OAI211_X1 U6220 ( .C1(n5014), .C2(n6697), .A(n5002), .B(n5001), .ZN(U3081)
         );
  OAI22_X1 U6221 ( .A1(n5222), .A2(n6852), .B1(n5009), .B2(n6850), .ZN(n5003)
         );
  AOI21_X1 U6222 ( .B1(n6855), .B2(n6723), .A(n5003), .ZN(n5005) );
  NAND2_X1 U6223 ( .A1(n5011), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5004) );
  OAI211_X1 U6224 ( .C1(n5014), .C2(n6860), .A(n5005), .B(n5004), .ZN(U3080)
         );
  INV_X1 U6225 ( .A(n6808), .ZN(n6755) );
  OAI22_X1 U6226 ( .A1(n5222), .A2(n6800), .B1(n5009), .B2(n6799), .ZN(n5006)
         );
  AOI21_X1 U6227 ( .B1(n6755), .B2(n6723), .A(n5006), .ZN(n5008) );
  NAND2_X1 U6228 ( .A1(n5011), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5007) );
  OAI211_X1 U6229 ( .C1(n5014), .C2(n6702), .A(n5008), .B(n5007), .ZN(U3082)
         );
  OAI22_X1 U6230 ( .A1(n5222), .A2(n6769), .B1(n5009), .B2(n6704), .ZN(n5010)
         );
  AOI21_X1 U6231 ( .B1(n6764), .B2(n6723), .A(n5010), .ZN(n5013) );
  NAND2_X1 U6232 ( .A1(n5011), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5012) );
  OAI211_X1 U6233 ( .C1(n5014), .C2(n6758), .A(n5013), .B(n5012), .ZN(U3083)
         );
  AOI21_X1 U6234 ( .B1(n6660), .B2(STATEBS16_REG_SCAN_IN), .A(n6722), .ZN(
        n6664) );
  NAND2_X1 U6235 ( .A1(n5149), .A2(n5017), .ZN(n6658) );
  OAI211_X1 U6236 ( .C1(n6725), .C2(n5134), .A(n6664), .B(n6658), .ZN(n5021)
         );
  NOR2_X1 U6237 ( .A1(n5018), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6665)
         );
  NAND2_X1 U6238 ( .A1(n6665), .A2(n6718), .ZN(n5045) );
  NOR2_X1 U6239 ( .A1(n5022), .A2(n6345), .ZN(n6303) );
  INV_X1 U6240 ( .A(n5145), .ZN(n5148) );
  AOI21_X1 U6241 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6301), .A(n5019), .ZN(
        n5144) );
  OAI21_X1 U6242 ( .B1(n6345), .B2(n5148), .A(n5144), .ZN(n5064) );
  AOI211_X1 U6243 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5045), .A(n6303), .B(
        n5064), .ZN(n5020) );
  NAND2_X1 U6244 ( .A1(n5044), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5025) );
  NOR2_X1 U6245 ( .A1(n4832), .A2(n6722), .ZN(n6715) );
  NOR2_X1 U6246 ( .A1(n5145), .A2(n6301), .ZN(n5068) );
  AOI22_X1 U6247 ( .A1(n6715), .A2(n5149), .B1(n6713), .B2(n5068), .ZN(n5046)
         );
  OAI22_X1 U6248 ( .A1(n5046), .A2(n6717), .B1(n6661), .B2(n5045), .ZN(n5023)
         );
  AOI21_X1 U6249 ( .B1(n5048), .B2(n6731), .A(n5023), .ZN(n5024) );
  OAI211_X1 U6250 ( .C1(n6734), .C2(n6671), .A(n5025), .B(n5024), .ZN(U3052)
         );
  NAND2_X1 U6251 ( .A1(n5044), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5028) );
  OAI22_X1 U6252 ( .A1(n5046), .A2(n6688), .B1(n6784), .B2(n5045), .ZN(n5026)
         );
  AOI21_X1 U6253 ( .B1(n5048), .B2(n6744), .A(n5026), .ZN(n5027) );
  OAI211_X1 U6254 ( .C1(n6671), .C2(n6785), .A(n5028), .B(n5027), .ZN(U3055)
         );
  NAND2_X1 U6255 ( .A1(n5044), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5031) );
  OAI22_X1 U6256 ( .A1(n5046), .A2(n6678), .B1(n6770), .B2(n5045), .ZN(n5029)
         );
  AOI21_X1 U6257 ( .B1(n5048), .B2(n6736), .A(n5029), .ZN(n5030) );
  OAI211_X1 U6258 ( .C1(n6671), .C2(n6771), .A(n5031), .B(n5030), .ZN(U3053)
         );
  NAND2_X1 U6259 ( .A1(n5044), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5034) );
  OAI22_X1 U6260 ( .A1(n5046), .A2(n6758), .B1(n6704), .B2(n5045), .ZN(n5032)
         );
  AOI21_X1 U6261 ( .B1(n5048), .B2(n6764), .A(n5032), .ZN(n5033) );
  OAI211_X1 U6262 ( .C1(n6671), .C2(n6769), .A(n5034), .B(n5033), .ZN(U3059)
         );
  NAND2_X1 U6263 ( .A1(n5044), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5037) );
  OAI22_X1 U6264 ( .A1(n5046), .A2(n6683), .B1(n6777), .B2(n5045), .ZN(n5035)
         );
  AOI21_X1 U6265 ( .B1(n5048), .B2(n6740), .A(n5035), .ZN(n5036) );
  OAI211_X1 U6266 ( .C1(n6671), .C2(n6778), .A(n5037), .B(n5036), .ZN(U3054)
         );
  NAND2_X1 U6267 ( .A1(n5044), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5040) );
  OAI22_X1 U6268 ( .A1(n5046), .A2(n6697), .B1(n6791), .B2(n5045), .ZN(n5038)
         );
  AOI21_X1 U6269 ( .B1(n5048), .B2(n6751), .A(n5038), .ZN(n5039) );
  OAI211_X1 U6270 ( .C1(n6671), .C2(n6792), .A(n5040), .B(n5039), .ZN(U3057)
         );
  NAND2_X1 U6271 ( .A1(n5044), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5043) );
  OAI22_X1 U6272 ( .A1(n5046), .A2(n6860), .B1(n6850), .B2(n5045), .ZN(n5041)
         );
  AOI21_X1 U6273 ( .B1(n5048), .B2(n6855), .A(n5041), .ZN(n5042) );
  OAI211_X1 U6274 ( .C1(n6671), .C2(n6852), .A(n5043), .B(n5042), .ZN(U3056)
         );
  NAND2_X1 U6275 ( .A1(n5044), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5050) );
  OAI22_X1 U6276 ( .A1(n5046), .A2(n6702), .B1(n6799), .B2(n5045), .ZN(n5047)
         );
  AOI21_X1 U6277 ( .B1(n5048), .B2(n6755), .A(n5047), .ZN(n5049) );
  OAI211_X1 U6278 ( .C1(n6671), .C2(n6800), .A(n5050), .B(n5049), .ZN(U3058)
         );
  OAI21_X1 U6279 ( .B1(n5053), .B2(n5052), .A(n5051), .ZN(n5376) );
  INV_X1 U6280 ( .A(n5054), .ZN(n5057) );
  INV_X1 U6281 ( .A(n5055), .ZN(n5056) );
  AND2_X1 U6282 ( .A1(n5055), .A2(n5054), .ZN(n5298) );
  AOI21_X1 U6283 ( .B1(n5057), .B2(n5056), .A(n5298), .ZN(n5443) );
  INV_X1 U6284 ( .A(n5058), .ZN(n5453) );
  AOI22_X1 U6285 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6566), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n5059) );
  OAI21_X1 U6286 ( .B1(n5453), .B2(n6586), .A(n5059), .ZN(n5060) );
  AOI21_X1 U6287 ( .B1(n5443), .B2(n6571), .A(n5060), .ZN(n5061) );
  OAI21_X1 U6288 ( .B1(n6372), .B2(n5376), .A(n5061), .ZN(U2981) );
  INV_X1 U6289 ( .A(n5183), .ZN(n5062) );
  AOI21_X1 U6290 ( .B1(n5183), .B2(n6304), .A(n6725), .ZN(n5188) );
  INV_X1 U6291 ( .A(n5188), .ZN(n5182) );
  INV_X1 U6292 ( .A(n4728), .ZN(n6284) );
  NAND2_X1 U6293 ( .A1(n6284), .A2(n6280), .ZN(n5254) );
  OAI211_X1 U6294 ( .C1(n6725), .C2(n5063), .A(n5182), .B(n5180), .ZN(n5066)
         );
  NOR2_X1 U6295 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6296 ( .A1(n5217), .A2(n5345), .ZN(n5185) );
  OR2_X1 U6297 ( .A1(n5185), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5093)
         );
  AOI211_X1 U6298 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5093), .A(n6713), .B(
        n5064), .ZN(n5065) );
  NAND2_X1 U6299 ( .A1(n5092), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5073) );
  INV_X1 U6300 ( .A(n5180), .ZN(n5067) );
  NAND2_X1 U6301 ( .A1(n5067), .A2(n6304), .ZN(n5070) );
  NAND2_X1 U6302 ( .A1(n5068), .A2(n6303), .ZN(n5069) );
  OAI22_X1 U6303 ( .A1(n5094), .A2(n6678), .B1(n6770), .B2(n5093), .ZN(n5071)
         );
  AOI21_X1 U6304 ( .B1(n5096), .B2(n6736), .A(n5071), .ZN(n5072) );
  OAI211_X1 U6305 ( .C1(n5210), .C2(n6771), .A(n5073), .B(n5072), .ZN(U3021)
         );
  NAND2_X1 U6306 ( .A1(n5092), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5076) );
  OAI22_X1 U6307 ( .A1(n5094), .A2(n6688), .B1(n6784), .B2(n5093), .ZN(n5074)
         );
  AOI21_X1 U6308 ( .B1(n5096), .B2(n6744), .A(n5074), .ZN(n5075) );
  OAI211_X1 U6309 ( .C1(n5210), .C2(n6785), .A(n5076), .B(n5075), .ZN(U3023)
         );
  NAND2_X1 U6310 ( .A1(n5092), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5079) );
  OAI22_X1 U6311 ( .A1(n5094), .A2(n6697), .B1(n6791), .B2(n5093), .ZN(n5077)
         );
  AOI21_X1 U6312 ( .B1(n5096), .B2(n6751), .A(n5077), .ZN(n5078) );
  OAI211_X1 U6313 ( .C1(n5210), .C2(n6792), .A(n5079), .B(n5078), .ZN(U3025)
         );
  NAND2_X1 U6314 ( .A1(n5092), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5082) );
  OAI22_X1 U6315 ( .A1(n5094), .A2(n6860), .B1(n6850), .B2(n5093), .ZN(n5080)
         );
  AOI21_X1 U6316 ( .B1(n5096), .B2(n6855), .A(n5080), .ZN(n5081) );
  OAI211_X1 U6317 ( .C1(n5210), .C2(n6852), .A(n5082), .B(n5081), .ZN(U3024)
         );
  NAND2_X1 U6318 ( .A1(n5092), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5085) );
  OAI22_X1 U6319 ( .A1(n5094), .A2(n6702), .B1(n6799), .B2(n5093), .ZN(n5083)
         );
  AOI21_X1 U6320 ( .B1(n5096), .B2(n6755), .A(n5083), .ZN(n5084) );
  OAI211_X1 U6321 ( .C1(n5210), .C2(n6800), .A(n5085), .B(n5084), .ZN(U3026)
         );
  NAND2_X1 U6322 ( .A1(n5092), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5088) );
  OAI22_X1 U6323 ( .A1(n5094), .A2(n6683), .B1(n6777), .B2(n5093), .ZN(n5086)
         );
  AOI21_X1 U6324 ( .B1(n5096), .B2(n6740), .A(n5086), .ZN(n5087) );
  OAI211_X1 U6325 ( .C1(n5210), .C2(n6778), .A(n5088), .B(n5087), .ZN(U3022)
         );
  NAND2_X1 U6326 ( .A1(n5092), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5091) );
  OAI22_X1 U6327 ( .A1(n5094), .A2(n6717), .B1(n6661), .B2(n5093), .ZN(n5089)
         );
  AOI21_X1 U6328 ( .B1(n5096), .B2(n6731), .A(n5089), .ZN(n5090) );
  OAI211_X1 U6329 ( .C1(n5210), .C2(n6734), .A(n5091), .B(n5090), .ZN(U3020)
         );
  NAND2_X1 U6330 ( .A1(n5092), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5098) );
  OAI22_X1 U6331 ( .A1(n5094), .A2(n6758), .B1(n6704), .B2(n5093), .ZN(n5095)
         );
  AOI21_X1 U6332 ( .B1(n5096), .B2(n6764), .A(n5095), .ZN(n5097) );
  OAI211_X1 U6333 ( .C1(n5210), .C2(n6769), .A(n5098), .B(n5097), .ZN(U3027)
         );
  INV_X1 U6334 ( .A(n5443), .ZN(n5296) );
  INV_X1 U6335 ( .A(DATAI_5_), .ZN(n5099) );
  INV_X1 U6336 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6546) );
  OAI222_X1 U6337 ( .A1(n5296), .A2(n5859), .B1(n5860), .B2(n5099), .C1(n5856), 
        .C2(n6546), .ZN(U2886) );
  AOI21_X1 U6338 ( .B1(n5100), .B2(n6282), .A(n6722), .ZN(n5109) );
  NAND2_X1 U6339 ( .A1(n6453), .A2(n5101), .ZN(n6310) );
  OR2_X1 U6340 ( .A1(n6310), .A2(n6657), .ZN(n5103) );
  OR2_X1 U6341 ( .A1(n5102), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6306)
         );
  INV_X1 U6342 ( .A(n6306), .ZN(n5104) );
  NAND2_X1 U6343 ( .A1(n5104), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6344 ( .A1(n5103), .A2(n5133), .ZN(n5111) );
  INV_X1 U6345 ( .A(n5105), .ZN(n5106) );
  OAI22_X1 U6346 ( .A1(n5134), .A2(n6771), .B1(n6770), .B2(n5133), .ZN(n5108)
         );
  AOI21_X1 U6347 ( .B1(n6736), .B2(n6341), .A(n5108), .ZN(n5114) );
  INV_X1 U6348 ( .A(n5109), .ZN(n5112) );
  NAND2_X1 U6349 ( .A1(n6306), .A2(n6722), .ZN(n5110) );
  NAND2_X1 U6350 ( .A1(n5136), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5113) );
  OAI211_X1 U6351 ( .C1(n5139), .C2(n6678), .A(n5114), .B(n5113), .ZN(U3045)
         );
  OAI22_X1 U6352 ( .A1(n5134), .A2(n6792), .B1(n6791), .B2(n5133), .ZN(n5115)
         );
  AOI21_X1 U6353 ( .B1(n6751), .B2(n6341), .A(n5115), .ZN(n5117) );
  NAND2_X1 U6354 ( .A1(n5136), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5116) );
  OAI211_X1 U6355 ( .C1(n5139), .C2(n6697), .A(n5117), .B(n5116), .ZN(U3049)
         );
  OAI22_X1 U6356 ( .A1(n5134), .A2(n6734), .B1(n6661), .B2(n5133), .ZN(n5118)
         );
  AOI21_X1 U6357 ( .B1(n6731), .B2(n6341), .A(n5118), .ZN(n5120) );
  NAND2_X1 U6358 ( .A1(n5136), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5119) );
  OAI211_X1 U6359 ( .C1(n5139), .C2(n6717), .A(n5120), .B(n5119), .ZN(U3044)
         );
  OAI22_X1 U6360 ( .A1(n5134), .A2(n6769), .B1(n6704), .B2(n5133), .ZN(n5121)
         );
  AOI21_X1 U6361 ( .B1(n6764), .B2(n6341), .A(n5121), .ZN(n5123) );
  NAND2_X1 U6362 ( .A1(n5136), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5122) );
  OAI211_X1 U6363 ( .C1(n5139), .C2(n6758), .A(n5123), .B(n5122), .ZN(U3051)
         );
  OAI22_X1 U6364 ( .A1(n5134), .A2(n6800), .B1(n6799), .B2(n5133), .ZN(n5124)
         );
  AOI21_X1 U6365 ( .B1(n6755), .B2(n6341), .A(n5124), .ZN(n5126) );
  NAND2_X1 U6366 ( .A1(n5136), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5125) );
  OAI211_X1 U6367 ( .C1(n5139), .C2(n6702), .A(n5126), .B(n5125), .ZN(U3050)
         );
  OAI22_X1 U6368 ( .A1(n5134), .A2(n6785), .B1(n6784), .B2(n5133), .ZN(n5127)
         );
  AOI21_X1 U6369 ( .B1(n6744), .B2(n6341), .A(n5127), .ZN(n5129) );
  NAND2_X1 U6370 ( .A1(n5136), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5128) );
  OAI211_X1 U6371 ( .C1(n5139), .C2(n6688), .A(n5129), .B(n5128), .ZN(U3047)
         );
  OAI22_X1 U6372 ( .A1(n5134), .A2(n6778), .B1(n6777), .B2(n5133), .ZN(n5130)
         );
  AOI21_X1 U6373 ( .B1(n6740), .B2(n6341), .A(n5130), .ZN(n5132) );
  NAND2_X1 U6374 ( .A1(n5136), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5131) );
  OAI211_X1 U6375 ( .C1(n5139), .C2(n6683), .A(n5132), .B(n5131), .ZN(U3046)
         );
  OAI22_X1 U6376 ( .A1(n5134), .A2(n6852), .B1(n6850), .B2(n5133), .ZN(n5135)
         );
  AOI21_X1 U6377 ( .B1(n6855), .B2(n6341), .A(n5135), .ZN(n5138) );
  NAND2_X1 U6378 ( .A1(n5136), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5137) );
  OAI211_X1 U6379 ( .C1(n5139), .C2(n6860), .A(n5138), .B(n5137), .ZN(U3048)
         );
  INV_X1 U6380 ( .A(n6801), .ZN(n5140) );
  NOR3_X1 U6381 ( .A1(n5140), .A2(n5175), .A3(n6722), .ZN(n5142) );
  OAI22_X1 U6382 ( .A1(n5142), .A2(n6725), .B1(n6453), .B2(n5141), .ZN(n5147)
         );
  NAND2_X1 U6383 ( .A1(n5143), .A2(n6718), .ZN(n5172) );
  OAI21_X1 U6384 ( .B1(n5145), .B2(n6345), .A(n5144), .ZN(n5218) );
  AOI211_X1 U6385 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5172), .A(n6303), .B(
        n5218), .ZN(n5146) );
  NAND2_X1 U6386 ( .A1(n5171), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5152)
         );
  AND2_X1 U6387 ( .A1(n4832), .A2(n6304), .ZN(n5391) );
  NOR2_X1 U6388 ( .A1(n5148), .A2(n6301), .ZN(n5223) );
  AOI22_X1 U6389 ( .A1(n5391), .A2(n5149), .B1(n6713), .B2(n5223), .ZN(n5173)
         );
  OAI22_X1 U6390 ( .A1(n5173), .A2(n6758), .B1(n6704), .B2(n5172), .ZN(n5150)
         );
  AOI21_X1 U6391 ( .B1(n5175), .B2(n6706), .A(n5150), .ZN(n5151) );
  OAI211_X1 U6392 ( .C1(n6801), .C2(n6343), .A(n5152), .B(n5151), .ZN(U3123)
         );
  NAND2_X1 U6393 ( .A1(n5171), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5155)
         );
  OAI22_X1 U6394 ( .A1(n5173), .A2(n6688), .B1(n6784), .B2(n5172), .ZN(n5153)
         );
  AOI21_X1 U6395 ( .B1(n5175), .B2(n6685), .A(n5153), .ZN(n5154) );
  OAI211_X1 U6396 ( .C1(n6801), .C2(n6790), .A(n5155), .B(n5154), .ZN(U3119)
         );
  NAND2_X1 U6397 ( .A1(n5171), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5158)
         );
  OAI22_X1 U6398 ( .A1(n5173), .A2(n6702), .B1(n6799), .B2(n5172), .ZN(n5156)
         );
  AOI21_X1 U6399 ( .B1(n5175), .B2(n6699), .A(n5156), .ZN(n5157) );
  OAI211_X1 U6400 ( .C1(n6801), .C2(n6808), .A(n5158), .B(n5157), .ZN(U3122)
         );
  NAND2_X1 U6401 ( .A1(n5171), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5161)
         );
  OAI22_X1 U6402 ( .A1(n5173), .A2(n6697), .B1(n6791), .B2(n5172), .ZN(n5159)
         );
  AOI21_X1 U6403 ( .B1(n5175), .B2(n6694), .A(n5159), .ZN(n5160) );
  OAI211_X1 U6404 ( .C1(n6801), .C2(n6797), .A(n5161), .B(n5160), .ZN(U3121)
         );
  NAND2_X1 U6405 ( .A1(n5171), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5164)
         );
  OAI22_X1 U6406 ( .A1(n5173), .A2(n6860), .B1(n6850), .B2(n5172), .ZN(n5162)
         );
  AOI21_X1 U6407 ( .B1(n5175), .B2(n6690), .A(n5162), .ZN(n5163) );
  OAI211_X1 U6408 ( .C1(n6801), .C2(n6329), .A(n5164), .B(n5163), .ZN(U3120)
         );
  NAND2_X1 U6409 ( .A1(n5171), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5167)
         );
  OAI22_X1 U6410 ( .A1(n5173), .A2(n6683), .B1(n6777), .B2(n5172), .ZN(n5165)
         );
  AOI21_X1 U6411 ( .B1(n5175), .B2(n6680), .A(n5165), .ZN(n5166) );
  OAI211_X1 U6412 ( .C1(n6801), .C2(n6783), .A(n5167), .B(n5166), .ZN(U3118)
         );
  NAND2_X1 U6413 ( .A1(n5171), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5170)
         );
  OAI22_X1 U6414 ( .A1(n5173), .A2(n6678), .B1(n6770), .B2(n5172), .ZN(n5168)
         );
  AOI21_X1 U6415 ( .B1(n5175), .B2(n6675), .A(n5168), .ZN(n5169) );
  OAI211_X1 U6416 ( .C1(n6801), .C2(n6776), .A(n5170), .B(n5169), .ZN(U3117)
         );
  NAND2_X1 U6417 ( .A1(n5171), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5177)
         );
  OAI22_X1 U6418 ( .A1(n5173), .A2(n6717), .B1(n6661), .B2(n5172), .ZN(n5174)
         );
  AOI21_X1 U6419 ( .B1(n5175), .B2(n6663), .A(n5174), .ZN(n5176) );
  OAI211_X1 U6420 ( .C1(n6801), .C2(n6316), .A(n5177), .B(n5176), .ZN(U3116)
         );
  INV_X1 U6421 ( .A(DATAI_4_), .ZN(n6511) );
  XOR2_X1 U6422 ( .A(n5178), .B(n4951), .Z(n6572) );
  INV_X1 U6423 ( .A(n6572), .ZN(n5179) );
  INV_X1 U6424 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6975) );
  OAI222_X1 U6425 ( .A1(n5860), .A2(n6511), .B1(n5859), .B2(n5179), .C1(n6975), 
        .C2(n5856), .ZN(U2887) );
  OR2_X1 U6426 ( .A1(n5185), .A2(n6718), .ZN(n5209) );
  OAI21_X1 U6427 ( .B1(n5180), .B2(n6657), .A(n5209), .ZN(n5187) );
  INV_X1 U6428 ( .A(n5185), .ZN(n5181) );
  OAI22_X1 U6429 ( .A1(n5210), .A2(n6343), .B1(n6704), .B2(n5209), .ZN(n5184)
         );
  AOI21_X1 U6430 ( .B1(n6706), .B2(n6308), .A(n5184), .ZN(n5190) );
  NAND2_X1 U6431 ( .A1(n5185), .A2(n6722), .ZN(n5186) );
  NAND2_X1 U6432 ( .A1(n5212), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5189) );
  OAI211_X1 U6433 ( .C1(n5215), .C2(n6758), .A(n5190), .B(n5189), .ZN(U3035)
         );
  OAI22_X1 U6434 ( .A1(n5210), .A2(n6797), .B1(n6791), .B2(n5209), .ZN(n5191)
         );
  AOI21_X1 U6435 ( .B1(n6694), .B2(n6308), .A(n5191), .ZN(n5193) );
  NAND2_X1 U6436 ( .A1(n5212), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5192) );
  OAI211_X1 U6437 ( .C1(n5215), .C2(n6697), .A(n5193), .B(n5192), .ZN(U3033)
         );
  OAI22_X1 U6438 ( .A1(n5210), .A2(n6776), .B1(n6770), .B2(n5209), .ZN(n5194)
         );
  AOI21_X1 U6439 ( .B1(n6675), .B2(n6308), .A(n5194), .ZN(n5196) );
  NAND2_X1 U6440 ( .A1(n5212), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n5195) );
  OAI211_X1 U6441 ( .C1(n5215), .C2(n6678), .A(n5196), .B(n5195), .ZN(U3029)
         );
  OAI22_X1 U6442 ( .A1(n5210), .A2(n6790), .B1(n6784), .B2(n5209), .ZN(n5197)
         );
  AOI21_X1 U6443 ( .B1(n6685), .B2(n6308), .A(n5197), .ZN(n5199) );
  NAND2_X1 U6444 ( .A1(n5212), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5198) );
  OAI211_X1 U6445 ( .C1(n5215), .C2(n6688), .A(n5199), .B(n5198), .ZN(U3031)
         );
  OAI22_X1 U6446 ( .A1(n5210), .A2(n6316), .B1(n6661), .B2(n5209), .ZN(n5200)
         );
  AOI21_X1 U6447 ( .B1(n6663), .B2(n6308), .A(n5200), .ZN(n5202) );
  NAND2_X1 U6448 ( .A1(n5212), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5201) );
  OAI211_X1 U6449 ( .C1(n5215), .C2(n6717), .A(n5202), .B(n5201), .ZN(U3028)
         );
  OAI22_X1 U6450 ( .A1(n5210), .A2(n6783), .B1(n6777), .B2(n5209), .ZN(n5203)
         );
  AOI21_X1 U6451 ( .B1(n6680), .B2(n6308), .A(n5203), .ZN(n5205) );
  NAND2_X1 U6452 ( .A1(n5212), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5204) );
  OAI211_X1 U6453 ( .C1(n5215), .C2(n6683), .A(n5205), .B(n5204), .ZN(U3030)
         );
  OAI22_X1 U6454 ( .A1(n5210), .A2(n6329), .B1(n6850), .B2(n5209), .ZN(n5206)
         );
  AOI21_X1 U6455 ( .B1(n6690), .B2(n6308), .A(n5206), .ZN(n5208) );
  NAND2_X1 U6456 ( .A1(n5212), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5207) );
  OAI211_X1 U6457 ( .C1(n5215), .C2(n6860), .A(n5208), .B(n5207), .ZN(U3032)
         );
  OAI22_X1 U6458 ( .A1(n5210), .A2(n6808), .B1(n6799), .B2(n5209), .ZN(n5211)
         );
  AOI21_X1 U6459 ( .B1(n6699), .B2(n6308), .A(n5211), .ZN(n5214) );
  NAND2_X1 U6460 ( .A1(n5212), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5213) );
  OAI211_X1 U6461 ( .C1(n5215), .C2(n6702), .A(n5214), .B(n5213), .ZN(U3034)
         );
  AOI21_X1 U6462 ( .B1(n5287), .B2(n5222), .A(n6371), .ZN(n5221) );
  OAI21_X1 U6463 ( .B1(n6453), .B2(n5254), .A(n6304), .ZN(n5220) );
  NAND2_X1 U6464 ( .A1(n5217), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5259) );
  OR2_X1 U6465 ( .A1(n5259), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5247)
         );
  AOI211_X1 U6466 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5247), .A(n6713), .B(
        n5218), .ZN(n5219) );
  NAND2_X1 U6467 ( .A1(n5246), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5227) );
  INV_X1 U6468 ( .A(n5254), .ZN(n5224) );
  AOI22_X1 U6469 ( .A1(n5391), .A2(n5224), .B1(n6303), .B2(n5223), .ZN(n5248)
         );
  OAI22_X1 U6470 ( .A1(n5248), .A2(n6688), .B1(n6784), .B2(n5247), .ZN(n5225)
         );
  AOI21_X1 U6471 ( .B1(n5250), .B2(n6744), .A(n5225), .ZN(n5226) );
  OAI211_X1 U6472 ( .C1(n5287), .C2(n6785), .A(n5227), .B(n5226), .ZN(U3087)
         );
  NAND2_X1 U6473 ( .A1(n5246), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5230) );
  OAI22_X1 U6474 ( .A1(n5248), .A2(n6758), .B1(n6704), .B2(n5247), .ZN(n5228)
         );
  AOI21_X1 U6475 ( .B1(n5250), .B2(n6764), .A(n5228), .ZN(n5229) );
  OAI211_X1 U6476 ( .C1(n5287), .C2(n6769), .A(n5230), .B(n5229), .ZN(U3091)
         );
  NAND2_X1 U6477 ( .A1(n5246), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5233) );
  OAI22_X1 U6478 ( .A1(n5248), .A2(n6697), .B1(n6791), .B2(n5247), .ZN(n5231)
         );
  AOI21_X1 U6479 ( .B1(n5250), .B2(n6751), .A(n5231), .ZN(n5232) );
  OAI211_X1 U6480 ( .C1(n5287), .C2(n6792), .A(n5233), .B(n5232), .ZN(U3089)
         );
  NAND2_X1 U6481 ( .A1(n5246), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5236) );
  OAI22_X1 U6482 ( .A1(n5248), .A2(n6717), .B1(n6661), .B2(n5247), .ZN(n5234)
         );
  AOI21_X1 U6483 ( .B1(n5250), .B2(n6731), .A(n5234), .ZN(n5235) );
  OAI211_X1 U6484 ( .C1(n5287), .C2(n6734), .A(n5236), .B(n5235), .ZN(U3084)
         );
  NAND2_X1 U6485 ( .A1(n5246), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5239) );
  OAI22_X1 U6486 ( .A1(n5248), .A2(n6860), .B1(n6850), .B2(n5247), .ZN(n5237)
         );
  AOI21_X1 U6487 ( .B1(n5250), .B2(n6855), .A(n5237), .ZN(n5238) );
  OAI211_X1 U6488 ( .C1(n5287), .C2(n6852), .A(n5239), .B(n5238), .ZN(U3088)
         );
  NAND2_X1 U6489 ( .A1(n5246), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5242) );
  OAI22_X1 U6490 ( .A1(n5248), .A2(n6683), .B1(n6777), .B2(n5247), .ZN(n5240)
         );
  AOI21_X1 U6491 ( .B1(n5250), .B2(n6740), .A(n5240), .ZN(n5241) );
  OAI211_X1 U6492 ( .C1(n5287), .C2(n6778), .A(n5242), .B(n5241), .ZN(U3086)
         );
  NAND2_X1 U6493 ( .A1(n5246), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5245) );
  OAI22_X1 U6494 ( .A1(n5248), .A2(n6678), .B1(n6770), .B2(n5247), .ZN(n5243)
         );
  AOI21_X1 U6495 ( .B1(n5250), .B2(n6736), .A(n5243), .ZN(n5244) );
  OAI211_X1 U6496 ( .C1(n5287), .C2(n6771), .A(n5245), .B(n5244), .ZN(U3085)
         );
  NAND2_X1 U6497 ( .A1(n5246), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5252) );
  OAI22_X1 U6498 ( .A1(n5248), .A2(n6702), .B1(n6799), .B2(n5247), .ZN(n5249)
         );
  AOI21_X1 U6499 ( .B1(n5250), .B2(n6755), .A(n5249), .ZN(n5251) );
  OAI211_X1 U6500 ( .C1(n5287), .C2(n6800), .A(n5252), .B(n5251), .ZN(U3090)
         );
  INV_X1 U6501 ( .A(n5263), .ZN(n5253) );
  AOI21_X1 U6502 ( .B1(n5253), .B2(n6304), .A(n6725), .ZN(n5262) );
  INV_X1 U6503 ( .A(n5262), .ZN(n5258) );
  OR2_X1 U6504 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  OR2_X1 U6505 ( .A1(n5259), .A2(n6718), .ZN(n5286) );
  NAND2_X1 U6506 ( .A1(n5256), .A2(n5286), .ZN(n5261) );
  INV_X1 U6507 ( .A(n5259), .ZN(n5257) );
  NAND2_X1 U6508 ( .A1(n5259), .A2(n6722), .ZN(n5260) );
  NAND2_X1 U6509 ( .A1(n5285), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6510 ( .A1(n5263), .A2(n6659), .ZN(n5301) );
  OAI22_X1 U6511 ( .A1(n5287), .A2(n6316), .B1(n6661), .B2(n5286), .ZN(n5264)
         );
  AOI21_X1 U6512 ( .B1(n6856), .B2(n6663), .A(n5264), .ZN(n5265) );
  OAI211_X1 U6513 ( .C1(n5291), .C2(n6717), .A(n5266), .B(n5265), .ZN(U3092)
         );
  NAND2_X1 U6514 ( .A1(n5285), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n5269) );
  OAI22_X1 U6515 ( .A1(n5287), .A2(n6783), .B1(n6777), .B2(n5286), .ZN(n5267)
         );
  AOI21_X1 U6516 ( .B1(n6856), .B2(n6680), .A(n5267), .ZN(n5268) );
  OAI211_X1 U6517 ( .C1(n5291), .C2(n6683), .A(n5269), .B(n5268), .ZN(U3094)
         );
  NAND2_X1 U6518 ( .A1(n5285), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n5272) );
  OAI22_X1 U6519 ( .A1(n5287), .A2(n6343), .B1(n6704), .B2(n5286), .ZN(n5270)
         );
  AOI21_X1 U6520 ( .B1(n6856), .B2(n6706), .A(n5270), .ZN(n5271) );
  OAI211_X1 U6521 ( .C1(n5291), .C2(n6758), .A(n5272), .B(n5271), .ZN(U3099)
         );
  NAND2_X1 U6522 ( .A1(n5285), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n5275) );
  OAI22_X1 U6523 ( .A1(n5287), .A2(n6776), .B1(n6770), .B2(n5286), .ZN(n5273)
         );
  AOI21_X1 U6524 ( .B1(n6856), .B2(n6675), .A(n5273), .ZN(n5274) );
  OAI211_X1 U6525 ( .C1(n5291), .C2(n6678), .A(n5275), .B(n5274), .ZN(U3093)
         );
  NAND2_X1 U6526 ( .A1(n5285), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n5278) );
  OAI22_X1 U6527 ( .A1(n5287), .A2(n6808), .B1(n6799), .B2(n5286), .ZN(n5276)
         );
  AOI21_X1 U6528 ( .B1(n6856), .B2(n6699), .A(n5276), .ZN(n5277) );
  OAI211_X1 U6529 ( .C1(n5291), .C2(n6702), .A(n5278), .B(n5277), .ZN(U3098)
         );
  NAND2_X1 U6530 ( .A1(n5285), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n5281) );
  OAI22_X1 U6531 ( .A1(n5287), .A2(n6790), .B1(n6784), .B2(n5286), .ZN(n5279)
         );
  AOI21_X1 U6532 ( .B1(n6856), .B2(n6685), .A(n5279), .ZN(n5280) );
  OAI211_X1 U6533 ( .C1(n5291), .C2(n6688), .A(n5281), .B(n5280), .ZN(U3095)
         );
  NAND2_X1 U6534 ( .A1(n5285), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n5284) );
  OAI22_X1 U6535 ( .A1(n5287), .A2(n6329), .B1(n6850), .B2(n5286), .ZN(n5282)
         );
  AOI21_X1 U6536 ( .B1(n6856), .B2(n6690), .A(n5282), .ZN(n5283) );
  OAI211_X1 U6537 ( .C1(n5291), .C2(n6860), .A(n5284), .B(n5283), .ZN(U3096)
         );
  NAND2_X1 U6538 ( .A1(n5285), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n5290) );
  OAI22_X1 U6539 ( .A1(n5287), .A2(n6797), .B1(n6791), .B2(n5286), .ZN(n5288)
         );
  AOI21_X1 U6540 ( .B1(n6856), .B2(n6694), .A(n5288), .ZN(n5289) );
  OAI211_X1 U6541 ( .C1(n5291), .C2(n6697), .A(n5290), .B(n5289), .ZN(U3097)
         );
  INV_X1 U6542 ( .A(n6429), .ZN(n5293) );
  AOI21_X1 U6543 ( .B1(n5293), .B2(n6428), .A(n5292), .ZN(n5295) );
  OR2_X1 U6544 ( .A1(n5295), .A2(n5294), .ZN(n5447) );
  OAI222_X1 U6545 ( .A1(n5447), .A2(n5802), .B1(n6481), .B2(n4372), .C1(n6474), 
        .C2(n5296), .ZN(U2854) );
  NOR2_X1 U6546 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  INV_X1 U6547 ( .A(DATAI_6_), .ZN(n5300) );
  OAI222_X1 U6548 ( .A1(n6561), .A2(n5859), .B1(n5856), .B2(n6494), .C1(n5860), 
        .C2(n5300), .ZN(U2885) );
  AOI21_X1 U6549 ( .B1(n5301), .B2(n6853), .A(n6371), .ZN(n5302) );
  AND2_X1 U6550 ( .A1(n6301), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5392)
         );
  NAND2_X1 U6551 ( .A1(n5303), .A2(n6718), .ZN(n6851) );
  OAI22_X1 U6552 ( .A1(n6853), .A2(n6734), .B1(n6851), .B2(n6661), .ZN(n5304)
         );
  AOI21_X1 U6553 ( .B1(n6856), .B2(n6731), .A(n5304), .ZN(n5311) );
  INV_X1 U6554 ( .A(n5305), .ZN(n5309) );
  OAI21_X1 U6555 ( .B1(n6301), .B2(n6345), .A(n5306), .ZN(n5386) );
  NOR2_X1 U6556 ( .A1(n5386), .A2(n6713), .ZN(n6311) );
  AND2_X1 U6557 ( .A1(n5345), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5388) );
  AOI21_X1 U6558 ( .B1(n6851), .B2(STATE2_REG_3__SCAN_IN), .A(n5388), .ZN(
        n5307) );
  NAND2_X1 U6559 ( .A1(n6857), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5310)
         );
  OAI211_X1 U6560 ( .C1(n6861), .C2(n6717), .A(n5311), .B(n5310), .ZN(U3100)
         );
  OAI22_X1 U6561 ( .A1(n6853), .A2(n6800), .B1(n6851), .B2(n6799), .ZN(n5312)
         );
  AOI21_X1 U6562 ( .B1(n6856), .B2(n6755), .A(n5312), .ZN(n5314) );
  NAND2_X1 U6563 ( .A1(n6857), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5313)
         );
  OAI211_X1 U6564 ( .C1(n6861), .C2(n6702), .A(n5314), .B(n5313), .ZN(U3106)
         );
  OAI22_X1 U6565 ( .A1(n6853), .A2(n6778), .B1(n6851), .B2(n6777), .ZN(n5315)
         );
  AOI21_X1 U6566 ( .B1(n6856), .B2(n6740), .A(n5315), .ZN(n5317) );
  NAND2_X1 U6567 ( .A1(n6857), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5316)
         );
  OAI211_X1 U6568 ( .C1(n6861), .C2(n6683), .A(n5317), .B(n5316), .ZN(U3102)
         );
  OAI22_X1 U6569 ( .A1(n6853), .A2(n6769), .B1(n6851), .B2(n6704), .ZN(n5318)
         );
  AOI21_X1 U6570 ( .B1(n6856), .B2(n6764), .A(n5318), .ZN(n5320) );
  NAND2_X1 U6571 ( .A1(n6857), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5319)
         );
  OAI211_X1 U6572 ( .C1(n6861), .C2(n6758), .A(n5320), .B(n5319), .ZN(U3107)
         );
  OAI22_X1 U6573 ( .A1(n6853), .A2(n6771), .B1(n6851), .B2(n6770), .ZN(n5321)
         );
  AOI21_X1 U6574 ( .B1(n6856), .B2(n6736), .A(n5321), .ZN(n5323) );
  NAND2_X1 U6575 ( .A1(n6857), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5322)
         );
  OAI211_X1 U6576 ( .C1(n6861), .C2(n6678), .A(n5323), .B(n5322), .ZN(U3101)
         );
  OAI22_X1 U6577 ( .A1(n6853), .A2(n6792), .B1(n6851), .B2(n6791), .ZN(n5324)
         );
  AOI21_X1 U6578 ( .B1(n6856), .B2(n6751), .A(n5324), .ZN(n5326) );
  NAND2_X1 U6579 ( .A1(n6857), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5325)
         );
  OAI211_X1 U6580 ( .C1(n6861), .C2(n6697), .A(n5326), .B(n5325), .ZN(U3105)
         );
  OAI22_X1 U6581 ( .A1(n6853), .A2(n6785), .B1(n6851), .B2(n6784), .ZN(n5327)
         );
  AOI21_X1 U6582 ( .B1(n6856), .B2(n6744), .A(n5327), .ZN(n5329) );
  NAND2_X1 U6583 ( .A1(n6857), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5328)
         );
  OAI211_X1 U6584 ( .C1(n6861), .C2(n6688), .A(n5329), .B(n5328), .ZN(U3103)
         );
  NAND2_X1 U6585 ( .A1(n5330), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5331) );
  OR2_X1 U6586 ( .A1(n5332), .A2(n5331), .ZN(n5336) );
  INV_X1 U6587 ( .A(n5336), .ZN(n5340) );
  NAND2_X1 U6588 ( .A1(n5341), .A2(n5333), .ZN(n5339) );
  OAI211_X1 U6589 ( .C1(n5337), .C2(n5336), .A(n5335), .B(n5334), .ZN(n5338)
         );
  OAI211_X1 U6590 ( .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n5340), .A(n5339), .B(n5338), .ZN(n5344) );
  INV_X1 U6591 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U6592 ( .A1(n5342), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5343) );
  INV_X1 U6593 ( .A(n5347), .ZN(n5350) );
  INV_X1 U6594 ( .A(n5346), .ZN(n5349) );
  OAI21_X1 U6595 ( .B1(n5347), .B2(n5346), .A(n5345), .ZN(n5348) );
  OAI21_X1 U6596 ( .B1(n5350), .B2(n5349), .A(n5348), .ZN(n5359) );
  NOR2_X1 U6597 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n5352) );
  OAI21_X1 U6598 ( .B1(n5353), .B2(n5352), .A(n5351), .ZN(n5354) );
  AOI21_X1 U6599 ( .B1(n5359), .B2(n7116), .A(n5358), .ZN(n6354) );
  AOI21_X1 U6600 ( .B1(n6354), .B2(n6359), .A(n6938), .ZN(n5364) );
  NAND2_X1 U6601 ( .A1(STATE2_REG_1__SCAN_IN), .A2(READY_N), .ZN(n5360) );
  AOI21_X1 U6602 ( .B1(n6938), .B2(n5360), .A(n6345), .ZN(n5361) );
  OAI21_X1 U6603 ( .B1(n5363), .B2(n5362), .A(n5361), .ZN(n6347) );
  NOR2_X1 U6604 ( .A1(n5364), .A2(n6347), .ZN(n6364) );
  OAI21_X1 U6605 ( .B1(n6364), .B2(n6938), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5366) );
  NAND2_X1 U6606 ( .A1(n5366), .A2(n5365), .ZN(U3453) );
  NAND2_X1 U6607 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5367), .ZN(n6261)
         );
  INV_X1 U6608 ( .A(n5368), .ZN(n5369) );
  OAI22_X1 U6609 ( .A1(n6645), .A2(n5369), .B1(n6646), .B2(n6266), .ZN(n6650)
         );
  AOI21_X1 U6610 ( .B1(n6269), .B2(n6261), .A(n6650), .ZN(n6621) );
  AOI21_X1 U6611 ( .B1(n7150), .B2(n5370), .A(n6621), .ZN(n5374) );
  AND3_X1 U6612 ( .A1(n5371), .A2(n7150), .A3(n6651), .ZN(n5373) );
  OAI22_X1 U6613 ( .A1(n6252), .A2(n5447), .B1(n5444), .B2(n6577), .ZN(n5372)
         );
  NOR3_X1 U6614 ( .A1(n5374), .A2(n5373), .A3(n5372), .ZN(n5375) );
  OAI21_X1 U6615 ( .B1(n6275), .B2(n5376), .A(n5375), .ZN(U3013) );
  NAND2_X1 U6616 ( .A1(n5378), .A2(n5379), .ZN(n5380) );
  NAND2_X1 U6617 ( .A1(n5377), .A2(n5380), .ZN(n6046) );
  AOI22_X1 U6618 ( .A1(n5851), .A2(DATAI_10_), .B1(n5850), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5381) );
  OAI21_X1 U6619 ( .B1(n6046), .B2(n5859), .A(n5381), .ZN(U2881) );
  NOR3_X1 U6620 ( .A1(n5383), .A2(n5420), .A3(n6722), .ZN(n5385) );
  OAI22_X1 U6621 ( .A1(n5385), .A2(n6725), .B1(n6453), .B2(n5384), .ZN(n5390)
         );
  NOR2_X1 U6622 ( .A1(n5386), .A2(n6303), .ZN(n6729) );
  NAND2_X1 U6623 ( .A1(n5387), .A2(n6718), .ZN(n5417) );
  AOI21_X1 U6624 ( .B1(n5417), .B2(STATE2_REG_3__SCAN_IN), .A(n5388), .ZN(
        n5389) );
  NAND3_X1 U6625 ( .A1(n5390), .A2(n6729), .A3(n5389), .ZN(n5416) );
  NAND2_X1 U6626 ( .A1(n5416), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5397)
         );
  NAND2_X1 U6627 ( .A1(n5391), .A2(n6714), .ZN(n5394) );
  NAND2_X1 U6628 ( .A1(n6713), .A2(n5392), .ZN(n5393) );
  OAI22_X1 U6629 ( .A1(n5418), .A2(n6688), .B1(n6784), .B2(n5417), .ZN(n5395)
         );
  AOI21_X1 U6630 ( .B1(n5420), .B2(n6685), .A(n5395), .ZN(n5396) );
  OAI211_X1 U6631 ( .C1(n5423), .C2(n6790), .A(n5397), .B(n5396), .ZN(U3135)
         );
  NAND2_X1 U6632 ( .A1(n5416), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5400)
         );
  OAI22_X1 U6633 ( .A1(n5418), .A2(n6717), .B1(n6661), .B2(n5417), .ZN(n5398)
         );
  AOI21_X1 U6634 ( .B1(n5420), .B2(n6663), .A(n5398), .ZN(n5399) );
  OAI211_X1 U6635 ( .C1(n5423), .C2(n6316), .A(n5400), .B(n5399), .ZN(U3132)
         );
  NAND2_X1 U6636 ( .A1(n5416), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5403)
         );
  OAI22_X1 U6637 ( .A1(n5418), .A2(n6758), .B1(n6704), .B2(n5417), .ZN(n5401)
         );
  AOI21_X1 U6638 ( .B1(n5420), .B2(n6706), .A(n5401), .ZN(n5402) );
  OAI211_X1 U6639 ( .C1(n5423), .C2(n6343), .A(n5403), .B(n5402), .ZN(U3139)
         );
  NAND2_X1 U6640 ( .A1(n5416), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5406)
         );
  OAI22_X1 U6641 ( .A1(n5418), .A2(n6702), .B1(n6799), .B2(n5417), .ZN(n5404)
         );
  AOI21_X1 U6642 ( .B1(n5420), .B2(n6699), .A(n5404), .ZN(n5405) );
  OAI211_X1 U6643 ( .C1(n5423), .C2(n6808), .A(n5406), .B(n5405), .ZN(U3138)
         );
  NAND2_X1 U6644 ( .A1(n5416), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5409)
         );
  OAI22_X1 U6645 ( .A1(n5418), .A2(n6697), .B1(n6791), .B2(n5417), .ZN(n5407)
         );
  AOI21_X1 U6646 ( .B1(n5420), .B2(n6694), .A(n5407), .ZN(n5408) );
  OAI211_X1 U6647 ( .C1(n5423), .C2(n6797), .A(n5409), .B(n5408), .ZN(U3137)
         );
  NAND2_X1 U6648 ( .A1(n5416), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5412)
         );
  OAI22_X1 U6649 ( .A1(n5418), .A2(n6683), .B1(n6777), .B2(n5417), .ZN(n5410)
         );
  AOI21_X1 U6650 ( .B1(n5420), .B2(n6680), .A(n5410), .ZN(n5411) );
  OAI211_X1 U6651 ( .C1(n5423), .C2(n6783), .A(n5412), .B(n5411), .ZN(U3134)
         );
  NAND2_X1 U6652 ( .A1(n5416), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5415)
         );
  OAI22_X1 U6653 ( .A1(n5418), .A2(n6678), .B1(n6770), .B2(n5417), .ZN(n5413)
         );
  AOI21_X1 U6654 ( .B1(n5420), .B2(n6675), .A(n5413), .ZN(n5414) );
  OAI211_X1 U6655 ( .C1(n5423), .C2(n6776), .A(n5415), .B(n5414), .ZN(U3133)
         );
  NAND2_X1 U6656 ( .A1(n5416), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5422)
         );
  OAI22_X1 U6657 ( .A1(n5418), .A2(n6860), .B1(n6850), .B2(n5417), .ZN(n5419)
         );
  AOI21_X1 U6658 ( .B1(n5420), .B2(n6690), .A(n5419), .ZN(n5421) );
  OAI211_X1 U6659 ( .C1(n5423), .C2(n6329), .A(n5422), .B(n5421), .ZN(U3136)
         );
  INV_X1 U6660 ( .A(n5424), .ZN(n5425) );
  AND2_X4 U6661 ( .A1(n5426), .A2(n5425), .ZN(n6463) );
  INV_X1 U6662 ( .A(n6042), .ZN(n5440) );
  NAND2_X1 U6663 ( .A1(n5797), .A2(n5427), .ZN(n5428) );
  NAND2_X1 U6664 ( .A1(n6248), .A2(n5428), .ZN(n6260) );
  INV_X1 U6665 ( .A(n6401), .ZN(n5429) );
  OAI211_X1 U6666 ( .C1(REIP_REG_10__SCAN_IN), .C2(REIP_REG_9__SCAN_IN), .A(
        n5430), .B(n5429), .ZN(n5431) );
  OAI22_X1 U6667 ( .A1(n6452), .A2(n6260), .B1(n6402), .B2(n5431), .ZN(n5439)
         );
  INV_X1 U6668 ( .A(n6433), .ZN(n5459) );
  OAI21_X1 U6669 ( .B1(n5459), .B2(n6401), .A(n6435), .ZN(n6405) );
  INV_X1 U6670 ( .A(EBX_REG_31__SCAN_IN), .ZN(n7090) );
  NAND2_X1 U6671 ( .A1(n5432), .A2(n7090), .ZN(n5433) );
  NOR2_X1 U6672 ( .A1(n5456), .A2(n5433), .ZN(n5434) );
  NOR2_X1 U6673 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  AOI22_X1 U6674 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6458), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n6419), .ZN(n5437) );
  NAND2_X1 U6675 ( .A1(n6433), .A2(n5509), .ZN(n6430) );
  OAI211_X1 U6676 ( .C1(n6405), .C2(n6041), .A(n5437), .B(n6430), .ZN(n5438)
         );
  AOI211_X1 U6677 ( .C1(n6463), .C2(n5440), .A(n5439), .B(n5438), .ZN(n5441)
         );
  OAI21_X1 U6678 ( .B1(n6424), .B2(n6046), .A(n5441), .ZN(U2817) );
  INV_X1 U6679 ( .A(EBX_REG_10__SCAN_IN), .ZN(n7019) );
  OAI222_X1 U6680 ( .A1(n6260), .A2(n5802), .B1(n6481), .B2(n7019), .C1(n6474), 
        .C2(n6046), .ZN(U2849) );
  OR2_X1 U6681 ( .A1(n5458), .A2(n5510), .ZN(n5442) );
  NAND2_X1 U6682 ( .A1(n6424), .A2(n5442), .ZN(n6446) );
  NAND2_X1 U6683 ( .A1(n5443), .A2(n6446), .ZN(n5452) );
  OAI21_X1 U6684 ( .B1(n6402), .B2(n5771), .A(n6433), .ZN(n6417) );
  OAI21_X1 U6685 ( .B1(n6402), .B2(n5445), .A(n5444), .ZN(n5450) );
  NOR2_X1 U6686 ( .A1(n6443), .A2(n4372), .ZN(n5449) );
  NAND2_X1 U6687 ( .A1(n6419), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5446)
         );
  OAI211_X1 U6688 ( .C1(n6452), .C2(n5447), .A(n6430), .B(n5446), .ZN(n5448)
         );
  AOI211_X1 U6689 ( .C1(n6417), .C2(n5450), .A(n5449), .B(n5448), .ZN(n5451)
         );
  OAI211_X1 U6690 ( .C1(n6449), .C2(n5453), .A(n5452), .B(n5451), .ZN(U2822)
         );
  OAI22_X1 U6691 ( .A1(n5454), .A2(n6452), .B1(n6402), .B2(REIP_REG_1__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6692 ( .A1(n5456), .A2(n5455), .ZN(n5457) );
  OR2_X1 U6693 ( .A1(n5458), .A2(n5457), .ZN(n6454) );
  NAND2_X1 U6694 ( .A1(n6458), .A2(EBX_REG_1__SCAN_IN), .ZN(n5461) );
  AOI22_X1 U6695 ( .A1(n6419), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5459), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5460) );
  OAI211_X1 U6696 ( .C1(n6454), .C2(n6280), .A(n5461), .B(n5460), .ZN(n5462)
         );
  AOI211_X1 U6697 ( .C1(n6463), .C2(n4785), .A(n5463), .B(n5462), .ZN(n5464)
         );
  OAI21_X1 U6698 ( .B1(n6460), .B2(n5465), .A(n5464), .ZN(U2826) );
  NOR2_X1 U6699 ( .A1(n6443), .A2(n7050), .ZN(n5468) );
  OAI22_X1 U6700 ( .A1(n6657), .A2(n6454), .B1(n6452), .B2(n5466), .ZN(n5467)
         );
  AOI211_X1 U6701 ( .C1(REIP_REG_0__SCAN_IN), .C2(n6435), .A(n5468), .B(n5467), 
        .ZN(n5470) );
  OAI21_X1 U6702 ( .B1(n6463), .B2(n6419), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5469) );
  OAI211_X1 U6703 ( .C1(n6460), .C2(n5471), .A(n5470), .B(n5469), .ZN(U2827)
         );
  AND2_X1 U6704 ( .A1(n5377), .A2(n5472), .ZN(n5474) );
  OR2_X1 U6705 ( .A1(n5474), .A2(n5473), .ZN(n6470) );
  AOI22_X1 U6706 ( .A1(n5851), .A2(DATAI_11_), .B1(n5850), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5475) );
  OAI21_X1 U6707 ( .B1(n6470), .B2(n5859), .A(n5475), .ZN(U2880) );
  OAI21_X1 U6708 ( .B1(n6402), .B2(REIP_REG_1__SCAN_IN), .A(n6433), .ZN(n6450)
         );
  NAND2_X1 U6709 ( .A1(n6389), .A2(REIP_REG_1__SCAN_IN), .ZN(n6441) );
  XNOR2_X1 U6710 ( .A(n5477), .B(n5476), .ZN(n6643) );
  AOI22_X1 U6711 ( .A1(n6458), .A2(EBX_REG_2__SCAN_IN), .B1(n6439), .B2(n6643), 
        .ZN(n5480) );
  INV_X1 U6712 ( .A(n6454), .ZN(n5478) );
  AOI22_X1 U6713 ( .A1(n5478), .A2(n4728), .B1(n6419), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5479) );
  OAI211_X1 U6714 ( .C1(REIP_REG_2__SCAN_IN), .C2(n6441), .A(n5480), .B(n5479), 
        .ZN(n5481) );
  AOI21_X1 U6715 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6450), .A(n5481), .ZN(n5484)
         );
  INV_X1 U6716 ( .A(n6585), .ZN(n5482) );
  NAND2_X1 U6717 ( .A1(n6463), .A2(n5482), .ZN(n5483) );
  OAI211_X1 U6718 ( .C1(n5485), .C2(n6460), .A(n5484), .B(n5483), .ZN(U2825)
         );
  INV_X1 U6719 ( .A(n6073), .ZN(n5492) );
  OAI22_X1 U6720 ( .A1(n6455), .A2(n6918), .B1(n6443), .B2(n5486), .ZN(n5489)
         );
  OAI21_X1 U6721 ( .B1(n4577), .B2(n6424), .A(n5493), .ZN(U2797) );
  OAI21_X1 U6722 ( .B1(n5494), .B2(n5496), .A(n5495), .ZN(n6004) );
  AOI22_X1 U6723 ( .A1(n5851), .A2(DATAI_14_), .B1(n5850), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5497) );
  OAI21_X1 U6724 ( .B1(n6004), .B2(n5859), .A(n5497), .ZN(U2877) );
  INV_X1 U6725 ( .A(n5498), .ZN(n5721) );
  AND2_X1 U6726 ( .A1(n5721), .A2(n5499), .ZN(n5500) );
  NOR2_X1 U6727 ( .A1(n5703), .A2(n5500), .ZN(n6215) );
  INV_X1 U6728 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U6729 ( .A1(n6419), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5501)
         );
  OAI211_X1 U6730 ( .C1(n6443), .C2(n6977), .A(n6430), .B(n5501), .ZN(n5502)
         );
  AOI21_X1 U6731 ( .B1(n6215), .B2(n6439), .A(n5502), .ZN(n5508) );
  INV_X1 U6732 ( .A(n6006), .ZN(n5506) );
  NAND2_X1 U6733 ( .A1(n5504), .A2(n5503), .ZN(n5505) );
  AOI22_X1 U6734 ( .A1(n6463), .A2(n5506), .B1(n5706), .B2(n5505), .ZN(n5507)
         );
  OAI211_X1 U6735 ( .C1(n6004), .C2(n6424), .A(n5508), .B(n5507), .ZN(U2813)
         );
  OR2_X1 U6736 ( .A1(n5509), .A2(READREQUEST_REG_SCAN_IN), .ZN(n5512) );
  NAND2_X1 U6737 ( .A1(n4360), .A2(n5510), .ZN(n5511) );
  MUX2_X1 U6738 ( .A(n5512), .B(n5511), .S(n6842), .Z(U3474) );
  NAND2_X1 U6739 ( .A1(n5804), .A2(n6411), .ZN(n5522) );
  INV_X1 U6740 ( .A(n5513), .ZN(n5514) );
  NAND2_X1 U6741 ( .A1(n6463), .A2(n5514), .ZN(n5516) );
  NAND2_X1 U6742 ( .A1(n6458), .A2(EBX_REG_29__SCAN_IN), .ZN(n5515) );
  OAI211_X1 U6743 ( .C1(n6455), .C2(n5517), .A(n5516), .B(n5515), .ZN(n5520)
         );
  AND3_X1 U6744 ( .A1(n5533), .A2(REIP_REG_28__SCAN_IN), .A3(n5518), .ZN(n5519) );
  AOI211_X1 U6745 ( .C1(n5532), .C2(REIP_REG_29__SCAN_IN), .A(n5520), .B(n5519), .ZN(n5521) );
  OAI211_X1 U6746 ( .C1(n6452), .C2(n6080), .A(n5522), .B(n5521), .ZN(U2798)
         );
  OR2_X1 U6747 ( .A1(n5526), .A2(n5525), .ZN(n5527) );
  NAND2_X1 U6748 ( .A1(n5528), .A2(n5527), .ZN(n6086) );
  INV_X1 U6749 ( .A(n5862), .ZN(n5531) );
  NAND2_X1 U6750 ( .A1(n6419), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5529)
         );
  OAI21_X1 U6751 ( .B1(n6443), .B2(n5778), .A(n5529), .ZN(n5530) );
  AOI21_X1 U6752 ( .B1(n6463), .B2(n5531), .A(n5530), .ZN(n5535) );
  OAI21_X1 U6753 ( .B1(n5533), .B2(REIP_REG_28__SCAN_IN), .A(n5532), .ZN(n5534) );
  OAI211_X1 U6754 ( .C1(n6086), .C2(n6452), .A(n5535), .B(n5534), .ZN(n5536)
         );
  INV_X1 U6755 ( .A(n5536), .ZN(n5537) );
  OAI21_X1 U6756 ( .B1(n5869), .B2(n6424), .A(n5537), .ZN(U2799) );
  INV_X1 U6757 ( .A(n5538), .ZN(n5554) );
  INV_X1 U6758 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U6759 ( .A1(n6463), .A2(n5873), .ZN(n5540) );
  NAND2_X1 U6760 ( .A1(n6458), .A2(EBX_REG_27__SCAN_IN), .ZN(n5539) );
  OAI211_X1 U6761 ( .C1(n6455), .C2(n5875), .A(n5540), .B(n5539), .ZN(n5541)
         );
  AOI21_X1 U6762 ( .B1(n5554), .B2(REIP_REG_27__SCAN_IN), .A(n5541), .ZN(n5545) );
  INV_X1 U6763 ( .A(n5542), .ZN(n5555) );
  NAND3_X1 U6764 ( .A1(n5555), .A2(REIP_REG_26__SCAN_IN), .A3(n5543), .ZN(
        n5544) );
  OAI211_X1 U6765 ( .C1(n6096), .C2(n6452), .A(n5545), .B(n5544), .ZN(n5546)
         );
  AOI21_X1 U6766 ( .B1(n5877), .B2(n6411), .A(n5546), .ZN(n5547) );
  INV_X1 U6767 ( .A(n5547), .ZN(U2800) );
  INV_X1 U6768 ( .A(n4458), .ZN(n5549) );
  INV_X1 U6769 ( .A(n5883), .ZN(n5815) );
  NAND2_X1 U6770 ( .A1(n5562), .A2(n5551), .ZN(n5552) );
  AND2_X1 U6771 ( .A1(n5553), .A2(n5552), .ZN(n6103) );
  OAI21_X1 U6772 ( .B1(n5555), .B2(REIP_REG_26__SCAN_IN), .A(n5554), .ZN(n5557) );
  AOI22_X1 U6773 ( .A1(n6458), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6419), .ZN(n5556) );
  OAI211_X1 U6774 ( .C1(n6449), .C2(n5881), .A(n5557), .B(n5556), .ZN(n5558)
         );
  AOI21_X1 U6775 ( .B1(n6103), .B2(n6439), .A(n5558), .ZN(n5559) );
  OAI21_X1 U6776 ( .B1(n5815), .B2(n6424), .A(n5559), .ZN(U2801) );
  OAI21_X1 U6777 ( .B1(n5574), .B2(n5563), .A(n5562), .ZN(n6114) );
  INV_X1 U6778 ( .A(n6114), .ZN(n5570) );
  INV_X1 U6779 ( .A(n5588), .ZN(n5605) );
  NOR3_X1 U6780 ( .A1(n5605), .A2(REIP_REG_24__SCAN_IN), .A3(n5564), .ZN(n5580) );
  INV_X1 U6781 ( .A(n5589), .ZN(n5576) );
  OAI21_X1 U6782 ( .B1(n5580), .B2(n5576), .A(REIP_REG_25__SCAN_IN), .ZN(n5567) );
  INV_X1 U6783 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5889) );
  INV_X1 U6784 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5780) );
  OAI22_X1 U6785 ( .A1(n6455), .A2(n5889), .B1(n6443), .B2(n5780), .ZN(n5565)
         );
  AOI21_X1 U6786 ( .B1(n6463), .B2(n5893), .A(n5565), .ZN(n5566) );
  OAI211_X1 U6787 ( .C1(REIP_REG_25__SCAN_IN), .C2(n5568), .A(n5567), .B(n5566), .ZN(n5569) );
  AOI21_X1 U6788 ( .B1(n5570), .B2(n6439), .A(n5569), .ZN(n5571) );
  OAI21_X1 U6789 ( .B1(n5890), .B2(n6424), .A(n5571), .ZN(U2802) );
  NOR2_X1 U6790 ( .A1(n3116), .A2(n5572), .ZN(n5573) );
  AOI21_X1 U6791 ( .B1(n5575), .B2(n5587), .A(n5574), .ZN(n6121) );
  NAND2_X1 U6792 ( .A1(n5576), .A2(REIP_REG_24__SCAN_IN), .ZN(n5578) );
  AOI22_X1 U6793 ( .A1(n6458), .A2(EBX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6419), .ZN(n5577) );
  OAI211_X1 U6794 ( .C1(n6449), .C2(n5912), .A(n5578), .B(n5577), .ZN(n5579)
         );
  AOI211_X1 U6795 ( .C1(n6121), .C2(n6439), .A(n5580), .B(n5579), .ZN(n5581)
         );
  OAI21_X1 U6796 ( .B1(n5915), .B2(n6424), .A(n5581), .ZN(U2803) );
  INV_X1 U6797 ( .A(n5582), .ZN(n5584) );
  AOI21_X1 U6798 ( .B1(n5584), .B2(n3279), .A(n3116), .ZN(n5923) );
  INV_X1 U6799 ( .A(n5923), .ZN(n5822) );
  NAND2_X1 U6800 ( .A1(n3121), .A2(n5585), .ZN(n5586) );
  NAND2_X1 U6801 ( .A1(n5587), .A2(n5586), .ZN(n6129) );
  INV_X1 U6802 ( .A(n6129), .ZN(n5594) );
  AOI21_X1 U6803 ( .B1(n5588), .B2(REIP_REG_22__SCAN_IN), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5590) );
  NOR2_X1 U6804 ( .A1(n5590), .A2(n5589), .ZN(n5593) );
  AOI22_X1 U6805 ( .A1(n6458), .A2(EBX_REG_23__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6419), .ZN(n5591) );
  OAI21_X1 U6806 ( .B1(n6449), .B2(n5921), .A(n5591), .ZN(n5592) );
  AOI211_X1 U6807 ( .C1(n5594), .C2(n6439), .A(n5593), .B(n5592), .ZN(n5595)
         );
  OAI21_X1 U6808 ( .B1(n5822), .B2(n6424), .A(n5595), .ZN(U2804) );
  AOI21_X1 U6809 ( .B1(n5597), .B2(n5596), .A(n5583), .ZN(n5933) );
  INV_X1 U6810 ( .A(n5933), .ZN(n5825) );
  NAND2_X1 U6811 ( .A1(n5598), .A2(n5599), .ZN(n5600) );
  NAND2_X1 U6812 ( .A1(n3121), .A2(n5600), .ZN(n6139) );
  INV_X1 U6813 ( .A(n6139), .ZN(n5607) );
  INV_X1 U6814 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5783) );
  OAI22_X1 U6815 ( .A1(n6455), .A2(n6980), .B1(n6443), .B2(n5783), .ZN(n5601)
         );
  AOI21_X1 U6816 ( .B1(n6463), .B2(n5930), .A(n5601), .ZN(n5604) );
  NOR3_X1 U6817 ( .A1(n5667), .A2(REIP_REG_21__SCAN_IN), .A3(n5602), .ZN(n5613) );
  OAI21_X1 U6818 ( .B1(n5613), .B2(n3164), .A(REIP_REG_22__SCAN_IN), .ZN(n5603) );
  OAI211_X1 U6819 ( .C1(n5605), .C2(REIP_REG_22__SCAN_IN), .A(n5604), .B(n5603), .ZN(n5606) );
  AOI21_X1 U6820 ( .B1(n5607), .B2(n6439), .A(n5606), .ZN(n5608) );
  OAI21_X1 U6821 ( .B1(n5825), .B2(n6424), .A(n5608), .ZN(U2805) );
  INV_X1 U6822 ( .A(n5609), .ZN(n5622) );
  OAI21_X1 U6823 ( .B1(n5622), .B2(n3138), .A(n5596), .ZN(n5943) );
  OR2_X1 U6824 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  NAND2_X1 U6825 ( .A1(n5598), .A2(n5612), .ZN(n6149) );
  INV_X1 U6826 ( .A(n6149), .ZN(n5619) );
  INV_X1 U6827 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5784) );
  OAI22_X1 U6828 ( .A1(n6455), .A2(n5938), .B1(n6443), .B2(n5784), .ZN(n5614)
         );
  AOI211_X1 U6829 ( .C1(n6463), .C2(n5940), .A(n5614), .B(n5613), .ZN(n5615)
         );
  OAI21_X1 U6830 ( .B1(n5617), .B2(n5616), .A(n5615), .ZN(n5618) );
  AOI21_X1 U6831 ( .B1(n5619), .B2(n6439), .A(n5618), .ZN(n5620) );
  OAI21_X1 U6832 ( .B1(n5943), .B2(n6424), .A(n5620), .ZN(U2806) );
  AOI21_X1 U6833 ( .B1(n5623), .B2(n5621), .A(n5622), .ZN(n5949) );
  INV_X1 U6834 ( .A(n5949), .ZN(n5830) );
  MUX2_X1 U6835 ( .A(n5626), .B(n5625), .S(n5624), .Z(n5628) );
  XNOR2_X1 U6836 ( .A(n5628), .B(n5627), .ZN(n6162) );
  INV_X1 U6837 ( .A(n6162), .ZN(n5633) );
  OAI21_X1 U6838 ( .B1(n5629), .B2(REIP_REG_20__SCAN_IN), .A(n3164), .ZN(n5631) );
  AOI22_X1 U6839 ( .A1(n6458), .A2(EBX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6419), .ZN(n5630) );
  OAI211_X1 U6840 ( .C1(n6449), .C2(n5947), .A(n5631), .B(n5630), .ZN(n5632)
         );
  AOI21_X1 U6841 ( .B1(n5633), .B2(n6439), .A(n5632), .ZN(n5634) );
  OAI21_X1 U6842 ( .B1(n5830), .B2(n6424), .A(n5634), .ZN(U2807) );
  OAI21_X1 U6843 ( .B1(n5635), .B2(n5636), .A(n5621), .ZN(n5956) );
  INV_X1 U6844 ( .A(n5674), .ZN(n5641) );
  INV_X1 U6845 ( .A(n5637), .ZN(n5639) );
  MUX2_X1 U6846 ( .A(n5640), .B(n5639), .S(n5638), .Z(n5658) );
  NAND2_X1 U6847 ( .A1(n5641), .A2(n5658), .ZN(n5661) );
  XOR2_X1 U6848 ( .A(n5642), .B(n5661), .Z(n6169) );
  INV_X1 U6849 ( .A(n5678), .ZN(n5651) );
  NAND2_X1 U6850 ( .A1(n6419), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5643)
         );
  OAI211_X1 U6851 ( .C1(n6443), .C2(n5644), .A(n6430), .B(n5643), .ZN(n5645)
         );
  AOI21_X1 U6852 ( .B1(n6463), .B2(n5959), .A(n5645), .ZN(n5649) );
  INV_X1 U6853 ( .A(n5667), .ZN(n5647) );
  OAI211_X1 U6854 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5647), .B(n5646), .ZN(n5648) );
  OAI211_X1 U6855 ( .C1(n5651), .C2(n5650), .A(n5649), .B(n5648), .ZN(n5652)
         );
  AOI21_X1 U6856 ( .B1(n6169), .B2(n6439), .A(n5652), .ZN(n5653) );
  OAI21_X1 U6857 ( .B1(n5956), .B2(n6424), .A(n5653), .ZN(U2808) );
  INV_X1 U6858 ( .A(n5654), .ZN(n5701) );
  NAND2_X1 U6859 ( .A1(n5700), .A2(n5696), .ZN(n5695) );
  INV_X1 U6860 ( .A(n5655), .ZN(n5671) );
  NOR2_X1 U6861 ( .A1(n5695), .A2(n5671), .ZN(n5670) );
  INV_X1 U6862 ( .A(n5635), .ZN(n5656) );
  OAI21_X1 U6863 ( .B1(n5670), .B2(n5657), .A(n5656), .ZN(n5970) );
  INV_X1 U6864 ( .A(n5658), .ZN(n5659) );
  NAND2_X1 U6865 ( .A1(n5674), .A2(n5659), .ZN(n5660) );
  INV_X1 U6866 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U6867 ( .A1(n6419), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5662)
         );
  OAI211_X1 U6868 ( .C1(n6443), .C2(n5663), .A(n5662), .B(n6430), .ZN(n5664)
         );
  AOI21_X1 U6869 ( .B1(n6463), .B2(n5967), .A(n5664), .ZN(n5666) );
  NAND2_X1 U6870 ( .A1(n5678), .A2(REIP_REG_18__SCAN_IN), .ZN(n5665) );
  OAI211_X1 U6871 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5667), .A(n5666), .B(n5665), .ZN(n5668) );
  AOI21_X1 U6872 ( .B1(n6181), .B2(n6439), .A(n5668), .ZN(n5669) );
  OAI21_X1 U6873 ( .B1(n5970), .B2(n6424), .A(n5669), .ZN(U2809) );
  AOI21_X1 U6874 ( .B1(n5671), .B2(n5695), .A(n5670), .ZN(n5983) );
  NAND2_X1 U6875 ( .A1(n5686), .A2(n5672), .ZN(n5673) );
  NAND2_X1 U6876 ( .A1(n5674), .A2(n5673), .ZN(n6189) );
  INV_X1 U6877 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U6878 ( .A1(n6419), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5675)
         );
  OAI211_X1 U6879 ( .C1(n6443), .C2(n5787), .A(n6430), .B(n5675), .ZN(n5676)
         );
  AOI21_X1 U6880 ( .B1(n6463), .B2(n5978), .A(n5676), .ZN(n5681) );
  NAND2_X1 U6881 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5687) );
  OAI21_X1 U6882 ( .B1(n5709), .B2(n5687), .A(n5677), .ZN(n5679) );
  NAND2_X1 U6883 ( .A1(n5679), .A2(n5678), .ZN(n5680) );
  OAI211_X1 U6884 ( .C1(n6189), .C2(n6452), .A(n5681), .B(n5680), .ZN(n5682)
         );
  AOI21_X1 U6885 ( .B1(n5983), .B2(n6411), .A(n5682), .ZN(n5683) );
  INV_X1 U6886 ( .A(n5683), .ZN(U2810) );
  OR2_X1 U6887 ( .A1(n5705), .A2(n5684), .ZN(n5685) );
  AND2_X1 U6888 ( .A1(n5686), .A2(n5685), .ZN(n6198) );
  OAI21_X1 U6889 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n5687), .ZN(n5694) );
  INV_X1 U6890 ( .A(n5988), .ZN(n5688) );
  NAND2_X1 U6891 ( .A1(n6463), .A2(n5688), .ZN(n5693) );
  INV_X1 U6892 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U6893 ( .A1(n6419), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5689)
         );
  OAI211_X1 U6894 ( .C1(n6443), .C2(n5690), .A(n6430), .B(n5689), .ZN(n5691)
         );
  AOI21_X1 U6895 ( .B1(n5706), .B2(REIP_REG_16__SCAN_IN), .A(n5691), .ZN(n5692) );
  OAI211_X1 U6896 ( .C1(n5709), .C2(n5694), .A(n5693), .B(n5692), .ZN(n5698)
         );
  OAI21_X1 U6897 ( .B1(n5700), .B2(n5696), .A(n5695), .ZN(n5992) );
  NOR2_X1 U6898 ( .A1(n5992), .A2(n6424), .ZN(n5697) );
  AOI211_X1 U6899 ( .C1(n6198), .C2(n6439), .A(n5698), .B(n5697), .ZN(n5699)
         );
  INV_X1 U6900 ( .A(n5699), .ZN(U2811) );
  AOI21_X1 U6901 ( .B1(n5701), .B2(n5495), .A(n5700), .ZN(n5999) );
  INV_X1 U6902 ( .A(n5999), .ZN(n5843) );
  NOR2_X1 U6903 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  OR2_X1 U6904 ( .A1(n5705), .A2(n5704), .ZN(n6206) );
  INV_X1 U6905 ( .A(n6206), .ZN(n5712) );
  NAND2_X1 U6906 ( .A1(n5706), .A2(REIP_REG_15__SCAN_IN), .ZN(n5708) );
  INV_X1 U6907 ( .A(n6430), .ZN(n6407) );
  AOI21_X1 U6908 ( .B1(n6419), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6407), 
        .ZN(n5707) );
  OAI211_X1 U6909 ( .C1(n5789), .C2(n6443), .A(n5708), .B(n5707), .ZN(n5711)
         );
  OAI22_X1 U6910 ( .A1(n6449), .A2(n5997), .B1(REIP_REG_15__SCAN_IN), .B2(
        n5709), .ZN(n5710) );
  AOI211_X1 U6911 ( .C1(n6439), .C2(n5712), .A(n5711), .B(n5710), .ZN(n5713)
         );
  OAI21_X1 U6912 ( .B1(n5843), .B2(n6424), .A(n5713), .ZN(U2812) );
  INV_X1 U6913 ( .A(n5716), .ZN(n5717) );
  AOI21_X1 U6914 ( .B1(n5718), .B2(n5714), .A(n5717), .ZN(n6015) );
  INV_X1 U6915 ( .A(n6015), .ZN(n5846) );
  AOI22_X1 U6916 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6458), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n6419), .ZN(n5730) );
  INV_X1 U6917 ( .A(n6013), .ZN(n5728) );
  NAND2_X1 U6918 ( .A1(n5737), .A2(n5719), .ZN(n5720) );
  NAND2_X1 U6919 ( .A1(n5721), .A2(n5720), .ZN(n6228) );
  INV_X1 U6920 ( .A(n6228), .ZN(n5722) );
  NAND2_X1 U6921 ( .A1(n5722), .A2(n6439), .ZN(n5726) );
  NAND2_X1 U6922 ( .A1(n6394), .A2(REIP_REG_13__SCAN_IN), .ZN(n5725) );
  OAI211_X1 U6923 ( .C1(REIP_REG_13__SCAN_IN), .C2(REIP_REG_12__SCAN_IN), .A(
        n5740), .B(n5723), .ZN(n5724) );
  NAND4_X1 U6924 ( .A1(n5726), .A2(n6430), .A3(n5725), .A4(n5724), .ZN(n5727)
         );
  AOI21_X1 U6925 ( .B1(n6463), .B2(n5728), .A(n5727), .ZN(n5729) );
  OAI211_X1 U6926 ( .C1(n5846), .C2(n6424), .A(n5730), .B(n5729), .ZN(U2814)
         );
  XOR2_X1 U6927 ( .A(n5731), .B(n5473), .Z(n6029) );
  INV_X1 U6928 ( .A(n5732), .ZN(n6027) );
  AOI22_X1 U6929 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6458), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6394), .ZN(n5733) );
  OAI211_X1 U6930 ( .C1(n6455), .C2(n5734), .A(n5733), .B(n6430), .ZN(n5735)
         );
  INV_X1 U6931 ( .A(n5735), .ZN(n5742) );
  OR2_X1 U6932 ( .A1(n6246), .A2(n5736), .ZN(n5738) );
  AND2_X1 U6933 ( .A1(n5738), .A2(n5737), .ZN(n6236) );
  AOI22_X1 U6934 ( .A1(n5740), .A2(n5739), .B1(n6236), .B2(n6439), .ZN(n5741)
         );
  OAI211_X1 U6935 ( .C1(n6449), .C2(n6027), .A(n5742), .B(n5741), .ZN(n5743)
         );
  AOI21_X1 U6936 ( .B1(n6411), .B2(n6029), .A(n5743), .ZN(n5744) );
  INV_X1 U6937 ( .A(n5744), .ZN(U2815) );
  INV_X1 U6938 ( .A(n5745), .ZN(n5747) );
  NAND2_X1 U6939 ( .A1(n5760), .A2(n5761), .ZN(n5746) );
  NOR2_X1 U6940 ( .A1(n5746), .A2(n5747), .ZN(n5796) );
  AOI21_X1 U6941 ( .B1(n5747), .B2(n5746), .A(n5796), .ZN(n6061) );
  INV_X1 U6942 ( .A(n6061), .ZN(n5855) );
  INV_X1 U6943 ( .A(n6059), .ZN(n5758) );
  OR2_X1 U6944 ( .A1(n5749), .A2(n5750), .ZN(n5751) );
  NAND2_X1 U6945 ( .A1(n5748), .A2(n5751), .ZN(n5799) );
  NAND3_X1 U6946 ( .A1(n6389), .A2(n6401), .A3(n5752), .ZN(n5753) );
  OAI21_X1 U6947 ( .B1(n5799), .B2(n6452), .A(n5753), .ZN(n5757) );
  AOI22_X1 U6948 ( .A1(EBX_REG_8__SCAN_IN), .A2(n6458), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n6419), .ZN(n5754) );
  OAI211_X1 U6949 ( .C1(n6405), .C2(n5755), .A(n5754), .B(n6430), .ZN(n5756)
         );
  AOI211_X1 U6950 ( .C1(n6463), .C2(n5758), .A(n5757), .B(n5756), .ZN(n5759)
         );
  OAI21_X1 U6951 ( .B1(n6424), .B2(n5855), .A(n5759), .ZN(U2819) );
  XOR2_X1 U6952 ( .A(n5761), .B(n5760), .Z(n6069) );
  NAND2_X1 U6953 ( .A1(n6069), .A2(n6411), .ZN(n5776) );
  NOR2_X1 U6954 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5762), .ZN(n5769) );
  INV_X1 U6955 ( .A(n5763), .ZN(n6418) );
  INV_X1 U6956 ( .A(n5764), .ZN(n5765) );
  AOI21_X1 U6957 ( .B1(n5294), .B2(n6418), .A(n5765), .ZN(n5766) );
  OR2_X1 U6958 ( .A1(n5749), .A2(n5766), .ZN(n5803) );
  INV_X1 U6959 ( .A(n5803), .ZN(n6606) );
  AOI22_X1 U6960 ( .A1(n6439), .A2(n6606), .B1(n6458), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5767) );
  OAI211_X1 U6961 ( .C1(n6455), .C2(n7159), .A(n5767), .B(n6430), .ZN(n5768)
         );
  AOI21_X1 U6962 ( .B1(n6389), .B2(n5769), .A(n5768), .ZN(n5775) );
  INV_X1 U6963 ( .A(n6067), .ZN(n5770) );
  NAND2_X1 U6964 ( .A1(n6463), .A2(n5770), .ZN(n5774) );
  NAND2_X1 U6965 ( .A1(n6556), .A2(n5771), .ZN(n5772) );
  NOR2_X1 U6966 ( .A1(n6402), .A2(n5772), .ZN(n6416) );
  OAI21_X1 U6967 ( .B1(n6417), .B2(n6416), .A(REIP_REG_7__SCAN_IN), .ZN(n5773)
         );
  NAND4_X1 U6968 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(U2820)
         );
  OAI22_X1 U6969 ( .A1(n5777), .A2(n5802), .B1(n7090), .B2(n6481), .ZN(U2828)
         );
  OAI222_X1 U6970 ( .A1(n5778), .A2(n6481), .B1(n5802), .B2(n6086), .C1(n5869), 
        .C2(n6474), .ZN(U2831) );
  AOI22_X1 U6971 ( .A1(n6103), .A2(n6478), .B1(n4564), .B2(EBX_REG_26__SCAN_IN), .ZN(n5779) );
  OAI21_X1 U6972 ( .B1(n5815), .B2(n6474), .A(n5779), .ZN(U2833) );
  OAI222_X1 U6973 ( .A1(n5780), .A2(n6481), .B1(n5802), .B2(n6114), .C1(n5890), 
        .C2(n6474), .ZN(U2834) );
  INV_X1 U6974 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6924) );
  INV_X1 U6975 ( .A(n6121), .ZN(n5781) );
  OAI222_X1 U6976 ( .A1(n6924), .A2(n6481), .B1(n5802), .B2(n5781), .C1(n5915), 
        .C2(n6474), .ZN(U2835) );
  INV_X1 U6977 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5782) );
  OAI222_X1 U6978 ( .A1(n5782), .A2(n6481), .B1(n5802), .B2(n6129), .C1(n5822), 
        .C2(n6474), .ZN(U2836) );
  OAI222_X1 U6979 ( .A1(n5783), .A2(n6481), .B1(n5802), .B2(n6139), .C1(n5825), 
        .C2(n6474), .ZN(U2837) );
  OAI222_X1 U6980 ( .A1(n5784), .A2(n6481), .B1(n5802), .B2(n6149), .C1(n5943), 
        .C2(n6474), .ZN(U2838) );
  OAI222_X1 U6981 ( .A1(n5802), .A2(n6162), .B1(n6481), .B2(n7141), .C1(n6474), 
        .C2(n5830), .ZN(U2839) );
  AOI22_X1 U6982 ( .A1(n6169), .A2(n6478), .B1(EBX_REG_19__SCAN_IN), .B2(n4564), .ZN(n5785) );
  OAI21_X1 U6983 ( .B1(n5956), .B2(n6474), .A(n5785), .ZN(U2840) );
  AOI22_X1 U6984 ( .A1(n6181), .A2(n6478), .B1(n4564), .B2(EBX_REG_18__SCAN_IN), .ZN(n5786) );
  OAI21_X1 U6985 ( .B1(n5970), .B2(n6474), .A(n5786), .ZN(U2841) );
  INV_X1 U6986 ( .A(n5983), .ZN(n5837) );
  OAI222_X1 U6987 ( .A1(n5787), .A2(n6481), .B1(n5802), .B2(n6189), .C1(n5837), 
        .C2(n6474), .ZN(U2842) );
  AOI22_X1 U6988 ( .A1(n6198), .A2(n6478), .B1(n4564), .B2(EBX_REG_16__SCAN_IN), .ZN(n5788) );
  OAI21_X1 U6989 ( .B1(n5992), .B2(n6474), .A(n5788), .ZN(U2843) );
  OAI222_X1 U6990 ( .A1(n6206), .A2(n5802), .B1(n5789), .B2(n6481), .C1(n5843), 
        .C2(n6474), .ZN(U2844) );
  INV_X1 U6991 ( .A(n6215), .ZN(n5790) );
  OAI222_X1 U6992 ( .A1(n5790), .A2(n5802), .B1(n6977), .B2(n6481), .C1(n6004), 
        .C2(n6474), .ZN(U2845) );
  INV_X1 U6993 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5791) );
  OAI22_X1 U6994 ( .A1(n6228), .A2(n5802), .B1(n5791), .B2(n6481), .ZN(n5792)
         );
  INV_X1 U6995 ( .A(n5792), .ZN(n5793) );
  OAI21_X1 U6996 ( .B1(n5846), .B2(n6474), .A(n5793), .ZN(U2846) );
  INV_X1 U6997 ( .A(n6236), .ZN(n5794) );
  INV_X1 U6998 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6973) );
  INV_X1 U6999 ( .A(n6029), .ZN(n5848) );
  OAI222_X1 U7000 ( .A1(n5794), .A2(n5802), .B1(n6481), .B2(n6973), .C1(n6474), 
        .C2(n5848), .ZN(U2847) );
  OAI21_X1 U7001 ( .B1(n5796), .B2(n5795), .A(n5378), .ZN(n6408) );
  INV_X1 U7002 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5798) );
  OAI21_X1 U7003 ( .B1(n4394), .B2(n3294), .A(n5797), .ZN(n6400) );
  OAI222_X1 U7004 ( .A1(n6408), .A2(n6474), .B1(n6481), .B2(n5798), .C1(n5802), 
        .C2(n6400), .ZN(U2850) );
  INV_X1 U7005 ( .A(n5799), .ZN(n6598) );
  AOI22_X1 U7006 ( .A1(n6478), .A2(n6598), .B1(n4564), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5800) );
  OAI21_X1 U7007 ( .B1(n5855), .B2(n6474), .A(n5800), .ZN(U2851) );
  INV_X1 U7008 ( .A(n6069), .ZN(n5858) );
  INV_X1 U7009 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5801) );
  OAI222_X1 U7010 ( .A1(n5803), .A2(n5802), .B1(n6474), .B2(n5858), .C1(n6481), 
        .C2(n5801), .ZN(U2852) );
  AOI22_X1 U7011 ( .A1(n5838), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n5850), .ZN(n5806) );
  NAND2_X1 U7012 ( .A1(n5839), .A2(DATAI_13_), .ZN(n5805) );
  OAI211_X1 U7013 ( .C1(n5807), .C2(n5859), .A(n5806), .B(n5805), .ZN(U2862)
         );
  AOI22_X1 U7014 ( .A1(n5838), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n5850), .ZN(n5809) );
  NAND2_X1 U7015 ( .A1(n5839), .A2(DATAI_12_), .ZN(n5808) );
  OAI211_X1 U7016 ( .C1(n5869), .C2(n5859), .A(n5809), .B(n5808), .ZN(U2863)
         );
  AOI22_X1 U7017 ( .A1(n5838), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5850), .ZN(n5811) );
  NAND2_X1 U7018 ( .A1(n5839), .A2(DATAI_11_), .ZN(n5810) );
  OAI211_X1 U7019 ( .C1(n5812), .C2(n5859), .A(n5811), .B(n5810), .ZN(U2864)
         );
  AOI22_X1 U7020 ( .A1(n5838), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5850), .ZN(n5814) );
  NAND2_X1 U7021 ( .A1(n5839), .A2(DATAI_10_), .ZN(n5813) );
  OAI211_X1 U7022 ( .C1(n5815), .C2(n5859), .A(n5814), .B(n5813), .ZN(U2865)
         );
  AOI22_X1 U7023 ( .A1(n5838), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n5850), .ZN(n5817) );
  NAND2_X1 U7024 ( .A1(n5839), .A2(DATAI_9_), .ZN(n5816) );
  OAI211_X1 U7025 ( .C1(n5890), .C2(n5859), .A(n5817), .B(n5816), .ZN(U2866)
         );
  AOI22_X1 U7026 ( .A1(n5838), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n5850), .ZN(n5819) );
  NAND2_X1 U7027 ( .A1(n5839), .A2(DATAI_8_), .ZN(n5818) );
  OAI211_X1 U7028 ( .C1(n5915), .C2(n5859), .A(n5819), .B(n5818), .ZN(U2867)
         );
  AOI22_X1 U7029 ( .A1(n5838), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n5850), .ZN(n5821) );
  NAND2_X1 U7030 ( .A1(n5839), .A2(DATAI_7_), .ZN(n5820) );
  OAI211_X1 U7031 ( .C1(n5822), .C2(n5859), .A(n5821), .B(n5820), .ZN(U2868)
         );
  AOI22_X1 U7032 ( .A1(n5838), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n5850), .ZN(n5824) );
  NAND2_X1 U7033 ( .A1(n5839), .A2(DATAI_6_), .ZN(n5823) );
  OAI211_X1 U7034 ( .C1(n5825), .C2(n5859), .A(n5824), .B(n5823), .ZN(U2869)
         );
  AOI22_X1 U7035 ( .A1(n5838), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n5850), .ZN(n5827) );
  NAND2_X1 U7036 ( .A1(n5839), .A2(DATAI_5_), .ZN(n5826) );
  OAI211_X1 U7037 ( .C1(n5943), .C2(n5859), .A(n5827), .B(n5826), .ZN(U2870)
         );
  AOI22_X1 U7038 ( .A1(n5838), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n5850), .ZN(n5829) );
  NAND2_X1 U7039 ( .A1(n5839), .A2(DATAI_4_), .ZN(n5828) );
  OAI211_X1 U7040 ( .C1(n5830), .C2(n5859), .A(n5829), .B(n5828), .ZN(U2871)
         );
  AOI22_X1 U7041 ( .A1(n5838), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n5850), .ZN(n5832) );
  NAND2_X1 U7042 ( .A1(n5839), .A2(DATAI_3_), .ZN(n5831) );
  OAI211_X1 U7043 ( .C1(n5956), .C2(n5859), .A(n5832), .B(n5831), .ZN(U2872)
         );
  AOI22_X1 U7044 ( .A1(n5838), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n5850), .ZN(n5834) );
  NAND2_X1 U7045 ( .A1(n5839), .A2(DATAI_2_), .ZN(n5833) );
  OAI211_X1 U7046 ( .C1(n5970), .C2(n5859), .A(n5834), .B(n5833), .ZN(U2873)
         );
  AOI22_X1 U7047 ( .A1(n5838), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n5850), .ZN(n5836) );
  NAND2_X1 U7048 ( .A1(n5839), .A2(DATAI_1_), .ZN(n5835) );
  OAI211_X1 U7049 ( .C1(n5837), .C2(n5859), .A(n5836), .B(n5835), .ZN(U2874)
         );
  AOI22_X1 U7050 ( .A1(n5838), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n5850), .ZN(n5841) );
  NAND2_X1 U7051 ( .A1(n5839), .A2(DATAI_0_), .ZN(n5840) );
  OAI211_X1 U7052 ( .C1(n5992), .C2(n5859), .A(n5841), .B(n5840), .ZN(U2875)
         );
  AOI22_X1 U7053 ( .A1(n5851), .A2(DATAI_15_), .B1(n5850), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5842) );
  OAI21_X1 U7054 ( .B1(n5843), .B2(n5859), .A(n5842), .ZN(U2876) );
  INV_X1 U7055 ( .A(DATAI_13_), .ZN(n5844) );
  OAI222_X1 U7056 ( .A1(n5846), .A2(n5859), .B1(n5856), .B2(n5845), .C1(n5844), 
        .C2(n5860), .ZN(U2878) );
  OAI222_X1 U7057 ( .A1(n5860), .A2(n5849), .B1(n5859), .B2(n5848), .C1(n5847), 
        .C2(n5856), .ZN(U2879) );
  AOI22_X1 U7058 ( .A1(n5851), .A2(DATAI_9_), .B1(n5850), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5852) );
  OAI21_X1 U7059 ( .B1(n6408), .B2(n5859), .A(n5852), .ZN(U2882) );
  OAI222_X1 U7060 ( .A1(n5855), .A2(n5859), .B1(n5856), .B2(n5854), .C1(n5853), 
        .C2(n5860), .ZN(U2883) );
  OAI222_X1 U7061 ( .A1(n5860), .A2(n4705), .B1(n5859), .B2(n5858), .C1(n5857), 
        .C2(n5856), .ZN(U2884) );
  NOR2_X1 U7062 ( .A1(n6577), .A2(n5861), .ZN(n6088) );
  NOR2_X1 U7063 ( .A1(n5862), .A2(n6586), .ZN(n5863) );
  AOI211_X1 U7064 ( .C1(PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n6578), .A(n6088), 
        .B(n5863), .ZN(n5868) );
  NAND2_X1 U7065 ( .A1(n6116), .A2(n5865), .ZN(n6107) );
  NAND2_X1 U7066 ( .A1(n5885), .A2(n3136), .ZN(n5871) );
  NAND2_X1 U7067 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  XNOR2_X1 U7068 ( .A(n5872), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6102)
         );
  NAND2_X1 U7069 ( .A1(n5873), .A2(n5979), .ZN(n5874) );
  NAND2_X1 U7070 ( .A1(n6566), .A2(REIP_REG_27__SCAN_IN), .ZN(n6095) );
  OAI211_X1 U7071 ( .C1(n5875), .C2(n5981), .A(n5874), .B(n6095), .ZN(n5876)
         );
  AOI21_X1 U7072 ( .B1(n5877), .B2(n6571), .A(n5876), .ZN(n5878) );
  OAI21_X1 U7073 ( .B1(n6102), .B2(n6372), .A(n5878), .ZN(U2959) );
  XNOR2_X1 U7074 ( .A(n6020), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5879)
         );
  NAND2_X1 U7075 ( .A1(n6566), .A2(REIP_REG_26__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7076 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5880)
         );
  OAI211_X1 U7077 ( .C1(n6586), .C2(n5881), .A(n6104), .B(n5880), .ZN(n5882)
         );
  AOI21_X1 U7078 ( .B1(n5883), .B2(n6571), .A(n5882), .ZN(n5884) );
  OAI21_X1 U7079 ( .B1(n6372), .B2(n6111), .A(n5884), .ZN(U2960) );
  INV_X1 U7080 ( .A(n5885), .ZN(n5888) );
  AOI21_X1 U7081 ( .B1(n5888), .B2(n5887), .A(n5886), .ZN(n6119) );
  NAND2_X1 U7082 ( .A1(n6566), .A2(REIP_REG_25__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7083 ( .B1(n5981), .B2(n5889), .A(n6112), .ZN(n5892) );
  NOR2_X1 U7084 ( .A1(n5890), .A2(n6054), .ZN(n5891) );
  AOI211_X1 U7085 ( .C1(n5893), .C2(n5979), .A(n5892), .B(n5891), .ZN(n5894)
         );
  OAI21_X1 U7086 ( .B1(n6119), .B2(n6372), .A(n5894), .ZN(U2961) );
  XNOR2_X1 U7087 ( .A(n6018), .B(n5897), .ZN(n5953) );
  NAND2_X1 U7088 ( .A1(n5896), .A2(n5895), .ZN(n5951) );
  NAND2_X1 U7089 ( .A1(n6020), .A2(n5897), .ZN(n5898) );
  AND2_X2 U7090 ( .A1(n5951), .A2(n5898), .ZN(n5918) );
  XNOR2_X1 U7091 ( .A(n3113), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5944)
         );
  XNOR2_X1 U7092 ( .A(n6018), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5936)
         );
  INV_X1 U7093 ( .A(n5935), .ZN(n5902) );
  INV_X1 U7094 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7095 ( .A1(n3113), .A2(n5926), .ZN(n5925) );
  NOR2_X1 U7096 ( .A1(n5925), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5907)
         );
  INV_X1 U7097 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n7110) );
  AOI21_X1 U7098 ( .B1(n5907), .B2(n7110), .A(n5899), .ZN(n5900) );
  INV_X1 U7099 ( .A(n5900), .ZN(n5901) );
  INV_X1 U7100 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n7048) );
  NOR2_X1 U7101 ( .A1(n3113), .A2(n7048), .ZN(n5905) );
  NAND4_X1 U7102 ( .A1(n5905), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .A4(n7110), .ZN(n5903) );
  OAI21_X1 U7103 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n7110), .A(n5903), 
        .ZN(n5904) );
  NAND3_X1 U7104 ( .A1(n5905), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7105 ( .A1(n5906), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5908) );
  OR2_X1 U7106 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  AND3_X2 U7107 ( .A1(n5911), .A2(n5910), .A3(n5909), .ZN(n6127) );
  AND2_X1 U7108 ( .A1(n6566), .A2(REIP_REG_24__SCAN_IN), .ZN(n6120) );
  AOI21_X1 U7109 ( .B1(n6578), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n6120), 
        .ZN(n5914) );
  OR2_X1 U7110 ( .A1(n6586), .A2(n5912), .ZN(n5913) );
  OAI211_X1 U7111 ( .C1(n5915), .C2(n6054), .A(n5914), .B(n5913), .ZN(n5916)
         );
  INV_X1 U7112 ( .A(n5916), .ZN(n5917) );
  OAI21_X1 U7113 ( .B1(n6127), .B2(n6372), .A(n5917), .ZN(U2962) );
  NAND3_X1 U7114 ( .A1(n6018), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n6142), .ZN(n5919) );
  NAND2_X1 U7115 ( .A1(n6566), .A2(REIP_REG_23__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7116 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5920)
         );
  OAI211_X1 U7117 ( .C1(n6586), .C2(n5921), .A(n6128), .B(n5920), .ZN(n5922)
         );
  AOI21_X1 U7118 ( .B1(n5923), .B2(n6571), .A(n5922), .ZN(n5924) );
  OAI21_X1 U7119 ( .B1(n6136), .B2(n6372), .A(n5924), .ZN(U2963) );
  OAI21_X1 U7120 ( .B1(n3113), .B2(n5926), .A(n5925), .ZN(n5927) );
  NAND2_X1 U7121 ( .A1(n5979), .A2(n5930), .ZN(n5931) );
  NAND2_X1 U7122 ( .A1(n6566), .A2(REIP_REG_22__SCAN_IN), .ZN(n6138) );
  OAI211_X1 U7123 ( .C1(n5981), .C2(n6980), .A(n5931), .B(n6138), .ZN(n5932)
         );
  AOI21_X1 U7124 ( .B1(n5933), .B2(n6571), .A(n5932), .ZN(n5934) );
  OAI21_X1 U7125 ( .B1(n6146), .B2(n6372), .A(n5934), .ZN(U2964) );
  OAI21_X1 U7126 ( .B1(n5937), .B2(n5936), .A(n5935), .ZN(n6147) );
  NAND2_X1 U7127 ( .A1(n6147), .A2(n3784), .ZN(n5942) );
  NAND2_X1 U7128 ( .A1(n6566), .A2(REIP_REG_21__SCAN_IN), .ZN(n6148) );
  OAI21_X1 U7129 ( .B1(n5981), .B2(n5938), .A(n6148), .ZN(n5939) );
  AOI21_X1 U7130 ( .B1(n5979), .B2(n5940), .A(n5939), .ZN(n5941) );
  OAI211_X1 U7131 ( .C1(n6054), .C2(n5943), .A(n5942), .B(n5941), .ZN(U2965)
         );
  XNOR2_X1 U7132 ( .A(n5945), .B(n5944), .ZN(n6168) );
  NAND2_X1 U7133 ( .A1(n6566), .A2(REIP_REG_20__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7134 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5946)
         );
  OAI211_X1 U7135 ( .C1(n6586), .C2(n5947), .A(n6161), .B(n5946), .ZN(n5948)
         );
  AOI21_X1 U7136 ( .B1(n5949), .B2(n6571), .A(n5948), .ZN(n5950) );
  OAI21_X1 U7137 ( .B1(n6168), .B2(n6372), .A(n5950), .ZN(U2966) );
  INV_X1 U7138 ( .A(n5951), .ZN(n5952) );
  AOI21_X1 U7139 ( .B1(n5954), .B2(n5953), .A(n5952), .ZN(n6176) );
  INV_X1 U7140 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7141 ( .A1(n6566), .A2(REIP_REG_19__SCAN_IN), .ZN(n6170) );
  OAI21_X1 U7142 ( .B1(n5981), .B2(n5955), .A(n6170), .ZN(n5958) );
  NOR2_X1 U7143 ( .A1(n5956), .A2(n6054), .ZN(n5957) );
  AOI211_X1 U7144 ( .C1(n5979), .C2(n5959), .A(n5958), .B(n5957), .ZN(n5960)
         );
  OAI21_X1 U7145 ( .B1(n6176), .B2(n6372), .A(n5960), .ZN(U2967) );
  INV_X1 U7146 ( .A(n5961), .ZN(n5962) );
  OAI21_X1 U7147 ( .B1(n3113), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5962), 
        .ZN(n5974) );
  OR2_X1 U7148 ( .A1(n6018), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5985)
         );
  NOR3_X1 U7149 ( .A1(n5963), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5985), 
        .ZN(n5975) );
  NOR2_X1 U7150 ( .A1(n6577), .A2(n5964), .ZN(n6180) );
  NOR2_X1 U7151 ( .A1(n5981), .A2(n5965), .ZN(n5966) );
  AOI211_X1 U7152 ( .C1(n5979), .C2(n5967), .A(n6180), .B(n5966), .ZN(n5968)
         );
  OAI211_X1 U7153 ( .C1(n6054), .C2(n5970), .A(n5969), .B(n5968), .ZN(U2968)
         );
  INV_X1 U7154 ( .A(n5971), .ZN(n5977) );
  NOR2_X1 U7155 ( .A1(n6020), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5973)
         );
  INV_X1 U7156 ( .A(n5985), .ZN(n5972) );
  OAI22_X1 U7157 ( .A1(n5974), .A2(n5973), .B1(n5972), .B2(n6937), .ZN(n5976)
         );
  AOI21_X1 U7158 ( .B1(n5977), .B2(n5976), .A(n5975), .ZN(n6193) );
  NAND2_X1 U7159 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  NAND2_X1 U7160 ( .A1(n6566), .A2(REIP_REG_17__SCAN_IN), .ZN(n6187) );
  OAI211_X1 U7161 ( .C1(n5981), .C2(n7046), .A(n5980), .B(n6187), .ZN(n5982)
         );
  AOI21_X1 U7162 ( .B1(n5983), .B2(n6571), .A(n5982), .ZN(n5984) );
  OAI21_X1 U7163 ( .B1(n6193), .B2(n6372), .A(n5984), .ZN(U2969) );
  OAI21_X1 U7164 ( .B1(n3113), .B2(n7144), .A(n5985), .ZN(n5986) );
  XNOR2_X1 U7165 ( .A(n5961), .B(n5986), .ZN(n6194) );
  NAND2_X1 U7166 ( .A1(n6194), .A2(n3784), .ZN(n5991) );
  NOR2_X1 U7167 ( .A1(n6577), .A2(n5987), .ZN(n6197) );
  NOR2_X1 U7168 ( .A1(n6586), .A2(n5988), .ZN(n5989) );
  AOI211_X1 U7169 ( .C1(n6578), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6197), 
        .B(n5989), .ZN(n5990) );
  OAI211_X1 U7170 ( .C1(n6054), .C2(n5992), .A(n5991), .B(n5990), .ZN(U2970)
         );
  INV_X1 U7171 ( .A(n5963), .ZN(n5994) );
  AOI21_X1 U7172 ( .B1(n5995), .B2(n5993), .A(n5994), .ZN(n6211) );
  NAND2_X1 U7173 ( .A1(n6566), .A2(REIP_REG_15__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7174 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5996)
         );
  OAI211_X1 U7175 ( .C1(n6586), .C2(n5997), .A(n6205), .B(n5996), .ZN(n5998)
         );
  AOI21_X1 U7176 ( .B1(n5999), .B2(n6571), .A(n5998), .ZN(n6000) );
  OAI21_X1 U7177 ( .B1(n6211), .B2(n6372), .A(n6000), .ZN(U2971) );
  XNOR2_X1 U7178 ( .A(n6018), .B(n6002), .ZN(n6003) );
  XNOR2_X1 U7179 ( .A(n6001), .B(n6003), .ZN(n6226) );
  INV_X1 U7180 ( .A(n6004), .ZN(n6008) );
  AND2_X1 U7181 ( .A1(n6566), .A2(REIP_REG_14__SCAN_IN), .ZN(n6214) );
  AOI21_X1 U7182 ( .B1(n6578), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6214), 
        .ZN(n6005) );
  OAI21_X1 U7183 ( .B1(n6006), .B2(n6586), .A(n6005), .ZN(n6007) );
  AOI21_X1 U7184 ( .B1(n6008), .B2(n6571), .A(n6007), .ZN(n6009) );
  OAI21_X1 U7185 ( .B1(n6226), .B2(n6372), .A(n6009), .ZN(U2972) );
  XOR2_X1 U7186 ( .A(n6010), .B(n6011), .Z(n6234) );
  NAND2_X1 U7187 ( .A1(n6566), .A2(REIP_REG_13__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7188 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6012)
         );
  OAI211_X1 U7189 ( .C1(n6586), .C2(n6013), .A(n6227), .B(n6012), .ZN(n6014)
         );
  AOI21_X1 U7190 ( .B1(n6015), .B2(n6571), .A(n6014), .ZN(n6016) );
  OAI21_X1 U7191 ( .B1(n6234), .B2(n6372), .A(n6016), .ZN(U2973) );
  OAI21_X1 U7192 ( .B1(n6018), .B2(n7018), .A(n6017), .ZN(n6025) );
  NOR2_X1 U7193 ( .A1(n6020), .A2(n6593), .ZN(n6049) );
  AOI21_X1 U7194 ( .B1(n6019), .B2(n6047), .A(n6049), .ZN(n6040) );
  NAND2_X1 U7195 ( .A1(n6040), .A2(n6021), .ZN(n6032) );
  OAI21_X1 U7196 ( .B1(n6032), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n3113), 
        .ZN(n6022) );
  OAI21_X1 U7197 ( .B1(n6040), .B2(n6023), .A(n6022), .ZN(n6024) );
  XOR2_X1 U7198 ( .A(n6025), .B(n6024), .Z(n6245) );
  AND2_X1 U7199 ( .A1(n6566), .A2(REIP_REG_12__SCAN_IN), .ZN(n6235) );
  AOI21_X1 U7200 ( .B1(n6578), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6235), 
        .ZN(n6026) );
  OAI21_X1 U7201 ( .B1(n6027), .B2(n6586), .A(n6026), .ZN(n6028) );
  AOI21_X1 U7202 ( .B1(n6029), .B2(n6571), .A(n6028), .ZN(n6030) );
  OAI21_X1 U7203 ( .B1(n6245), .B2(n6372), .A(n6030), .ZN(U2974) );
  INV_X1 U7204 ( .A(n6040), .ZN(n6031) );
  AOI22_X1 U7205 ( .A1(n3113), .A2(n6032), .B1(n6031), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6034) );
  XNOR2_X1 U7206 ( .A(n3710), .B(n6240), .ZN(n6033) );
  XNOR2_X1 U7207 ( .A(n6034), .B(n6033), .ZN(n6258) );
  INV_X1 U7208 ( .A(n6470), .ZN(n6037) );
  NAND2_X1 U7209 ( .A1(n6566), .A2(REIP_REG_11__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7210 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6035)
         );
  OAI211_X1 U7211 ( .C1(n6586), .C2(n6395), .A(n6251), .B(n6035), .ZN(n6036)
         );
  AOI21_X1 U7212 ( .B1(n6037), .B2(n6571), .A(n6036), .ZN(n6038) );
  OAI21_X1 U7213 ( .B1(n6258), .B2(n6372), .A(n6038), .ZN(U2975) );
  XNOR2_X1 U7214 ( .A(n6020), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6039)
         );
  XNOR2_X1 U7215 ( .A(n6040), .B(n6039), .ZN(n6259) );
  NAND2_X1 U7216 ( .A1(n6259), .A2(n3784), .ZN(n6045) );
  NOR2_X1 U7217 ( .A1(n6577), .A2(n6041), .ZN(n6263) );
  NOR2_X1 U7218 ( .A1(n6586), .A2(n6042), .ZN(n6043) );
  AOI211_X1 U7219 ( .C1(n6578), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6263), 
        .B(n6043), .ZN(n6044) );
  OAI211_X1 U7220 ( .C1(n6054), .C2(n6046), .A(n6045), .B(n6044), .ZN(U2976)
         );
  INV_X1 U7221 ( .A(n6047), .ZN(n6048) );
  NOR2_X1 U7222 ( .A1(n6049), .A2(n6048), .ZN(n6050) );
  XOR2_X1 U7223 ( .A(n6050), .B(n6019), .Z(n6590) );
  NAND2_X1 U7224 ( .A1(n6590), .A2(n3784), .ZN(n6053) );
  AND2_X1 U7225 ( .A1(n6566), .A2(REIP_REG_9__SCAN_IN), .ZN(n6587) );
  NOR2_X1 U7226 ( .A1(n6586), .A2(n6409), .ZN(n6051) );
  AOI211_X1 U7227 ( .C1(n6578), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6587), 
        .B(n6051), .ZN(n6052) );
  OAI211_X1 U7228 ( .C1(n6054), .C2(n6408), .A(n6053), .B(n6052), .ZN(U2977)
         );
  OAI21_X1 U7229 ( .B1(n6057), .B2(n6056), .A(n6055), .ZN(n6599) );
  NAND2_X1 U7230 ( .A1(n6566), .A2(REIP_REG_8__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U7231 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6058)
         );
  OAI211_X1 U7232 ( .C1(n6586), .C2(n6059), .A(n6596), .B(n6058), .ZN(n6060)
         );
  AOI21_X1 U7233 ( .B1(n6061), .B2(n6571), .A(n6060), .ZN(n6062) );
  OAI21_X1 U7234 ( .B1(n6599), .B2(n6372), .A(n6062), .ZN(U2978) );
  OAI21_X1 U7235 ( .B1(n6065), .B2(n6064), .A(n6063), .ZN(n6607) );
  NAND2_X1 U7236 ( .A1(n6566), .A2(REIP_REG_7__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U7237 ( .A1(n6578), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6066)
         );
  OAI211_X1 U7238 ( .C1(n6586), .C2(n6067), .A(n6604), .B(n6066), .ZN(n6068)
         );
  AOI21_X1 U7239 ( .B1(n6069), .B2(n6571), .A(n6068), .ZN(n6070) );
  OAI21_X1 U7240 ( .B1(n6372), .B2(n6607), .A(n6070), .ZN(U2979) );
  INV_X1 U7241 ( .A(n6074), .ZN(n6075) );
  OAI21_X1 U7242 ( .B1(n6076), .B2(n6275), .A(n6075), .ZN(U2988) );
  INV_X1 U7243 ( .A(n6077), .ZN(n6083) );
  NOR2_X1 U7244 ( .A1(n6078), .A2(n6082), .ZN(n6081) );
  INV_X1 U7245 ( .A(n6085), .ZN(n6094) );
  NOR2_X1 U7246 ( .A1(n6086), .A2(n6252), .ZN(n6087) );
  AOI211_X1 U7247 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n6100), .A(n6088), .B(n6087), .ZN(n6093) );
  INV_X1 U7248 ( .A(n6097), .ZN(n6091) );
  NAND3_X1 U7249 ( .A1(n6091), .A2(n6090), .A3(n6089), .ZN(n6092) );
  OAI211_X1 U7250 ( .C1(n6094), .C2(n6275), .A(n6093), .B(n6092), .ZN(U2990)
         );
  OAI21_X1 U7251 ( .B1(n6096), .B2(n6252), .A(n6095), .ZN(n6099) );
  NOR2_X1 U7252 ( .A1(n6097), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6098)
         );
  AOI211_X1 U7253 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n6100), .A(n6099), .B(n6098), .ZN(n6101) );
  OAI21_X1 U7254 ( .B1(n6102), .B2(n6275), .A(n6101), .ZN(U2991) );
  INV_X1 U7255 ( .A(n6103), .ZN(n6105) );
  OAI21_X1 U7256 ( .B1(n6105), .B2(n6252), .A(n6104), .ZN(n6106) );
  AOI21_X1 U7257 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n6124), .A(n6106), 
        .ZN(n6110) );
  NAND3_X1 U7258 ( .A1(n6117), .A2(n6108), .A3(n6107), .ZN(n6109) );
  OAI211_X1 U7259 ( .C1(n6111), .C2(n6275), .A(n6110), .B(n6109), .ZN(U2992)
         );
  NAND2_X1 U7260 ( .A1(n6124), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6113) );
  OAI211_X1 U7261 ( .C1(n6114), .C2(n6252), .A(n6113), .B(n6112), .ZN(n6115)
         );
  AOI21_X1 U7262 ( .B1(n6117), .B2(n6116), .A(n6115), .ZN(n6118) );
  OAI21_X1 U7263 ( .B1(n6119), .B2(n6275), .A(n6118), .ZN(U2993) );
  AOI21_X1 U7264 ( .B1(n6121), .B2(n6644), .A(n6120), .ZN(n6126) );
  INV_X1 U7265 ( .A(n6122), .ZN(n6123) );
  OAI211_X1 U7266 ( .C1(n6134), .C2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n6124), .B(n6123), .ZN(n6125) );
  OAI211_X1 U7267 ( .C1(n6127), .C2(n6275), .A(n6126), .B(n6125), .ZN(U2994)
         );
  INV_X1 U7268 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6133) );
  OAI21_X1 U7269 ( .B1(n6129), .B2(n6252), .A(n6128), .ZN(n6132) );
  NOR2_X1 U7270 ( .A1(n6130), .A2(n6133), .ZN(n6131) );
  AOI211_X1 U7271 ( .C1(n6134), .C2(n6133), .A(n6132), .B(n6131), .ZN(n6135)
         );
  OAI21_X1 U7272 ( .B1(n6136), .B2(n6275), .A(n6135), .ZN(U2995) );
  INV_X1 U7273 ( .A(n6137), .ZN(n6151) );
  OAI21_X1 U7274 ( .B1(n6139), .B2(n6252), .A(n6138), .ZN(n6144) );
  INV_X1 U7275 ( .A(n6140), .ZN(n6154) );
  NOR3_X1 U7276 ( .A1(n6154), .A2(n6142), .A3(n6141), .ZN(n6143) );
  AOI211_X1 U7277 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n6151), .A(n6144), .B(n6143), .ZN(n6145) );
  OAI21_X1 U7278 ( .B1(n6146), .B2(n6275), .A(n6145), .ZN(U2996) );
  NAND2_X1 U7279 ( .A1(n6147), .A2(n6649), .ZN(n6153) );
  OAI21_X1 U7280 ( .B1(n6149), .B2(n6252), .A(n6148), .ZN(n6150) );
  AOI21_X1 U7281 ( .B1(n6151), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6150), 
        .ZN(n6152) );
  OAI211_X1 U7282 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n6154), .A(n6153), .B(n6152), .ZN(U2997) );
  INV_X1 U7283 ( .A(n6269), .ZN(n6160) );
  OAI21_X1 U7284 ( .B1(n6156), .B2(n6937), .A(n6155), .ZN(n6158) );
  NAND2_X1 U7285 ( .A1(n6158), .A2(n6157), .ZN(n6191) );
  NOR2_X1 U7286 ( .A1(n6239), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6159)
         );
  NOR2_X1 U7287 ( .A1(n6191), .A2(n6159), .ZN(n6185) );
  OAI21_X1 U7288 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6160), .A(n6185), 
        .ZN(n6174) );
  OAI21_X1 U7289 ( .B1(n6162), .B2(n6252), .A(n6161), .ZN(n6166) );
  NOR3_X1 U7290 ( .A1(n6172), .A2(n6164), .A3(n6163), .ZN(n6165) );
  AOI211_X1 U7291 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n6174), .A(n6166), .B(n6165), .ZN(n6167) );
  OAI21_X1 U7292 ( .B1(n6168), .B2(n6275), .A(n6167), .ZN(U2998) );
  NAND2_X1 U7293 ( .A1(n6169), .A2(n6644), .ZN(n6171) );
  OAI211_X1 U7294 ( .C1(n6172), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n6171), .B(n6170), .ZN(n6173) );
  AOI21_X1 U7295 ( .B1(n6174), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n6173), 
        .ZN(n6175) );
  OAI21_X1 U7296 ( .B1(n6176), .B2(n6275), .A(n6175), .ZN(U2999) );
  NAND2_X1 U7297 ( .A1(n6177), .A2(n6649), .ZN(n6183) );
  NOR2_X1 U7298 ( .A1(n6178), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6179)
         );
  AOI211_X1 U7299 ( .C1(n6644), .C2(n6181), .A(n6180), .B(n6179), .ZN(n6182)
         );
  OAI211_X1 U7300 ( .C1(n6185), .C2(n6184), .A(n6183), .B(n6182), .ZN(U3000)
         );
  NAND2_X1 U7301 ( .A1(n6186), .A2(n6937), .ZN(n6188) );
  OAI211_X1 U7302 ( .C1(n6252), .C2(n6189), .A(n6188), .B(n6187), .ZN(n6190)
         );
  AOI21_X1 U7303 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6191), .A(n6190), 
        .ZN(n6192) );
  OAI21_X1 U7304 ( .B1(n6193), .B2(n6275), .A(n6192), .ZN(U3001) );
  INV_X1 U7305 ( .A(n6194), .ZN(n6204) );
  INV_X1 U7306 ( .A(n6239), .ZN(n6195) );
  NOR4_X1 U7307 ( .A1(n6253), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6200), 
        .A4(n7117), .ZN(n6196) );
  AOI211_X1 U7308 ( .C1(n6644), .C2(n6198), .A(n6197), .B(n6196), .ZN(n6203)
         );
  NOR3_X1 U7309 ( .A1(n6253), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n6200), 
        .ZN(n6207) );
  OAI22_X1 U7310 ( .A1(n6220), .A2(n6267), .B1(n6199), .B2(n6266), .ZN(n6256)
         );
  AND2_X1 U7311 ( .A1(n6269), .A2(n6200), .ZN(n6201) );
  OR2_X1 U7312 ( .A1(n6256), .A2(n6201), .ZN(n6209) );
  OAI21_X1 U7313 ( .B1(n6207), .B2(n6209), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n6202) );
  OAI211_X1 U7314 ( .C1(n6204), .C2(n6275), .A(n6203), .B(n6202), .ZN(U3002)
         );
  OAI21_X1 U7315 ( .B1(n6206), .B2(n6252), .A(n6205), .ZN(n6208) );
  AOI211_X1 U7316 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n6209), .A(n6208), .B(n6207), .ZN(n6210) );
  OAI21_X1 U7317 ( .B1(n6211), .B2(n6275), .A(n6210), .ZN(U3003) );
  INV_X1 U7318 ( .A(n6217), .ZN(n6212) );
  NOR3_X1 U7319 ( .A1(n6253), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n6212), 
        .ZN(n6213) );
  AOI211_X1 U7320 ( .C1(n6644), .C2(n6215), .A(n6214), .B(n6213), .ZN(n6225)
         );
  OAI22_X1 U7321 ( .A1(n6218), .A2(n6217), .B1(n6237), .B2(n6216), .ZN(n6219)
         );
  OR2_X1 U7322 ( .A1(n6256), .A2(n6219), .ZN(n6232) );
  INV_X1 U7323 ( .A(n6220), .ZN(n6222) );
  NAND2_X1 U7324 ( .A1(n6237), .A2(n7166), .ZN(n6229) );
  AOI21_X1 U7325 ( .B1(n6222), .B2(n6221), .A(n6229), .ZN(n6223) );
  OAI21_X1 U7326 ( .B1(n6232), .B2(n6223), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n6224) );
  OAI211_X1 U7327 ( .C1(n6226), .C2(n6275), .A(n6225), .B(n6224), .ZN(U3004)
         );
  OAI21_X1 U7328 ( .B1(n6228), .B2(n6252), .A(n6227), .ZN(n6231) );
  NOR2_X1 U7329 ( .A1(n6253), .A2(n6229), .ZN(n6230) );
  AOI211_X1 U7330 ( .C1(INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n6232), .A(n6231), .B(n6230), .ZN(n6233) );
  OAI21_X1 U7331 ( .B1(n6234), .B2(n6275), .A(n6233), .ZN(U3005) );
  AOI21_X1 U7332 ( .B1(n6236), .B2(n6644), .A(n6235), .ZN(n6244) );
  AOI21_X1 U7333 ( .B1(n6239), .B2(n6238), .A(n6237), .ZN(n6242) );
  OAI21_X1 U7334 ( .B1(n6253), .B2(n6240), .A(n7018), .ZN(n6241) );
  OAI21_X1 U7335 ( .B1(n6242), .B2(n6256), .A(n6241), .ZN(n6243) );
  OAI211_X1 U7336 ( .C1(n6245), .C2(n6275), .A(n6244), .B(n6243), .ZN(U3006)
         );
  INV_X1 U7337 ( .A(n6246), .ZN(n6250) );
  NAND2_X1 U7338 ( .A1(n6248), .A2(n6247), .ZN(n6249) );
  NAND2_X1 U7339 ( .A1(n6250), .A2(n6249), .ZN(n6469) );
  OAI21_X1 U7340 ( .B1(n6469), .B2(n6252), .A(n6251), .ZN(n6255) );
  NOR2_X1 U7341 ( .A1(n6253), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6254)
         );
  AOI211_X1 U7342 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6256), .A(n6255), .B(n6254), .ZN(n6257) );
  OAI21_X1 U7343 ( .B1(n6258), .B2(n6275), .A(n6257), .ZN(U3007) );
  INV_X1 U7344 ( .A(n6259), .ZN(n6276) );
  INV_X1 U7345 ( .A(n6260), .ZN(n6264) );
  AOI21_X1 U7346 ( .B1(n6646), .B2(n6651), .A(n6645), .ZN(n6634) );
  NOR2_X1 U7347 ( .A1(n6634), .A2(n6261), .ZN(n6616) );
  NAND2_X1 U7348 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6616), .ZN(n6612)
         );
  NOR4_X1 U7349 ( .A1(n6595), .A2(n6593), .A3(INSTADDRPOINTER_REG_10__SCAN_IN), 
        .A4(n6612), .ZN(n6262) );
  AOI211_X1 U7350 ( .C1(n6644), .C2(n6264), .A(n6263), .B(n6262), .ZN(n6274)
         );
  OAI22_X1 U7351 ( .A1(n6268), .A2(n6267), .B1(n6266), .B2(n6265), .ZN(n6608)
         );
  AOI21_X1 U7352 ( .B1(n6595), .B2(n6269), .A(n6608), .ZN(n6594) );
  INV_X1 U7353 ( .A(n6594), .ZN(n6272) );
  INV_X1 U7354 ( .A(n6612), .ZN(n6270) );
  NAND2_X1 U7355 ( .A1(n6593), .A2(n6270), .ZN(n6271) );
  NOR2_X1 U7356 ( .A1(n6271), .A2(n6595), .ZN(n6589) );
  OAI21_X1 U7357 ( .B1(n6272), .B2(n6589), .A(INSTADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n6273) );
  OAI211_X1 U7358 ( .C1(n6276), .C2(n6275), .A(n6274), .B(n6273), .ZN(U3008)
         );
  OAI211_X1 U7359 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6278), .A(n6277), .B(
        n6304), .ZN(n6279) );
  OAI21_X1 U7360 ( .B1(n6291), .B2(n6280), .A(n6279), .ZN(n6281) );
  MUX2_X1 U7361 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n6281), .S(n6656), 
        .Z(U3464) );
  XNOR2_X1 U7362 ( .A(n6283), .B(n6282), .ZN(n6285) );
  OAI22_X1 U7363 ( .A1(n6285), .A2(n6722), .B1(n6284), .B2(n6291), .ZN(n6286)
         );
  MUX2_X1 U7364 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n6286), .S(n6656), 
        .Z(U3463) );
  INV_X1 U7365 ( .A(n6287), .ZN(n6293) );
  NOR3_X1 U7366 ( .A1(n6290), .A2(n6289), .A3(n6288), .ZN(n6292) );
  OAI222_X1 U7367 ( .A1(n6307), .A2(n6293), .B1(n6722), .B2(n6292), .C1(n6291), 
        .C2(n6453), .ZN(n6294) );
  MUX2_X1 U7368 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n6294), .S(n6656), 
        .Z(U3462) );
  INV_X1 U7369 ( .A(n6295), .ZN(n6298) );
  OAI22_X1 U7370 ( .A1(n6298), .A2(n6297), .B1(n6296), .B2(n6349), .ZN(n6300)
         );
  MUX2_X1 U7371 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6300), .S(n6299), 
        .Z(U3456) );
  INV_X1 U7372 ( .A(n6310), .ZN(n6305) );
  INV_X1 U7373 ( .A(n6301), .ZN(n6302) );
  NOR2_X1 U7374 ( .A1(n6302), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6712)
         );
  AOI22_X1 U7375 ( .A1(n6305), .A2(n6304), .B1(n6303), .B2(n6712), .ZN(n6339)
         );
  INV_X1 U7376 ( .A(n6661), .ZN(n6720) );
  NOR2_X1 U7377 ( .A1(n6306), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6337)
         );
  OAI21_X1 U7378 ( .B1(n6308), .B2(n6341), .A(n6307), .ZN(n6309) );
  AOI21_X1 U7379 ( .B1(n6310), .B2(n6309), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6312) );
  AOI22_X1 U7380 ( .A1(n6720), .A2(n6337), .B1(INSTQUEUE_REG_2__0__SCAN_IN), 
        .B2(n6336), .ZN(n6313) );
  OAI21_X1 U7381 ( .B1(n6339), .B2(n6717), .A(n6313), .ZN(n6314) );
  AOI21_X1 U7382 ( .B1(n6341), .B2(n6663), .A(n6314), .ZN(n6315) );
  OAI21_X1 U7383 ( .B1(n6344), .B2(n6316), .A(n6315), .ZN(U3036) );
  INV_X1 U7384 ( .A(n6770), .ZN(n6735) );
  AOI22_X1 U7385 ( .A1(n6735), .A2(n6337), .B1(INSTQUEUE_REG_2__1__SCAN_IN), 
        .B2(n6336), .ZN(n6317) );
  OAI21_X1 U7386 ( .B1(n6339), .B2(n6678), .A(n6317), .ZN(n6318) );
  AOI21_X1 U7387 ( .B1(n6341), .B2(n6675), .A(n6318), .ZN(n6319) );
  OAI21_X1 U7388 ( .B1(n6344), .B2(n6776), .A(n6319), .ZN(U3037) );
  INV_X1 U7389 ( .A(n6777), .ZN(n6739) );
  AOI22_X1 U7390 ( .A1(n6739), .A2(n6337), .B1(INSTQUEUE_REG_2__2__SCAN_IN), 
        .B2(n6336), .ZN(n6320) );
  OAI21_X1 U7391 ( .B1(n6339), .B2(n6683), .A(n6320), .ZN(n6321) );
  AOI21_X1 U7392 ( .B1(n6341), .B2(n6680), .A(n6321), .ZN(n6322) );
  OAI21_X1 U7393 ( .B1(n6344), .B2(n6783), .A(n6322), .ZN(U3038) );
  INV_X1 U7394 ( .A(n6784), .ZN(n6743) );
  AOI22_X1 U7395 ( .A1(n6743), .A2(n6337), .B1(INSTQUEUE_REG_2__3__SCAN_IN), 
        .B2(n6336), .ZN(n6323) );
  OAI21_X1 U7396 ( .B1(n6339), .B2(n6688), .A(n6323), .ZN(n6324) );
  AOI21_X1 U7397 ( .B1(n6341), .B2(n6685), .A(n6324), .ZN(n6325) );
  OAI21_X1 U7398 ( .B1(n6344), .B2(n6790), .A(n6325), .ZN(U3039) );
  AOI22_X1 U7399 ( .A1(n3191), .A2(n6337), .B1(INSTQUEUE_REG_2__4__SCAN_IN), 
        .B2(n6336), .ZN(n6326) );
  OAI21_X1 U7400 ( .B1(n6339), .B2(n6860), .A(n6326), .ZN(n6327) );
  AOI21_X1 U7401 ( .B1(n6341), .B2(n6690), .A(n6327), .ZN(n6328) );
  OAI21_X1 U7402 ( .B1(n6344), .B2(n6329), .A(n6328), .ZN(U3040) );
  INV_X1 U7403 ( .A(n6791), .ZN(n6750) );
  AOI22_X1 U7404 ( .A1(n6750), .A2(n6337), .B1(INSTQUEUE_REG_2__5__SCAN_IN), 
        .B2(n6336), .ZN(n6330) );
  OAI21_X1 U7405 ( .B1(n6339), .B2(n6697), .A(n6330), .ZN(n6331) );
  AOI21_X1 U7406 ( .B1(n6341), .B2(n6694), .A(n6331), .ZN(n6332) );
  OAI21_X1 U7407 ( .B1(n6344), .B2(n6797), .A(n6332), .ZN(U3041) );
  INV_X1 U7408 ( .A(n6799), .ZN(n6754) );
  AOI22_X1 U7409 ( .A1(n6754), .A2(n6337), .B1(INSTQUEUE_REG_2__6__SCAN_IN), 
        .B2(n6336), .ZN(n6333) );
  OAI21_X1 U7410 ( .B1(n6339), .B2(n6702), .A(n6333), .ZN(n6334) );
  AOI21_X1 U7411 ( .B1(n6341), .B2(n6699), .A(n6334), .ZN(n6335) );
  OAI21_X1 U7412 ( .B1(n6344), .B2(n6808), .A(n6335), .ZN(U3042) );
  INV_X1 U7413 ( .A(n6704), .ZN(n6760) );
  AOI22_X1 U7414 ( .A1(n6760), .A2(n6337), .B1(INSTQUEUE_REG_2__7__SCAN_IN), 
        .B2(n6336), .ZN(n6338) );
  OAI21_X1 U7415 ( .B1(n6339), .B2(n6758), .A(n6338), .ZN(n6340) );
  AOI21_X1 U7416 ( .B1(n6341), .B2(n6706), .A(n6340), .ZN(n6342) );
  OAI21_X1 U7417 ( .B1(n6344), .B2(n6343), .A(n6342), .ZN(U3043) );
  AOI21_X1 U7418 ( .B1(READY_N), .B2(n6345), .A(n6364), .ZN(n6358) );
  AND2_X1 U7419 ( .A1(n6346), .A2(n6358), .ZN(n6351) );
  OAI21_X1 U7420 ( .B1(n6349), .B2(n6348), .A(n6347), .ZN(n6350) );
  MUX2_X1 U7421 ( .A(n6351), .B(n6350), .S(n6938), .Z(n6353) );
  OAI211_X1 U7422 ( .C1(n6354), .C2(n6365), .A(n6353), .B(n6352), .ZN(U3148)
         );
  NOR2_X1 U7423 ( .A1(n6938), .A2(READY_N), .ZN(n6356) );
  AOI21_X1 U7424 ( .B1(n6357), .B2(n6356), .A(n6355), .ZN(n6363) );
  OR3_X1 U7425 ( .A1(n6360), .A2(n6359), .A3(n6358), .ZN(n6361) );
  OAI211_X1 U7426 ( .C1(n6364), .C2(n6363), .A(n6362), .B(n6361), .ZN(U3149)
         );
  AND2_X1 U7427 ( .A1(n6497), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NAND2_X1 U7428 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6844), .ZN(n6368) );
  OAI21_X1 U7429 ( .B1(n6366), .B2(n6365), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6367) );
  OAI21_X1 U7430 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6368), .A(n6367), .ZN(
        U2790) );
  NOR2_X1 U7431 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6370) );
  OAI21_X1 U7432 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6370), .A(n6849), .ZN(n6369)
         );
  OAI21_X1 U7433 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6849), .A(n6369), .ZN(
        U2791) );
  OAI21_X1 U7434 ( .B1(n6370), .B2(BS16_N), .A(n6829), .ZN(n6827) );
  OAI21_X1 U7435 ( .B1(n6829), .B2(n6371), .A(n6827), .ZN(U2792) );
  OAI21_X1 U7436 ( .B1(n6374), .B2(n6373), .A(n6372), .ZN(U2793) );
  NOR4_X1 U7437 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6375) );
  INV_X1 U7438 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n7045) );
  NAND2_X1 U7439 ( .A1(n6375), .A2(n7045), .ZN(n6997) );
  INV_X1 U7440 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n7080) );
  INV_X1 U7441 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n7084) );
  NAND2_X1 U7442 ( .A1(n7080), .A2(n7084), .ZN(n6995) );
  AOI211_X1 U7443 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_9__SCAN_IN), .B(n6995), 
        .ZN(n6376) );
  INV_X1 U7444 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6978) );
  INV_X1 U7445 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6915) );
  NAND3_X1 U7446 ( .A1(n6376), .A2(n6978), .A3(n6915), .ZN(n6383) );
  OR4_X1 U7447 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(
        n6382) );
  NOR4_X1 U7448 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n6380) );
  NOR4_X1 U7449 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(
        DATAWIDTH_REG_6__SCAN_IN), .ZN(n6379) );
  NOR4_X1 U7450 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n6378) );
  NOR4_X1 U7451 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6377) );
  NAND4_X1 U7452 ( .A1(n6380), .A2(n6379), .A3(n6378), .A4(n6377), .ZN(n6381)
         );
  INV_X1 U7453 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6824) );
  NOR3_X1 U7454 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6385) );
  OAI21_X1 U7455 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6385), .A(n6833), .ZN(n6384)
         );
  OAI21_X1 U7456 ( .B1(n6833), .B2(n6824), .A(n6384), .ZN(U2794) );
  INV_X1 U7457 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6828) );
  AOI21_X1 U7458 ( .B1(n6926), .B2(n6828), .A(n6385), .ZN(n6386) );
  INV_X1 U7459 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6912) );
  INV_X1 U7460 ( .A(n6833), .ZN(n6835) );
  AOI22_X1 U7461 ( .A1(n6833), .A2(n6386), .B1(n6912), .B2(n6835), .ZN(U2795)
         );
  INV_X1 U7462 ( .A(n6469), .ZN(n6391) );
  AND3_X1 U7463 ( .A1(n6389), .A2(n6388), .A3(n6387), .ZN(n6390) );
  AOI21_X1 U7464 ( .B1(n6391), .B2(n6439), .A(n6390), .ZN(n6399) );
  INV_X1 U7465 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6473) );
  OAI22_X1 U7466 ( .A1(n6473), .A2(n6443), .B1(n6392), .B2(n6455), .ZN(n6393)
         );
  AOI211_X1 U7467 ( .C1(REIP_REG_11__SCAN_IN), .C2(n6394), .A(n6407), .B(n6393), .ZN(n6398) );
  OAI22_X1 U7468 ( .A1(n6470), .A2(n6424), .B1(n6395), .B2(n6449), .ZN(n6396)
         );
  INV_X1 U7469 ( .A(n6396), .ZN(n6397) );
  NAND3_X1 U7470 ( .A1(n6399), .A2(n6398), .A3(n6397), .ZN(U2816) );
  INV_X1 U7471 ( .A(n6400), .ZN(n6588) );
  NOR3_X1 U7472 ( .A1(n6402), .A2(n6401), .A3(REIP_REG_9__SCAN_IN), .ZN(n6403)
         );
  AOI21_X1 U7473 ( .B1(n6588), .B2(n6439), .A(n6403), .ZN(n6415) );
  OAI22_X1 U7474 ( .A1(n6405), .A2(n6404), .B1(n7025), .B2(n6455), .ZN(n6406)
         );
  AOI211_X1 U7475 ( .C1(n6458), .C2(EBX_REG_9__SCAN_IN), .A(n6407), .B(n6406), 
        .ZN(n6414) );
  INV_X1 U7476 ( .A(n6408), .ZN(n6412) );
  INV_X1 U7477 ( .A(n6409), .ZN(n6410) );
  AOI22_X1 U7478 ( .A1(n6412), .A2(n6411), .B1(n6410), .B2(n6463), .ZN(n6413)
         );
  NAND3_X1 U7479 ( .A1(n6415), .A2(n6414), .A3(n6413), .ZN(U2818) );
  INV_X1 U7480 ( .A(EBX_REG_6__SCAN_IN), .ZN(n7130) );
  AOI21_X1 U7481 ( .B1(n6417), .B2(REIP_REG_6__SCAN_IN), .A(n6416), .ZN(n6427)
         );
  INV_X1 U7482 ( .A(n6565), .ZN(n6422) );
  XNOR2_X1 U7483 ( .A(n5294), .B(n6418), .ZN(n6613) );
  NAND2_X1 U7484 ( .A1(n6419), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6420)
         );
  OAI211_X1 U7485 ( .C1(n6452), .C2(n6613), .A(n6430), .B(n6420), .ZN(n6421)
         );
  AOI21_X1 U7486 ( .B1(n6463), .B2(n6422), .A(n6421), .ZN(n6423) );
  OAI21_X1 U7487 ( .B1(n6561), .B2(n6424), .A(n6423), .ZN(n6425) );
  INV_X1 U7488 ( .A(n6425), .ZN(n6426) );
  OAI211_X1 U7489 ( .C1(n7130), .C2(n6443), .A(n6427), .B(n6426), .ZN(U2821)
         );
  XNOR2_X1 U7490 ( .A(n6429), .B(n6428), .ZN(n6623) );
  OAI21_X1 U7491 ( .B1(n6455), .B2(n6431), .A(n6430), .ZN(n6438) );
  AND3_X1 U7492 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U7493 ( .A1(n6433), .A2(n6432), .ZN(n6434) );
  NAND2_X1 U7494 ( .A1(n6435), .A2(n6434), .ZN(n6468) );
  NOR2_X1 U7495 ( .A1(n6468), .A2(n6436), .ZN(n6437) );
  AOI211_X1 U7496 ( .C1(n6439), .C2(n6623), .A(n6438), .B(n6437), .ZN(n6448)
         );
  NAND2_X1 U7497 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n6440) );
  NOR3_X1 U7498 ( .A1(n6441), .A2(REIP_REG_4__SCAN_IN), .A3(n6440), .ZN(n6445)
         );
  INV_X1 U7499 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6952) );
  OAI22_X1 U7500 ( .A1(n6952), .A2(n6443), .B1(n6454), .B2(n6442), .ZN(n6444)
         );
  AOI211_X1 U7501 ( .C1(n6572), .C2(n6446), .A(n6445), .B(n6444), .ZN(n6447)
         );
  OAI211_X1 U7502 ( .C1(n6575), .C2(n6449), .A(n6448), .B(n6447), .ZN(U2823)
         );
  INV_X1 U7503 ( .A(n6450), .ZN(n6451) );
  NAND2_X1 U7504 ( .A1(n6451), .A2(REIP_REG_2__SCAN_IN), .ZN(n6466) );
  NOR2_X1 U7505 ( .A1(n6452), .A2(n6630), .ZN(n6457) );
  OAI22_X1 U7506 ( .A1(n6455), .A2(n7064), .B1(n6454), .B2(n6453), .ZN(n6456)
         );
  AOI211_X1 U7507 ( .C1(n6458), .C2(EBX_REG_3__SCAN_IN), .A(n6457), .B(n6456), 
        .ZN(n6459) );
  OAI21_X1 U7508 ( .B1(n6461), .B2(n6460), .A(n6459), .ZN(n6462) );
  AOI21_X1 U7509 ( .B1(n6464), .B2(n6463), .A(n6462), .ZN(n6465) );
  OAI221_X1 U7510 ( .B1(n6468), .B2(n6467), .C1(n6468), .C2(n6466), .A(n6465), 
        .ZN(U2824) );
  OAI22_X1 U7511 ( .A1(n6470), .A2(n6474), .B1(n5802), .B2(n6469), .ZN(n6471)
         );
  INV_X1 U7512 ( .A(n6471), .ZN(n6472) );
  OAI21_X1 U7513 ( .B1(n6473), .B2(n6481), .A(n6472), .ZN(U2848) );
  OAI22_X1 U7514 ( .A1(n6561), .A2(n6474), .B1(n6613), .B2(n5802), .ZN(n6475)
         );
  INV_X1 U7515 ( .A(n6475), .ZN(n6476) );
  OAI21_X1 U7516 ( .B1(n7130), .B2(n6481), .A(n6476), .ZN(U2853) );
  AOI22_X1 U7517 ( .A1(n6572), .A2(n6479), .B1(n6478), .B2(n6623), .ZN(n6477)
         );
  OAI21_X1 U7518 ( .B1(n6952), .B2(n6481), .A(n6477), .ZN(U2855) );
  AOI22_X1 U7519 ( .A1(n6582), .A2(n6479), .B1(n6478), .B2(n6643), .ZN(n6480)
         );
  OAI21_X1 U7520 ( .B1(n7066), .B2(n6481), .A(n6480), .ZN(U2857) );
  INV_X1 U7521 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n6891) );
  AOI22_X1 U7522 ( .A1(n6482), .A2(EAX_REG_29__SCAN_IN), .B1(n6839), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n6483) );
  OAI21_X1 U7523 ( .B1(n6891), .B2(n6492), .A(n6483), .ZN(U2894) );
  INV_X1 U7524 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6485) );
  AOI22_X1 U7525 ( .A1(n6497), .A2(DATAO_REG_15__SCAN_IN), .B1(n6839), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6484) );
  OAI21_X1 U7526 ( .B1(n6485), .B2(n6500), .A(n6484), .ZN(U2908) );
  AOI22_X1 U7527 ( .A1(n6497), .A2(DATAO_REG_13__SCAN_IN), .B1(n6839), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6486) );
  OAI21_X1 U7528 ( .B1(n5845), .B2(n6500), .A(n6486), .ZN(U2910) );
  INV_X1 U7529 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6488) );
  AOI22_X1 U7530 ( .A1(n6497), .A2(DATAO_REG_10__SCAN_IN), .B1(n6839), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6487) );
  OAI21_X1 U7531 ( .B1(n6488), .B2(n6500), .A(n6487), .ZN(U2913) );
  INV_X1 U7532 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n6896) );
  AOI22_X1 U7533 ( .A1(n6490), .A2(EAX_REG_9__SCAN_IN), .B1(n6839), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6489) );
  OAI21_X1 U7534 ( .B1(n6896), .B2(n6492), .A(n6489), .ZN(U2914) );
  INV_X1 U7535 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n7092) );
  AOI22_X1 U7536 ( .A1(n6490), .A2(EAX_REG_7__SCAN_IN), .B1(n6839), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n6491) );
  OAI21_X1 U7537 ( .B1(n7092), .B2(n6492), .A(n6491), .ZN(U2916) );
  AOI22_X1 U7538 ( .A1(n6497), .A2(DATAO_REG_6__SCAN_IN), .B1(n6839), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n6493) );
  OAI21_X1 U7539 ( .B1(n6494), .B2(n6500), .A(n6493), .ZN(U2917) );
  AOI22_X1 U7540 ( .A1(n6497), .A2(DATAO_REG_5__SCAN_IN), .B1(n6839), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n6495) );
  OAI21_X1 U7541 ( .B1(n6546), .B2(n6500), .A(n6495), .ZN(U2918) );
  AOI22_X1 U7542 ( .A1(n6497), .A2(DATAO_REG_4__SCAN_IN), .B1(n6839), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n6496) );
  OAI21_X1 U7543 ( .B1(n6975), .B2(n6500), .A(n6496), .ZN(U2919) );
  AOI22_X1 U7544 ( .A1(n6497), .A2(DATAO_REG_3__SCAN_IN), .B1(n6839), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n6498) );
  OAI21_X1 U7545 ( .B1(n7160), .B2(n6500), .A(n6498), .ZN(U2920) );
  INV_X1 U7546 ( .A(EAX_REG_0__SCAN_IN), .ZN(n7078) );
  AOI22_X1 U7547 ( .A1(n6497), .A2(DATAO_REG_0__SCAN_IN), .B1(n6839), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n6499) );
  OAI21_X1 U7548 ( .B1(n7078), .B2(n6500), .A(n6499), .ZN(U2923) );
  INV_X1 U7549 ( .A(DATAI_0_), .ZN(n6501) );
  NOR2_X1 U7550 ( .A1(n6516), .A2(n6501), .ZN(n6535) );
  AOI21_X1 U7551 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6549), .A(n6535), .ZN(n6502) );
  OAI21_X1 U7552 ( .B1(n4013), .B2(n6545), .A(n6502), .ZN(U2924) );
  INV_X1 U7553 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6506) );
  INV_X1 U7554 ( .A(DATAI_1_), .ZN(n6504) );
  NOR2_X1 U7555 ( .A1(n6516), .A2(n6504), .ZN(n6537) );
  AOI21_X1 U7556 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6553), .A(n6537), .ZN(n6505) );
  OAI21_X1 U7557 ( .B1(n6506), .B2(n6545), .A(n6505), .ZN(U2925) );
  AOI21_X1 U7558 ( .B1(UWORD_REG_2__SCAN_IN), .B2(n6553), .A(n6507), .ZN(n6508) );
  OAI21_X1 U7559 ( .B1(n6509), .B2(n6545), .A(n6508), .ZN(U2926) );
  NOR2_X1 U7560 ( .A1(n6516), .A2(n4975), .ZN(n6539) );
  AOI21_X1 U7561 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6553), .A(n6539), .ZN(n6510) );
  OAI21_X1 U7562 ( .B1(n4049), .B2(n6545), .A(n6510), .ZN(U2927) );
  NOR2_X1 U7563 ( .A1(n6516), .A2(n6511), .ZN(n6541) );
  AOI21_X1 U7564 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6553), .A(n6541), .ZN(n6512) );
  OAI21_X1 U7565 ( .B1(n6513), .B2(n6545), .A(n6512), .ZN(U2928) );
  INV_X1 U7566 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6515) );
  NOR2_X1 U7567 ( .A1(n6516), .A2(n5099), .ZN(n6543) );
  AOI21_X1 U7568 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6553), .A(n6543), .ZN(n6514) );
  OAI21_X1 U7569 ( .B1(n6515), .B2(n6545), .A(n6514), .ZN(U2929) );
  INV_X1 U7570 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6518) );
  INV_X1 U7571 ( .A(n6516), .ZN(n6531) );
  AOI22_X1 U7572 ( .A1(n6549), .A2(UWORD_REG_6__SCAN_IN), .B1(n6531), .B2(
        DATAI_6_), .ZN(n6517) );
  OAI21_X1 U7573 ( .B1(n6518), .B2(n6545), .A(n6517), .ZN(U2930) );
  INV_X1 U7574 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6976) );
  AOI22_X1 U7575 ( .A1(n6553), .A2(UWORD_REG_7__SCAN_IN), .B1(n6531), .B2(
        DATAI_7_), .ZN(n6519) );
  OAI21_X1 U7576 ( .B1(n6976), .B2(n6545), .A(n6519), .ZN(U2931) );
  AOI21_X1 U7577 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6553), .A(n6520), .ZN(n6521) );
  OAI21_X1 U7578 ( .B1(n4155), .B2(n6545), .A(n6521), .ZN(U2932) );
  NAND2_X1 U7579 ( .A1(n6531), .A2(DATAI_9_), .ZN(n6547) );
  INV_X1 U7580 ( .A(n6547), .ZN(n6522) );
  AOI21_X1 U7581 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6553), .A(n6522), .ZN(n6523) );
  OAI21_X1 U7582 ( .B1(n4172), .B2(n6545), .A(n6523), .ZN(U2933) );
  NAND2_X1 U7583 ( .A1(n6531), .A2(DATAI_10_), .ZN(n6550) );
  INV_X1 U7584 ( .A(n6550), .ZN(n6524) );
  AOI21_X1 U7585 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6553), .A(n6524), .ZN(
        n6525) );
  OAI21_X1 U7586 ( .B1(n6526), .B2(n6545), .A(n6525), .ZN(U2934) );
  INV_X1 U7587 ( .A(EAX_REG_27__SCAN_IN), .ZN(n7125) );
  AOI22_X1 U7588 ( .A1(n6553), .A2(UWORD_REG_11__SCAN_IN), .B1(n6531), .B2(
        DATAI_11_), .ZN(n6527) );
  OAI21_X1 U7589 ( .B1(n7125), .B2(n6545), .A(n6527), .ZN(U2935) );
  INV_X1 U7590 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6530) );
  AOI21_X1 U7591 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6553), .A(n6528), .ZN(
        n6529) );
  OAI21_X1 U7592 ( .B1(n6530), .B2(n6545), .A(n6529), .ZN(U2936) );
  INV_X1 U7593 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U7594 ( .A1(n6531), .A2(DATAI_13_), .ZN(n6554) );
  INV_X1 U7595 ( .A(n6554), .ZN(n6532) );
  AOI21_X1 U7596 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6553), .A(n6532), .ZN(
        n6533) );
  OAI21_X1 U7597 ( .B1(n6534), .B2(n6545), .A(n6533), .ZN(U2937) );
  AOI21_X1 U7598 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6553), .A(n6535), .ZN(n6536) );
  OAI21_X1 U7599 ( .B1(n7078), .B2(n6545), .A(n6536), .ZN(U2939) );
  INV_X1 U7600 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6972) );
  AOI21_X1 U7601 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6553), .A(n6537), .ZN(n6538) );
  OAI21_X1 U7602 ( .B1(n6972), .B2(n6545), .A(n6538), .ZN(U2940) );
  AOI21_X1 U7603 ( .B1(LWORD_REG_3__SCAN_IN), .B2(n6553), .A(n6539), .ZN(n6540) );
  OAI21_X1 U7604 ( .B1(n7160), .B2(n6545), .A(n6540), .ZN(U2942) );
  AOI21_X1 U7605 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6553), .A(n6541), .ZN(n6542) );
  OAI21_X1 U7606 ( .B1(n6975), .B2(n6545), .A(n6542), .ZN(U2943) );
  AOI21_X1 U7607 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6553), .A(n6543), .ZN(n6544) );
  OAI21_X1 U7608 ( .B1(n6546), .B2(n6545), .A(n6544), .ZN(U2944) );
  AOI22_X1 U7609 ( .A1(n6553), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n6552), .ZN(n6548) );
  NAND2_X1 U7610 ( .A1(n6548), .A2(n6547), .ZN(U2948) );
  AOI22_X1 U7611 ( .A1(n6549), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6552), .ZN(n6551) );
  NAND2_X1 U7612 ( .A1(n6551), .A2(n6550), .ZN(U2949) );
  AOI22_X1 U7613 ( .A1(n6553), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6552), .ZN(n6555) );
  NAND2_X1 U7614 ( .A1(n6555), .A2(n6554), .ZN(U2952) );
  NOR2_X1 U7615 ( .A1(n6577), .A2(n6556), .ZN(n6614) );
  AOI21_X1 U7616 ( .B1(n6578), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6614), 
        .ZN(n6564) );
  OAI21_X1 U7617 ( .B1(n6559), .B2(n6558), .A(n6557), .ZN(n6560) );
  INV_X1 U7618 ( .A(n6560), .ZN(n6617) );
  INV_X1 U7619 ( .A(n6561), .ZN(n6562) );
  AOI22_X1 U7620 ( .A1(n6617), .A2(n3784), .B1(n6571), .B2(n6562), .ZN(n6563)
         );
  OAI211_X1 U7621 ( .C1(n6586), .C2(n6565), .A(n6564), .B(n6563), .ZN(U2980)
         );
  AND2_X1 U7622 ( .A1(n6566), .A2(REIP_REG_4__SCAN_IN), .ZN(n6622) );
  AOI21_X1 U7623 ( .B1(n6578), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6622), 
        .ZN(n6574) );
  OAI21_X1 U7624 ( .B1(n6569), .B2(n6567), .A(n6568), .ZN(n6570) );
  INV_X1 U7625 ( .A(n6570), .ZN(n6624) );
  AOI22_X1 U7626 ( .A1(n6624), .A2(n3784), .B1(n6572), .B2(n6571), .ZN(n6573)
         );
  OAI211_X1 U7627 ( .C1(n6586), .C2(n6575), .A(n6574), .B(n6573), .ZN(U2982)
         );
  NOR2_X1 U7628 ( .A1(n6577), .A2(n6576), .ZN(n6642) );
  AOI21_X1 U7629 ( .B1(n6578), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n6642), 
        .ZN(n6584) );
  XNOR2_X1 U7630 ( .A(n6579), .B(n3616), .ZN(n6581) );
  XNOR2_X1 U7631 ( .A(n6581), .B(n6580), .ZN(n6648) );
  AOI22_X1 U7632 ( .A1(n6582), .A2(n6571), .B1(n3784), .B2(n6648), .ZN(n6583)
         );
  OAI211_X1 U7633 ( .C1(n6586), .C2(n6585), .A(n6584), .B(n6583), .ZN(U2984)
         );
  AOI21_X1 U7634 ( .B1(n6644), .B2(n6588), .A(n6587), .ZN(n6592) );
  AOI21_X1 U7635 ( .B1(n6590), .B2(n6649), .A(n6589), .ZN(n6591) );
  OAI211_X1 U7636 ( .C1(n6594), .C2(n6593), .A(n6592), .B(n6591), .ZN(U3009)
         );
  OAI21_X1 U7637 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6595), .ZN(n6603) );
  INV_X1 U7638 ( .A(n6596), .ZN(n6597) );
  AOI21_X1 U7639 ( .B1(n6644), .B2(n6598), .A(n6597), .ZN(n6602) );
  INV_X1 U7640 ( .A(n6599), .ZN(n6600) );
  AOI22_X1 U7641 ( .A1(n6600), .A2(n6649), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n6608), .ZN(n6601) );
  OAI211_X1 U7642 ( .C1(n6612), .C2(n6603), .A(n6602), .B(n6601), .ZN(U3010)
         );
  INV_X1 U7643 ( .A(n6604), .ZN(n6605) );
  AOI21_X1 U7644 ( .B1(n6644), .B2(n6606), .A(n6605), .ZN(n6611) );
  INV_X1 U7645 ( .A(n6607), .ZN(n6609) );
  AOI22_X1 U7646 ( .A1(n6609), .A2(n6649), .B1(INSTADDRPOINTER_REG_7__SCAN_IN), 
        .B2(n6608), .ZN(n6610) );
  OAI211_X1 U7647 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6612), .A(n6611), 
        .B(n6610), .ZN(U3011) );
  INV_X1 U7648 ( .A(n6613), .ZN(n6615) );
  AOI21_X1 U7649 ( .B1(n6644), .B2(n6615), .A(n6614), .ZN(n6619) );
  AOI22_X1 U7650 ( .A1(n6617), .A2(n6649), .B1(n6616), .B2(n6620), .ZN(n6618)
         );
  OAI211_X1 U7651 ( .C1(n6621), .C2(n6620), .A(n6619), .B(n6618), .ZN(U3012)
         );
  AOI21_X1 U7652 ( .B1(n6645), .B2(n6647), .A(n6650), .ZN(n6641) );
  AOI21_X1 U7653 ( .B1(n6644), .B2(n6623), .A(n6622), .ZN(n6628) );
  AOI211_X1 U7654 ( .C1(n6640), .C2(n6629), .A(n6634), .B(n6647), .ZN(n6626)
         );
  AOI22_X1 U7655 ( .A1(n6626), .A2(n6625), .B1(n6649), .B2(n6624), .ZN(n6627)
         );
  OAI211_X1 U7656 ( .C1(n6641), .C2(n6629), .A(n6628), .B(n6627), .ZN(U3014)
         );
  INV_X1 U7657 ( .A(n6630), .ZN(n6633) );
  INV_X1 U7658 ( .A(n6631), .ZN(n6632) );
  AOI21_X1 U7659 ( .B1(n6644), .B2(n6633), .A(n6632), .ZN(n6639) );
  NOR2_X1 U7660 ( .A1(n6647), .A2(n6634), .ZN(n6637) );
  INV_X1 U7661 ( .A(n6635), .ZN(n6636) );
  AOI22_X1 U7662 ( .A1(n6637), .A2(n6640), .B1(n6649), .B2(n6636), .ZN(n6638)
         );
  OAI211_X1 U7663 ( .C1(n6641), .C2(n6640), .A(n6639), .B(n6638), .ZN(U3015)
         );
  AOI21_X1 U7664 ( .B1(n6644), .B2(n6643), .A(n6642), .ZN(n6655) );
  OAI221_X1 U7665 ( .B1(n6647), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .C1(n6647), .C2(n6646), .A(n6645), .ZN(n6654) );
  AOI22_X1 U7666 ( .A1(n6650), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6649), 
        .B2(n6648), .ZN(n6653) );
  NAND3_X1 U7667 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n3616), .A3(n6651), 
        .ZN(n6652) );
  NAND4_X1 U7668 ( .A1(n6655), .A2(n6654), .A3(n6653), .A4(n6652), .ZN(U3016)
         );
  NOR2_X1 U7669 ( .A1(n7116), .A2(n6656), .ZN(U3019) );
  NAND2_X1 U7670 ( .A1(n6665), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6703) );
  OAI21_X1 U7671 ( .B1(n6658), .B2(n6657), .A(n6703), .ZN(n6669) );
  NOR2_X1 U7672 ( .A1(n6661), .A2(n6703), .ZN(n6662) );
  AOI21_X1 U7673 ( .B1(n6763), .B2(n6663), .A(n6662), .ZN(n6673) );
  INV_X1 U7674 ( .A(n6664), .ZN(n6670) );
  INV_X1 U7675 ( .A(n6665), .ZN(n6666) );
  NAND2_X1 U7676 ( .A1(n6666), .A2(n6722), .ZN(n6667) );
  OAI211_X1 U7677 ( .C1(n6670), .C2(n6669), .A(n6668), .B(n6667), .ZN(n6708)
         );
  AOI22_X1 U7678 ( .A1(n6708), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n6731), 
        .B2(n6707), .ZN(n6672) );
  OAI211_X1 U7679 ( .C1(n6711), .C2(n6717), .A(n6673), .B(n6672), .ZN(U3060)
         );
  NOR2_X1 U7680 ( .A1(n6770), .A2(n6703), .ZN(n6674) );
  AOI21_X1 U7681 ( .B1(n6763), .B2(n6675), .A(n6674), .ZN(n6677) );
  AOI22_X1 U7682 ( .A1(n6708), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n6736), 
        .B2(n6707), .ZN(n6676) );
  OAI211_X1 U7683 ( .C1(n6711), .C2(n6678), .A(n6677), .B(n6676), .ZN(U3061)
         );
  NOR2_X1 U7684 ( .A1(n6777), .A2(n6703), .ZN(n6679) );
  AOI21_X1 U7685 ( .B1(n6763), .B2(n6680), .A(n6679), .ZN(n6682) );
  AOI22_X1 U7686 ( .A1(n6708), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n6740), 
        .B2(n6707), .ZN(n6681) );
  OAI211_X1 U7687 ( .C1(n6711), .C2(n6683), .A(n6682), .B(n6681), .ZN(U3062)
         );
  NOR2_X1 U7688 ( .A1(n6784), .A2(n6703), .ZN(n6684) );
  AOI21_X1 U7689 ( .B1(n6763), .B2(n6685), .A(n6684), .ZN(n6687) );
  AOI22_X1 U7690 ( .A1(n6708), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n6744), 
        .B2(n6707), .ZN(n6686) );
  OAI211_X1 U7691 ( .C1(n6711), .C2(n6688), .A(n6687), .B(n6686), .ZN(U3063)
         );
  NOR2_X1 U7692 ( .A1(n6850), .A2(n6703), .ZN(n6689) );
  AOI21_X1 U7693 ( .B1(n6763), .B2(n6690), .A(n6689), .ZN(n6692) );
  AOI22_X1 U7694 ( .A1(n6708), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n6855), 
        .B2(n6707), .ZN(n6691) );
  OAI211_X1 U7695 ( .C1(n6711), .C2(n6860), .A(n6692), .B(n6691), .ZN(U3064)
         );
  NOR2_X1 U7696 ( .A1(n6791), .A2(n6703), .ZN(n6693) );
  AOI21_X1 U7697 ( .B1(n6763), .B2(n6694), .A(n6693), .ZN(n6696) );
  AOI22_X1 U7698 ( .A1(n6708), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n6751), 
        .B2(n6707), .ZN(n6695) );
  OAI211_X1 U7699 ( .C1(n6711), .C2(n6697), .A(n6696), .B(n6695), .ZN(U3065)
         );
  NOR2_X1 U7700 ( .A1(n6799), .A2(n6703), .ZN(n6698) );
  AOI21_X1 U7701 ( .B1(n6763), .B2(n6699), .A(n6698), .ZN(n6701) );
  AOI22_X1 U7702 ( .A1(n6708), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n6755), 
        .B2(n6707), .ZN(n6700) );
  OAI211_X1 U7703 ( .C1(n6711), .C2(n6702), .A(n6701), .B(n6700), .ZN(U3066)
         );
  NOR2_X1 U7704 ( .A1(n6704), .A2(n6703), .ZN(n6705) );
  AOI21_X1 U7705 ( .B1(n6763), .B2(n6706), .A(n6705), .ZN(n6710) );
  AOI22_X1 U7706 ( .A1(n6708), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n6764), 
        .B2(n6707), .ZN(n6709) );
  OAI211_X1 U7707 ( .C1(n6711), .C2(n6758), .A(n6710), .B(n6709), .ZN(U3067)
         );
  AOI22_X1 U7708 ( .A1(n6715), .A2(n6714), .B1(n6713), .B2(n6712), .ZN(n6716)
         );
  INV_X1 U7709 ( .A(n6717), .ZN(n6721) );
  NAND2_X1 U7710 ( .A1(n6719), .A2(n6718), .ZN(n6727) );
  INV_X1 U7711 ( .A(n6727), .ZN(n6759) );
  AOI22_X1 U7712 ( .A1(n6762), .A2(n6721), .B1(n6720), .B2(n6759), .ZN(n6733)
         );
  NOR3_X1 U7713 ( .A1(n6763), .A2(n6723), .A3(n6722), .ZN(n6726) );
  OAI21_X1 U7714 ( .B1(n6726), .B2(n6725), .A(n6724), .ZN(n6730) );
  AOI21_X1 U7715 ( .B1(n6727), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6728) );
  NAND3_X1 U7716 ( .A1(n6730), .A2(n6729), .A3(n6728), .ZN(n6765) );
  AOI22_X1 U7717 ( .A1(n6765), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6731), 
        .B2(n6763), .ZN(n6732) );
  OAI211_X1 U7718 ( .C1(n6734), .C2(n6768), .A(n6733), .B(n6732), .ZN(U3068)
         );
  AOI22_X1 U7719 ( .A1(n6762), .A2(n6773), .B1(n6735), .B2(n6759), .ZN(n6738)
         );
  AOI22_X1 U7720 ( .A1(n6765), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6736), 
        .B2(n6763), .ZN(n6737) );
  OAI211_X1 U7721 ( .C1(n6771), .C2(n6768), .A(n6738), .B(n6737), .ZN(U3069)
         );
  AOI22_X1 U7722 ( .A1(n6762), .A2(n6780), .B1(n6739), .B2(n6759), .ZN(n6742)
         );
  AOI22_X1 U7723 ( .A1(n6765), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6740), 
        .B2(n6763), .ZN(n6741) );
  OAI211_X1 U7724 ( .C1(n6778), .C2(n6768), .A(n6742), .B(n6741), .ZN(U3070)
         );
  AOI22_X1 U7725 ( .A1(n6762), .A2(n6787), .B1(n6743), .B2(n6759), .ZN(n6746)
         );
  AOI22_X1 U7726 ( .A1(n6765), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6744), 
        .B2(n6763), .ZN(n6745) );
  OAI211_X1 U7727 ( .C1(n6785), .C2(n6768), .A(n6746), .B(n6745), .ZN(U3071)
         );
  INV_X1 U7728 ( .A(n6860), .ZN(n6747) );
  AOI22_X1 U7729 ( .A1(n6762), .A2(n6747), .B1(n3191), .B2(n6759), .ZN(n6749)
         );
  AOI22_X1 U7730 ( .A1(n6765), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6855), 
        .B2(n6763), .ZN(n6748) );
  OAI211_X1 U7731 ( .C1(n6852), .C2(n6768), .A(n6749), .B(n6748), .ZN(U3072)
         );
  AOI22_X1 U7732 ( .A1(n6762), .A2(n6794), .B1(n6750), .B2(n6759), .ZN(n6753)
         );
  AOI22_X1 U7733 ( .A1(n6765), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6751), 
        .B2(n6763), .ZN(n6752) );
  OAI211_X1 U7734 ( .C1(n6792), .C2(n6768), .A(n6753), .B(n6752), .ZN(U3073)
         );
  AOI22_X1 U7735 ( .A1(n6762), .A2(n6804), .B1(n6754), .B2(n6759), .ZN(n6757)
         );
  AOI22_X1 U7736 ( .A1(n6765), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6755), 
        .B2(n6763), .ZN(n6756) );
  OAI211_X1 U7737 ( .C1(n6800), .C2(n6768), .A(n6757), .B(n6756), .ZN(U3074)
         );
  INV_X1 U7738 ( .A(n6758), .ZN(n6761) );
  AOI22_X1 U7739 ( .A1(n6762), .A2(n6761), .B1(n6760), .B2(n6759), .ZN(n6767)
         );
  AOI22_X1 U7740 ( .A1(n6765), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6764), 
        .B2(n6763), .ZN(n6766) );
  OAI211_X1 U7741 ( .C1(n6769), .C2(n6768), .A(n6767), .B(n6766), .ZN(U3075)
         );
  OAI22_X1 U7742 ( .A1(n6801), .A2(n6771), .B1(n6770), .B2(n6798), .ZN(n6772)
         );
  INV_X1 U7743 ( .A(n6772), .ZN(n6775) );
  AOI22_X1 U7744 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6805), .B1(n6773), 
        .B2(n6803), .ZN(n6774) );
  OAI211_X1 U7745 ( .C1(n6853), .C2(n6776), .A(n6775), .B(n6774), .ZN(U3109)
         );
  OAI22_X1 U7746 ( .A1(n6801), .A2(n6778), .B1(n6777), .B2(n6798), .ZN(n6779)
         );
  INV_X1 U7747 ( .A(n6779), .ZN(n6782) );
  AOI22_X1 U7748 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6805), .B1(n6780), 
        .B2(n6803), .ZN(n6781) );
  OAI211_X1 U7749 ( .C1(n6853), .C2(n6783), .A(n6782), .B(n6781), .ZN(U3110)
         );
  OAI22_X1 U7750 ( .A1(n6801), .A2(n6785), .B1(n6784), .B2(n6798), .ZN(n6786)
         );
  INV_X1 U7751 ( .A(n6786), .ZN(n6789) );
  AOI22_X1 U7752 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6805), .B1(n6787), 
        .B2(n6803), .ZN(n6788) );
  OAI211_X1 U7753 ( .C1(n6853), .C2(n6790), .A(n6789), .B(n6788), .ZN(U3111)
         );
  OAI22_X1 U7754 ( .A1(n6801), .A2(n6792), .B1(n6791), .B2(n6798), .ZN(n6793)
         );
  INV_X1 U7755 ( .A(n6793), .ZN(n6796) );
  AOI22_X1 U7756 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6805), .B1(n6794), 
        .B2(n6803), .ZN(n6795) );
  OAI211_X1 U7757 ( .C1(n6853), .C2(n6797), .A(n6796), .B(n6795), .ZN(U3113)
         );
  OAI22_X1 U7758 ( .A1(n6801), .A2(n6800), .B1(n6799), .B2(n6798), .ZN(n6802)
         );
  INV_X1 U7759 ( .A(n6802), .ZN(n6807) );
  AOI22_X1 U7760 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6805), .B1(n6804), 
        .B2(n6803), .ZN(n6806) );
  OAI211_X1 U7761 ( .C1(n6853), .C2(n6808), .A(n6807), .B(n6806), .ZN(U3114)
         );
  INV_X1 U7762 ( .A(DATAWIDTH_REG_31__SCAN_IN), .ZN(n7061) );
  NOR2_X1 U7763 ( .A1(n6829), .A2(n7061), .ZN(U3151) );
  INV_X1 U7764 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6863) );
  NOR2_X1 U7765 ( .A1(n6829), .A2(n6863), .ZN(U3152) );
  INV_X1 U7766 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n7077) );
  NOR2_X1 U7767 ( .A1(n6829), .A2(n7077), .ZN(U3153) );
  AND2_X1 U7768 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6809), .ZN(U3154) );
  AND2_X1 U7769 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6809), .ZN(U3155) );
  AND2_X1 U7770 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6809), .ZN(U3156) );
  INV_X1 U7771 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6914) );
  NOR2_X1 U7772 ( .A1(n6829), .A2(n6914), .ZN(U3157) );
  INV_X1 U7773 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n7147) );
  NOR2_X1 U7774 ( .A1(n6829), .A2(n7147), .ZN(U3158) );
  NOR2_X1 U7775 ( .A1(n6829), .A2(n6915), .ZN(U3159) );
  AND2_X1 U7776 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6809), .ZN(U3160) );
  NOR2_X1 U7777 ( .A1(n6829), .A2(n7045), .ZN(U3161) );
  AND2_X1 U7778 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6809), .ZN(U3162) );
  AND2_X1 U7779 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6809), .ZN(U3163) );
  AND2_X1 U7780 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6809), .ZN(U3164) );
  INV_X1 U7781 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n7083) );
  NOR2_X1 U7782 ( .A1(n6829), .A2(n7083), .ZN(U3165) );
  AND2_X1 U7783 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6809), .ZN(U3166) );
  NOR2_X1 U7784 ( .A1(n6829), .A2(n7080), .ZN(U3167) );
  AND2_X1 U7785 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6809), .ZN(U3168) );
  AND2_X1 U7786 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6809), .ZN(U3169) );
  NOR2_X1 U7787 ( .A1(n6829), .A2(n6978), .ZN(U3170) );
  AND2_X1 U7788 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6809), .ZN(U3171) );
  AND2_X1 U7789 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6809), .ZN(U3172) );
  AND2_X1 U7790 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6809), .ZN(U3173) );
  NOR2_X1 U7791 ( .A1(n6829), .A2(n7084), .ZN(U3174) );
  INV_X1 U7792 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n7097) );
  NOR2_X1 U7793 ( .A1(n6829), .A2(n7097), .ZN(U3175) );
  INV_X1 U7794 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n7091) );
  NOR2_X1 U7795 ( .A1(n6829), .A2(n7091), .ZN(U3176) );
  AND2_X1 U7796 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6809), .ZN(U3177) );
  AND2_X1 U7797 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6809), .ZN(U3178) );
  AND2_X1 U7798 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6809), .ZN(U3179) );
  AND2_X1 U7799 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6809), .ZN(U3180) );
  NAND2_X1 U7800 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6812) );
  NAND2_X1 U7801 ( .A1(n6810), .A2(n6817), .ZN(n6811) );
  INV_X1 U7802 ( .A(NA_N), .ZN(n6818) );
  AOI221_X1 U7803 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6818), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6822) );
  AOI21_X1 U7804 ( .B1(n6812), .B2(n6811), .A(n6822), .ZN(n6813) );
  OAI221_X1 U7805 ( .B1(n6825), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6825), 
        .C2(n6814), .A(n6813), .ZN(U3181) );
  AOI221_X1 U7806 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6838), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6816) );
  AOI221_X1 U7807 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6816), .C2(HOLD), .A(n6815), .ZN(n6823) );
  INV_X1 U7808 ( .A(n6817), .ZN(n6819) );
  NAND4_X1 U7809 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n6819), .A4(n6818), .ZN(n6821) );
  NAND3_X1 U7810 ( .A1(READY_N), .A2(STATE_REG_2__SCAN_IN), .A3(
        STATE_REG_1__SCAN_IN), .ZN(n6820) );
  OAI211_X1 U7811 ( .C1(n6823), .C2(n6822), .A(n6821), .B(n6820), .ZN(U3183)
         );
  INV_X1 U7812 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6974) );
  AOI22_X1 U7813 ( .A1(n6825), .A2(n6912), .B1(n6974), .B2(n6849), .ZN(U3445)
         );
  MUX2_X1 U7814 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6849), .Z(U3446) );
  INV_X1 U7815 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n7146) );
  AOI22_X1 U7816 ( .A1(n6825), .A2(n6824), .B1(n7146), .B2(n6849), .ZN(U3447)
         );
  INV_X1 U7817 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6836) );
  INV_X1 U7818 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n7065) );
  AOI22_X1 U7819 ( .A1(n6825), .A2(n6836), .B1(n7065), .B2(n6849), .ZN(U3448)
         );
  OAI21_X1 U7820 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6829), .A(n6827), .ZN(
        n6826) );
  INV_X1 U7821 ( .A(n6826), .ZN(U3451) );
  OAI21_X1 U7822 ( .B1(n6829), .B2(n6828), .A(n6827), .ZN(U3452) );
  AOI21_X1 U7823 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6830) );
  AOI22_X1 U7824 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6830), .B2(n6926), .ZN(n6832) );
  INV_X1 U7825 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6831) );
  AOI22_X1 U7826 ( .A1(n6833), .A2(n6832), .B1(n6831), .B2(n6835), .ZN(U3468)
         );
  NOR2_X1 U7827 ( .A1(n6835), .A2(REIP_REG_1__SCAN_IN), .ZN(n6834) );
  AOI22_X1 U7828 ( .A1(n6836), .A2(n6835), .B1(n6928), .B2(n6834), .ZN(U3469)
         );
  NAND2_X1 U7829 ( .A1(n6849), .A2(W_R_N_REG_SCAN_IN), .ZN(n6837) );
  OAI21_X1 U7830 ( .B1(n6849), .B2(READREQUEST_REG_SCAN_IN), .A(n6837), .ZN(
        U3470) );
  AND2_X1 U7831 ( .A1(n6839), .A2(n6838), .ZN(n6841) );
  NOR3_X1 U7832 ( .A1(n6842), .A2(n6841), .A3(n6840), .ZN(n6848) );
  OAI211_X1 U7833 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n3590), .A(n6843), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6845) );
  AOI21_X1 U7834 ( .B1(n6845), .B2(STATE2_REG_0__SCAN_IN), .A(n6844), .ZN(
        n6847) );
  NAND2_X1 U7835 ( .A1(n6848), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6846) );
  OAI21_X1 U7836 ( .B1(n6848), .B2(n6847), .A(n6846), .ZN(U3472) );
  MUX2_X1 U7837 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6849), .Z(U3473) );
  OAI22_X1 U7838 ( .A1(n6853), .A2(n6852), .B1(n6851), .B2(n6850), .ZN(n6854)
         );
  AOI21_X1 U7839 ( .B1(n6856), .B2(n6855), .A(n6854), .ZN(n6859) );
  NAND2_X1 U7840 ( .A1(n6857), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6858)
         );
  OAI211_X1 U7841 ( .C1(n6861), .C2(n6860), .A(n6859), .B(n6858), .ZN(n7183)
         );
  INV_X1 U7842 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n7010) );
  AOI22_X1 U7843 ( .A1(n7010), .A2(keyinput3), .B1(keyinput89), .B2(n6863), 
        .ZN(n6862) );
  OAI221_X1 U7844 ( .B1(n7010), .B2(keyinput3), .C1(n6863), .C2(keyinput89), 
        .A(n6862), .ZN(n6873) );
  INV_X1 U7845 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6865) );
  AOI22_X1 U7846 ( .A1(n6865), .A2(keyinput106), .B1(n6972), .B2(keyinput46), 
        .ZN(n6864) );
  OAI221_X1 U7847 ( .B1(n6865), .B2(keyinput106), .C1(n6972), .C2(keyinput46), 
        .A(n6864), .ZN(n6872) );
  INV_X1 U7848 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6979) );
  AOI22_X1 U7849 ( .A1(n6973), .A2(keyinput59), .B1(keyinput4), .B2(n6979), 
        .ZN(n6866) );
  OAI221_X1 U7850 ( .B1(n6973), .B2(keyinput59), .C1(n6979), .C2(keyinput4), 
        .A(n6866), .ZN(n6871) );
  INV_X1 U7851 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6869) );
  INV_X1 U7852 ( .A(DATAI_30_), .ZN(n6868) );
  AOI22_X1 U7853 ( .A1(n6869), .A2(keyinput24), .B1(keyinput83), .B2(n6868), 
        .ZN(n6867) );
  OAI221_X1 U7854 ( .B1(n6869), .B2(keyinput24), .C1(n6868), .C2(keyinput83), 
        .A(n6867), .ZN(n6870) );
  NOR4_X1 U7855 ( .A1(n6873), .A2(n6872), .A3(n6871), .A4(n6870), .ZN(n7181)
         );
  INV_X1 U7856 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6876) );
  AOI22_X1 U7857 ( .A1(n6876), .A2(keyinput122), .B1(keyinput103), .B2(n6875), 
        .ZN(n6874) );
  OAI221_X1 U7858 ( .B1(n6876), .B2(keyinput122), .C1(n6875), .C2(keyinput103), 
        .A(n6874), .ZN(n6885) );
  INV_X1 U7859 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6988) );
  AOI22_X1 U7860 ( .A1(n6988), .A2(keyinput81), .B1(keyinput75), .B2(n6878), 
        .ZN(n6877) );
  OAI221_X1 U7861 ( .B1(n6988), .B2(keyinput81), .C1(n6878), .C2(keyinput75), 
        .A(n6877), .ZN(n6884) );
  AOI22_X1 U7862 ( .A1(n6974), .A2(keyinput68), .B1(n6975), .B2(keyinput69), 
        .ZN(n6879) );
  OAI221_X1 U7863 ( .B1(n6974), .B2(keyinput68), .C1(n6975), .C2(keyinput69), 
        .A(n6879), .ZN(n6883) );
  XNOR2_X1 U7864 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .B(keyinput14), .ZN(n6880)
         );
  OAI21_X1 U7865 ( .B1(n6881), .B2(keyinput7), .A(n6880), .ZN(n6882) );
  NOR4_X1 U7866 ( .A1(n6885), .A2(n6884), .A3(n6883), .A4(n6882), .ZN(n7180)
         );
  INV_X1 U7867 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n7011) );
  AOI22_X1 U7868 ( .A1(n7011), .A2(keyinput102), .B1(keyinput127), .B2(n6980), 
        .ZN(n6886) );
  OAI221_X1 U7869 ( .B1(n7011), .B2(keyinput102), .C1(n6980), .C2(keyinput127), 
        .A(n6886), .ZN(n6971) );
  INV_X1 U7870 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6888) );
  AOI22_X1 U7871 ( .A1(n7009), .A2(keyinput23), .B1(n6888), .B2(keyinput2), 
        .ZN(n6887) );
  OAI221_X1 U7872 ( .B1(n7009), .B2(keyinput23), .C1(n6888), .C2(keyinput2), 
        .A(n6887), .ZN(n6970) );
  OAI22_X1 U7873 ( .A1(n6977), .A2(keyinput44), .B1(n7023), .B2(keyinput80), 
        .ZN(n6889) );
  AOI221_X1 U7874 ( .B1(n6977), .B2(keyinput44), .C1(keyinput80), .C2(n7023), 
        .A(n6889), .ZN(n6908) );
  OAI22_X1 U7875 ( .A1(n6987), .A2(keyinput116), .B1(n6891), .B2(keyinput90), 
        .ZN(n6890) );
  AOI221_X1 U7876 ( .B1(n6987), .B2(keyinput116), .C1(keyinput90), .C2(n6891), 
        .A(n6890), .ZN(n6907) );
  INV_X1 U7877 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6893) );
  AOI22_X1 U7878 ( .A1(n6978), .A2(keyinput124), .B1(n6893), .B2(keyinput8), 
        .ZN(n6892) );
  OAI221_X1 U7879 ( .B1(n6978), .B2(keyinput124), .C1(n6893), .C2(keyinput8), 
        .A(n6892), .ZN(n6905) );
  INV_X1 U7880 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U7881 ( .A1(n6896), .A2(keyinput94), .B1(n6895), .B2(keyinput56), 
        .ZN(n6894) );
  OAI221_X1 U7882 ( .B1(n6896), .B2(keyinput94), .C1(n6895), .C2(keyinput56), 
        .A(n6894), .ZN(n6904) );
  INV_X1 U7883 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6899) );
  INV_X1 U7884 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6898) );
  AOI22_X1 U7885 ( .A1(n6899), .A2(keyinput35), .B1(keyinput112), .B2(n6898), 
        .ZN(n6897) );
  OAI221_X1 U7886 ( .B1(n6899), .B2(keyinput35), .C1(n6898), .C2(keyinput112), 
        .A(n6897), .ZN(n6903) );
  AOI22_X1 U7887 ( .A1(n6976), .A2(keyinput86), .B1(n6901), .B2(keyinput65), 
        .ZN(n6900) );
  OAI221_X1 U7888 ( .B1(n6976), .B2(keyinput86), .C1(n6901), .C2(keyinput65), 
        .A(n6900), .ZN(n6902) );
  NOR4_X1 U7889 ( .A1(n6905), .A2(n6904), .A3(n6903), .A4(n6902), .ZN(n6906)
         );
  NAND3_X1 U7890 ( .A1(n6908), .A2(n6907), .A3(n6906), .ZN(n6969) );
  AOI22_X1 U7891 ( .A1(n7026), .A2(keyinput15), .B1(keyinput99), .B2(n6910), 
        .ZN(n6909) );
  OAI221_X1 U7892 ( .B1(n7026), .B2(keyinput15), .C1(n6910), .C2(keyinput99), 
        .A(n6909), .ZN(n6922) );
  AOI22_X1 U7893 ( .A1(n6912), .A2(keyinput18), .B1(n7018), .B2(keyinput98), 
        .ZN(n6911) );
  OAI221_X1 U7894 ( .B1(n6912), .B2(keyinput18), .C1(n7018), .C2(keyinput98), 
        .A(n6911), .ZN(n6921) );
  AOI22_X1 U7895 ( .A1(n6915), .A2(keyinput34), .B1(keyinput20), .B2(n6914), 
        .ZN(n6913) );
  OAI221_X1 U7896 ( .B1(n6915), .B2(keyinput34), .C1(n6914), .C2(keyinput20), 
        .A(n6913), .ZN(n6920) );
  INV_X1 U7897 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n6917) );
  AOI22_X1 U7898 ( .A1(n6918), .A2(keyinput40), .B1(n6917), .B2(keyinput71), 
        .ZN(n6916) );
  OAI221_X1 U7899 ( .B1(n6918), .B2(keyinput40), .C1(n6917), .C2(keyinput71), 
        .A(n6916), .ZN(n6919) );
  NOR4_X1 U7900 ( .A1(n6922), .A2(n6921), .A3(n6920), .A4(n6919), .ZN(n6967)
         );
  INV_X1 U7901 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n7008) );
  AOI22_X1 U7902 ( .A1(n7008), .A2(keyinput121), .B1(keyinput57), .B2(n6924), 
        .ZN(n6923) );
  OAI221_X1 U7903 ( .B1(n7008), .B2(keyinput121), .C1(n6924), .C2(keyinput57), 
        .A(n6923), .ZN(n6934) );
  AOI22_X1 U7904 ( .A1(n6926), .A2(keyinput38), .B1(keyinput123), .B2(n7024), 
        .ZN(n6925) );
  OAI221_X1 U7905 ( .B1(n6926), .B2(keyinput38), .C1(n7024), .C2(keyinput123), 
        .A(n6925), .ZN(n6933) );
  AOI22_X1 U7906 ( .A1(n6985), .A2(keyinput36), .B1(keyinput26), .B2(n6928), 
        .ZN(n6927) );
  OAI221_X1 U7907 ( .B1(n6985), .B2(keyinput36), .C1(n6928), .C2(keyinput26), 
        .A(n6927), .ZN(n6932) );
  INV_X1 U7908 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n7022) );
  INV_X1 U7909 ( .A(EAX_REG_31__SCAN_IN), .ZN(n6930) );
  AOI22_X1 U7910 ( .A1(n7022), .A2(keyinput27), .B1(n6930), .B2(keyinput49), 
        .ZN(n6929) );
  OAI221_X1 U7911 ( .B1(n7022), .B2(keyinput27), .C1(n6930), .C2(keyinput49), 
        .A(n6929), .ZN(n6931) );
  NOR4_X1 U7912 ( .A1(n6934), .A2(n6933), .A3(n6932), .A4(n6931), .ZN(n6966)
         );
  INV_X1 U7913 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6936) );
  AOI22_X1 U7914 ( .A1(n6937), .A2(keyinput73), .B1(n6936), .B2(keyinput105), 
        .ZN(n6935) );
  OAI221_X1 U7915 ( .B1(n6937), .B2(keyinput73), .C1(n6936), .C2(keyinput105), 
        .A(n6935), .ZN(n6942) );
  XNOR2_X1 U7916 ( .A(n6938), .B(keyinput53), .ZN(n6941) );
  XNOR2_X1 U7917 ( .A(n6939), .B(keyinput48), .ZN(n6940) );
  OR3_X1 U7918 ( .A1(n6942), .A2(n6941), .A3(n6940), .ZN(n6950) );
  AOI22_X1 U7919 ( .A1(n6945), .A2(keyinput109), .B1(keyinput125), .B2(n6944), 
        .ZN(n6943) );
  OAI221_X1 U7920 ( .B1(n6945), .B2(keyinput109), .C1(n6944), .C2(keyinput125), 
        .A(n6943), .ZN(n6949) );
  AOI22_X1 U7921 ( .A1(n6947), .A2(keyinput61), .B1(n7019), .B2(keyinput70), 
        .ZN(n6946) );
  OAI221_X1 U7922 ( .B1(n6947), .B2(keyinput61), .C1(n7019), .C2(keyinput70), 
        .A(n6946), .ZN(n6948) );
  NOR3_X1 U7923 ( .A1(n6950), .A2(n6949), .A3(n6948), .ZN(n6965) );
  INV_X1 U7924 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6953) );
  AOI22_X1 U7925 ( .A1(n6953), .A2(keyinput118), .B1(keyinput9), .B2(n6952), 
        .ZN(n6951) );
  OAI221_X1 U7926 ( .B1(n6953), .B2(keyinput118), .C1(n6952), .C2(keyinput9), 
        .A(n6951), .ZN(n6963) );
  INV_X1 U7927 ( .A(DATAI_29_), .ZN(n6956) );
  AOI22_X1 U7928 ( .A1(n6956), .A2(keyinput82), .B1(n6955), .B2(keyinput17), 
        .ZN(n6954) );
  OAI221_X1 U7929 ( .B1(n6956), .B2(keyinput82), .C1(n6955), .C2(keyinput17), 
        .A(n6954), .ZN(n6962) );
  INV_X1 U7930 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n6986) );
  AOI22_X1 U7931 ( .A1(n6986), .A2(keyinput95), .B1(keyinput13), .B2(n6958), 
        .ZN(n6957) );
  OAI221_X1 U7932 ( .B1(n6986), .B2(keyinput95), .C1(n6958), .C2(keyinput13), 
        .A(n6957), .ZN(n6961) );
  INV_X1 U7933 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n7007) );
  AOI22_X1 U7934 ( .A1(n7007), .A2(keyinput126), .B1(keyinput31), .B2(n7025), 
        .ZN(n6959) );
  OAI221_X1 U7935 ( .B1(n7007), .B2(keyinput126), .C1(n7025), .C2(keyinput31), 
        .A(n6959), .ZN(n6960) );
  NOR4_X1 U7936 ( .A1(n6963), .A2(n6962), .A3(n6961), .A4(n6960), .ZN(n6964)
         );
  NAND4_X1 U7937 ( .A1(n6967), .A2(n6966), .A3(n6965), .A4(n6964), .ZN(n6968)
         );
  NOR4_X1 U7938 ( .A1(n6971), .A2(n6970), .A3(n6969), .A4(n6968), .ZN(n7179)
         );
  NAND4_X1 U7939 ( .A1(DATAI_30_), .A2(DATAO_REG_1__SCAN_IN), .A3(n6973), .A4(
        n6972), .ZN(n6984) );
  NAND4_X1 U7940 ( .A1(REIP_REG_13__SCAN_IN), .A2(LWORD_REG_14__SCAN_IN), .A3(
        n6975), .A4(n6974), .ZN(n6983) );
  NAND4_X1 U7941 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        DATAO_REG_29__SCAN_IN), .A3(n6977), .A4(n6976), .ZN(n6982) );
  NAND4_X1 U7942 ( .A1(DATAO_REG_9__SCAN_IN), .A2(n6980), .A3(n6979), .A4(
        n6978), .ZN(n6981) );
  NOR4_X1 U7943 ( .A1(n6984), .A2(n6983), .A3(n6982), .A4(n6981), .ZN(n7006)
         );
  INV_X1 U7944 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n7131) );
  NAND4_X1 U7945 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(
        INSTQUEUE_REG_12__3__SCAN_IN), .A3(n7131), .A4(n6985), .ZN(n6993) );
  INV_X1 U7946 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n7114) );
  NAND4_X1 U7947 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n7114), .A3(n6987), 
        .A4(n6986), .ZN(n6992) );
  INV_X1 U7948 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n7049) );
  NAND4_X1 U7949 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        INSTQUEUE_REG_8__2__SCAN_IN), .A3(n6988), .A4(n7049), .ZN(n6991) );
  INV_X1 U7950 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6989) );
  INV_X1 U7951 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n7143) );
  NAND4_X1 U7952 ( .A1(n6989), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .A3(
        INSTQUEUE_REG_14__6__SCAN_IN), .A4(n7143), .ZN(n6990) );
  NOR4_X1 U7953 ( .A1(n6993), .A2(n6992), .A3(n6991), .A4(n6990), .ZN(n7005)
         );
  NAND4_X1 U7954 ( .A1(ADDRESS_REG_20__SCAN_IN), .A2(DATAWIDTH_REG_29__SCAN_IN), .A3(LWORD_REG_2__SCAN_IN), .A4(n7078), .ZN(n6994) );
  NOR4_X1 U7955 ( .A1(DATAO_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(n6995), .A4(n6994), .ZN(n7004) );
  NOR4_X1 U7956 ( .A1(EAX_REG_27__SCAN_IN), .A2(UWORD_REG_2__SCAN_IN), .A3(
        n3829), .A4(n7130), .ZN(n6996) );
  NAND3_X1 U7957 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        BE_N_REG_1__SCAN_IN), .A3(n6996), .ZN(n7002) );
  NOR4_X1 U7958 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(EBX_REG_5__SCAN_IN), .A3(INSTADDRPOINTER_REG_15__SCAN_IN), .A4(ADDRESS_REG_3__SCAN_IN), .ZN(n7000) );
  NOR4_X1 U7959 ( .A1(ADDRESS_REG_9__SCAN_IN), .A2(n7090), .A3(n7101), .A4(
        n7091), .ZN(n6999) );
  NOR4_X1 U7960 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(DATAI_11_), .A3(
        ADDRESS_REG_11__SCAN_IN), .A4(n6997), .ZN(n6998) );
  NAND4_X1 U7961 ( .A1(n7000), .A2(n6999), .A3(n6998), .A4(n7160), .ZN(n7001)
         );
  NOR4_X1 U7962 ( .A1(EBX_REG_29__SCAN_IN), .A2(n7141), .A3(n7002), .A4(n7001), 
        .ZN(n7003) );
  NAND4_X1 U7963 ( .A1(n7006), .A2(n7005), .A3(n7004), .A4(n7003), .ZN(n7040)
         );
  INV_X1 U7964 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n7042) );
  NOR4_X1 U7965 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(
        INSTQUEUE_REG_0__0__SCAN_IN), .A3(n7007), .A4(n7042), .ZN(n7038) );
  INV_X1 U7966 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n7162) );
  NOR4_X1 U7967 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(
        INSTQUEUE_REG_1__4__SCAN_IN), .A3(n7008), .A4(n7162), .ZN(n7037) );
  NAND4_X1 U7968 ( .A1(STATE2_REG_0__SCAN_IN), .A2(
        INSTQUEUE_REG_13__4__SCAN_IN), .A3(PHYADDRPOINTER_REG_7__SCAN_IN), 
        .A4(DATAI_17_), .ZN(n7017) );
  INV_X1 U7969 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n7074) );
  NOR4_X1 U7970 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(
        INSTQUEUE_REG_8__7__SCAN_IN), .A3(n7009), .A4(n7074), .ZN(n7015) );
  NOR4_X1 U7971 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(
        INSTQUEUE_REG_8__0__SCAN_IN), .A3(INSTQUEUE_REG_13__0__SCAN_IN), .A4(
        n7010), .ZN(n7014) );
  INV_X1 U7972 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n7126) );
  NOR4_X1 U7973 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(
        INSTQUEUE_REG_13__1__SCAN_IN), .A3(INSTQUEUE_REG_5__7__SCAN_IN), .A4(
        n7126), .ZN(n7013) );
  INV_X1 U7974 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n7163) );
  NOR4_X1 U7975 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(
        INSTQUEUE_REG_12__7__SCAN_IN), .A3(n7011), .A4(n7163), .ZN(n7012) );
  NAND4_X1 U7976 ( .A1(n7015), .A2(n7014), .A3(n7013), .A4(n7012), .ZN(n7016)
         );
  NOR4_X1 U7977 ( .A1(n7018), .A2(n7166), .A3(n7017), .A4(n7016), .ZN(n7036)
         );
  NOR4_X1 U7978 ( .A1(ADDRESS_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(LWORD_REG_12__SCAN_IN), .A4(
        n7019), .ZN(n7020) );
  NAND3_X1 U7979 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        DATAO_REG_18__SCAN_IN), .A3(n7020), .ZN(n7034) );
  NAND4_X1 U7980 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(BE_N_REG_0__SCAN_IN), .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(n7059), .ZN(n7021) );
  NOR3_X1 U7981 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n7048), .A3(n7021), .ZN(
        n7032) );
  NAND4_X1 U7982 ( .A1(EAX_REG_31__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .A3(
        BYTEENABLE_REG_3__SCAN_IN), .A4(n7022), .ZN(n7030) );
  NAND4_X1 U7983 ( .A1(n7024), .A2(n7023), .A3(REIP_REG_1__SCAN_IN), .A4(
        EBX_REG_24__SCAN_IN), .ZN(n7029) );
  NAND4_X1 U7984 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(EBX_REG_4__SCAN_IN), .A3(DATAI_29_), .A4(n7025), .ZN(n7028) );
  NAND4_X1 U7985 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(
        ADDRESS_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(n7026), 
        .ZN(n7027) );
  NOR4_X1 U7986 ( .A1(n7030), .A2(n7029), .A3(n7028), .A4(n7027), .ZN(n7031)
         );
  NAND4_X1 U7987 ( .A1(EBX_REG_0__SCAN_IN), .A2(n7032), .A3(n7031), .A4(n7066), 
        .ZN(n7033) );
  NOR4_X1 U7988 ( .A1(EBX_REG_27__SCAN_IN), .A2(UWORD_REG_4__SCAN_IN), .A3(
        n7034), .A4(n7033), .ZN(n7035) );
  NAND4_X1 U7989 ( .A1(n7038), .A2(n7037), .A3(n7036), .A4(n7035), .ZN(n7039)
         );
  OAI21_X1 U7990 ( .B1(n7040), .B2(n7039), .A(DATAO_REG_2__SCAN_IN), .ZN(n7177) );
  AOI22_X1 U7991 ( .A1(n7043), .A2(keyinput58), .B1(n7042), .B2(keyinput77), 
        .ZN(n7041) );
  OAI221_X1 U7992 ( .B1(n7043), .B2(keyinput58), .C1(n7042), .C2(keyinput77), 
        .A(n7041), .ZN(n7056) );
  AOI22_X1 U7993 ( .A1(n7046), .A2(keyinput92), .B1(keyinput51), .B2(n7045), 
        .ZN(n7044) );
  OAI221_X1 U7994 ( .B1(n7046), .B2(keyinput92), .C1(n7045), .C2(keyinput51), 
        .A(n7044), .ZN(n7055) );
  AOI22_X1 U7995 ( .A1(n7049), .A2(keyinput60), .B1(keyinput74), .B2(n7048), 
        .ZN(n7047) );
  OAI221_X1 U7996 ( .B1(n7049), .B2(keyinput60), .C1(n7048), .C2(keyinput74), 
        .A(n7047), .ZN(n7054) );
  XOR2_X1 U7997 ( .A(n7050), .B(keyinput85), .Z(n7052) );
  XNOR2_X1 U7998 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .B(keyinput29), .ZN(n7051) );
  NAND2_X1 U7999 ( .A1(n7052), .A2(n7051), .ZN(n7053) );
  NOR4_X1 U8000 ( .A1(n7056), .A2(n7055), .A3(n7054), .A4(n7053), .ZN(n7108)
         );
  INV_X1 U8001 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n7058) );
  AOI22_X1 U8002 ( .A1(n7059), .A2(keyinput30), .B1(n7058), .B2(keyinput84), 
        .ZN(n7057) );
  OAI221_X1 U8003 ( .B1(n7059), .B2(keyinput30), .C1(n7058), .C2(keyinput84), 
        .A(n7057), .ZN(n7072) );
  INV_X1 U8004 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n7062) );
  AOI22_X1 U8005 ( .A1(n7062), .A2(keyinput87), .B1(keyinput96), .B2(n7061), 
        .ZN(n7060) );
  OAI221_X1 U8006 ( .B1(n7062), .B2(keyinput87), .C1(n7061), .C2(keyinput96), 
        .A(n7060), .ZN(n7071) );
  AOI22_X1 U8007 ( .A1(n7065), .A2(keyinput25), .B1(n7064), .B2(keyinput66), 
        .ZN(n7063) );
  OAI221_X1 U8008 ( .B1(n7065), .B2(keyinput25), .C1(n7064), .C2(keyinput66), 
        .A(n7063), .ZN(n7070) );
  XOR2_X1 U8009 ( .A(n7066), .B(keyinput101), .Z(n7068) );
  XNOR2_X1 U8010 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .B(keyinput79), .ZN(n7067) );
  NAND2_X1 U8011 ( .A1(n7068), .A2(n7067), .ZN(n7069) );
  NOR4_X1 U8012 ( .A1(n7072), .A2(n7071), .A3(n7070), .A4(n7069), .ZN(n7107)
         );
  AOI22_X1 U8013 ( .A1(n7075), .A2(keyinput111), .B1(n7074), .B2(keyinput91), 
        .ZN(n7073) );
  OAI221_X1 U8014 ( .B1(n7075), .B2(keyinput111), .C1(n7074), .C2(keyinput91), 
        .A(n7073), .ZN(n7088) );
  AOI22_X1 U8015 ( .A1(n7078), .A2(keyinput22), .B1(keyinput113), .B2(n7077), 
        .ZN(n7076) );
  OAI221_X1 U8016 ( .B1(n7078), .B2(keyinput22), .C1(n7077), .C2(keyinput113), 
        .A(n7076), .ZN(n7087) );
  AOI22_X1 U8017 ( .A1(n7081), .A2(keyinput117), .B1(keyinput100), .B2(n7080), 
        .ZN(n7079) );
  OAI221_X1 U8018 ( .B1(n7081), .B2(keyinput117), .C1(n7080), .C2(keyinput100), 
        .A(n7079), .ZN(n7086) );
  AOI22_X1 U8019 ( .A1(n7084), .A2(keyinput6), .B1(keyinput54), .B2(n7083), 
        .ZN(n7082) );
  OAI221_X1 U8020 ( .B1(n7084), .B2(keyinput6), .C1(n7083), .C2(keyinput54), 
        .A(n7082), .ZN(n7085) );
  NOR4_X1 U8021 ( .A1(n7088), .A2(n7087), .A3(n7086), .A4(n7085), .ZN(n7106)
         );
  AOI22_X1 U8022 ( .A1(n7091), .A2(keyinput78), .B1(n7090), .B2(keyinput50), 
        .ZN(n7089) );
  OAI221_X1 U8023 ( .B1(n7091), .B2(keyinput78), .C1(n7090), .C2(keyinput50), 
        .A(n7089), .ZN(n7095) );
  XNOR2_X1 U8024 ( .A(n7092), .B(keyinput37), .ZN(n7094) );
  XOR2_X1 U8025 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .B(keyinput67), .Z(n7093)
         );
  OR3_X1 U8026 ( .A1(n7095), .A2(n7094), .A3(n7093), .ZN(n7104) );
  INV_X1 U8027 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n7098) );
  AOI22_X1 U8028 ( .A1(n7098), .A2(keyinput104), .B1(keyinput28), .B2(n7097), 
        .ZN(n7096) );
  OAI221_X1 U8029 ( .B1(n7098), .B2(keyinput104), .C1(n7097), .C2(keyinput28), 
        .A(n7096), .ZN(n7103) );
  AOI22_X1 U8030 ( .A1(n7101), .A2(keyinput93), .B1(keyinput115), .B2(n7100), 
        .ZN(n7099) );
  OAI221_X1 U8031 ( .B1(n7101), .B2(keyinput93), .C1(n7100), .C2(keyinput115), 
        .A(n7099), .ZN(n7102) );
  NOR3_X1 U8032 ( .A1(n7104), .A2(n7103), .A3(n7102), .ZN(n7105) );
  NAND4_X1 U8033 ( .A1(n7108), .A2(n7107), .A3(n7106), .A4(n7105), .ZN(n7176)
         );
  INV_X1 U8034 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n7111) );
  AOI22_X1 U8035 ( .A1(n7111), .A2(keyinput43), .B1(keyinput110), .B2(n7110), 
        .ZN(n7109) );
  OAI221_X1 U8036 ( .B1(n7111), .B2(keyinput43), .C1(n7110), .C2(keyinput110), 
        .A(n7109), .ZN(n7123) );
  AOI22_X1 U8037 ( .A1(n7114), .A2(keyinput5), .B1(keyinput114), .B2(n7113), 
        .ZN(n7112) );
  OAI221_X1 U8038 ( .B1(n7114), .B2(keyinput5), .C1(n7113), .C2(keyinput114), 
        .A(n7112), .ZN(n7122) );
  AOI22_X1 U8039 ( .A1(n7117), .A2(keyinput76), .B1(n7116), .B2(keyinput108), 
        .ZN(n7115) );
  OAI221_X1 U8040 ( .B1(n7117), .B2(keyinput76), .C1(n7116), .C2(keyinput108), 
        .A(n7115), .ZN(n7121) );
  INV_X1 U8041 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n7119) );
  AOI22_X1 U8042 ( .A1(n7119), .A2(keyinput62), .B1(keyinput119), .B2(n4372), 
        .ZN(n7118) );
  OAI221_X1 U8043 ( .B1(n7119), .B2(keyinput62), .C1(n4372), .C2(keyinput119), 
        .A(n7118), .ZN(n7120) );
  NOR4_X1 U8044 ( .A1(n7123), .A2(n7122), .A3(n7121), .A4(n7120), .ZN(n7174)
         );
  AOI22_X1 U8045 ( .A1(n7126), .A2(keyinput45), .B1(keyinput11), .B2(n7125), 
        .ZN(n7124) );
  OAI221_X1 U8046 ( .B1(n7126), .B2(keyinput45), .C1(n7125), .C2(keyinput11), 
        .A(n7124), .ZN(n7138) );
  INV_X1 U8047 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n7128) );
  AOI22_X1 U8048 ( .A1(n7128), .A2(keyinput42), .B1(keyinput41), .B2(n3829), 
        .ZN(n7127) );
  OAI221_X1 U8049 ( .B1(n7128), .B2(keyinput42), .C1(n3829), .C2(keyinput41), 
        .A(n7127), .ZN(n7137) );
  AOI22_X1 U8050 ( .A1(n7131), .A2(keyinput72), .B1(keyinput52), .B2(n7130), 
        .ZN(n7129) );
  OAI221_X1 U8051 ( .B1(n7131), .B2(keyinput72), .C1(n7130), .C2(keyinput52), 
        .A(n7129), .ZN(n7136) );
  INV_X1 U8052 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n7133) );
  AOI22_X1 U8053 ( .A1(n7134), .A2(keyinput39), .B1(n7133), .B2(keyinput88), 
        .ZN(n7132) );
  OAI221_X1 U8054 ( .B1(n7134), .B2(keyinput39), .C1(n7133), .C2(keyinput88), 
        .A(n7132), .ZN(n7135) );
  NOR4_X1 U8055 ( .A1(n7138), .A2(n7137), .A3(n7136), .A4(n7135), .ZN(n7173)
         );
  AOI22_X1 U8056 ( .A1(n7141), .A2(keyinput107), .B1(n7140), .B2(keyinput12), 
        .ZN(n7139) );
  OAI221_X1 U8057 ( .B1(n7141), .B2(keyinput107), .C1(n7140), .C2(keyinput12), 
        .A(n7139), .ZN(n7154) );
  AOI22_X1 U8058 ( .A1(n7144), .A2(keyinput21), .B1(n7143), .B2(keyinput63), 
        .ZN(n7142) );
  OAI221_X1 U8059 ( .B1(n7144), .B2(keyinput21), .C1(n7143), .C2(keyinput63), 
        .A(n7142), .ZN(n7153) );
  AOI22_X1 U8060 ( .A1(n7147), .A2(keyinput64), .B1(n7146), .B2(keyinput10), 
        .ZN(n7145) );
  OAI221_X1 U8061 ( .B1(n7147), .B2(keyinput64), .C1(n7146), .C2(keyinput10), 
        .A(n7145), .ZN(n7152) );
  INV_X1 U8062 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n7149) );
  AOI22_X1 U8063 ( .A1(n7150), .A2(keyinput16), .B1(n7149), .B2(keyinput1), 
        .ZN(n7148) );
  OAI221_X1 U8064 ( .B1(n7150), .B2(keyinput16), .C1(n7149), .C2(keyinput1), 
        .A(n7148), .ZN(n7151) );
  NOR4_X1 U8065 ( .A1(n7154), .A2(n7153), .A3(n7152), .A4(n7151), .ZN(n7172)
         );
  INV_X1 U8066 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n7156) );
  AOI22_X1 U8067 ( .A1(n7157), .A2(keyinput19), .B1(keyinput97), .B2(n7156), 
        .ZN(n7155) );
  OAI221_X1 U8068 ( .B1(n7157), .B2(keyinput19), .C1(n7156), .C2(keyinput97), 
        .A(n7155), .ZN(n7170) );
  AOI22_X1 U8069 ( .A1(n7160), .A2(keyinput55), .B1(n7159), .B2(keyinput120), 
        .ZN(n7158) );
  OAI221_X1 U8070 ( .B1(n7160), .B2(keyinput55), .C1(n7159), .C2(keyinput120), 
        .A(n7158), .ZN(n7169) );
  AOI22_X1 U8071 ( .A1(n7163), .A2(keyinput33), .B1(n7162), .B2(keyinput47), 
        .ZN(n7161) );
  OAI221_X1 U8072 ( .B1(n7163), .B2(keyinput33), .C1(n7162), .C2(keyinput47), 
        .A(n7161), .ZN(n7168) );
  INV_X1 U8073 ( .A(DATAI_17_), .ZN(n7165) );
  AOI22_X1 U8074 ( .A1(n7166), .A2(keyinput0), .B1(keyinput32), .B2(n7165), 
        .ZN(n7164) );
  OAI221_X1 U8075 ( .B1(n7166), .B2(keyinput0), .C1(n7165), .C2(keyinput32), 
        .A(n7164), .ZN(n7167) );
  NOR4_X1 U8076 ( .A1(n7170), .A2(n7169), .A3(n7168), .A4(n7167), .ZN(n7171)
         );
  NAND4_X1 U8077 ( .A1(n7174), .A2(n7173), .A3(n7172), .A4(n7171), .ZN(n7175)
         );
  AOI211_X1 U8078 ( .C1(keyinput7), .C2(n7177), .A(n7176), .B(n7175), .ZN(
        n7178) );
  NAND4_X1 U8079 ( .A1(n7181), .A2(n7180), .A3(n7179), .A4(n7178), .ZN(n7182)
         );
  XNOR2_X1 U8080 ( .A(n7183), .B(n7182), .ZN(U3104) );
  INV_X2 U3569 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6938) );
  CLKBUF_X1 U3588 ( .A(n4279), .Z(n4225) );
  CLKBUF_X1 U3591 ( .A(n3406), .Z(n4188) );
  CLKBUF_X1 U3691 ( .A(n3448), .Z(n4328) );
  CLKBUF_X2 U3702 ( .A(n3434), .Z(n4698) );
  CLKBUF_X1 U3703 ( .A(n4271), .Z(n4252) );
endmodule

