

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, 
        DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, 
        DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, 
        DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, 
        DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, 
        DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, 
        DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_,
         DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_,
         DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_,
         DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_,
         DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_,
         DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
         HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN,
         P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN,
         P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN,
         P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN,
         P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN,
         P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN,
         P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN,
         P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN,
         P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN,
         P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
         P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
         P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
         P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
         P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
         P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
         P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
         P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
         P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
         P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
         P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN,
         P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
         P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
         P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
         P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN,
         P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
         P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
         P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN,
         P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
         P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
         P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN,
         P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
         P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
         P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN,
         P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN,
         P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN,
         P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN,
         P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN,
         P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
         P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
         P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN,
         P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
         P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
         P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN,
         P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
         P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
         P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN,
         P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
         P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
         P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
         P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
         P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n10951, n10952, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
         n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484,
         n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492,
         n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500,
         n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508,
         n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516,
         n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
         n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
         n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540,
         n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
         n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556,
         n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564,
         n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572,
         n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580,
         n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588,
         n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
         n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
         n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612,
         n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
         n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628,
         n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636,
         n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644,
         n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652,
         n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660,
         n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
         n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
         n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684,
         n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
         n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700,
         n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708,
         n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716,
         n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724,
         n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732,
         n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
         n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
         n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756,
         n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
         n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772,
         n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780,
         n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788,
         n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796,
         n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804,
         n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
         n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
         n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828,
         n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
         n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844,
         n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852,
         n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860,
         n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868,
         n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876,
         n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884,
         n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
         n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900,
         n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
         n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916,
         n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924,
         n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932,
         n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940,
         n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
         n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956,
         n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
         n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972,
         n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
         n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988,
         n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996,
         n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004,
         n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012,
         n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
         n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028,
         n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
         n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044,
         n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
         n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060,
         n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068,
         n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076,
         n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084,
         n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092,
         n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100,
         n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
         n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116,
         n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
         n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
         n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140,
         n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148,
         n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156,
         n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164,
         n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172,
         n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
         n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188,
         n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
         n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
         n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212,
         n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220,
         n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228,
         n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
         n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244,
         n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252,
         n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260,
         n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268,
         n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276,
         n22277, n22278, n22279;

  AOI221_X1 U11058 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17974), .C1(
        n17973), .C2(n17974), .A(n17972), .ZN(n21175) );
  INV_X2 U11059 ( .A(n21419), .ZN(n14073) );
  NAND2_X1 U11060 ( .A1(n12312), .A2(n12311), .ZN(n15605) );
  OR3_X1 U11061 ( .A1(n13858), .A2(n14073), .A3(n11584), .ZN(n21483) );
  OAI211_X1 U11062 ( .C1(n12657), .C2(n12656), .A(n21206), .B(n21205), .ZN(
        n20786) );
  NAND2_X1 U11063 ( .A1(n12721), .A2(n12651), .ZN(n12660) );
  NAND2_X1 U11064 ( .A1(n11363), .A2(n11805), .ZN(n11832) );
  NAND2_X1 U11065 ( .A1(n11755), .A2(n11813), .ZN(n11366) );
  OR2_X1 U11066 ( .A1(n11793), .A2(n11792), .ZN(n11794) );
  INV_X2 U11067 ( .A(n15490), .ZN(n19381) );
  CLKBUF_X2 U11068 ( .A(n13305), .Z(n10958) );
  XNOR2_X1 U11069 ( .A(n11110), .B(n11781), .ZN(n14382) );
  INV_X1 U11070 ( .A(n14320), .ZN(n10965) );
  CLKBUF_X3 U11071 ( .A(n12482), .Z(n17656) );
  INV_X2 U11072 ( .A(n17406), .ZN(n10970) );
  INV_X2 U11073 ( .A(n12572), .ZN(n17489) );
  CLKBUF_X2 U11074 ( .A(n12512), .Z(n17599) );
  CLKBUF_X2 U11075 ( .A(n12517), .Z(n17536) );
  AND2_X1 U11076 ( .A1(n14502), .A2(n13145), .ZN(n13706) );
  AND2_X1 U11077 ( .A1(n13134), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13605) );
  CLKBUF_X2 U11078 ( .A(n11515), .Z(n12049) );
  INV_X2 U11079 ( .A(n11395), .ZN(n13301) );
  CLKBUF_X2 U11080 ( .A(n11460), .Z(n12360) );
  AND2_X1 U11081 ( .A1(n13127), .A2(n13335), .ZN(n13598) );
  AND2_X1 U11082 ( .A1(n13335), .A2(n13125), .ZN(n13155) );
  AND2_X1 U11083 ( .A1(n13335), .A2(n13124), .ZN(n13599) );
  BUF_X1 U11084 ( .A(n12557), .Z(n17510) );
  NOR2_X1 U11085 ( .A1(n12434), .A2(n12430), .ZN(n12475) );
  CLKBUF_X3 U11086 ( .A(n12518), .Z(n10960) );
  NAND2_X1 U11087 ( .A1(n20784), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12434) );
  INV_X1 U11088 ( .A(n11682), .ZN(n12400) );
  AND2_X1 U11089 ( .A1(n11709), .A2(n11680), .ZN(n11683) );
  NOR2_X1 U11090 ( .A1(n13015), .A2(n13014), .ZN(n13020) );
  INV_X1 U11092 ( .A(n11680), .ZN(n11700) );
  AND2_X1 U11093 ( .A1(n11491), .A2(n11490), .ZN(n11502) );
  AND2_X1 U11095 ( .A1(n11421), .A2(n11422), .ZN(n11503) );
  AND2_X1 U11096 ( .A1(n11417), .A2(n14270), .ZN(n11722) );
  BUF_X1 U11097 ( .A(n11840), .Z(n10976) );
  AND2_X1 U11098 ( .A1(n11166), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11418) );
  OAI22_X2 U11099 ( .A1(n20066), .A2(n14567), .B1(n17001), .B2(n14566), .ZN(
        n22040) );
  NAND2_X2 U11100 ( .A1(n20021), .A2(n15727), .ZN(n14566) );
  AND2_X1 U11101 ( .A1(n11411), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11420) );
  AND2_X1 U11102 ( .A1(n14286), .A2(n21655), .ZN(n11364) );
  INV_X1 U11103 ( .A(n15264), .ZN(n13108) );
  INV_X1 U11104 ( .A(n13462), .ZN(n13134) );
  CLKBUF_X3 U11105 ( .A(n13108), .Z(n15556) );
  CLKBUF_X3 U11106 ( .A(n13146), .Z(n13492) );
  AND2_X1 U11107 ( .A1(n13136), .A2(n13511), .ZN(n14512) );
  AND2_X1 U11108 ( .A1(n14986), .A2(n14984), .ZN(n14989) );
  NAND2_X1 U11109 ( .A1(n11680), .A2(n11682), .ZN(n11689) );
  AND3_X1 U11110 ( .A1(n13041), .A2(n14136), .A3(n13040), .ZN(n13965) );
  NOR2_X1 U11111 ( .A1(n16201), .A2(n13426), .ZN(n13469) );
  AND2_X2 U11112 ( .A1(n13492), .A2(n13511), .ZN(n13707) );
  OR2_X1 U11114 ( .A1(n20518), .A2(n11194), .ZN(n11192) );
  AND2_X1 U11115 ( .A1(n11686), .A2(n14410), .ZN(n11702) );
  NAND2_X1 U11116 ( .A1(n14250), .A2(n12787), .ZN(n12797) );
  AND4_X2 U11118 ( .A1(n11459), .A2(n11458), .A3(n11457), .A4(n11456), .ZN(
        n11686) );
  INV_X1 U11119 ( .A(n11573), .ZN(n14568) );
  NOR2_X1 U11120 ( .A1(n16203), .A2(n16202), .ZN(n16201) );
  AND2_X1 U11121 ( .A1(n15080), .A2(n15079), .ZN(n16651) );
  INV_X1 U11122 ( .A(n18087), .ZN(n18059) );
  INV_X1 U11124 ( .A(n11023), .ZN(n15578) );
  OR2_X1 U11125 ( .A1(n16284), .A2(n16283), .ZN(n16286) );
  NOR2_X1 U11126 ( .A1(n11006), .A2(n18371), .ZN(n18370) );
  AND2_X1 U11127 ( .A1(n14339), .A2(n10997), .ZN(n14681) );
  CLKBUF_X2 U11128 ( .A(n13024), .Z(n14142) );
  INV_X1 U11129 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13511) );
  NOR2_X1 U11130 ( .A1(n21240), .A2(n20161), .ZN(n20502) );
  INV_X1 U11131 ( .A(n17927), .ZN(n18061) );
  NAND2_X1 U11132 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20809) );
  AND2_X1 U11133 ( .A1(n11679), .A2(n11031), .ZN(n11179) );
  BUF_X1 U11134 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11531) );
  NAND2_X1 U11135 ( .A1(n14469), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13462) );
  OR2_X1 U11136 ( .A1(n15663), .A2(n21630), .ZN(n10951) );
  AND2_X1 U11138 ( .A1(n11685), .A2(n12777), .ZN(n10952) );
  NAND2_X2 U11139 ( .A1(n14306), .A2(n14305), .ZN(n14304) );
  OAI21_X2 U11140 ( .B1(n16450), .B2(n16401), .A(n16400), .ZN(n16634) );
  NOR2_X2 U11141 ( .A1(n10984), .A2(n16254), .ZN(n16247) );
  AND2_X1 U11142 ( .A1(n11418), .A2(n11420), .ZN(n11515) );
  NOR2_X2 U11143 ( .A1(n17997), .A2(n12542), .ZN(n17973) );
  AOI211_X2 U11144 ( .C1(n12747), .C2(n21119), .A(n21065), .B(n21079), .ZN(
        n21066) );
  NOR2_X2 U11145 ( .A1(n14998), .A2(n18244), .ZN(n15006) );
  XNOR2_X2 U11146 ( .A(n14324), .B(n11202), .ZN(n14998) );
  AND2_X2 U11147 ( .A1(n14989), .A2(n14988), .ZN(n19185) );
  NOR3_X2 U11148 ( .A1(n16120), .A2(n10966), .A3(n15517), .ZN(n15535) );
  AND2_X2 U11149 ( .A1(n14989), .A2(n17101), .ZN(n15095) );
  AND2_X2 U11150 ( .A1(n14987), .A2(n14988), .ZN(n15096) );
  NOR2_X2 U11151 ( .A1(n16369), .A2(n16370), .ZN(n16368) );
  NOR2_X2 U11152 ( .A1(n21032), .A2(n12897), .ZN(n21062) );
  XNOR2_X2 U11153 ( .A(n15134), .B(n15135), .ZN(n15133) );
  NOR2_X2 U11154 ( .A1(n20798), .A2(n20786), .ZN(n12695) );
  NOR2_X2 U11155 ( .A1(n12876), .A2(n11387), .ZN(n15818) );
  NOR2_X2 U11156 ( .A1(n15838), .A2(n12874), .ZN(n12876) );
  INV_X2 U11158 ( .A(n10952), .ZN(n10954) );
  AOI211_X2 U11159 ( .C1(n17163), .C2(n16107), .A(n15484), .B(n15483), .ZN(
        n15485) );
  XNOR2_X1 U11160 ( .A(n17896), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10956) );
  NAND2_X2 U11161 ( .A1(n11772), .A2(n11771), .ZN(n11822) );
  NOR2_X2 U11162 ( .A1(n15207), .A2(n16265), .ZN(n16255) );
  AND2_X1 U11164 ( .A1(n13495), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13305) );
  XNOR2_X2 U11165 ( .A(n12540), .B(n17718), .ZN(n18018) );
  AND3_X4 U11166 ( .A1(n11250), .A2(n11035), .A3(n11249), .ZN(n17718) );
  AND2_X4 U11167 ( .A1(n13143), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13525) );
  OAI22_X1 U11168 ( .A1(n15822), .A2(n15821), .B1(n15820), .B2(n15819), .ZN(
        n15967) );
  AND2_X1 U11169 ( .A1(n11379), .A2(n12867), .ZN(n11378) );
  OR2_X1 U11170 ( .A1(n11381), .A2(n11380), .ZN(n11379) );
  AND2_X1 U11171 ( .A1(n15890), .A2(n12859), .ZN(n11381) );
  NOR2_X1 U11172 ( .A1(n19984), .A2(n12858), .ZN(n15890) );
  NOR3_X1 U11173 ( .A1(n15310), .A2(n10966), .A3(n16491), .ZN(n15534) );
  INV_X4 U11174 ( .A(n19993), .ZN(n20015) );
  NOR2_X1 U11175 ( .A1(n17785), .A2(n12553), .ZN(n17834) );
  AND2_X1 U11176 ( .A1(n12548), .A2(n11246), .ZN(n11245) );
  INV_X1 U11177 ( .A(n21111), .ZN(n21202) );
  NAND2_X1 U11178 ( .A1(n11366), .A2(n11779), .ZN(n11831) );
  INV_X2 U11179 ( .A(n21185), .ZN(n20874) );
  NAND2_X1 U11180 ( .A1(n19946), .A2(n15576), .ZN(n15726) );
  NAND2_X1 U11181 ( .A1(n10964), .A2(n11109), .ZN(n11784) );
  NAND2_X2 U11183 ( .A1(n13965), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15264) );
  INV_X1 U11184 ( .A(n12730), .ZN(n18811) );
  INV_X2 U11185 ( .A(n13837), .ZN(n11085) );
  CLKBUF_X2 U11186 ( .A(n12991), .Z(n13968) );
  INV_X2 U11188 ( .A(n11686), .ZN(n11688) );
  AND4_X1 U11189 ( .A1(n11485), .A2(n11484), .A3(n11483), .A4(n11482), .ZN(
        n11491) );
  INV_X4 U11190 ( .A(n20184), .ZN(n17628) );
  CLKBUF_X2 U11191 ( .A(n12517), .Z(n17665) );
  CLKBUF_X2 U11192 ( .A(n12518), .Z(n10980) );
  CLKBUF_X2 U11193 ( .A(n11722), .Z(n12315) );
  CLKBUF_X2 U11194 ( .A(n11503), .Z(n12268) );
  CLKBUF_X2 U11195 ( .A(n11741), .Z(n11981) );
  INV_X2 U11196 ( .A(n11428), .ZN(n10971) );
  CLKBUF_X1 U11197 ( .A(n13134), .Z(n10959) );
  NOR2_X2 U11198 ( .A1(n12431), .A2(n11244), .ZN(n12465) );
  NOR2_X1 U11199 ( .A1(n12434), .A2(n12432), .ZN(n12481) );
  INV_X2 U11200 ( .A(n21161), .ZN(n10961) );
  NOR2_X1 U11201 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12909) );
  INV_X4 U11202 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20808) );
  INV_X1 U11203 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12698) );
  NAND2_X1 U11204 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20821) );
  INV_X1 U11205 ( .A(n20809), .ZN(n10962) );
  OR2_X1 U11206 ( .A1(n16347), .A2(n16767), .ZN(n11284) );
  NOR2_X1 U11207 ( .A1(n15805), .A2(n15804), .ZN(n15806) );
  INV_X1 U11208 ( .A(n15200), .ZN(n12077) );
  OR2_X1 U11209 ( .A1(n15914), .A2(n12857), .ZN(n19984) );
  OAI21_X1 U11210 ( .B1(n15139), .B2(n11050), .A(n18250), .ZN(n15318) );
  NAND2_X1 U11211 ( .A1(n11125), .A2(n11348), .ZN(n17099) );
  OR2_X1 U11212 ( .A1(n15888), .A2(n12863), .ZN(n15902) );
  NAND2_X1 U11213 ( .A1(n11026), .A2(n11117), .ZN(n14687) );
  AND2_X1 U11214 ( .A1(n11671), .A2(n11670), .ZN(n15931) );
  OR2_X1 U11215 ( .A1(n20015), .A2(n12860), .ZN(n15909) );
  OR2_X1 U11216 ( .A1(n20015), .A2(n21282), .ZN(n19983) );
  AND2_X1 U11217 ( .A1(n11192), .A2(n11064), .ZN(n20555) );
  AND2_X1 U11218 ( .A1(n11196), .A2(n11195), .ZN(n10988) );
  NAND2_X1 U11219 ( .A1(n17834), .A2(n21101), .ZN(n17833) );
  NAND2_X1 U11220 ( .A1(n11333), .A2(n11321), .ZN(n11325) );
  OAI21_X1 U11221 ( .B1(n12820), .B2(n11371), .A(n11914), .ZN(n14657) );
  AND2_X1 U11222 ( .A1(n15422), .A2(n15421), .ZN(n11333) );
  NAND2_X1 U11223 ( .A1(n12549), .A2(n11245), .ZN(n11247) );
  NAND2_X1 U11224 ( .A1(n20626), .A2(n18081), .ZN(n18002) );
  NAND2_X1 U11225 ( .A1(n14243), .A2(n13122), .ZN(n14339) );
  OR2_X1 U11226 ( .A1(n12661), .A2(n21270), .ZN(n17951) );
  OAI21_X2 U11227 ( .B1(n20096), .B2(P3_STATE2_REG_0__SCAN_IN), .A(n21270), 
        .ZN(n18087) );
  INV_X1 U11228 ( .A(n11906), .ZN(n11904) );
  XNOR2_X1 U11229 ( .A(n11880), .B(n11888), .ZN(n12808) );
  INV_X1 U11230 ( .A(n19308), .ZN(n15109) );
  CLKBUF_X1 U11231 ( .A(n14298), .Z(n16073) );
  NAND2_X1 U11232 ( .A1(n14215), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14250) );
  AND2_X1 U11233 ( .A1(n14987), .A2(n17101), .ZN(n19265) );
  NAND2_X1 U11234 ( .A1(n14999), .A2(n11010), .ZN(n15328) );
  XNOR2_X1 U11235 ( .A(n14170), .B(n14169), .ZN(n19142) );
  AND2_X1 U11236 ( .A1(n14982), .A2(n17101), .ZN(n19232) );
  XNOR2_X1 U11237 ( .A(n11831), .B(n11832), .ZN(n12788) );
  AND2_X1 U11238 ( .A1(n15005), .A2(n14984), .ZN(n14982) );
  NAND2_X1 U11239 ( .A1(n16723), .A2(n16724), .ZN(n16725) );
  AND2_X1 U11240 ( .A1(n15005), .A2(n14985), .ZN(n14983) );
  AND2_X1 U11241 ( .A1(n14986), .A2(n14985), .ZN(n14987) );
  AND2_X1 U11242 ( .A1(n14368), .A2(n11888), .ZN(n11106) );
  NAND2_X1 U11243 ( .A1(n11010), .A2(n15000), .ZN(n15103) );
  NAND2_X1 U11244 ( .A1(n14047), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14049) );
  OR2_X1 U11245 ( .A1(n17999), .A2(n17998), .ZN(n11268) );
  NAND2_X1 U11246 ( .A1(n16738), .A2(n16737), .ZN(n16739) );
  NAND2_X1 U11247 ( .A1(n11794), .A2(n11364), .ZN(n11363) );
  NAND2_X1 U11248 ( .A1(n13724), .A2(n13723), .ZN(n16738) );
  NOR2_X1 U11249 ( .A1(n12541), .A2(n18017), .ZN(n17999) );
  OR2_X1 U11250 ( .A1(n14660), .A2(n11139), .ZN(n21484) );
  NAND3_X1 U11251 ( .A1(n13104), .A2(n13103), .A3(n13102), .ZN(n14324) );
  AND2_X1 U11252 ( .A1(n11189), .A2(n20396), .ZN(n20433) );
  NAND2_X1 U11253 ( .A1(n11784), .A2(n11783), .ZN(n11793) );
  NAND2_X2 U11255 ( .A1(n15794), .A2(n14218), .ZN(n15801) );
  AND2_X1 U11256 ( .A1(n13098), .A2(n14980), .ZN(n18244) );
  NAND2_X1 U11257 ( .A1(n12405), .A2(n12404), .ZN(n15794) );
  NAND2_X1 U11258 ( .A1(n14942), .A2(n11613), .ZN(n19922) );
  NOR2_X2 U11259 ( .A1(n19941), .A2(n11606), .ZN(n14942) );
  NOR2_X2 U11260 ( .A1(n19585), .A2(n19641), .ZN(n19586) );
  NOR2_X2 U11261 ( .A1(n19429), .A2(n19639), .ZN(n19430) );
  NOR2_X2 U11262 ( .A1(n19379), .A2(n19639), .ZN(n19380) );
  NOR2_X2 U11263 ( .A1(n19381), .A2(n19641), .ZN(n19382) );
  OR2_X1 U11264 ( .A1(n18035), .A2(n11251), .ZN(n11250) );
  NOR2_X2 U11265 ( .A1(n19329), .A2(n19639), .ZN(n19330) );
  NOR2_X2 U11266 ( .A1(n19113), .A2(n19639), .ZN(n19114) );
  NAND2_X1 U11267 ( .A1(n11791), .A2(n11790), .ZN(n11792) );
  INV_X2 U11268 ( .A(n11059), .ZN(n10963) );
  OR2_X1 U11269 ( .A1(n15533), .A2(n14873), .ZN(n15358) );
  INV_X1 U11270 ( .A(n14382), .ZN(n10964) );
  NAND2_X1 U11271 ( .A1(n13071), .A2(n13070), .ZN(n13075) );
  NOR2_X1 U11272 ( .A1(n11187), .A2(n20421), .ZN(n11186) );
  OR2_X1 U11273 ( .A1(n13659), .A2(n13653), .ZN(n14927) );
  AOI21_X1 U11274 ( .B1(n14149), .B2(n13652), .A(n13651), .ZN(n13659) );
  OR2_X1 U11275 ( .A1(n13056), .A2(n14714), .ZN(n13057) );
  AND2_X1 U11276 ( .A1(n11720), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11781) );
  AND2_X1 U11277 ( .A1(n13048), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13045) );
  AND2_X1 U11278 ( .A1(n13061), .A2(n13062), .ZN(n13063) );
  AND2_X1 U11279 ( .A1(n11694), .A2(n11108), .ZN(n11107) );
  AND2_X1 U11280 ( .A1(n17880), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17915) );
  AND2_X1 U11281 ( .A1(n11691), .A2(n11692), .ZN(n11713) );
  AND2_X1 U11282 ( .A1(n13021), .A2(n14555), .ZN(n13896) );
  CLKBUF_X1 U11283 ( .A(n12696), .Z(n10972) );
  AND2_X1 U11284 ( .A1(n14160), .A2(n14159), .ZN(n14158) );
  AND2_X1 U11285 ( .A1(n14843), .A2(n15123), .ZN(n11150) );
  NOR2_X2 U11286 ( .A1(n12728), .A2(n12620), .ZN(n12652) );
  AND2_X1 U11287 ( .A1(n15579), .A2(n13950), .ZN(n13861) );
  OR2_X1 U11288 ( .A1(n15578), .A2(n13950), .ZN(n11662) );
  INV_X2 U11289 ( .A(n15264), .ZN(n15285) );
  NAND2_X1 U11290 ( .A1(n13032), .A2(n13031), .ZN(n13812) );
  OR2_X1 U11291 ( .A1(n14101), .A2(n13018), .ZN(n13021) );
  AOI21_X1 U11292 ( .B1(n20156), .B2(n18891), .A(n20602), .ZN(n12728) );
  CLKBUF_X1 U11293 ( .A(n13030), .Z(n14555) );
  NOR2_X1 U11294 ( .A1(n18076), .A2(n12491), .ZN(n18069) );
  NAND3_X1 U11295 ( .A1(n11575), .A2(n11711), .A3(n11574), .ZN(n11697) );
  OR2_X1 U11296 ( .A1(n11385), .A2(n14129), .ZN(n11204) );
  NOR2_X1 U11297 ( .A1(n18077), .A2(n18084), .ZN(n18076) );
  INV_X2 U11298 ( .A(n20693), .ZN(n20667) );
  AND2_X1 U11299 ( .A1(n11701), .A2(n15576), .ZN(n12418) );
  CLKBUF_X1 U11300 ( .A(n12776), .Z(n21274) );
  INV_X2 U11301 ( .A(n11050), .ZN(n10966) );
  CLKBUF_X1 U11302 ( .A(n11709), .Z(n14404) );
  OR2_X2 U11303 ( .A1(n20088), .A2(n20027), .ZN(n20074) );
  OR2_X1 U11304 ( .A1(n13614), .A2(n13613), .ZN(n13867) );
  NAND2_X1 U11305 ( .A1(n13035), .A2(n13579), .ZN(n13011) );
  NAND3_X1 U11306 ( .A1(n12631), .A2(n12630), .A3(n12629), .ZN(n20693) );
  INV_X2 U11307 ( .A(n14727), .ZN(n19642) );
  INV_X2 U11308 ( .A(n13024), .ZN(n19585) );
  NAND2_X1 U11309 ( .A1(n13024), .A2(n14727), .ZN(n13837) );
  INV_X1 U11310 ( .A(n12964), .ZN(n13035) );
  CLKBUF_X2 U11311 ( .A(n13579), .Z(n15490) );
  INV_X1 U11312 ( .A(n13024), .ZN(n10967) );
  NAND2_X1 U11313 ( .A1(n11075), .A2(n11074), .ZN(n12964) );
  INV_X2 U11314 ( .A(U214), .ZN(n20088) );
  NAND2_X1 U11315 ( .A1(n12951), .A2(n12950), .ZN(n12991) );
  AND3_X1 U11316 ( .A1(n10985), .A2(n17743), .A3(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17713) );
  NAND2_X1 U11317 ( .A1(n11079), .A2(n13511), .ZN(n11078) );
  NAND2_X1 U11318 ( .A1(n11077), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11076) );
  MUX2_X1 U11319 ( .A(n12963), .B(n12962), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14129) );
  AND4_X1 U11320 ( .A1(n11495), .A2(n11494), .A3(n11493), .A4(n11492), .ZN(
        n11501) );
  AND4_X1 U11321 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n11500) );
  AND4_X1 U11322 ( .A1(n11442), .A2(n11441), .A3(n11440), .A4(n11439), .ZN(
        n11459) );
  AND4_X1 U11323 ( .A1(n11446), .A2(n11445), .A3(n11444), .A4(n11443), .ZN(
        n11458) );
  AND4_X1 U11324 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(
        n11457) );
  AND4_X1 U11325 ( .A1(n11474), .A2(n11473), .A3(n11472), .A4(n11471), .ZN(
        n11481) );
  CLKBUF_X2 U11326 ( .A(n12452), .Z(n17640) );
  AND4_X1 U11327 ( .A1(n11479), .A2(n11478), .A3(n11477), .A4(n11476), .ZN(
        n11480) );
  AND4_X1 U11328 ( .A1(n13001), .A2(n13000), .A3(n12999), .A4(n12998), .ZN(
        n13002) );
  AND2_X1 U11329 ( .A1(n11197), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10985) );
  AND2_X1 U11330 ( .A1(n11517), .A2(n11522), .ZN(n11118) );
  AND4_X1 U11331 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n11456) );
  INV_X2 U11333 ( .A(n18977), .ZN(U215) );
  CLKBUF_X1 U11334 ( .A(n14088), .Z(n19108) );
  INV_X2 U11335 ( .A(n21704), .ZN(n10969) );
  AND2_X1 U11336 ( .A1(n11199), .A2(n11198), .ZN(n11197) );
  INV_X1 U11337 ( .A(n12451), .ZN(n12572) );
  INV_X1 U11338 ( .A(n11428), .ZN(n12366) );
  NOR2_X1 U11339 ( .A1(n12433), .A2(n12432), .ZN(n12482) );
  NOR2_X1 U11340 ( .A1(n12433), .A2(n20821), .ZN(n12451) );
  BUF_X2 U11341 ( .A(n13141), .Z(n13495) );
  INV_X2 U11342 ( .A(n19756), .ZN(n19816) );
  AND2_X2 U11343 ( .A1(n11421), .A2(n11419), .ZN(n11840) );
  AND3_X1 U11344 ( .A1(n10962), .A2(n20808), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12557) );
  AND2_X1 U11345 ( .A1(n14270), .A2(n11418), .ZN(n11460) );
  OR2_X2 U11346 ( .A1(n12431), .A2(n20821), .ZN(n17598) );
  NOR2_X2 U11347 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17691), .ZN(n21161) );
  INV_X2 U11348 ( .A(n22276), .ZN(n22279) );
  OAI21_X1 U11349 ( .B1(n13793), .B2(n13792), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14088) );
  AND3_X2 U11350 ( .A1(n14487), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13146) );
  CLKBUF_X1 U11351 ( .A(n12698), .Z(n20794) );
  NAND2_X1 U11352 ( .A1(n14469), .A2(n14490), .ZN(n13334) );
  AND2_X2 U11353 ( .A1(n13127), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13128) );
  AND2_X2 U11354 ( .A1(n12909), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13142) );
  AND2_X2 U11355 ( .A1(n13144), .A2(n14490), .ZN(n13141) );
  NAND2_X1 U11356 ( .A1(n12698), .A2(n20784), .ZN(n12433) );
  AND2_X1 U11357 ( .A1(n11376), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11419) );
  AND2_X1 U11358 ( .A1(n11412), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11417) );
  NOR2_X1 U11359 ( .A1(n20221), .A2(n11183), .ZN(n11182) );
  AND2_X1 U11360 ( .A1(n11531), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14269) );
  NAND2_X1 U11361 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21214), .ZN(
        n12432) );
  CLKBUF_X1 U11362 ( .A(n13144), .Z(n14502) );
  NAND2_X2 U11363 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12698), .ZN(
        n12431) );
  INV_X2 U11364 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20784) );
  NOR2_X2 U11365 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21900) );
  INV_X2 U11366 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21214) );
  NOR2_X2 U11367 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14270) );
  AND2_X2 U11368 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16085) );
  AND2_X1 U11369 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13144) );
  NOR2_X2 U11370 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14469) );
  XNOR2_X1 U11372 ( .A(n14049), .B(n12785), .ZN(n14215) );
  NAND2_X2 U11373 ( .A1(n12077), .A2(n12076), .ZN(n15232) );
  NAND2_X1 U11374 ( .A1(n15818), .A2(n15816), .ZN(n15817) );
  NOR2_X2 U11375 ( .A1(n12450), .A2(n12449), .ZN(n20774) );
  OAI211_X1 U11376 ( .C1(n11328), .C2(n11325), .A(n16568), .B(n11323), .ZN(
        n16396) );
  OAI22_X2 U11377 ( .A1(n15882), .A2(n15881), .B1(n19971), .B2(n16041), .ZN(
        n20001) );
  AOI21_X4 U11378 ( .B1(n16635), .B2(n16403), .A(n16402), .ZN(n17176) );
  XNOR2_X2 U11379 ( .A(n16406), .B(n11096), .ZN(n11164) );
  OAI21_X2 U11380 ( .B1(n17176), .B2(n16405), .A(n16404), .ZN(n16406) );
  AOI21_X1 U11381 ( .B1(n18535), .B2(n17202), .A(n11160), .ZN(n17187) );
  OAI21_X2 U11382 ( .B1(n14661), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11733), 
        .ZN(n11754) );
  XNOR2_X1 U11383 ( .A(n14978), .B(n13098), .ZN(n14994) );
  AOI211_X1 U11384 ( .C1(n12799), .C2(n21929), .A(n14373), .B(n14378), .ZN(
        n14375) );
  XNOR2_X2 U11385 ( .A(n11865), .B(n14368), .ZN(n12799) );
  INV_X1 U11386 ( .A(n12788), .ZN(n10974) );
  INV_X1 U11387 ( .A(n10974), .ZN(n10975) );
  BUF_X8 U11388 ( .A(n11840), .Z(n10977) );
  NAND2_X1 U11389 ( .A1(n11419), .A2(n16085), .ZN(n11428) );
  INV_X1 U11390 ( .A(n13457), .ZN(n10979) );
  NOR2_X4 U11391 ( .A1(n20770), .A2(n20769), .ZN(n20767) );
  NOR2_X1 U11392 ( .A1(n12430), .A2(n20809), .ZN(n12518) );
  INV_X1 U11393 ( .A(n17951), .ZN(n10981) );
  INV_X1 U11394 ( .A(n17951), .ZN(n10982) );
  OAI21_X1 U11395 ( .B1(n13583), .B2(n13029), .A(n13028), .ZN(n13038) );
  OR2_X1 U11396 ( .A1(n12400), .A2(n21655), .ZN(n11777) );
  NAND2_X1 U11397 ( .A1(n11087), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13022) );
  NAND2_X1 U11398 ( .A1(n13055), .A2(n11084), .ZN(n11087) );
  NAND2_X1 U11399 ( .A1(n11086), .A2(n11019), .ZN(n11084) );
  NAND2_X1 U11400 ( .A1(n11377), .A2(n12866), .ZN(n15868) );
  NAND2_X1 U11401 ( .A1(n11570), .A2(n11408), .ZN(n11137) );
  NAND2_X1 U11402 ( .A1(n11106), .A2(n11889), .ZN(n11906) );
  BUF_X1 U11403 ( .A(n11447), .Z(n12367) );
  AOI21_X1 U11404 ( .B1(n11822), .B2(n11821), .A(n12842), .ZN(n11813) );
  NOR2_X1 U11405 ( .A1(n11693), .A2(n14268), .ZN(n11108) );
  INV_X1 U11406 ( .A(n11093), .ZN(n11091) );
  NAND2_X1 U11407 ( .A1(n11081), .A2(n12992), .ZN(n11080) );
  AOI21_X1 U11408 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19255), .A(
        n13513), .ZN(n13515) );
  NOR2_X1 U11409 ( .A1(n13512), .A2(n13557), .ZN(n13513) );
  INV_X1 U11410 ( .A(n14136), .ZN(n13903) );
  NOR2_X1 U11411 ( .A1(n20639), .A2(n12508), .ZN(n12525) );
  NAND2_X1 U11412 ( .A1(n16079), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12381) );
  XNOR2_X1 U11413 ( .A(n12823), .B(n11945), .ZN(n12833) );
  OR2_X1 U11414 ( .A1(n20015), .A2(n15933), .ZN(n12854) );
  INV_X1 U11415 ( .A(n12846), .ZN(n11778) );
  NOR2_X1 U11416 ( .A1(n11121), .A2(n11120), .ZN(n11119) );
  NAND2_X1 U11417 ( .A1(n15488), .A2(n15489), .ZN(n15531) );
  INV_X1 U11418 ( .A(n16348), .ZN(n11340) );
  NAND2_X1 U11419 ( .A1(n10986), .A2(n11322), .ZN(n11324) );
  NOR2_X1 U11420 ( .A1(n16709), .A2(n11290), .ZN(n11289) );
  INV_X1 U11421 ( .A(n16690), .ZN(n11290) );
  AND2_X1 U11422 ( .A1(n15147), .A2(n11279), .ZN(n11278) );
  INV_X1 U11423 ( .A(n14845), .ZN(n11279) );
  NAND2_X1 U11424 ( .A1(n13116), .A2(n13115), .ZN(n11304) );
  OR2_X1 U11425 ( .A1(n17101), .A2(n14557), .ZN(n13116) );
  INV_X1 U11426 ( .A(n13682), .ZN(n13775) );
  AND2_X1 U11427 ( .A1(n11021), .A2(n19585), .ZN(n13748) );
  AND2_X1 U11428 ( .A1(n13591), .A2(n13968), .ZN(n13025) );
  NOR2_X1 U11429 ( .A1(n20631), .A2(n12527), .ZN(n12539) );
  OAI21_X1 U11430 ( .B1(n18012), .B2(n18011), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12688) );
  NAND2_X1 U11431 ( .A1(n11143), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n11142) );
  INV_X2 U11432 ( .A(n12330), .ZN(n12386) );
  AND2_X1 U11433 ( .A1(n21922), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12385) );
  INV_X1 U11434 ( .A(n11136), .ZN(n11135) );
  NAND2_X1 U11435 ( .A1(n14687), .A2(n11382), .ZN(n19957) );
  NOR2_X1 U11436 ( .A1(n19960), .A2(n11383), .ZN(n11382) );
  INV_X1 U11437 ( .A(n12822), .ZN(n11383) );
  CLKBUF_X2 U11438 ( .A(n13654), .Z(n15550) );
  NAND2_X1 U11439 ( .A1(n20396), .A2(n11001), .ZN(n11193) );
  CLKBUF_X1 U11441 ( .A(n12463), .Z(n20196) );
  NAND2_X1 U11442 ( .A1(n11142), .A2(n21627), .ZN(n15590) );
  AND2_X1 U11443 ( .A1(n17151), .A2(n16832), .ZN(n17190) );
  OR2_X1 U11444 ( .A1(n11732), .A2(n11731), .ZN(n12789) );
  NAND2_X1 U11445 ( .A1(n14410), .A2(n11699), .ZN(n11703) );
  AND2_X1 U11446 ( .A1(n14270), .A2(n11421), .ZN(n11475) );
  AND4_X1 U11447 ( .A1(n15324), .A2(n15323), .A3(n15322), .A4(n15321), .ZN(
        n15335) );
  NAND2_X1 U11448 ( .A1(n13061), .A2(n13039), .ZN(n13048) );
  NOR2_X1 U11449 ( .A1(n13038), .A2(n13037), .ZN(n13039) );
  NAND2_X1 U11450 ( .A1(n13054), .A2(n19642), .ZN(n11088) );
  NAND2_X1 U11451 ( .A1(n13896), .A2(n13031), .ZN(n13051) );
  AND2_X1 U11452 ( .A1(n11902), .A2(n11901), .ZN(n11905) );
  CLKBUF_X1 U11453 ( .A(n11516), .Z(n12296) );
  NOR2_X1 U11454 ( .A1(n15576), .A2(n21922), .ZN(n11824) );
  AND2_X1 U11455 ( .A1(n11927), .A2(n11926), .ZN(n11939) );
  INV_X1 U11456 ( .A(n11905), .ZN(n11903) );
  CLKBUF_X3 U11457 ( .A(n11475), .Z(n12340) );
  AOI21_X1 U11458 ( .B1(n11701), .B2(n11700), .A(n11681), .ZN(n12766) );
  NAND2_X1 U11459 ( .A1(n11272), .A2(n16315), .ZN(n11271) );
  INV_X1 U11460 ( .A(n16577), .ZN(n11272) );
  NAND2_X1 U11461 ( .A1(n15474), .A2(n15473), .ZN(n15478) );
  INV_X1 U11462 ( .A(n15472), .ZN(n15474) );
  AND2_X1 U11463 ( .A1(n15117), .A2(n15116), .ZN(n15120) );
  INV_X1 U11464 ( .A(n13075), .ZN(n13072) );
  NOR2_X1 U11465 ( .A1(n19478), .A2(n11083), .ZN(n11082) );
  NAND2_X1 U11466 ( .A1(n12952), .A2(n12953), .ZN(n13899) );
  INV_X2 U11467 ( .A(n13334), .ZN(n13476) );
  NAND2_X1 U11468 ( .A1(n14129), .A2(n19534), .ZN(n13015) );
  NAND2_X1 U11469 ( .A1(n12473), .A2(n20644), .ZN(n12508) );
  NAND2_X1 U11470 ( .A1(n15596), .A2(n11360), .ZN(n11359) );
  INV_X1 U11471 ( .A(n15606), .ZN(n11360) );
  AND2_X1 U11472 ( .A1(n11362), .A2(n15630), .ZN(n11361) );
  INV_X1 U11473 ( .A(n12381), .ZN(n12353) );
  AND2_X1 U11474 ( .A1(n15670), .A2(n12247), .ZN(n11362) );
  NOR2_X1 U11475 ( .A1(n11357), .A2(n11356), .ZN(n11355) );
  INV_X1 U11476 ( .A(n15711), .ZN(n11356) );
  NAND2_X1 U11477 ( .A1(n11350), .A2(n15201), .ZN(n11349) );
  INV_X1 U11478 ( .A(n11351), .ZN(n11350) );
  NAND2_X1 U11479 ( .A1(n19928), .A2(n15672), .ZN(n11172) );
  NAND2_X1 U11480 ( .A1(n12871), .A2(n20009), .ZN(n15826) );
  INV_X1 U11481 ( .A(n12866), .ZN(n11380) );
  INV_X1 U11482 ( .A(n15225), .ZN(n12853) );
  NOR2_X1 U11483 ( .A1(n11170), .A2(n14649), .ZN(n11169) );
  INV_X1 U11484 ( .A(n14653), .ZN(n11170) );
  INV_X1 U11485 ( .A(n14426), .ZN(n11168) );
  OR2_X1 U11486 ( .A1(n11768), .A2(n11767), .ZN(n12790) );
  OR2_X1 U11487 ( .A1(n11747), .A2(n11746), .ZN(n12846) );
  INV_X1 U11488 ( .A(n11721), .ZN(n11109) );
  XNOR2_X1 U11489 ( .A(n11758), .B(n11757), .ZN(n11374) );
  AOI21_X1 U11490 ( .B1(n11408), .B2(n11569), .A(n11051), .ZN(n11138) );
  NOR2_X1 U11491 ( .A1(n15444), .A2(n15309), .ZN(n15488) );
  NAND2_X1 U11492 ( .A1(n15344), .A2(n15345), .ZN(n15533) );
  NAND2_X1 U11493 ( .A1(n13409), .A2(n16206), .ZN(n13425) );
  NAND2_X1 U11494 ( .A1(n11311), .A2(n16219), .ZN(n11310) );
  NAND2_X1 U11495 ( .A1(n11313), .A2(n13408), .ZN(n11312) );
  AND2_X1 U11496 ( .A1(n16255), .A2(n11065), .ZN(n16223) );
  INV_X1 U11497 ( .A(n16235), .ZN(n11314) );
  OAI21_X1 U11498 ( .B1(n11278), .B2(n11277), .A(n14880), .ZN(n11276) );
  INV_X1 U11499 ( .A(n14712), .ZN(n11241) );
  XNOR2_X1 U11500 ( .A(n14326), .B(n11203), .ZN(n14325) );
  INV_X1 U11501 ( .A(n14327), .ZN(n11203) );
  INV_X1 U11502 ( .A(n16570), .ZN(n11321) );
  NAND2_X1 U11503 ( .A1(n11295), .A2(n16334), .ZN(n11294) );
  INV_X1 U11504 ( .A(n15192), .ZN(n11295) );
  NAND2_X1 U11505 ( .A1(n11209), .A2(n15179), .ZN(n11208) );
  INV_X1 U11506 ( .A(n14971), .ZN(n11209) );
  NOR2_X1 U11507 ( .A1(n14905), .A2(n14906), .ZN(n14915) );
  INV_X1 U11508 ( .A(n14831), .ZN(n11214) );
  INV_X1 U11509 ( .A(n15351), .ZN(n11092) );
  INV_X1 U11510 ( .A(n11332), .ZN(n11331) );
  NAND2_X1 U11511 ( .A1(n11091), .A2(n15351), .ZN(n11090) );
  INV_X1 U11512 ( .A(n15372), .ZN(n11330) );
  AND2_X1 U11513 ( .A1(n11289), .A2(n11287), .ZN(n11286) );
  INV_X1 U11514 ( .A(n16136), .ZN(n11287) );
  INV_X1 U11515 ( .A(n16725), .ZN(n11288) );
  NOR2_X1 U11516 ( .A1(n14706), .A2(n11216), .ZN(n11215) );
  INV_X1 U11517 ( .A(n14853), .ZN(n11216) );
  NOR2_X1 U11518 ( .A1(n15468), .A2(n11129), .ZN(n11128) );
  INV_X1 U11519 ( .A(n15300), .ZN(n15294) );
  NAND2_X1 U11520 ( .A1(n17099), .A2(n15051), .ZN(n15134) );
  AOI221_X1 U11521 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n13515), 
        .C1(n13917), .C2(n13515), .A(n13514), .ZN(n13844) );
  NAND2_X1 U11522 ( .A1(n14986), .A2(n11010), .ZN(n15007) );
  AND4_X1 U11523 ( .A1(n12936), .A2(n12935), .A3(n12934), .A4(n12933), .ZN(
        n12937) );
  NAND2_X1 U11524 ( .A1(n12914), .A2(n13511), .ZN(n11075) );
  NAND2_X1 U11525 ( .A1(n12919), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11074) );
  INV_X1 U11526 ( .A(n17847), .ZN(n11256) );
  NAND2_X1 U11527 ( .A1(n17833), .A2(n12554), .ZN(n12555) );
  NAND2_X1 U11528 ( .A1(n18031), .A2(n12682), .ZN(n12684) );
  XNOR2_X1 U11529 ( .A(n12671), .B(n11097), .ZN(n12670) );
  INV_X1 U11530 ( .A(n20644), .ZN(n11097) );
  NOR2_X1 U11531 ( .A1(n20667), .A2(n18851), .ZN(n12721) );
  NOR2_X1 U11532 ( .A1(n12660), .A2(n20796), .ZN(n16807) );
  NOR2_X1 U11533 ( .A1(n20784), .A2(n20817), .ZN(n12425) );
  NOR4_X1 U11534 ( .A1(n12730), .A2(n12649), .A3(n12657), .A4(n12734), .ZN(
        n12696) );
  NAND2_X1 U11535 ( .A1(n11676), .A2(n11140), .ZN(n11139) );
  INV_X1 U11536 ( .A(n11141), .ZN(n11140) );
  AND2_X1 U11537 ( .A1(n12359), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12388) );
  AND2_X1 U11538 ( .A1(n12199), .A2(n12198), .ZN(n15683) );
  CLKBUF_X1 U11539 ( .A(n15684), .Z(n15685) );
  INV_X1 U11540 ( .A(n15703), .ZN(n15766) );
  CLKBUF_X1 U11541 ( .A(n15702), .Z(n15703) );
  OR2_X1 U11542 ( .A1(n14080), .A2(n14077), .ZN(n15942) );
  INV_X1 U11543 ( .A(n14684), .ZN(n11117) );
  OR2_X1 U11544 ( .A1(n14080), .A2(n15575), .ZN(n21368) );
  NAND2_X1 U11545 ( .A1(n11365), .A2(n11779), .ZN(n11816) );
  INV_X1 U11546 ( .A(n11366), .ZN(n11365) );
  NAND2_X1 U11547 ( .A1(n21829), .A2(n21655), .ZN(n11855) );
  INV_X1 U11548 ( .A(n14570), .ZN(n21783) );
  NAND2_X1 U11549 ( .A1(n11683), .A2(n11389), .ZN(n13956) );
  INV_X1 U11550 ( .A(n13956), .ZN(n16079) );
  NOR2_X1 U11551 ( .A1(n21907), .A2(n21783), .ZN(n21858) );
  NOR2_X1 U11552 ( .A1(n21850), .A2(n21783), .ZN(n21914) );
  NAND2_X1 U11553 ( .A1(n16073), .A2(n14379), .ZN(n21868) );
  NAND2_X1 U11554 ( .A1(n15311), .A2(n15312), .ZN(n15444) );
  NOR2_X1 U11555 ( .A1(n15433), .A2(n15306), .ZN(n15307) );
  NAND2_X1 U11556 ( .A1(n15427), .A2(n15428), .ZN(n15433) );
  NAND2_X1 U11557 ( .A1(n15398), .A2(n15399), .ZN(n15424) );
  NAND2_X1 U11558 ( .A1(n15353), .A2(n15354), .ZN(n15374) );
  NAND2_X1 U11559 ( .A1(n18370), .A2(n16321), .ZN(n16576) );
  AND3_X1 U11560 ( .A1(n13737), .A2(n13736), .A3(n13735), .ZN(n16709) );
  AND2_X2 U11561 ( .A1(n13023), .A2(n19534), .ZN(n14136) );
  NOR2_X1 U11562 ( .A1(n15496), .A2(n16111), .ZN(n14713) );
  NAND2_X1 U11563 ( .A1(n15452), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15496) );
  NAND2_X1 U11564 ( .A1(n16096), .A2(n11000), .ZN(n16097) );
  XNOR2_X1 U11565 ( .A(n15479), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17129) );
  INV_X1 U11566 ( .A(n15477), .ZN(n11347) );
  INV_X1 U11567 ( .A(n11346), .ZN(n11345) );
  OAI21_X1 U11568 ( .B1(n16482), .B2(n11347), .A(n17129), .ZN(n11346) );
  NOR2_X1 U11569 ( .A1(n14865), .A2(n16485), .ZN(n14866) );
  AND2_X1 U11570 ( .A1(n16293), .A2(n11296), .ZN(n13778) );
  NOR2_X1 U11571 ( .A1(n11299), .A2(n11297), .ZN(n11296) );
  NAND2_X1 U11572 ( .A1(n11298), .A2(n16294), .ZN(n11297) );
  INV_X1 U11573 ( .A(n11069), .ZN(n11298) );
  NAND2_X1 U11574 ( .A1(n13778), .A2(n13779), .ZN(n15553) );
  AND2_X1 U11575 ( .A1(n16198), .A2(n11217), .ZN(n15555) );
  AND2_X1 U11576 ( .A1(n11218), .A2(n15455), .ZN(n11217) );
  NAND2_X1 U11577 ( .A1(n11029), .A2(n11340), .ZN(n11338) );
  AND2_X1 U11578 ( .A1(n15438), .A2(n15435), .ZN(n11341) );
  NAND2_X1 U11579 ( .A1(n11328), .A2(n11327), .ZN(n11326) );
  INV_X1 U11580 ( .A(n11324), .ZN(n11327) );
  AND2_X2 U11581 ( .A1(n16416), .A2(n15481), .ZN(n16567) );
  INV_X1 U11582 ( .A(n11164), .ZN(n11165) );
  NAND2_X1 U11583 ( .A1(n11089), .A2(n15351), .ZN(n16460) );
  NAND2_X1 U11584 ( .A1(n11095), .A2(n11093), .ZN(n11089) );
  NAND2_X1 U11585 ( .A1(n11288), .A2(n11289), .ZN(n16689) );
  AND2_X1 U11586 ( .A1(n16416), .A2(n11130), .ZN(n16704) );
  INV_X1 U11587 ( .A(n16692), .ZN(n11130) );
  NAND2_X1 U11588 ( .A1(n16704), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17142) );
  NAND2_X1 U11589 ( .A1(n16755), .A2(n15471), .ZN(n16483) );
  AND3_X1 U11590 ( .A1(n13666), .A2(n13665), .A3(n13664), .ZN(n14845) );
  NAND2_X1 U11591 ( .A1(n11280), .A2(n11278), .ZN(n15146) );
  INV_X1 U11592 ( .A(n14846), .ZN(n11280) );
  NAND2_X1 U11593 ( .A1(n11319), .A2(n15054), .ZN(n16774) );
  INV_X1 U11594 ( .A(n11304), .ZN(n13118) );
  NAND2_X1 U11595 ( .A1(n11304), .A2(n11303), .ZN(n13121) );
  INV_X1 U11596 ( .A(n13117), .ZN(n11303) );
  NAND2_X1 U11597 ( .A1(n14255), .A2(n11306), .ZN(n11302) );
  NAND4_X1 U11598 ( .A1(n13121), .A2(n11302), .A3(n13119), .A4(n11305), .ZN(
        n14243) );
  NAND2_X1 U11599 ( .A1(n18244), .A2(n13087), .ZN(n13089) );
  AND2_X1 U11600 ( .A1(n13092), .A2(n13091), .ZN(n14168) );
  OR2_X1 U11601 ( .A1(n14994), .A2(n14557), .ZN(n13092) );
  OR2_X1 U11602 ( .A1(n13084), .A2(n13083), .ZN(n11305) );
  AND2_X1 U11603 ( .A1(n19239), .A2(n19238), .ZN(n19258) );
  AND2_X1 U11604 ( .A1(n19239), .A2(n19525), .ZN(n19225) );
  INV_X1 U11605 ( .A(n19125), .ZN(n19254) );
  NOR2_X1 U11606 ( .A1(n19239), .A2(n19525), .ZN(n19178) );
  NAND2_X1 U11607 ( .A1(n15000), .A2(n15006), .ZN(n19154) );
  OAI21_X2 U11608 ( .B1(n18606), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n19116), 
        .ZN(n19281) );
  OR2_X1 U11609 ( .A1(n19142), .A2(n19141), .ZN(n19147) );
  INV_X1 U11610 ( .A(n19281), .ZN(n19639) );
  NAND2_X1 U11611 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19281), .ZN(n19641) );
  OR2_X1 U11612 ( .A1(n19142), .A2(n19123), .ZN(n19125) );
  NAND2_X1 U11613 ( .A1(n19110), .A2(n19525), .ZN(n19143) );
  INV_X1 U11614 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19214) );
  INV_X1 U11615 ( .A(n20549), .ZN(n11191) );
  INV_X1 U11616 ( .A(n12471), .ZN(n11099) );
  INV_X1 U11617 ( .A(n12467), .ZN(n11100) );
  INV_X1 U11618 ( .A(n12470), .ZN(n11101) );
  AOI21_X1 U11619 ( .B1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n17640), .A(
        n11103), .ZN(n11102) );
  INV_X1 U11620 ( .A(n12469), .ZN(n11103) );
  NAND2_X1 U11621 ( .A1(n17815), .A2(n11049), .ZN(n17907) );
  NAND2_X1 U11622 ( .A1(n12690), .A2(n18000), .ZN(n17957) );
  INV_X1 U11623 ( .A(n12688), .ZN(n12686) );
  NAND2_X1 U11624 ( .A1(n11263), .A2(n11262), .ZN(n12751) );
  AND2_X1 U11625 ( .A1(n11264), .A2(n21057), .ZN(n11262) );
  NOR2_X1 U11626 ( .A1(n17762), .A2(n12555), .ZN(n17813) );
  NAND2_X1 U11627 ( .A1(n11252), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11251) );
  NAND2_X1 U11628 ( .A1(n12511), .A2(n11252), .ZN(n11249) );
  OR2_X1 U11629 ( .A1(n18035), .A2(n20903), .ZN(n11254) );
  INV_X1 U11630 ( .A(n21233), .ZN(n21224) );
  NAND2_X1 U11631 ( .A1(n11678), .A2(n19891), .ZN(n11180) );
  INV_X1 U11632 ( .A(n11142), .ZN(n11678) );
  INV_X1 U11633 ( .A(n11143), .ZN(n15591) );
  OR2_X1 U11634 ( .A1(n11676), .A2(n11675), .ZN(n21623) );
  AND2_X1 U11635 ( .A1(n21483), .A2(n12391), .ZN(n21618) );
  INV_X1 U11636 ( .A(n21634), .ZN(n21613) );
  INV_X1 U11637 ( .A(n21623), .ZN(n21597) );
  AND2_X1 U11638 ( .A1(n14227), .A2(n14226), .ZN(n19820) );
  XNOR2_X1 U11639 ( .A(n12756), .B(n12387), .ZN(n12774) );
  AOI21_X1 U11640 ( .B1(n20014), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n21376), .ZN(n11114) );
  XNOR2_X1 U11641 ( .A(n11115), .B(n11614), .ZN(n21383) );
  NOR2_X1 U11642 ( .A1(n19970), .A2(n11116), .ZN(n11115) );
  AND2_X1 U11643 ( .A1(n19972), .A2(n19971), .ZN(n11116) );
  CLKBUF_X1 U11644 ( .A(n14661), .Z(n14662) );
  XNOR2_X1 U11645 ( .A(n15555), .B(n15554), .ZN(n16110) );
  NOR2_X1 U11646 ( .A1(n17198), .A2(n16343), .ZN(n11229) );
  INV_X1 U11647 ( .A(n11228), .ZN(n11227) );
  AOI21_X1 U11648 ( .B1(n17200), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16342), .ZN(n11228) );
  NAND2_X1 U11649 ( .A1(n18534), .A2(n17203), .ZN(n11162) );
  NAND2_X1 U11650 ( .A1(n18533), .A2(n17190), .ZN(n11161) );
  NOR2_X1 U11651 ( .A1(n17183), .A2(n11163), .ZN(n18535) );
  NOR2_X1 U11652 ( .A1(n11164), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11163) );
  INV_X1 U11653 ( .A(n17152), .ZN(n17203) );
  NAND2_X1 U11654 ( .A1(n18623), .A2(n13848), .ZN(n17151) );
  INV_X1 U11655 ( .A(n17190), .ZN(n17207) );
  INV_X1 U11656 ( .A(n17151), .ZN(n17200) );
  AOI21_X1 U11657 ( .B1(n16345), .B2(n18556), .A(n11283), .ZN(n11282) );
  NAND2_X1 U11658 ( .A1(n15565), .A2(n11013), .ZN(n11283) );
  INV_X1 U11659 ( .A(n18579), .ZN(n18553) );
  INV_X1 U11660 ( .A(n19290), .ZN(n19304) );
  INV_X1 U11661 ( .A(n19525), .ZN(n19238) );
  INV_X1 U11662 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n17222) );
  NAND2_X1 U11663 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n20588), .ZN(n20572) );
  INV_X1 U11664 ( .A(n20570), .ZN(n20587) );
  NAND2_X1 U11665 ( .A1(n17845), .A2(n21209), .ZN(n12745) );
  AOI21_X1 U11666 ( .B1(n11259), .B2(n17910), .A(n12691), .ZN(n12740) );
  INV_X1 U11667 ( .A(n21086), .ZN(n21092) );
  INV_X1 U11668 ( .A(n11690), .ZN(n11691) );
  OAI21_X1 U11669 ( .B1(n11689), .B2(n10954), .A(n13946), .ZN(n11690) );
  AND4_X1 U11670 ( .A1(n15100), .A2(n15099), .A3(n15098), .A4(n15097), .ZN(
        n15114) );
  AND2_X1 U11671 ( .A1(n19288), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13563) );
  OAI211_X1 U11672 ( .C1(n15300), .C2(n13869), .A(n13043), .B(n13042), .ZN(
        n13044) );
  NAND2_X1 U11673 ( .A1(n10965), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13071) );
  NAND2_X1 U11674 ( .A1(n11546), .A2(n11529), .ZN(n11535) );
  NOR2_X1 U11675 ( .A1(n11680), .A2(n21655), .ZN(n11538) );
  INV_X1 U11676 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11166) );
  OR2_X1 U11677 ( .A1(n11900), .A2(n11899), .ZN(n12826) );
  OR2_X1 U11678 ( .A1(n11877), .A2(n11876), .ZN(n12815) );
  NAND2_X1 U11679 ( .A1(n11758), .A2(n11756), .ZN(n11721) );
  INV_X1 U11680 ( .A(n11518), .ZN(n11120) );
  NAND2_X1 U11681 ( .A1(n11447), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11122) );
  NAND2_X1 U11682 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11124) );
  AOI22_X1 U11683 ( .A1(n11503), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11123) );
  NOR2_X1 U11684 ( .A1(n15358), .A2(n15357), .ZN(n15356) );
  NAND2_X1 U11685 ( .A1(n15371), .A2(n11060), .ZN(n11332) );
  AND2_X1 U11686 ( .A1(n15338), .A2(n15337), .ZN(n15473) );
  AND4_X1 U11687 ( .A1(n13524), .A2(n13523), .A3(n13522), .A4(n13521), .ZN(
        n13533) );
  INV_X1 U11688 ( .A(n15119), .ZN(n15121) );
  NAND2_X1 U11689 ( .A1(n13011), .A2(n14129), .ZN(n11126) );
  NAND2_X1 U11690 ( .A1(n13510), .A2(n13509), .ZN(n13558) );
  NOR2_X1 U11691 ( .A1(n13024), .A2(n13579), .ZN(n13591) );
  INV_X1 U11692 ( .A(n13387), .ZN(n13445) );
  AND2_X1 U11693 ( .A1(n15005), .A2(n16170), .ZN(n14999) );
  AOI22_X1 U11694 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U11695 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12910) );
  AOI22_X1 U11696 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12916) );
  INV_X1 U11697 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14481) );
  NAND2_X1 U11698 ( .A1(n20789), .A2(n20810), .ZN(n12579) );
  OR2_X1 U11699 ( .A1(n12676), .A2(n20647), .ZN(n12671) );
  NAND2_X1 U11700 ( .A1(n11537), .A2(n11853), .ZN(n11568) );
  NAND2_X1 U11701 ( .A1(n11688), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11141) );
  MUX2_X1 U11702 ( .A(n11659), .B(n13950), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n11589) );
  NAND2_X1 U11703 ( .A1(n11355), .A2(n11062), .ZN(n11354) );
  NAND2_X1 U11704 ( .A1(n15716), .A2(n11358), .ZN(n11357) );
  INV_X1 U11705 ( .A(n15642), .ZN(n11358) );
  OR2_X1 U11706 ( .A1(n12043), .A2(n11352), .ZN(n11351) );
  AND2_X1 U11707 ( .A1(n15161), .A2(n15169), .ZN(n11352) );
  AND3_X1 U11708 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(n11908), .ZN(n11928) );
  OR2_X1 U11709 ( .A1(n15719), .A2(n15714), .ZN(n11177) );
  AND2_X1 U11710 ( .A1(n20015), .A2(n21287), .ZN(n12858) );
  AND2_X1 U11711 ( .A1(n11940), .A2(n11903), .ZN(n11367) );
  OR2_X1 U11712 ( .A1(n20015), .A2(n12861), .ZN(n15912) );
  INV_X1 U11713 ( .A(n11696), .ZN(n11653) );
  NAND2_X1 U11714 ( .A1(n11023), .A2(n10954), .ZN(n11659) );
  NAND2_X1 U11715 ( .A1(n11524), .A2(n12400), .ZN(n11944) );
  NOR2_X1 U11716 ( .A1(n11686), .A2(n21655), .ZN(n11524) );
  OR2_X1 U11717 ( .A1(n11804), .A2(n11803), .ZN(n12791) );
  OAI21_X1 U11718 ( .B1(n11531), .B2(n11782), .A(n11781), .ZN(n11783) );
  OR2_X1 U11719 ( .A1(n11785), .A2(n13979), .ZN(n11791) );
  NAND2_X1 U11720 ( .A1(n11749), .A2(n11777), .ZN(n11941) );
  INV_X1 U11721 ( .A(n11944), .ZN(n11853) );
  OR2_X1 U11722 ( .A1(n11689), .A2(n11688), .ZN(n11576) );
  OR2_X1 U11723 ( .A1(n11785), .A2(n11376), .ZN(n11839) );
  INV_X1 U11724 ( .A(n11806), .ZN(n11709) );
  AOI21_X1 U11725 ( .B1(n21275), .B2(n21654), .A(n21658), .ZN(n14380) );
  NOR2_X1 U11726 ( .A1(n11154), .A2(n15185), .ZN(n11153) );
  INV_X1 U11727 ( .A(n15391), .ZN(n11154) );
  NOR2_X1 U11728 ( .A1(n11158), .A2(n15373), .ZN(n11157) );
  INV_X1 U11729 ( .A(n15354), .ZN(n11158) );
  AND2_X1 U11730 ( .A1(n15356), .A2(n15361), .ZN(n15353) );
  AND3_X1 U11731 ( .A1(n11150), .A2(n11149), .A3(n11148), .ZN(n15344) );
  NAND2_X1 U11732 ( .A1(n11150), .A2(n11149), .ZN(n15126) );
  INV_X1 U11733 ( .A(n14721), .ZN(n14724) );
  NOR2_X1 U11734 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13335) );
  AND2_X1 U11735 ( .A1(n11061), .A2(n16239), .ZN(n11315) );
  AND2_X1 U11736 ( .A1(n10994), .A2(n13258), .ZN(n11316) );
  NOR2_X1 U11737 ( .A1(n16104), .A2(n16355), .ZN(n15452) );
  NOR2_X1 U11738 ( .A1(n16091), .A2(n11238), .ZN(n11237) );
  INV_X1 U11739 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11238) );
  NOR2_X1 U11740 ( .A1(n16426), .A2(n11232), .ZN(n11231) );
  INV_X1 U11741 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11232) );
  NOR2_X1 U11742 ( .A1(n18297), .A2(n11235), .ZN(n11234) );
  INV_X1 U11743 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11235) );
  NAND2_X1 U11744 ( .A1(n13107), .A2(n13106), .ZN(n14327) );
  NAND2_X1 U11745 ( .A1(n11301), .A2(n11300), .ZN(n11299) );
  INV_X1 U11746 ( .A(n16276), .ZN(n11300) );
  INV_X1 U11747 ( .A(n16283), .ZN(n11301) );
  AND2_X1 U11748 ( .A1(n11338), .A2(n11337), .ZN(n11336) );
  INV_X1 U11749 ( .A(n15486), .ZN(n11337) );
  AND2_X1 U11750 ( .A1(n11220), .A2(n11219), .ZN(n11218) );
  INV_X1 U11751 ( .A(n16180), .ZN(n11219) );
  NOR2_X1 U11752 ( .A1(n11221), .A2(n16193), .ZN(n11220) );
  INV_X1 U11753 ( .A(n16199), .ZN(n11221) );
  OR2_X1 U11754 ( .A1(n16368), .A2(n16348), .ZN(n16350) );
  INV_X1 U11755 ( .A(n16308), .ZN(n11273) );
  NOR2_X1 U11756 ( .A1(n16233), .A2(n16225), .ZN(n16216) );
  OR2_X1 U11757 ( .A1(n15382), .A2(n10966), .ZN(n15410) );
  NOR2_X1 U11758 ( .A1(n11094), .A2(n15352), .ZN(n11093) );
  AND2_X1 U11759 ( .A1(n14332), .A2(n14323), .ZN(n11224) );
  INV_X1 U11760 ( .A(n14341), .ZN(n11225) );
  INV_X1 U11761 ( .A(n15115), .ZN(n14871) );
  NAND2_X1 U11762 ( .A1(n13097), .A2(n13099), .ZN(n13090) );
  INV_X1 U11763 ( .A(n13016), .ZN(n13017) );
  OR2_X1 U11764 ( .A1(n13632), .A2(n13631), .ZN(n13884) );
  OR2_X1 U11765 ( .A1(n14158), .A2(n13636), .ZN(n13652) );
  NAND2_X1 U11766 ( .A1(n11052), .A2(n13899), .ZN(n14126) );
  INV_X1 U11767 ( .A(n15328), .ZN(n19212) );
  NOR2_X1 U11768 ( .A1(n13799), .A2(n13579), .ZN(n13019) );
  INV_X1 U11769 ( .A(n12579), .ZN(n12452) );
  INV_X1 U11770 ( .A(n17735), .ZN(n11198) );
  XOR2_X1 U11771 ( .A(n20647), .B(n20774), .Z(n12492) );
  NOR2_X1 U11772 ( .A1(n12555), .A2(n11070), .ZN(n11261) );
  NAND2_X1 U11773 ( .A1(n21038), .A2(n21016), .ZN(n11265) );
  NOR2_X1 U11774 ( .A1(n17732), .A2(n21132), .ZN(n17706) );
  NAND2_X1 U11775 ( .A1(n11270), .A2(n12543), .ZN(n11269) );
  INV_X1 U11776 ( .A(n12542), .ZN(n11270) );
  AND2_X1 U11777 ( .A1(n17869), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12542) );
  NAND2_X1 U11778 ( .A1(n12490), .A2(n20647), .ZN(n12672) );
  INV_X1 U11779 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21217) );
  NAND2_X1 U11780 ( .A1(n11138), .A2(n15582), .ZN(n11136) );
  CLKBUF_X1 U11781 ( .A(n11705), .Z(n11577) );
  NOR2_X1 U11782 ( .A1(n15597), .A2(n19888), .ZN(n11143) );
  NAND2_X1 U11783 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n11147) );
  NOR2_X1 U11784 ( .A1(n19870), .A2(n11132), .ZN(n11131) );
  INV_X1 U11785 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n11132) );
  NAND2_X1 U11786 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n11145) );
  AND2_X1 U11787 ( .A1(n14050), .A2(n11672), .ZN(n11676) );
  INV_X1 U11788 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14754) );
  OR2_X1 U11789 ( .A1(n14660), .A2(n21922), .ZN(n14597) );
  MUX2_X1 U11790 ( .A(n15587), .B(n13950), .S(n15598), .Z(n11666) );
  OR2_X1 U11791 ( .A1(n11172), .A2(n15632), .ZN(n11171) );
  AND2_X1 U11792 ( .A1(n11622), .A2(n11621), .ZN(n15219) );
  NOR2_X1 U11793 ( .A1(n19923), .A2(n15219), .ZN(n15220) );
  NOR2_X1 U11794 ( .A1(n12333), .A2(n15841), .ZN(n12334) );
  OR2_X1 U11795 ( .A1(n12339), .A2(n12338), .ZN(n15606) );
  CLKBUF_X1 U11796 ( .A(n15618), .Z(n15619) );
  AND2_X1 U11797 ( .A1(n12378), .A2(n21635), .ZN(n12263) );
  NOR2_X1 U11798 ( .A1(n12227), .A2(n21609), .ZN(n12228) );
  NAND2_X1 U11799 ( .A1(n12228), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12283) );
  NAND2_X1 U11800 ( .A1(n12197), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12227) );
  NOR2_X1 U11801 ( .A1(n12147), .A2(n12146), .ZN(n12148) );
  NAND2_X1 U11802 ( .A1(n12148), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12196) );
  CLKBUF_X1 U11803 ( .A(n15693), .Z(n15694) );
  NOR2_X1 U11804 ( .A1(n12124), .A2(n21535), .ZN(n12125) );
  NAND2_X1 U11805 ( .A1(n12125), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12147) );
  AND2_X1 U11806 ( .A1(n12127), .A2(n12126), .ZN(n15711) );
  NOR2_X1 U11807 ( .A1(n12078), .A2(n12060), .ZN(n12079) );
  NAND2_X1 U11808 ( .A1(n12059), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12078) );
  CLKBUF_X1 U11809 ( .A(n15200), .Z(n15233) );
  NOR2_X1 U11810 ( .A1(n12038), .A2(n12024), .ZN(n12044) );
  CLKBUF_X1 U11811 ( .A(n14808), .Z(n14809) );
  NAND2_X1 U11812 ( .A1(n11946), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11966) );
  AND2_X1 U11813 ( .A1(n11928), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11946) );
  AOI21_X1 U11814 ( .B1(n12808), .B2(n12069), .A(n11887), .ZN(n14647) );
  NOR2_X1 U11815 ( .A1(n11856), .A2(n14606), .ZN(n11908) );
  NAND2_X1 U11816 ( .A1(n11864), .A2(n11863), .ZN(n14425) );
  CLKBUF_X1 U11817 ( .A(n14424), .Z(n14648) );
  NOR3_X1 U11818 ( .A1(n15634), .A2(n15622), .A3(n15610), .ZN(n15608) );
  NAND2_X1 U11819 ( .A1(n15849), .A2(n12873), .ZN(n15838) );
  NOR2_X1 U11820 ( .A1(n15689), .A2(n15678), .ZN(n19929) );
  OAI21_X1 U11821 ( .B1(n15887), .B2(n11380), .A(n11378), .ZN(n12868) );
  OR2_X1 U11822 ( .A1(n15698), .A2(n15691), .ZN(n15689) );
  NOR3_X1 U11823 ( .A1(n15720), .A2(n11177), .A3(n11175), .ZN(n19936) );
  OR2_X1 U11824 ( .A1(n11178), .A2(n11176), .ZN(n11175) );
  INV_X1 U11825 ( .A(n19934), .ZN(n11176) );
  NAND2_X1 U11826 ( .A1(n19936), .A2(n15696), .ZN(n15698) );
  NOR2_X1 U11827 ( .A1(n15720), .A2(n11177), .ZN(n15713) );
  OR2_X1 U11828 ( .A1(n15644), .A2(n15645), .ZN(n15720) );
  AND2_X1 U11829 ( .A1(n15220), .A2(n15203), .ZN(n15238) );
  NAND2_X1 U11830 ( .A1(n15238), .A2(n15237), .ZN(n15644) );
  OR2_X1 U11831 ( .A1(n19922), .A2(n11181), .ZN(n19923) );
  OR2_X1 U11832 ( .A1(n19921), .A2(n19920), .ZN(n11181) );
  NOR2_X1 U11833 ( .A1(n15922), .A2(n15932), .ZN(n19972) );
  AND2_X1 U11834 ( .A1(n11610), .A2(n11609), .ZN(n14940) );
  NAND2_X1 U11835 ( .A1(n11168), .A2(n10989), .ZN(n19941) );
  INV_X1 U11836 ( .A(n14799), .ZN(n11167) );
  NAND2_X1 U11837 ( .A1(n11168), .A2(n11169), .ZN(n14798) );
  NOR2_X1 U11838 ( .A1(n14426), .A2(n14649), .ZN(n14654) );
  AND2_X1 U11839 ( .A1(n14416), .A2(n14415), .ZN(n14428) );
  NAND2_X1 U11840 ( .A1(n14304), .A2(n11020), .ZN(n14611) );
  NOR2_X1 U11841 ( .A1(n16063), .A2(n14614), .ZN(n15941) );
  AND2_X1 U11842 ( .A1(n14062), .A2(n14061), .ZN(n14080) );
  NAND2_X1 U11843 ( .A1(n11374), .A2(n21655), .ZN(n11772) );
  NAND2_X1 U11844 ( .A1(n11784), .A2(n14438), .ZN(n14661) );
  OR2_X1 U11845 ( .A1(n12799), .A2(n10975), .ZN(n21807) );
  INV_X1 U11846 ( .A(n14368), .ZN(n14371) );
  NAND2_X1 U11847 ( .A1(n12799), .A2(n10974), .ZN(n21869) );
  OR3_X1 U11848 ( .A1(n21837), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14380), 
        .ZN(n14569) );
  AND3_X1 U11849 ( .A1(n13951), .A2(n12767), .A3(n13934), .ZN(n16868) );
  XNOR2_X1 U11850 ( .A(n15531), .B(n11068), .ZN(n15491) );
  AND2_X1 U11851 ( .A1(n15308), .A2(n15439), .ZN(n15311) );
  NOR2_X1 U11852 ( .A1(n15424), .A2(n15305), .ZN(n15427) );
  NOR2_X1 U11853 ( .A1(n15397), .A2(n15304), .ZN(n15398) );
  NAND2_X1 U11854 ( .A1(n12983), .A2(n13511), .ZN(n12990) );
  AND2_X1 U11855 ( .A1(n18423), .A2(n11033), .ZN(n18384) );
  NAND2_X1 U11856 ( .A1(n15380), .A2(n15379), .ZN(n15397) );
  NOR2_X1 U11857 ( .A1(n13579), .A2(n18347), .ZN(n15377) );
  NOR2_X1 U11858 ( .A1(n15385), .A2(n15377), .ZN(n15380) );
  NAND2_X1 U11859 ( .A1(n15392), .A2(n11151), .ZN(n15385) );
  NOR2_X1 U11860 ( .A1(n11152), .A2(n15383), .ZN(n11151) );
  INV_X1 U11861 ( .A(n11153), .ZN(n11152) );
  NAND2_X1 U11862 ( .A1(n15392), .A2(n15391), .ZN(n15394) );
  AND2_X1 U11863 ( .A1(n15389), .A2(n15069), .ZN(n15392) );
  NAND2_X1 U11864 ( .A1(n15353), .A2(n11157), .ZN(n15388) );
  AND2_X1 U11865 ( .A1(n15353), .A2(n11155), .ZN(n15389) );
  NOR2_X1 U11866 ( .A1(n11156), .A2(n15387), .ZN(n11155) );
  INV_X1 U11867 ( .A(n11157), .ZN(n11156) );
  OR2_X1 U11868 ( .A1(n13086), .A2(n13085), .ZN(n14980) );
  AND2_X1 U11869 ( .A1(n13184), .A2(n13183), .ZN(n13734) );
  NAND2_X1 U11870 ( .A1(n13169), .A2(n11406), .ZN(n14701) );
  NOR2_X1 U11871 ( .A1(n16284), .A2(n11299), .ZN(n16278) );
  NOR2_X1 U11872 ( .A1(n13469), .A2(n13468), .ZN(n16187) );
  NAND2_X1 U11873 ( .A1(n11308), .A2(n11307), .ZN(n16208) );
  OAI21_X1 U11874 ( .B1(n16220), .B2(n11312), .A(n11310), .ZN(n11309) );
  NAND2_X1 U11875 ( .A1(n16208), .A2(n16207), .ZN(n16206) );
  AOI22_X1 U11876 ( .A1(n16223), .A2(n16224), .B1(n13384), .B2(n19585), .ZN(
        n16220) );
  CLKBUF_X1 U11877 ( .A(n16223), .Z(n16234) );
  AND2_X1 U11878 ( .A1(n16255), .A2(n11061), .ZN(n16246) );
  NAND2_X1 U11879 ( .A1(n16255), .A2(n11315), .ZN(n16238) );
  AND2_X1 U11880 ( .A1(n13752), .A2(n13751), .ZN(n15192) );
  AND2_X1 U11881 ( .A1(n14825), .A2(n11316), .ZN(n15209) );
  NAND2_X1 U11882 ( .A1(n11286), .A2(n16126), .ZN(n11285) );
  INV_X1 U11883 ( .A(n11276), .ZN(n11275) );
  AND2_X1 U11884 ( .A1(n13121), .A2(n13120), .ZN(n13122) );
  INV_X1 U11885 ( .A(n14088), .ZN(n19109) );
  NAND2_X1 U11886 ( .A1(n16099), .A2(n11236), .ZN(n16104) );
  AND2_X1 U11887 ( .A1(n10999), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11236) );
  NAND2_X1 U11888 ( .A1(n16099), .A2(n10999), .ZN(n16102) );
  NAND2_X1 U11889 ( .A1(n16099), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16092) );
  NOR2_X1 U11890 ( .A1(n16100), .A2(n16390), .ZN(n16099) );
  NAND2_X1 U11891 ( .A1(n16098), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16100) );
  AND2_X1 U11892 ( .A1(n16096), .A2(n11230), .ZN(n16098) );
  AND2_X1 U11893 ( .A1(n11000), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11230) );
  INV_X1 U11894 ( .A(n16407), .ZN(n11096) );
  NAND2_X1 U11895 ( .A1(n16096), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16095) );
  NOR2_X1 U11896 ( .A1(n16093), .A2(n16094), .ZN(n16096) );
  NAND2_X1 U11897 ( .A1(n15188), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16093) );
  NOR2_X1 U11898 ( .A1(n15187), .A2(n18330), .ZN(n15188) );
  AND2_X1 U11899 ( .A1(n15074), .A2(n11233), .ZN(n15076) );
  AND2_X1 U11900 ( .A1(n10993), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11233) );
  NAND2_X1 U11901 ( .A1(n15076), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15187) );
  NAND2_X1 U11902 ( .A1(n15074), .A2(n10993), .ZN(n15075) );
  NOR2_X1 U11903 ( .A1(n15071), .A2(n18275), .ZN(n15074) );
  NAND2_X1 U11904 ( .A1(n15074), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15073) );
  INV_X1 U11905 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18275) );
  NAND2_X1 U11906 ( .A1(n14866), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15071) );
  NOR2_X1 U11907 ( .A1(n18249), .A2(n11240), .ZN(n11239) );
  NOR2_X1 U11908 ( .A1(n14712), .A2(n17106), .ZN(n14834) );
  INV_X1 U11909 ( .A(n14325), .ZN(n11202) );
  NAND2_X1 U11910 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14712) );
  INV_X1 U11911 ( .A(n15534), .ZN(n11335) );
  NAND2_X1 U11912 ( .A1(n16198), .A2(n11220), .ZN(n16195) );
  NOR2_X1 U11913 ( .A1(n18459), .A2(n10966), .ZN(n16351) );
  NAND2_X1 U11914 ( .A1(n16293), .A2(n16294), .ZN(n16284) );
  NOR2_X1 U11915 ( .A1(n16350), .A2(n16349), .ZN(n16362) );
  NAND2_X1 U11916 ( .A1(n16548), .A2(n16547), .ZN(n11342) );
  NAND2_X1 U11917 ( .A1(n11320), .A2(n11324), .ZN(n11323) );
  NAND2_X1 U11918 ( .A1(n16567), .A2(n15512), .ZN(n16549) );
  AND2_X1 U11919 ( .A1(n13758), .A2(n13757), .ZN(n18371) );
  INV_X1 U11920 ( .A(n18351), .ZN(n11292) );
  INV_X1 U11921 ( .A(n11294), .ZN(n11293) );
  NAND2_X1 U11922 ( .A1(n11207), .A2(n16261), .ZN(n11206) );
  INV_X1 U11923 ( .A(n11208), .ZN(n11207) );
  NOR3_X1 U11924 ( .A1(n14972), .A2(n15213), .A3(n11208), .ZN(n16260) );
  NOR3_X1 U11925 ( .A1(n16652), .A2(n11294), .A3(n18351), .ZN(n18350) );
  NOR2_X1 U11926 ( .A1(n11213), .A2(n11212), .ZN(n11211) );
  INV_X1 U11927 ( .A(n14946), .ZN(n11212) );
  NAND2_X1 U11928 ( .A1(n11328), .A2(n11322), .ZN(n16450) );
  NAND2_X1 U11929 ( .A1(n11210), .A2(n11215), .ZN(n14855) );
  NOR2_X1 U11930 ( .A1(n14707), .A2(n14706), .ZN(n14854) );
  AOI21_X1 U11931 ( .B1(n11345), .B2(n11347), .A(n11028), .ZN(n11343) );
  INV_X1 U11932 ( .A(n16416), .ZN(n17167) );
  NOR2_X1 U11933 ( .A1(n14341), .A2(n11222), .ZN(n14642) );
  NAND2_X1 U11934 ( .A1(n11224), .A2(n11223), .ZN(n11222) );
  INV_X1 U11935 ( .A(n14587), .ZN(n11223) );
  NAND2_X1 U11936 ( .A1(n15467), .A2(n11127), .ZN(n16754) );
  NAND2_X1 U11937 ( .A1(n15459), .A2(n11128), .ZN(n11127) );
  OAI21_X1 U11938 ( .B1(n15460), .B2(n15465), .A(n15464), .ZN(n15466) );
  NAND2_X1 U11939 ( .A1(n11225), .A2(n11224), .ZN(n14588) );
  NAND2_X1 U11940 ( .A1(n11225), .A2(n14332), .ZN(n14333) );
  AND2_X1 U11941 ( .A1(n14150), .A2(n14523), .ZN(n18573) );
  XNOR2_X1 U11942 ( .A(n14158), .B(n13619), .ZN(n14145) );
  NOR2_X2 U11943 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13127) );
  INV_X1 U11944 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14487) );
  OR2_X1 U11945 ( .A1(n14098), .A2(n13577), .ZN(n14561) );
  NAND2_X1 U11946 ( .A1(n15008), .A2(n10973), .ZN(n19308) );
  NAND2_X1 U11947 ( .A1(n19281), .A2(n19304), .ZN(n19306) );
  AND2_X1 U11948 ( .A1(n19126), .A2(n19304), .ZN(n19130) );
  NAND2_X2 U11949 ( .A1(n13004), .A2(n13003), .ZN(n19534) );
  NAND2_X1 U11950 ( .A1(n12997), .A2(n13511), .ZN(n13004) );
  AND4_X1 U11951 ( .A1(n12996), .A2(n12995), .A3(n12994), .A4(n12993), .ZN(
        n12997) );
  INV_X1 U11952 ( .A(n14129), .ZN(n19478) );
  NAND2_X1 U11953 ( .A1(n12932), .A2(n13511), .ZN(n12939) );
  NAND2_X1 U11954 ( .A1(n12937), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12938) );
  AND4_X1 U11955 ( .A1(n12931), .A2(n12930), .A3(n12929), .A4(n12928), .ZN(
        n12932) );
  NAND2_X1 U11956 ( .A1(n21205), .A2(n21204), .ZN(n20593) );
  INV_X1 U11957 ( .A(n16825), .ZN(n21206) );
  NOR2_X1 U11958 ( .A1(n12731), .A2(n12733), .ZN(n21207) );
  OR2_X1 U11959 ( .A1(n20518), .A2(n11194), .ZN(n11196) );
  NOR2_X1 U11960 ( .A1(n20508), .A2(n11194), .ZN(n20509) );
  NOR2_X1 U11961 ( .A1(n11194), .A2(n20403), .ZN(n11187) );
  OR2_X1 U11962 ( .A1(n20406), .A2(n20407), .ZN(n11190) );
  INV_X1 U11963 ( .A(n20502), .ZN(n20517) );
  AOI21_X1 U11964 ( .B1(n17293), .B2(n17292), .A(n21263), .ZN(n20595) );
  NOR2_X1 U11965 ( .A1(n12433), .A2(n11244), .ZN(n12512) );
  AOI22_X1 U11966 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12425), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12480) );
  NAND2_X1 U11967 ( .A1(n12482), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12483) );
  INV_X1 U11968 ( .A(n18144), .ZN(n18145) );
  NOR2_X1 U11969 ( .A1(n21263), .A2(n21207), .ZN(n17688) );
  NOR2_X1 U11970 ( .A1(n21679), .A2(n20108), .ZN(n20594) );
  NAND2_X1 U11971 ( .A1(n17915), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17896) );
  NAND2_X1 U11972 ( .A1(n17768), .A2(n11403), .ZN(n17802) );
  AND2_X1 U11973 ( .A1(n17743), .A2(n11197), .ZN(n17929) );
  NAND2_X1 U11974 ( .A1(n10985), .A2(n17743), .ZN(n17925) );
  NAND2_X1 U11975 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n20988), .ZN(
        n20989) );
  NAND2_X1 U11976 ( .A1(n17743), .A2(n11199), .ZN(n17723) );
  INV_X1 U11977 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20323) );
  NAND2_X1 U11978 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11183) );
  NOR2_X1 U11979 ( .A1(n20221), .A2(n11185), .ZN(n11184) );
  XNOR2_X1 U11980 ( .A(n20871), .B(n12492), .ZN(n18068) );
  NOR2_X1 U11981 ( .A1(n12490), .A2(n12489), .ZN(n12491) );
  INV_X1 U11982 ( .A(n11258), .ZN(n11257) );
  AOI21_X1 U11983 ( .B1(n11258), .B2(n11256), .A(n12747), .ZN(n11255) );
  NOR2_X1 U11984 ( .A1(n20626), .A2(n17697), .ZN(n11258) );
  NAND2_X1 U11985 ( .A1(n17823), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n21032) );
  NOR2_X1 U11986 ( .A1(n17824), .A2(n21016), .ZN(n17823) );
  NOR2_X1 U11987 ( .A1(n11398), .A2(n20989), .ZN(n21084) );
  NOR2_X1 U11988 ( .A1(n21129), .A2(n11398), .ZN(n21087) );
  NAND2_X1 U11989 ( .A1(n17955), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n21130) );
  AND2_X1 U11990 ( .A1(n12549), .A2(n11248), .ZN(n17732) );
  INV_X1 U11991 ( .A(n12550), .ZN(n11248) );
  NAND2_X1 U11992 ( .A1(n20998), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21129) );
  NAND2_X1 U11993 ( .A1(n17957), .A2(n20969), .ZN(n17949) );
  AND2_X1 U11994 ( .A1(n11268), .A2(n11267), .ZN(n17756) );
  NOR2_X1 U11995 ( .A1(n11269), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11267) );
  INV_X1 U11996 ( .A(n11269), .ZN(n11266) );
  NAND2_X1 U11997 ( .A1(n18022), .A2(n12685), .ZN(n18012) );
  XNOR2_X1 U11998 ( .A(n12684), .B(n11105), .ZN(n18023) );
  INV_X1 U11999 ( .A(n12683), .ZN(n11105) );
  NAND2_X1 U12000 ( .A1(n18041), .A2(n12681), .ZN(n18032) );
  NAND2_X1 U12001 ( .A1(n18032), .A2(n18033), .ZN(n18031) );
  NAND2_X1 U12002 ( .A1(n20775), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18084) );
  NOR2_X1 U12003 ( .A1(n20814), .A2(n10972), .ZN(n20812) );
  NAND3_X1 U12004 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n21214), .ZN(n20817) );
  NAND2_X1 U12005 ( .A1(n20102), .A2(n16807), .ZN(n21203) );
  NOR2_X1 U12006 ( .A1(n12641), .A2(n12640), .ZN(n18851) );
  NOR2_X1 U12007 ( .A1(n12578), .A2(n12577), .ZN(n18772) );
  NAND2_X1 U12008 ( .A1(n12416), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15727)
         );
  NAND2_X1 U12009 ( .A1(n11137), .A2(n11133), .ZN(n14259) );
  NOR2_X1 U12010 ( .A1(n11136), .A2(n11134), .ZN(n11133) );
  NAND2_X1 U12011 ( .A1(n21629), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15638) );
  NOR2_X1 U12012 ( .A1(n21599), .A2(n11146), .ZN(n21629) );
  OR2_X1 U12013 ( .A1(n11147), .A2(n19881), .ZN(n11146) );
  NOR2_X1 U12014 ( .A1(n21599), .A2(n11147), .ZN(n11390) );
  NOR2_X1 U12015 ( .A1(n21599), .A2(n21600), .ZN(n21610) );
  AND2_X1 U12016 ( .A1(n21538), .A2(n11072), .ZN(n21588) );
  NAND2_X1 U12017 ( .A1(n21538), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n21558) );
  INV_X1 U12018 ( .A(n21627), .ZN(n21601) );
  NOR2_X1 U12019 ( .A1(n21510), .A2(n11144), .ZN(n21529) );
  OR2_X1 U12020 ( .A1(n11145), .A2(n19861), .ZN(n11144) );
  OR2_X1 U12021 ( .A1(n21510), .A2(n11145), .ZN(n15657) );
  NOR2_X1 U12022 ( .A1(n21510), .A2(n19969), .ZN(n21517) );
  INV_X1 U12023 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14606) );
  INV_X1 U12024 ( .A(n21615), .ZN(n21626) );
  INV_X1 U12025 ( .A(n21484), .ZN(n21493) );
  AND2_X1 U12026 ( .A1(n21483), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21615) );
  AND2_X1 U12027 ( .A1(n19946), .A2(n12394), .ZN(n19925) );
  NAND2_X1 U12028 ( .A1(n13991), .A2(n13990), .ZN(n19946) );
  INV_X1 U12029 ( .A(n19925), .ZN(n19942) );
  INV_X1 U12030 ( .A(n15786), .ZN(n15776) );
  INV_X1 U12031 ( .A(n15794), .ZN(n15798) );
  NOR2_X1 U12032 ( .A1(n15798), .A2(n14218), .ZN(n15799) );
  INV_X1 U12033 ( .A(n15799), .ZN(n15796) );
  BUF_X1 U12034 ( .A(n14630), .Z(n21278) );
  BUF_X1 U12035 ( .A(n14629), .Z(n19841) );
  NAND2_X1 U12036 ( .A1(n12393), .A2(n14223), .ZN(n21777) );
  OR2_X1 U12037 ( .A1(n21775), .A2(n14410), .ZN(n21772) );
  OAI21_X1 U12038 ( .B1(n15595), .B2(n15596), .A(n12755), .ZN(n15825) );
  AOI21_X1 U12039 ( .B1(n15688), .B2(n15687), .A(n15686), .ZN(n21591) );
  AND2_X1 U12040 ( .A1(n15898), .A2(n12771), .ZN(n19989) );
  NAND2_X1 U12041 ( .A1(n15088), .A2(n12851), .ZN(n15224) );
  NAND2_X1 U12042 ( .A1(n14687), .A2(n12822), .ZN(n19959) );
  NAND2_X1 U12043 ( .A1(n19947), .A2(n12814), .ZN(n14685) );
  OR2_X1 U12044 ( .A1(n12768), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21419) );
  INV_X1 U12045 ( .A(n21382), .ZN(n21422) );
  INV_X1 U12046 ( .A(n21414), .ZN(n21421) );
  INV_X1 U12047 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21892) );
  INV_X1 U12048 ( .A(n11368), .ZN(n14315) );
  AND2_X1 U12049 ( .A1(n14300), .A2(n21900), .ZN(n21862) );
  NAND2_X1 U12050 ( .A1(n11794), .A2(n14286), .ZN(n21877) );
  INV_X1 U12051 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13961) );
  NOR2_X1 U12052 ( .A1(n21807), .A2(n21868), .ZN(n22202) );
  OR2_X1 U12053 ( .A1(n14441), .A2(n21844), .ZN(n22208) );
  OAI211_X1 U12054 ( .C1(n22215), .C2(n21837), .A(n21836), .B(n21858), .ZN(
        n22218) );
  OR2_X1 U12055 ( .A1(n21869), .A2(n21844), .ZN(n22157) );
  AND2_X1 U12056 ( .A1(n21905), .A2(n21872), .ZN(n22251) );
  OAI211_X1 U12057 ( .C1(n22257), .C2(n21915), .A(n21914), .B(n21913), .ZN(
        n22260) );
  NAND2_X1 U12058 ( .A1(n21905), .A2(n21779), .ZN(n22270) );
  AND2_X1 U12059 ( .A1(n21932), .A2(n21931), .ZN(n22268) );
  NOR2_X1 U12060 ( .A1(n13821), .A2(n21837), .ZN(n21658) );
  INV_X1 U12061 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16886) );
  AND2_X1 U12062 ( .A1(n16886), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21649) );
  INV_X1 U12063 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21690) );
  NAND2_X1 U12064 ( .A1(n21690), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21684) );
  AND2_X1 U12065 ( .A1(n14551), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18619) );
  INV_X1 U12066 ( .A(n15491), .ZN(n16120) );
  NAND2_X1 U12067 ( .A1(n18484), .A2(n18483), .ZN(n18481) );
  NAND2_X1 U12068 ( .A1(n18465), .A2(n18464), .ZN(n18463) );
  OR2_X1 U12069 ( .A1(n18452), .A2(n18451), .ZN(n18454) );
  INV_X1 U12070 ( .A(n15307), .ZN(n15437) );
  NAND2_X1 U12071 ( .A1(n18407), .A2(n18406), .ZN(n18405) );
  NAND2_X1 U12072 ( .A1(n18396), .A2(n18395), .ZN(n18394) );
  NOR2_X1 U12073 ( .A1(n18473), .A2(n17222), .ZN(n18474) );
  INV_X1 U12074 ( .A(n18490), .ZN(n18470) );
  OR2_X1 U12075 ( .A1(n18384), .A2(n18385), .ZN(n18387) );
  INV_X1 U12076 ( .A(n18423), .ZN(n18436) );
  INV_X1 U12077 ( .A(n18494), .ZN(n18471) );
  OR3_X1 U12078 ( .A1(n14737), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n21699), 
        .ZN(n18478) );
  AND2_X1 U12079 ( .A1(n11243), .A2(n11242), .ZN(n18423) );
  NAND2_X1 U12080 ( .A1(n15561), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11242) );
  NAND2_X1 U12081 ( .A1(n16343), .A2(n14714), .ZN(n11243) );
  CLKBUF_X1 U12082 ( .A(n14716), .Z(n18482) );
  INV_X1 U12083 ( .A(n18329), .ZN(n18498) );
  INV_X1 U12084 ( .A(n18478), .ZN(n18501) );
  INV_X1 U12085 ( .A(n16341), .ZN(n18502) );
  OR2_X1 U12086 ( .A1(n13151), .A2(n13150), .ZN(n14680) );
  INV_X1 U12087 ( .A(n16253), .ZN(n16266) );
  NAND2_X1 U12088 ( .A1(n14339), .A2(n10991), .ZN(n14638) );
  INV_X1 U12089 ( .A(n19123), .ZN(n19141) );
  NOR2_X1 U12090 ( .A1(n16725), .A2(n16709), .ZN(n16691) );
  AND2_X1 U12091 ( .A1(n19531), .A2(n11083), .ZN(n19633) );
  INV_X1 U12092 ( .A(n19579), .ZN(n19634) );
  INV_X1 U12093 ( .A(n19524), .ZN(n19583) );
  BUF_X1 U12095 ( .A(n17256), .Z(n17265) );
  NOR2_X1 U12096 ( .A1(n17241), .A2(n17265), .ZN(n17254) );
  AND2_X1 U12097 ( .A1(n14974), .A2(n14973), .ZN(n18318) );
  NAND2_X1 U12098 ( .A1(n16484), .A2(n15477), .ZN(n17130) );
  INV_X1 U12099 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16485) );
  CLKBUF_X1 U12100 ( .A(n14986), .Z(n16157) );
  AND2_X1 U12101 ( .A1(n15553), .A2(n13782), .ZN(n16113) );
  OR2_X1 U12102 ( .A1(n15555), .A2(n15456), .ZN(n18479) );
  NAND2_X1 U12103 ( .A1(n11339), .A2(n11338), .ZN(n15487) );
  NAND2_X1 U12104 ( .A1(n11326), .A2(n11333), .ZN(n16572) );
  XNOR2_X1 U12105 ( .A(n17142), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18525) );
  OAI21_X1 U12106 ( .B1(n16460), .B2(n15372), .A(n15371), .ZN(n17141) );
  INV_X1 U12107 ( .A(n16728), .ZN(n16694) );
  NAND2_X1 U12108 ( .A1(n15146), .A2(n13702), .ZN(n14882) );
  NOR2_X1 U12109 ( .A1(n14846), .A2(n14845), .ZN(n15148) );
  NAND2_X1 U12110 ( .A1(n15469), .A2(n15140), .ZN(n15141) );
  INV_X1 U12111 ( .A(n18512), .ZN(n18584) );
  INV_X1 U12112 ( .A(n16773), .ZN(n11348) );
  AND2_X1 U12113 ( .A1(n14150), .A2(n14138), .ZN(n18568) );
  INV_X1 U12114 ( .A(n16767), .ZN(n18582) );
  INV_X1 U12115 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19288) );
  INV_X1 U12116 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19260) );
  INV_X1 U12117 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19256) );
  AND2_X1 U12118 ( .A1(n11302), .A2(n11305), .ZN(n14245) );
  AND2_X1 U12119 ( .A1(n13121), .A2(n13119), .ZN(n14244) );
  INV_X1 U12120 ( .A(n14168), .ZN(n14170) );
  XNOR2_X1 U12121 ( .A(n14254), .B(n14256), .ZN(n19525) );
  INV_X1 U12122 ( .A(n14255), .ZN(n14256) );
  INV_X1 U12123 ( .A(n19239), .ZN(n19110) );
  INV_X1 U12124 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13917) );
  OAI22_X1 U12125 ( .A1(n19251), .A2(n19247), .B1(n19246), .B2(n19245), .ZN(
        n19718) );
  INV_X1 U12126 ( .A(n19714), .ZN(n19704) );
  OAI21_X1 U12127 ( .B1(n19157), .B2(n19156), .A(n19155), .ZN(n19668) );
  INV_X1 U12128 ( .A(n19411), .ZN(n19416) );
  INV_X1 U12129 ( .A(n19657), .ZN(n19660) );
  INV_X1 U12130 ( .A(n19363), .ZN(n19365) );
  INV_X1 U12131 ( .A(n19567), .ZN(n19569) );
  INV_X1 U12132 ( .A(n19507), .ZN(n19514) );
  INV_X1 U12133 ( .A(n19460), .ZN(n19466) );
  INV_X1 U12134 ( .A(n19650), .ZN(n19652) );
  INV_X1 U12135 ( .A(n19414), .ZN(n19415) );
  INV_X1 U12136 ( .A(n19537), .ZN(n19745) );
  INV_X1 U12137 ( .A(n19286), .ZN(n19317) );
  OR2_X1 U12138 ( .A1(n19143), .A2(n19125), .ZN(n19650) );
  NAND2_X1 U12139 ( .A1(n11192), .A2(n11193), .ZN(n20548) );
  AND2_X1 U12140 ( .A1(n11190), .A2(n20396), .ZN(n20420) );
  AND2_X1 U12141 ( .A1(n17438), .A2(n17675), .ZN(n17626) );
  AND2_X1 U12142 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17626), .ZN(n17654) );
  INV_X1 U12143 ( .A(n17684), .ZN(n17438) );
  NOR2_X1 U12144 ( .A1(n20717), .A2(n20711), .ZN(n20710) );
  NOR2_X1 U12145 ( .A1(n20729), .A2(n20694), .ZN(n20700) );
  NOR2_X1 U12146 ( .A1(n20693), .A2(n20736), .ZN(n20730) );
  NOR3_X1 U12147 ( .A1(n20744), .A2(n20692), .A3(n20691), .ZN(n20737) );
  NOR3_X1 U12148 ( .A1(n20693), .A2(n20744), .A3(n20654), .ZN(n20685) );
  NAND2_X1 U12149 ( .A1(n20755), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n20744) );
  NOR2_X1 U12150 ( .A1(n12440), .A2(n12439), .ZN(n20639) );
  NOR2_X1 U12151 ( .A1(n11100), .A2(n11099), .ZN(n11098) );
  NOR2_X1 U12152 ( .A1(n20667), .A2(n20601), .ZN(n20768) );
  NAND2_X1 U12153 ( .A1(n20602), .A2(n20779), .ZN(n20773) );
  INV_X1 U12154 ( .A(n20601), .ZN(n20779) );
  INV_X1 U12155 ( .A(n20773), .ZN(n20776) );
  CLKBUF_X1 U12156 ( .A(n18159), .Z(n18167) );
  CLKBUF_X1 U12157 ( .A(n20142), .Z(n20150) );
  AND2_X1 U12158 ( .A1(n17889), .A2(n10982), .ZN(n17890) );
  INV_X1 U12159 ( .A(n17880), .ZN(n17882) );
  NAND2_X1 U12160 ( .A1(n17815), .A2(n10992), .ZN(n17865) );
  NOR2_X1 U12161 ( .A1(n17950), .A2(n17948), .ZN(n20988) );
  INV_X1 U12162 ( .A(n18002), .ZN(n17952) );
  NOR3_X2 U12163 ( .A1(n18059), .A2(P3_STATEBS16_REG_SCAN_IN), .A3(n20785), 
        .ZN(n17917) );
  NOR2_X2 U12164 ( .A1(n20626), .A2(n18090), .ZN(n18004) );
  NAND2_X1 U12165 ( .A1(n11071), .A2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n20198) );
  NOR2_X1 U12166 ( .A1(n20183), .A2(n18058), .ZN(n18048) );
  INV_X2 U12167 ( .A(n10981), .ZN(n18091) );
  OAI21_X1 U12168 ( .B1(n21062), .B2(n21202), .A(n11104), .ZN(n21079) );
  OR2_X1 U12169 ( .A1(n21064), .A2(n21063), .ZN(n11104) );
  AND2_X1 U12170 ( .A1(n17813), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17870) );
  NAND2_X1 U12171 ( .A1(n12549), .A2(n12548), .ZN(n17924) );
  INV_X1 U12172 ( .A(n11247), .ZN(n17923) );
  NOR2_X1 U12173 ( .A1(n17949), .A2(n17950), .ZN(n20998) );
  NAND2_X1 U12174 ( .A1(n20812), .A2(n20795), .ZN(n21185) );
  OAI21_X1 U12175 ( .B1(n20987), .B2(n20945), .A(n21078), .ZN(n21197) );
  NAND2_X1 U12176 ( .A1(n11250), .A2(n11249), .ZN(n18024) );
  INV_X1 U12177 ( .A(n21078), .ZN(n21068) );
  CLKBUF_X1 U12178 ( .A(n21161), .Z(n21189) );
  INV_X1 U12179 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21216) );
  INV_X1 U12180 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16822) );
  INV_X1 U12181 ( .A(n12433), .ZN(n20789) );
  AOI211_X1 U12182 ( .C1(n21249), .C2(P3_FLUSH_REG_SCAN_IN), .A(n21248), .B(
        n16810), .ZN(n20828) );
  INV_X1 U12183 ( .A(n20828), .ZN(n20826) );
  NOR2_X1 U12184 ( .A1(n21726), .A2(n18214), .ZN(n18194) );
  AND2_X1 U12185 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n21678), .ZN(n21682) );
  INV_X1 U12186 ( .A(n15727), .ZN(n14377) );
  CLKBUF_X1 U12187 ( .A(n18649), .Z(n18977) );
  OAI21_X1 U12188 ( .B1(n15931), .B2(n21638), .A(n11179), .ZN(P1_U2809) );
  AOI21_X1 U12189 ( .B1(n21435), .B2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n11372), .ZN(n21436) );
  OAI21_X1 U12190 ( .B1(n21638), .B2(n11375), .A(n11373), .ZN(n11372) );
  INV_X1 U12191 ( .A(n11111), .ZN(n19973) );
  OAI21_X1 U12192 ( .B1(n21383), .B2(n21639), .A(n11112), .ZN(n11111) );
  INV_X1 U12193 ( .A(n11113), .ZN(n11112) );
  OAI21_X1 U12194 ( .B1(n16341), .B2(n17207), .A(n11226), .ZN(n16344) );
  NOR2_X1 U12195 ( .A1(n11229), .A2(n11227), .ZN(n11226) );
  AOI211_X1 U12196 ( .C1(n17200), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15520), .B(n15497), .ZN(n15498) );
  NAND2_X1 U12197 ( .A1(n11162), .A2(n11161), .ZN(n11160) );
  NAND2_X1 U12198 ( .A1(n11284), .A2(n11016), .ZN(P2_U3015) );
  NAND2_X1 U12199 ( .A1(n18499), .A2(n18553), .ZN(n11281) );
  AOI211_X1 U12200 ( .C1(n11011), .C2(n20560), .A(n20579), .B(n20559), .ZN(
        n20564) );
  OAI211_X1 U12201 ( .C1(n17888), .C2(n20921), .A(n12905), .B(n12904), .ZN(
        n12906) );
  NOR2_X1 U12202 ( .A1(n11008), .A2(n12752), .ZN(n12753) );
  AND4_X1 U12203 ( .A1(n11241), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10983) );
  AND2_X2 U12204 ( .A1(n13335), .A2(n13126), .ZN(n13600) );
  INV_X1 U12205 ( .A(n14994), .ZN(n16170) );
  OR3_X1 U12206 ( .A1(n14972), .A2(n15213), .A3(n11206), .ZN(n10984) );
  NAND3_X2 U12207 ( .A1(n11119), .A2(n11118), .A3(n11030), .ZN(n11685) );
  INV_X1 U12208 ( .A(n18025), .ZN(n11252) );
  INV_X1 U12209 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20183) );
  AND4_X1 U12210 ( .A1(n16404), .A2(n15405), .A3(n15404), .A4(n16409), .ZN(
        n10986) );
  OR2_X1 U12211 ( .A1(n16576), .A2(n11271), .ZN(n10987) );
  AND2_X1 U12212 ( .A1(n11169), .A2(n11167), .ZN(n10989) );
  OR2_X1 U12213 ( .A1(n11336), .A2(n15534), .ZN(n10990) );
  NOR2_X1 U12214 ( .A1(n16652), .A2(n15192), .ZN(n15191) );
  AND2_X1 U12215 ( .A1(n14338), .A2(n13123), .ZN(n10991) );
  AND2_X1 U12216 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10992) );
  INV_X1 U12217 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17106) );
  AND2_X1 U12218 ( .A1(n11234), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10993) );
  AND2_X1 U12219 ( .A1(n13233), .A2(n14965), .ZN(n10994) );
  AND2_X1 U12220 ( .A1(n15036), .A2(n15016), .ZN(n10995) );
  AND2_X1 U12221 ( .A1(n10992), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10996) );
  AND2_X1 U12222 ( .A1(n10991), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10997) );
  INV_X2 U12223 ( .A(n13340), .ZN(n13143) );
  AND2_X1 U12224 ( .A1(n10964), .A2(n11368), .ZN(n10998) );
  AND2_X1 U12225 ( .A1(n11237), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10999) );
  AND2_X1 U12226 ( .A1(n11231), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11000) );
  AND2_X1 U12227 ( .A1(n11045), .A2(n11673), .ZN(n21590) );
  NAND2_X1 U12228 ( .A1(n20547), .A2(n11195), .ZN(n11001) );
  AND2_X1 U12229 ( .A1(n12764), .A2(n21900), .ZN(n20021) );
  AND2_X1 U12230 ( .A1(n15512), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11002) );
  AND2_X1 U12231 ( .A1(n11131), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n11003) );
  AND2_X1 U12232 ( .A1(n11002), .A2(n15515), .ZN(n11004) );
  INV_X2 U12233 ( .A(n21702), .ZN(n17281) );
  NOR2_X2 U12234 ( .A1(n12434), .A2(n11244), .ZN(n12529) );
  AND2_X2 U12235 ( .A1(n13396), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13271) );
  OR3_X1 U12236 ( .A1(n16576), .A2(n11271), .A3(n11273), .ZN(n11005) );
  OR2_X1 U12237 ( .A1(n16652), .A2(n11291), .ZN(n11006) );
  NAND2_X2 U12238 ( .A1(n11656), .A2(n10954), .ZN(n11696) );
  NAND2_X1 U12239 ( .A1(n11095), .A2(n15342), .ZN(n16480) );
  AND2_X2 U12240 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11422) );
  NOR2_X1 U12241 ( .A1(n15232), .A2(n15642), .ZN(n15641) );
  AND2_X1 U12242 ( .A1(n15676), .A2(n12247), .ZN(n15668) );
  NAND2_X1 U12243 ( .A1(n16483), .A2(n16482), .ZN(n16484) );
  XNOR2_X1 U12244 ( .A(n15553), .B(n15552), .ZN(n18499) );
  OR2_X1 U12245 ( .A1(n14935), .A2(n15161), .ZN(n15160) );
  AND2_X1 U12246 ( .A1(n16198), .A2(n11218), .ZN(n11007) );
  NOR3_X1 U12247 ( .A1(n12751), .A2(n21150), .A3(n17847), .ZN(n11008) );
  NAND2_X1 U12248 ( .A1(n15392), .A2(n11153), .ZN(n11009) );
  NAND2_X1 U12249 ( .A1(n11215), .A2(n11214), .ZN(n11213) );
  AND2_X1 U12250 ( .A1(n18511), .A2(n14998), .ZN(n11010) );
  XOR2_X1 U12251 ( .A(n20566), .B(n20567), .Z(n11011) );
  OR2_X1 U12252 ( .A1(n11695), .A2(n11686), .ZN(n11012) );
  NAND2_X1 U12253 ( .A1(n11353), .A2(n11355), .ZN(n15701) );
  NOR2_X1 U12254 ( .A1(n15232), .A2(n11357), .ZN(n15710) );
  NAND2_X1 U12255 ( .A1(n15138), .A2(n15137), .ZN(n15460) );
  NAND2_X1 U12256 ( .A1(n15122), .A2(n15472), .ZN(n15139) );
  NOR2_X1 U12257 ( .A1(n16209), .A2(n16210), .ZN(n16198) );
  INV_X1 U12258 ( .A(n11369), .ZN(n11828) );
  OR3_X1 U12259 ( .A1(n16492), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15549), .ZN(n11013) );
  NAND2_X1 U12260 ( .A1(n11342), .A2(n15435), .ZN(n16384) );
  OR2_X1 U12261 ( .A1(n15605), .A2(n11359), .ZN(n12755) );
  NAND2_X1 U12262 ( .A1(n16567), .A2(n11004), .ZN(n15493) );
  XNOR2_X1 U12263 ( .A(n15472), .B(n15473), .ZN(n15458) );
  INV_X1 U12264 ( .A(n15458), .ZN(n11129) );
  OAI211_X1 U12265 ( .C1(n16187), .C2(n16191), .A(n16182), .B(n16188), .ZN(
        n16174) );
  INV_X1 U12266 ( .A(n14129), .ZN(n13023) );
  NAND2_X1 U12267 ( .A1(n11904), .A2(n11367), .ZN(n12823) );
  XNOR2_X1 U12268 ( .A(n15560), .B(n15559), .ZN(n16341) );
  AND2_X1 U12269 ( .A1(n15446), .A2(n11340), .ZN(n11014) );
  AND2_X1 U12270 ( .A1(n16567), .A2(n11002), .ZN(n16374) );
  NAND2_X1 U12271 ( .A1(n11305), .A2(n11306), .ZN(n14254) );
  AND2_X1 U12272 ( .A1(n15089), .A2(n12841), .ZN(n11015) );
  AND3_X1 U12273 ( .A1(n11384), .A2(n11282), .A3(n11281), .ZN(n11016) );
  NOR2_X1 U12274 ( .A1(n11005), .A2(n16301), .ZN(n16293) );
  AND2_X1 U12275 ( .A1(n11339), .A2(n11336), .ZN(n11017) );
  NOR2_X1 U12276 ( .A1(n16220), .A2(n16219), .ZN(n11018) );
  AND2_X1 U12277 ( .A1(n12966), .A2(n11085), .ZN(n11019) );
  AND2_X1 U12278 ( .A1(n12798), .A2(n11594), .ZN(n11020) );
  AND2_X1 U12279 ( .A1(n13579), .A2(n17222), .ZN(n11021) );
  AND2_X1 U12280 ( .A1(n12853), .A2(n12851), .ZN(n11022) );
  INV_X1 U12281 ( .A(n11683), .ZN(n12758) );
  INV_X1 U12282 ( .A(n12992), .ZN(n12953) );
  AND2_X1 U12283 ( .A1(n11688), .A2(n11685), .ZN(n11023) );
  AND2_X1 U12284 ( .A1(n11086), .A2(n12966), .ZN(n11024) );
  AND4_X1 U12285 ( .A1(n12468), .A2(n12472), .A3(n11102), .A4(n11101), .ZN(
        n11025) );
  AND2_X1 U12286 ( .A1(n19947), .A2(n12814), .ZN(n11026) );
  NAND2_X1 U12287 ( .A1(n11779), .A2(n11755), .ZN(n11027) );
  AND2_X1 U12288 ( .A1(n15480), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11028) );
  AND2_X1 U12289 ( .A1(n15448), .A2(n16508), .ZN(n11029) );
  NAND2_X1 U12290 ( .A1(n15121), .A2(n15120), .ZN(n15472) );
  NAND2_X1 U12291 ( .A1(n16198), .A2(n16199), .ZN(n16192) );
  AND3_X1 U12292 ( .A1(n11519), .A2(n11523), .A3(n11520), .ZN(n11030) );
  AND3_X1 U12293 ( .A1(n12392), .A2(n11180), .A3(n11677), .ZN(n11031) );
  AND2_X1 U12294 ( .A1(n15887), .A2(n15890), .ZN(n11032) );
  NAND2_X1 U12295 ( .A1(n18367), .A2(n18369), .ZN(n11033) );
  INV_X1 U12296 ( .A(n14843), .ZN(n14841) );
  NAND2_X1 U12297 ( .A1(n11014), .A2(n11335), .ZN(n11034) );
  NAND2_X1 U12298 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12526), .ZN(
        n11035) );
  NAND2_X1 U12299 ( .A1(n11137), .A2(n11138), .ZN(n13821) );
  NAND2_X1 U12300 ( .A1(n11481), .A2(n11480), .ZN(n11806) );
  BUF_X4 U12301 ( .A(n11475), .Z(n12365) );
  AND2_X1 U12302 ( .A1(n11137), .A2(n11135), .ZN(n12393) );
  AND2_X1 U12303 ( .A1(n11288), .A2(n11286), .ZN(n11036) );
  INV_X1 U12304 ( .A(n13727), .ZN(n13682) );
  NAND2_X1 U12305 ( .A1(n16754), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16755) );
  NOR2_X1 U12306 ( .A1(n14935), .A2(n11351), .ZN(n15199) );
  NAND2_X1 U12307 ( .A1(n11950), .A2(n11951), .ZN(n14696) );
  NAND2_X1 U12308 ( .A1(n14825), .A2(n10994), .ZN(n11037) );
  OR2_X1 U12309 ( .A1(n14842), .A2(n14841), .ZN(n11038) );
  AND2_X1 U12310 ( .A1(n16096), .A2(n11231), .ZN(n11039) );
  AND2_X1 U12311 ( .A1(n15074), .A2(n11234), .ZN(n11040) );
  NOR2_X2 U12312 ( .A1(n14701), .A2(n13734), .ZN(n14825) );
  INV_X1 U12313 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18058) );
  NOR3_X1 U12314 ( .A1(n15720), .A2(n11177), .A3(n11178), .ZN(n15705) );
  AND2_X1 U12315 ( .A1(n10996), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11041) );
  NOR2_X1 U12316 ( .A1(n16249), .A2(n16240), .ZN(n16230) );
  NOR2_X2 U12317 ( .A1(n11701), .A2(n21922), .ZN(n12069) );
  INV_X1 U12318 ( .A(n12069), .ZN(n11371) );
  INV_X1 U12319 ( .A(n12991), .ZN(n13783) );
  INV_X1 U12320 ( .A(n13968), .ZN(n11083) );
  NAND2_X1 U12321 ( .A1(n17839), .A2(n18087), .ZN(n17881) );
  NAND2_X1 U12322 ( .A1(n11937), .A2(n11936), .ZN(n14800) );
  NOR2_X1 U12323 ( .A1(n21540), .A2(n21539), .ZN(n21538) );
  NOR3_X1 U12324 ( .A1(n15689), .A2(n15678), .A3(n11171), .ZN(n11173) );
  NAND2_X1 U12325 ( .A1(n21538), .A2(n11003), .ZN(n21571) );
  NAND2_X1 U12326 ( .A1(n12661), .A2(n21103), .ZN(n17697) );
  NOR2_X1 U12327 ( .A1(n15638), .A2(n19884), .ZN(n15612) );
  AND2_X1 U12328 ( .A1(n15566), .A2(n15576), .ZN(n11704) );
  AND2_X1 U12329 ( .A1(n16255), .A2(n13296), .ZN(n16243) );
  NAND2_X1 U12330 ( .A1(n14825), .A2(n13233), .ZN(n14920) );
  OR2_X1 U12331 ( .A1(n14972), .A2(n11208), .ZN(n11042) );
  OR3_X1 U12332 ( .A1(n15689), .A2(n15678), .A3(n11172), .ZN(n11043) );
  NOR2_X1 U12333 ( .A1(n16576), .A2(n16577), .ZN(n16314) );
  OR2_X1 U12334 ( .A1(n16652), .A2(n11294), .ZN(n11044) );
  NOR2_X1 U12335 ( .A1(n14660), .A2(n11141), .ZN(n11045) );
  OAI21_X1 U12336 ( .B1(n11332), .B2(n11330), .A(n17139), .ZN(n11329) );
  INV_X1 U12337 ( .A(n11329), .ZN(n11322) );
  OR2_X1 U12338 ( .A1(n15720), .A2(n15719), .ZN(n11046) );
  AND2_X1 U12339 ( .A1(n11698), .A2(n11714), .ZN(n11047) );
  INV_X1 U12340 ( .A(n11268), .ZN(n17997) );
  OR2_X1 U12341 ( .A1(n11359), .A2(n12757), .ZN(n11048) );
  NAND2_X1 U12342 ( .A1(n14724), .A2(n14723), .ZN(n14842) );
  INV_X1 U12343 ( .A(n14842), .ZN(n11149) );
  AND2_X1 U12344 ( .A1(n11041), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11049) );
  INV_X1 U12345 ( .A(n15232), .ZN(n11353) );
  INV_X2 U12346 ( .A(n19993), .ZN(n19971) );
  INV_X2 U12347 ( .A(n12852), .ZN(n19993) );
  INV_X1 U12348 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11376) );
  NAND2_X2 U12349 ( .A1(n13722), .A2(n13721), .ZN(n11050) );
  AND2_X1 U12350 ( .A1(n11941), .A2(n11571), .ZN(n11051) );
  NOR3_X1 U12351 ( .A1(n15689), .A2(n15678), .A3(n11174), .ZN(n15671) );
  AND2_X1 U12352 ( .A1(n11080), .A2(n13968), .ZN(n11052) );
  AND2_X1 U12353 ( .A1(n19963), .A2(n12841), .ZN(n11053) );
  AND2_X1 U12354 ( .A1(n11268), .A2(n11266), .ZN(n11054) );
  INV_X1 U12355 ( .A(n13702), .ZN(n11277) );
  AND2_X1 U12356 ( .A1(n11316), .A2(n15208), .ZN(n11055) );
  AND2_X1 U12357 ( .A1(n10995), .A2(n15052), .ZN(n11056) );
  NAND2_X1 U12358 ( .A1(n14339), .A2(n14338), .ZN(n14319) );
  AND2_X1 U12359 ( .A1(n17815), .A2(n10996), .ZN(n11057) );
  AND3_X1 U12360 ( .A1(n11204), .A2(n13585), .A3(n11205), .ZN(n13578) );
  NOR2_X1 U12361 ( .A1(n15235), .A2(n19866), .ZN(n15236) );
  NAND2_X1 U12362 ( .A1(n21529), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15235) );
  NAND4_X1 U12363 ( .A1(n11204), .A2(n13585), .A3(n11205), .A4(n14136), .ZN(
        n14119) );
  NOR2_X1 U12364 ( .A1(n14707), .A2(n11213), .ZN(n14901) );
  NAND2_X1 U12365 ( .A1(n14999), .A2(n15006), .ZN(n15104) );
  AND2_X1 U12366 ( .A1(n16099), .A2(n11237), .ZN(n11058) );
  AND2_X1 U12367 ( .A1(n13967), .A2(n18619), .ZN(n11059) );
  NOR2_X1 U12368 ( .A1(n17766), .A2(n20424), .ZN(n17768) );
  NOR2_X1 U12369 ( .A1(n17802), .A2(n17818), .ZN(n17815) );
  OR2_X1 U12370 ( .A1(n16144), .A2(n15376), .ZN(n11060) );
  AND2_X1 U12371 ( .A1(n13296), .A2(n16244), .ZN(n11061) );
  INV_X1 U12372 ( .A(n15582), .ZN(n21664) );
  AND2_X1 U12373 ( .A1(n12145), .A2(n12144), .ZN(n11062) );
  INV_X1 U12374 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18249) );
  INV_X1 U12375 ( .A(n19928), .ZN(n11174) );
  NAND2_X1 U12376 ( .A1(n12539), .A2(n12663), .ZN(n17869) );
  INV_X1 U12377 ( .A(n17869), .ZN(n17971) );
  AND2_X1 U12378 ( .A1(n21538), .A2(n11131), .ZN(n11063) );
  AND2_X1 U12379 ( .A1(n11193), .A2(n11191), .ZN(n11064) );
  AND2_X1 U12380 ( .A1(n11315), .A2(n11314), .ZN(n11065) );
  AND2_X1 U12381 ( .A1(n11254), .A2(n11253), .ZN(n11066) );
  INV_X1 U12382 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21655) );
  INV_X1 U12383 ( .A(n20520), .ZN(n11195) );
  NAND2_X1 U12384 ( .A1(n14259), .A2(n13826), .ZN(n13858) );
  NAND2_X1 U12385 ( .A1(n12393), .A2(n16868), .ZN(n21639) );
  INV_X1 U12386 ( .A(n21639), .ZN(n20020) );
  NOR2_X1 U12387 ( .A1(n18014), .A2(n17944), .ZN(n17743) );
  AND2_X1 U12388 ( .A1(n17815), .A2(n11041), .ZN(n11067) );
  OR2_X1 U12389 ( .A1(n15490), .A2(n16112), .ZN(n11068) );
  AND2_X1 U12390 ( .A1(n13774), .A2(n13773), .ZN(n11069) );
  INV_X1 U12391 ( .A(n11704), .ZN(n11134) );
  INV_X1 U12392 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11201) );
  INV_X1 U12393 ( .A(n21434), .ZN(n11375) );
  AND3_X1 U12394 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(n11184), .ZN(n17943) );
  NAND2_X1 U12395 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11070) );
  AND2_X1 U12396 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11071) );
  AND2_X1 U12397 ( .A1(n11003), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n11072) );
  AND2_X1 U12398 ( .A1(n11004), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11073) );
  INV_X1 U12399 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11200) );
  INV_X1 U12400 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11185) );
  INV_X1 U12401 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11246) );
  NOR2_X1 U12402 ( .A1(n17706), .A2(n17785), .ZN(n17705) );
  OAI21_X1 U12403 ( .B1(n20024), .B2(n21515), .A(n11114), .ZN(n11113) );
  OAI22_X2 U12404 ( .A1(n20072), .A2(n14567), .B1(n16916), .B2(n14566), .ZN(
        n22164) );
  NAND2_X1 U12405 ( .A1(n20021), .A2(n14377), .ZN(n14567) );
  NOR4_X2 U12406 ( .A1(n20943), .A2(n20927), .A3(n17869), .A4(n17718), .ZN(
        n17984) );
  NOR2_X2 U12407 ( .A1(n20740), .A2(n18773), .ZN(n18724) );
  OAI22_X2 U12408 ( .A1(n20064), .A2(n14567), .B1(n17002), .B2(n14566), .ZN(
        n22001) );
  OAI22_X2 U12409 ( .A1(n20070), .A2(n14567), .B1(n17017), .B2(n14566), .ZN(
        n22121) );
  NOR4_X4 U12410 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n20785), .ZN(n20560) );
  NOR2_X2 U12411 ( .A1(n13982), .A2(n19585), .ZN(n14091) );
  NAND4_X1 U12412 ( .A1(n12923), .A2(n12921), .A3(n12922), .A4(n12920), .ZN(
        n11079) );
  NAND2_X4 U12413 ( .A1(n11078), .A2(n11076), .ZN(n13579) );
  NAND4_X1 U12414 ( .A1(n12925), .A2(n12927), .A3(n12924), .A4(n12926), .ZN(
        n11077) );
  NAND3_X1 U12415 ( .A1(n13899), .A2(n11082), .A3(n11080), .ZN(n11086) );
  INV_X1 U12416 ( .A(n13905), .ZN(n11081) );
  NAND2_X1 U12417 ( .A1(n13010), .A2(n13583), .ZN(n14132) );
  AND2_X2 U12418 ( .A1(n14132), .A2(n11088), .ZN(n13055) );
  NAND2_X1 U12419 ( .A1(n16752), .A2(n16753), .ZN(n11095) );
  INV_X1 U12420 ( .A(n15342), .ZN(n11094) );
  OAI211_X2 U12421 ( .C1(n11095), .C2(n11092), .A(n11090), .B(n11331), .ZN(
        n11328) );
  NAND3_X1 U12422 ( .A1(n15017), .A2(n15037), .A3(n10995), .ZN(n15054) );
  NAND3_X1 U12423 ( .A1(n15017), .A2(n15037), .A3(n11056), .ZN(n15119) );
  NAND3_X1 U12424 ( .A1(n11025), .A2(n12466), .A3(n11098), .ZN(n20644) );
  NAND2_X2 U12425 ( .A1(n19963), .A2(n11015), .ZN(n15088) );
  NAND2_X2 U12426 ( .A1(n15921), .A2(n12854), .ZN(n15887) );
  NAND2_X2 U12427 ( .A1(n15088), .A2(n11022), .ZN(n15921) );
  NAND4_X1 U12428 ( .A1(n11719), .A2(n11713), .A3(n11107), .A4(n11047), .ZN(
        n11707) );
  OAI21_X2 U12429 ( .B1(n11785), .B2(n11718), .A(n11717), .ZN(n11110) );
  INV_X2 U12430 ( .A(n11685), .ZN(n14410) );
  NAND3_X1 U12431 ( .A1(n11124), .A2(n11123), .A3(n11122), .ZN(n11121) );
  INV_X1 U12432 ( .A(n16774), .ZN(n11125) );
  AND2_X1 U12433 ( .A1(n11126), .A2(n13901), .ZN(n11205) );
  OAI21_X1 U12434 ( .B1(n13901), .B2(n11393), .A(n11126), .ZN(n13008) );
  INV_X2 U12435 ( .A(n13334), .ZN(n13396) );
  AOI22_X1 U12436 ( .A1(n13476), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12921) );
  INV_X2 U12437 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14490) );
  NAND2_X1 U12438 ( .A1(n15594), .A2(n10951), .ZN(P1_U2810) );
  AOI21_X1 U12439 ( .B1(n11680), .B2(n14410), .A(n11702), .ZN(n11546) );
  INV_X1 U12440 ( .A(n14597), .ZN(n14593) );
  INV_X1 U12441 ( .A(n14886), .ZN(n11148) );
  INV_X1 U12442 ( .A(n13128), .ZN(n13457) );
  AND2_X2 U12443 ( .A1(n10979), .A2(n13511), .ZN(n13156) );
  NAND2_X1 U12444 ( .A1(n11159), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13107) );
  OAI21_X1 U12445 ( .B1(n11159), .B2(n11409), .A(n13060), .ZN(n13064) );
  AOI21_X2 U12446 ( .B1(n11159), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13034), .ZN(n13047) );
  AOI21_X1 U12447 ( .B1(n11159), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13066), .ZN(n13073) );
  NAND2_X2 U12448 ( .A1(n13022), .A2(n13051), .ZN(n11159) );
  OAI21_X2 U12449 ( .B1(n16774), .B2(n11050), .A(n15038), .ZN(n15044) );
  NOR2_X2 U12450 ( .A1(n11165), .A2(n18538), .ZN(n17183) );
  OR2_X2 U12452 ( .A1(n11438), .A2(n11437), .ZN(n12777) );
  INV_X1 U12453 ( .A(n11173), .ZN(n15634) );
  INV_X1 U12454 ( .A(n15706), .ZN(n11178) );
  XNOR2_X2 U12455 ( .A(n17896), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n20396) );
  NAND3_X1 U12456 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(n11182), .ZN(n18014) );
  NAND2_X1 U12457 ( .A1(n20406), .A2(n20396), .ZN(n11188) );
  NAND2_X1 U12458 ( .A1(n11188), .A2(n11186), .ZN(n11189) );
  INV_X1 U12459 ( .A(n11190), .ZN(n20419) );
  INV_X1 U12460 ( .A(n11189), .ZN(n20432) );
  INV_X1 U12461 ( .A(n11196), .ZN(n20519) );
  AND2_X1 U12462 ( .A1(n20322), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11199) );
  INV_X1 U12463 ( .A(n14119), .ZN(n13036) );
  NOR2_X1 U12464 ( .A1(n14972), .A2(n14971), .ZN(n15180) );
  INV_X1 U12465 ( .A(n14707), .ZN(n11210) );
  NAND2_X1 U12466 ( .A1(n11210), .A2(n11211), .ZN(n14905) );
  NAND2_X1 U12467 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11240) );
  NAND3_X1 U12468 ( .A1(n11241), .A2(n11239), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14865) );
  NAND3_X1 U12469 ( .A1(n11241), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14863) );
  NAND2_X2 U12470 ( .A1(n20808), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11244) );
  AND2_X2 U12471 ( .A1(n11247), .A2(n17869), .ZN(n17785) );
  INV_X1 U12472 ( .A(n11254), .ZN(n18034) );
  INV_X1 U12473 ( .A(n12511), .ZN(n11253) );
  NAND2_X1 U12474 ( .A1(n17846), .A2(n17847), .ZN(n17845) );
  OAI21_X1 U12475 ( .B1(n17846), .B2(n11257), .A(n11255), .ZN(n11259) );
  INV_X1 U12476 ( .A(n17762), .ZN(n11260) );
  NAND2_X1 U12477 ( .A1(n11261), .A2(n11260), .ZN(n11263) );
  AND2_X1 U12478 ( .A1(n11263), .A2(n11264), .ZN(n12556) );
  OAI21_X1 U12479 ( .B1(n17833), .B2(n11265), .A(n17869), .ZN(n11264) );
  NAND3_X1 U12480 ( .A1(n13005), .A2(n13579), .A3(n14097), .ZN(n13006) );
  NAND2_X1 U12481 ( .A1(n14846), .A2(n13702), .ZN(n11274) );
  NAND2_X1 U12482 ( .A1(n11274), .A2(n11275), .ZN(n13724) );
  NOR2_X2 U12483 ( .A1(n16725), .A2(n11285), .ZN(n15080) );
  NAND3_X1 U12484 ( .A1(n11293), .A2(n16328), .A3(n11292), .ZN(n11291) );
  NAND2_X1 U12485 ( .A1(n13084), .A2(n13083), .ZN(n11306) );
  NAND2_X1 U12486 ( .A1(n16220), .A2(n11311), .ZN(n11307) );
  INV_X1 U12487 ( .A(n11309), .ZN(n11308) );
  INV_X1 U12488 ( .A(n13408), .ZN(n11311) );
  INV_X1 U12489 ( .A(n16219), .ZN(n11313) );
  NAND2_X1 U12490 ( .A1(n14825), .A2(n11055), .ZN(n15207) );
  NAND2_X1 U12491 ( .A1(n15037), .A2(n15036), .ZN(n11317) );
  NAND2_X1 U12492 ( .A1(n15017), .A2(n15016), .ZN(n11318) );
  NAND2_X1 U12493 ( .A1(n11318), .A2(n11317), .ZN(n11319) );
  INV_X1 U12494 ( .A(n11325), .ZN(n11320) );
  INV_X1 U12495 ( .A(n15447), .ZN(n11334) );
  OAI21_X1 U12496 ( .B1(n11334), .B2(n11034), .A(n10990), .ZN(n15492) );
  NAND2_X1 U12497 ( .A1(n15447), .A2(n11014), .ZN(n11339) );
  NAND2_X1 U12498 ( .A1(n11342), .A2(n11341), .ZN(n16369) );
  OAI21_X1 U12499 ( .B1(n16483), .B2(n11347), .A(n11345), .ZN(n17128) );
  NAND2_X2 U12500 ( .A1(n11344), .A2(n11343), .ZN(n16416) );
  NAND2_X1 U12501 ( .A1(n16483), .A2(n11345), .ZN(n11344) );
  NAND3_X2 U12502 ( .A1(n15469), .A2(n15140), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15459) );
  AND2_X2 U12503 ( .A1(n16567), .A2(n11073), .ZN(n16354) );
  OR2_X2 U12504 ( .A1(n14935), .A2(n11349), .ZN(n15200) );
  NOR2_X2 U12505 ( .A1(n15232), .A2(n11354), .ZN(n15702) );
  NAND3_X1 U12506 ( .A1(n11950), .A2(n11951), .A3(n11396), .ZN(n14743) );
  NOR2_X2 U12507 ( .A1(n14743), .A2(n14810), .ZN(n14808) );
  NOR2_X1 U12508 ( .A1(n15605), .A2(n15606), .ZN(n15595) );
  NOR2_X2 U12509 ( .A1(n15605), .A2(n11048), .ZN(n12756) );
  NAND2_X1 U12510 ( .A1(n15676), .A2(n11361), .ZN(n15618) );
  AND2_X1 U12511 ( .A1(n15676), .A2(n11362), .ZN(n15629) );
  INV_X1 U12512 ( .A(n15618), .ZN(n12312) );
  NAND2_X1 U12513 ( .A1(n11904), .A2(n11903), .ZN(n11938) );
  CLKBUF_X1 U12514 ( .A(n11374), .Z(n11368) );
  OAI21_X1 U12515 ( .B1(n14315), .B2(n11371), .A(n11370), .ZN(n11369) );
  INV_X1 U12516 ( .A(n11827), .ZN(n11370) );
  AOI21_X1 U12517 ( .B1(n11368), .B2(n16083), .A(n13957), .ZN(n16854) );
  NAND2_X1 U12518 ( .A1(n21456), .A2(n11368), .ZN(n11373) );
  AND2_X2 U12519 ( .A1(n11418), .A2(n11419), .ZN(n11846) );
  NAND2_X1 U12520 ( .A1(n14304), .A2(n12798), .ZN(n12806) );
  NAND2_X1 U12521 ( .A1(n14611), .A2(n14613), .ZN(n12807) );
  NAND2_X1 U12522 ( .A1(n15887), .A2(n11381), .ZN(n11377) );
  OAI21_X2 U12523 ( .B1(n15826), .B2(n15827), .A(n19993), .ZN(n15849) );
  OR3_X4 U12524 ( .A1(n17705), .A2(n21019), .A3(n17703), .ZN(n17762) );
  AOI21_X1 U12525 ( .B1(n16345), .B2(n17203), .A(n16344), .ZN(n16346) );
  CLKBUF_X1 U12526 ( .A(n15207), .Z(n16264) );
  NAND2_X1 U12527 ( .A1(n16216), .A2(n15279), .ZN(n16209) );
  NOR2_X1 U12528 ( .A1(n17973), .A2(n21139), .ZN(n12550) );
  AND2_X1 U12529 ( .A1(n14125), .A2(n13055), .ZN(n13056) );
  OR2_X2 U12530 ( .A1(n15869), .A2(n20002), .ZN(n15870) );
  INV_X1 U12531 ( .A(n16216), .ZN(n16227) );
  NOR2_X2 U12532 ( .A1(n18068), .A2(n18069), .ZN(n18067) );
  INV_X1 U12533 ( .A(n14679), .ZN(n13169) );
  INV_X1 U12534 ( .A(n13069), .ZN(n13070) );
  INV_X1 U12535 ( .A(n14698), .ZN(n11951) );
  NAND2_X1 U12536 ( .A1(n13562), .A2(n13837), .ZN(n13585) );
  INV_X1 U12537 ( .A(n11709), .ZN(n11701) );
  OR2_X1 U12538 ( .A1(n14245), .A2(n14244), .ZN(n14246) );
  AND2_X1 U12539 ( .A1(n13102), .A2(n13100), .ZN(n13076) );
  INV_X1 U12540 ( .A(n14998), .ZN(n14988) );
  BUF_X2 U12541 ( .A(n14998), .Z(n17101) );
  INV_X1 U12542 ( .A(n14064), .ZN(n14070) );
  NAND4_X1 U12543 ( .A1(n11702), .A2(n14268), .A3(n11700), .A4(n12418), .ZN(
        n14064) );
  NAND2_X1 U12544 ( .A1(n14676), .A2(n14675), .ZN(n14707) );
  NAND2_X1 U12545 ( .A1(n16230), .A2(n16231), .ZN(n16233) );
  INV_X1 U12546 ( .A(n14677), .ZN(n14676) );
  NAND2_X1 U12547 ( .A1(n10956), .A2(n11400), .ZN(n20381) );
  INV_X1 U12548 ( .A(n20396), .ZN(n11194) );
  NAND2_X1 U12549 ( .A1(n10967), .A2(n19642), .ZN(n13562) );
  NAND2_X1 U12550 ( .A1(n12774), .A2(n12406), .ZN(n12423) );
  INV_X1 U12551 ( .A(n11583), .ZN(n12384) );
  INV_X1 U12552 ( .A(n12384), .ZN(n12378) );
  OR2_X1 U12553 ( .A1(n16341), .A2(n18512), .ZN(n11384) );
  AND2_X1 U12554 ( .A1(n13591), .A2(n13035), .ZN(n11385) );
  NOR2_X1 U12555 ( .A1(n21831), .A2(n21849), .ZN(n11386) );
  AND2_X1 U12556 ( .A1(n19971), .A2(n12875), .ZN(n11387) );
  NOR2_X1 U12557 ( .A1(n21538), .A2(n21601), .ZN(n11388) );
  AND2_X1 U12558 ( .A1(n12400), .A2(n15576), .ZN(n11389) );
  INV_X1 U12559 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12489) );
  OR2_X1 U12560 ( .A1(n15535), .A2(n15542), .ZN(n11391) );
  OR2_X1 U12561 ( .A1(n11696), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11392) );
  NAND2_X1 U12562 ( .A1(n11938), .A2(n11939), .ZN(n12824) );
  AND2_X1 U12563 ( .A1(n12964), .A2(n12992), .ZN(n11393) );
  INV_X1 U12564 ( .A(n14598), .ZN(n11693) );
  AND2_X1 U12565 ( .A1(n13424), .A2(n13445), .ZN(n11394) );
  CLKBUF_X3 U12566 ( .A(n12465), .Z(n17498) );
  NAND2_X1 U12567 ( .A1(n13135), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11395) );
  INV_X1 U12568 ( .A(n13605), .ZN(n13692) );
  INV_X1 U12569 ( .A(n13597), .ZN(n12952) );
  NAND3_X1 U12570 ( .A1(n11965), .A2(n11964), .A3(n11963), .ZN(n11396) );
  AND4_X1 U12571 ( .A1(n15519), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15518), .A4(n15517), .ZN(n11397) );
  OR2_X1 U12572 ( .A1(n17827), .A2(n17765), .ZN(n11398) );
  OR2_X1 U12573 ( .A1(n11696), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11399) );
  INV_X1 U12574 ( .A(n12425), .ZN(n20184) );
  NOR2_X1 U12575 ( .A1(n12430), .A2(n12431), .ZN(n12517) );
  OR2_X1 U12576 ( .A1(n20380), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11400) );
  INV_X1 U12577 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12891) );
  AND4_X1 U12578 ( .A1(n12479), .A2(n12478), .A3(n12477), .A4(n12476), .ZN(
        n11401) );
  AND2_X1 U12579 ( .A1(n12386), .A2(P1_EAX_REG_5__SCAN_IN), .ZN(n11402) );
  INV_X1 U12580 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12747) );
  AND2_X1 U12581 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11403) );
  OR2_X1 U12582 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11404) );
  OR2_X1 U12583 ( .A1(n11696), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11405) );
  NAND2_X1 U12584 ( .A1(n13168), .A2(n13167), .ZN(n11406) );
  AND4_X1 U12585 ( .A1(n11416), .A2(n11415), .A3(n11414), .A4(n11413), .ZN(
        n11407) );
  OR2_X1 U12586 ( .A1(n11568), .A2(n11582), .ZN(n11408) );
  CLKBUF_X3 U12587 ( .A(n12529), .Z(n17520) );
  AND3_X1 U12588 ( .A1(n14136), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11085), 
        .ZN(n11409) );
  NAND2_X1 U12589 ( .A1(n14727), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18227) );
  BUF_X2 U12590 ( .A(n14995), .Z(n15005) );
  AND2_X2 U12591 ( .A1(n11420), .A2(n16085), .ZN(n11841) );
  AND4_X1 U12592 ( .A1(n11427), .A2(n11426), .A3(n11425), .A4(n11424), .ZN(
        n11410) );
  OAI21_X1 U12593 ( .B1(n11689), .B2(n11686), .A(n11527), .ZN(n11528) );
  INV_X1 U12594 ( .A(n11528), .ZN(n11529) );
  OR2_X1 U12595 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11834), .ZN(
        n11555) );
  OR2_X1 U12596 ( .A1(n11533), .A2(n11580), .ZN(n11534) );
  NAND2_X1 U12597 ( .A1(n13041), .A2(n19478), .ZN(n12966) );
  INV_X1 U12598 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11718) );
  OAI211_X1 U12599 ( .C1(n15300), .C2(n18577), .A(n13068), .B(n13067), .ZN(
        n13069) );
  AOI22_X1 U12600 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12961) );
  NOR2_X1 U12601 ( .A1(n11538), .A2(n14410), .ZN(n11537) );
  OR2_X1 U12602 ( .A1(n11925), .A2(n11924), .ZN(n12835) );
  NAND2_X1 U12603 ( .A1(n11696), .A2(n11695), .ZN(n11698) );
  AOI22_X1 U12604 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11477) );
  NOR2_X1 U12605 ( .A1(n13812), .A2(n14142), .ZN(n13037) );
  INV_X1 U12606 ( .A(n13558), .ZN(n13512) );
  OR2_X1 U12607 ( .A1(n12703), .A2(n12716), .ZN(n12699) );
  OR2_X1 U12608 ( .A1(n11565), .A2(n11564), .ZN(n11567) );
  NAND2_X1 U12609 ( .A1(n11687), .A2(n12776), .ZN(n11692) );
  INV_X1 U12610 ( .A(n15169), .ZN(n12013) );
  INV_X1 U12611 ( .A(n11939), .ZN(n11940) );
  INV_X1 U12612 ( .A(n15234), .ZN(n12076) );
  AND4_X1 U12613 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11490) );
  NOR2_X1 U12614 ( .A1(n13579), .A2(n12991), .ZN(n12965) );
  OAI21_X1 U12615 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n20794), .A(
        n12699), .ZN(n12705) );
  AND2_X1 U12616 ( .A1(n17976), .A2(n20956), .ZN(n12543) );
  NAND2_X1 U12617 ( .A1(n11567), .A2(n11566), .ZN(n11582) );
  INV_X1 U12618 ( .A(n15746), .ZN(n12247) );
  INV_X1 U12619 ( .A(n11935), .ZN(n11936) );
  INV_X1 U12620 ( .A(n15621), .ZN(n12311) );
  AND2_X1 U12621 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n12284), .ZN(
        n12285) );
  INV_X1 U12622 ( .A(n11824), .ZN(n12330) );
  INV_X1 U12623 ( .A(n11662), .ZN(n11642) );
  AND2_X1 U12624 ( .A1(n13700), .A2(n13699), .ZN(n15336) );
  AND2_X1 U12625 ( .A1(n13425), .A2(n11394), .ZN(n13426) );
  NAND2_X1 U12626 ( .A1(n11018), .A2(n11311), .ZN(n13409) );
  AND2_X1 U12627 ( .A1(n13681), .A2(n13680), .ZN(n15115) );
  INV_X1 U12628 ( .A(n18227), .ZN(n13031) );
  NAND2_X1 U12629 ( .A1(n13075), .A2(n13074), .ZN(n13100) );
  INV_X1 U12630 ( .A(n15479), .ZN(n15480) );
  OR2_X1 U12631 ( .A1(n15478), .A2(n10966), .ZN(n15479) );
  INV_X1 U12632 ( .A(n15466), .ZN(n15467) );
  INV_X1 U12633 ( .A(n19534), .ZN(n14097) );
  NAND2_X1 U12634 ( .A1(n12988), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12989) );
  INV_X1 U12635 ( .A(n17658), .ZN(n17406) );
  AND2_X1 U12636 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12496), .ZN(
        n12497) );
  INV_X1 U12637 ( .A(n12430), .ZN(n20810) );
  NAND2_X1 U12638 ( .A1(n20156), .A2(n20693), .ZN(n12657) );
  NOR2_X1 U12639 ( .A1(n11686), .A2(n11685), .ZN(n12776) );
  INV_X1 U12640 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11996) );
  NOR2_X1 U12641 ( .A1(n11402), .A2(n11913), .ZN(n11914) );
  NAND2_X1 U12642 ( .A1(n12285), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12333) );
  NAND2_X1 U12643 ( .A1(n11992), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11997) );
  AND2_X1 U12644 ( .A1(n11617), .A2(n11616), .ZN(n19921) );
  OR2_X1 U12645 ( .A1(n11852), .A2(n11851), .ZN(n12803) );
  INV_X1 U12646 ( .A(n15942), .ZN(n16063) );
  NAND2_X1 U12647 ( .A1(n11839), .A2(n11838), .ZN(n14381) );
  INV_X1 U12648 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21880) );
  INV_X1 U12649 ( .A(n15576), .ZN(n12394) );
  INV_X1 U12650 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n11585) );
  AND2_X1 U12651 ( .A1(n14142), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13082) );
  BUF_X1 U12652 ( .A(n10965), .Z(n15293) );
  INV_X1 U12653 ( .A(n16342), .ZN(n15563) );
  NOR2_X1 U12654 ( .A1(n18449), .A2(n10966), .ZN(n16349) );
  AND2_X1 U12655 ( .A1(n16611), .A2(n16612), .ZN(n16403) );
  XNOR2_X1 U12656 ( .A(n15478), .B(n10966), .ZN(n15475) );
  NAND2_X1 U12657 ( .A1(n13096), .A2(n13095), .ZN(n14255) );
  INV_X1 U12658 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15263) );
  INV_X1 U12659 ( .A(n20184), .ZN(n17612) );
  BUF_X2 U12660 ( .A(n12557), .Z(n17642) );
  INV_X1 U12661 ( .A(n12695), .ZN(n20814) );
  AND2_X1 U12662 ( .A1(n11630), .A2(n11629), .ZN(n15719) );
  NOR2_X1 U12663 ( .A1(n11997), .A2(n11996), .ZN(n11998) );
  AND2_X1 U12664 ( .A1(n12044), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12059) );
  NOR2_X1 U12665 ( .A1(n11966), .A2(n14754), .ZN(n11992) );
  NAND2_X1 U12666 ( .A1(n21639), .A2(n12769), .ZN(n15898) );
  OR2_X1 U12667 ( .A1(n14080), .A2(n16081), .ZN(n16062) );
  NAND2_X1 U12668 ( .A1(n14437), .A2(n12775), .ZN(n21827) );
  OR2_X1 U12669 ( .A1(n21869), .A2(n21868), .ZN(n21874) );
  OR2_X1 U12670 ( .A1(n14069), .A2(n14068), .ZN(n16880) );
  NAND2_X1 U12671 ( .A1(n15307), .A2(n15436), .ZN(n15440) );
  OR2_X1 U12672 ( .A1(n18221), .A2(n14731), .ZN(n18493) );
  NOR2_X1 U12673 ( .A1(n19369), .A2(n19419), .ZN(n13123) );
  INV_X1 U12674 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18297) );
  NOR2_X1 U12675 ( .A1(n15524), .A2(n15523), .ZN(n15525) );
  OR2_X1 U12676 ( .A1(n16694), .A2(n15511), .ZN(n16575) );
  AND2_X1 U12677 ( .A1(n13020), .A2(n13017), .ZN(n14101) );
  NAND2_X1 U12678 ( .A1(n13089), .A2(n13088), .ZN(n13964) );
  INV_X1 U12679 ( .A(n19258), .ZN(n19293) );
  INV_X1 U12680 ( .A(n19287), .ZN(n19224) );
  NAND2_X1 U12681 ( .A1(n19142), .A2(n19141), .ZN(n19287) );
  NAND2_X1 U12682 ( .A1(n19214), .A2(n17222), .ZN(n19290) );
  OAI21_X1 U12683 ( .B1(n12654), .B2(n21198), .A(n21239), .ZN(n16825) );
  INV_X1 U12684 ( .A(n20586), .ZN(n20562) );
  INV_X1 U12685 ( .A(n20159), .ZN(n20161) );
  AOI211_X1 U12686 ( .C1(n17656), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n12628), .B(n12627), .ZN(n12629) );
  INV_X1 U12687 ( .A(n18772), .ZN(n20655) );
  NAND2_X1 U12688 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n20779), .ZN(n20770) );
  NOR2_X1 U12689 ( .A1(n12486), .A2(n12485), .ZN(n12487) );
  NAND2_X1 U12690 ( .A1(n12661), .A2(n12655), .ZN(n21205) );
  INV_X1 U12691 ( .A(n17917), .ZN(n17897) );
  INV_X1 U12692 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20316) );
  INV_X1 U12693 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20221) );
  NAND2_X1 U12694 ( .A1(n12903), .A2(n21078), .ZN(n12905) );
  NOR2_X1 U12695 ( .A1(n12663), .A2(n17697), .ZN(n21131) );
  INV_X1 U12696 ( .A(n12547), .ZN(n12548) );
  INV_X1 U12697 ( .A(n21153), .ZN(n21103) );
  INV_X1 U12698 ( .A(n20955), .ZN(n21162) );
  NOR2_X1 U12699 ( .A1(n12599), .A2(n12598), .ZN(n20156) );
  NOR3_X1 U12700 ( .A1(n12660), .A2(n20655), .A3(n12652), .ZN(n12655) );
  OR2_X1 U12701 ( .A1(n13822), .A2(n21664), .ZN(n13826) );
  NAND2_X1 U12702 ( .A1(n11998), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12038) );
  AND2_X1 U12703 ( .A1(n21483), .A2(n14596), .ZN(n21634) );
  INV_X1 U12704 ( .A(n12419), .ZN(n12420) );
  NOR2_X1 U12705 ( .A1(n21278), .A2(n19820), .ZN(n14629) );
  INV_X1 U12706 ( .A(n21772), .ZN(n21740) );
  INV_X1 U12707 ( .A(n21777), .ZN(n21744) );
  OR2_X2 U12708 ( .A1(n14259), .A2(n14258), .ZN(n21775) );
  NOR2_X1 U12709 ( .A1(n12196), .A2(n21577), .ZN(n12197) );
  NAND2_X1 U12710 ( .A1(n12079), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12124) );
  NAND2_X1 U12711 ( .A1(n15817), .A2(n12880), .ZN(n12884) );
  NOR2_X1 U12712 ( .A1(n15941), .A2(n14618), .ZN(n21301) );
  INV_X1 U12713 ( .A(n16062), .ZN(n14614) );
  NOR2_X1 U12714 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16813) );
  NOR2_X2 U12715 ( .A1(n21807), .A2(n21827), .ZN(n22189) );
  OAI211_X1 U12716 ( .C1(n21803), .C2(n21802), .A(n21858), .B(n21801), .ZN(
        n22196) );
  NOR2_X2 U12717 ( .A1(n21807), .A2(n21903), .ZN(n22201) );
  OAI21_X1 U12718 ( .B1(n14764), .B2(n14765), .A(n21914), .ZN(n14789) );
  NOR2_X1 U12719 ( .A1(n14441), .A2(n21827), .ZN(n14793) );
  INV_X1 U12720 ( .A(n22208), .ZN(n22069) );
  INV_X1 U12721 ( .A(n22067), .ZN(n22210) );
  INV_X1 U12722 ( .A(n14422), .ZN(n22217) );
  INV_X1 U12723 ( .A(n21827), .ZN(n21872) );
  INV_X1 U12724 ( .A(n22157), .ZN(n22230) );
  NAND2_X1 U12725 ( .A1(n16073), .A2(n12775), .ZN(n21903) );
  INV_X1 U12726 ( .A(n21874), .ZN(n22243) );
  NOR2_X1 U12727 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14380), .ZN(n14570) );
  NOR2_X1 U12728 ( .A1(n16073), .A2(n12775), .ZN(n21890) );
  INV_X1 U12729 ( .A(n22255), .ZN(n22259) );
  AND2_X1 U12730 ( .A1(n10975), .A2(n14368), .ZN(n21905) );
  AND2_X1 U12731 ( .A1(n21649), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n15582) );
  AND2_X1 U12732 ( .A1(n21684), .A2(n11586), .ZN(n11699) );
  INV_X1 U12733 ( .A(n18493), .ZN(n18473) );
  AND2_X1 U12734 ( .A1(n18221), .A2(n14720), .ZN(n18500) );
  INV_X1 U12735 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n14714) );
  XNOR2_X1 U12736 ( .A(n13964), .B(n13093), .ZN(n14169) );
  INV_X1 U12737 ( .A(n19531), .ZN(n19627) );
  AND2_X1 U12738 ( .A1(n17151), .A2(n13870), .ZN(n17163) );
  INV_X1 U12739 ( .A(n17156), .ZN(n17202) );
  INV_X1 U12741 ( .A(n18576), .ZN(n18556) );
  AND2_X1 U12742 ( .A1(n14113), .A2(n18619), .ZN(n14150) );
  NOR2_X1 U12743 ( .A1(n13964), .A2(n13963), .ZN(n19123) );
  NAND2_X1 U12744 ( .A1(n14561), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18606) );
  OAI21_X1 U12745 ( .B1(n19316), .B2(n19315), .A(n19314), .ZN(n19748) );
  NOR2_X1 U12746 ( .A1(n19287), .A2(n19293), .ZN(n19750) );
  INV_X1 U12747 ( .A(n19721), .ZN(n19723) );
  OAI21_X1 U12748 ( .B1(n19251), .B2(n19250), .A(n19249), .ZN(n19717) );
  AND2_X1 U12749 ( .A1(n19225), .A2(n19224), .ZN(n19716) );
  INV_X1 U12750 ( .A(n19695), .ZN(n19698) );
  OAI21_X1 U12751 ( .B1(n19199), .B2(n19198), .A(n19197), .ZN(n19691) );
  AND2_X1 U12752 ( .A1(n19178), .A2(n19224), .ZN(n19690) );
  AND2_X1 U12753 ( .A1(n19142), .A2(n19123), .ZN(n19221) );
  INV_X1 U12754 ( .A(n19600), .ZN(n19678) );
  INV_X1 U12755 ( .A(n19147), .ZN(n19240) );
  INV_X1 U12756 ( .A(n19620), .ZN(n19621) );
  INV_X1 U12757 ( .A(n19734), .ZN(n19749) );
  INV_X1 U12758 ( .A(n19360), .ZN(n19366) );
  OAI21_X1 U12759 ( .B1(n16825), .B2(n20593), .A(n17688), .ZN(n20157) );
  INV_X1 U12760 ( .A(n17688), .ZN(n20108) );
  NOR2_X1 U12761 ( .A1(n20157), .A2(n20156), .ZN(n20159) );
  INV_X1 U12762 ( .A(n20572), .ZN(n20528) );
  NOR2_X1 U12763 ( .A1(n20423), .A2(n17653), .ZN(n17546) );
  INV_X1 U12764 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20190) );
  NOR2_X1 U12765 ( .A1(n20722), .A2(n20723), .ZN(n20721) );
  NAND2_X1 U12766 ( .A1(n20730), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n20729) );
  NOR2_X1 U12767 ( .A1(n20676), .A2(n20681), .ZN(n20675) );
  NOR2_X1 U12768 ( .A1(n20757), .A2(n20756), .ZN(n20755) );
  INV_X1 U12769 ( .A(n20768), .ZN(n20751) );
  AOI22_X1 U12770 ( .A1(n20596), .A2(n20595), .B1(n20594), .B2(n20593), .ZN(
        n20601) );
  INV_X1 U12771 ( .A(n20156), .ZN(n20592) );
  NOR2_X1 U12772 ( .A1(n20151), .A2(n20143), .ZN(n20142) );
  OAI21_X1 U12773 ( .B1(n20163), .B2(n17881), .A(n18773), .ZN(n17879) );
  INV_X1 U12774 ( .A(n17764), .ZN(n17928) );
  NOR2_X2 U12775 ( .A1(n20626), .A2(n20923), .ZN(n21194) );
  NAND2_X1 U12776 ( .A1(n20874), .A2(n21203), .ZN(n21153) );
  NOR2_X2 U12777 ( .A1(n12661), .A2(n21153), .ZN(n21111) );
  OAI22_X1 U12778 ( .A1(n21210), .A2(n17697), .B1(n21211), .B2(n21202), .ZN(
        n21236) );
  INV_X1 U12779 ( .A(n18207), .ZN(n18205) );
  INV_X1 U12780 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n21678) );
  AOI211_X1 U12781 ( .C1(n21590), .C2(n15963), .A(n15593), .B(n15592), .ZN(
        n15594) );
  INV_X1 U12782 ( .A(n21590), .ZN(n21638) );
  INV_X1 U12783 ( .A(n21618), .ZN(n21630) );
  OR2_X1 U12784 ( .A1(n14801), .A2(n14658), .ZN(n19953) );
  INV_X1 U12785 ( .A(n19820), .ZN(n19843) );
  INV_X1 U12786 ( .A(n21775), .ZN(n14264) );
  NAND2_X1 U12787 ( .A1(n12886), .A2(n20020), .ZN(n12887) );
  INV_X1 U12788 ( .A(n19989), .ZN(n20024) );
  INV_X1 U12789 ( .A(n20021), .ZN(n19975) );
  OR2_X1 U12790 ( .A1(n14080), .A2(n14072), .ZN(n21414) );
  OR2_X1 U12791 ( .A1(n14080), .A2(n14067), .ZN(n21382) );
  NAND2_X1 U12792 ( .A1(n21790), .A2(n21890), .ZN(n22193) );
  INV_X1 U12793 ( .A(n21808), .ZN(n22206) );
  INV_X1 U12794 ( .A(n22202), .ZN(n14796) );
  INV_X1 U12795 ( .A(n14793), .ZN(n14582) );
  AOI22_X1 U12796 ( .A1(n21819), .A2(n21823), .B1(n21907), .B2(n21818), .ZN(
        n22214) );
  OR2_X1 U12797 ( .A1(n14441), .A2(n21903), .ZN(n22067) );
  NAND2_X1 U12798 ( .A1(n21828), .A2(n21872), .ZN(n22226) );
  AOI22_X1 U12799 ( .A1(n21856), .A2(n21854), .B1(n21851), .B2(n21850), .ZN(
        n22234) );
  OR2_X1 U12800 ( .A1(n21869), .A2(n21903), .ZN(n22240) );
  AOI22_X1 U12801 ( .A1(n21879), .A2(n21885), .B1(n21907), .B2(n21878), .ZN(
        n22248) );
  NAND2_X1 U12802 ( .A1(n21905), .A2(n21890), .ZN(n22255) );
  NAND2_X1 U12803 ( .A1(n21905), .A2(n21904), .ZN(n22274) );
  NOR2_X1 U12804 ( .A1(n13817), .A2(n13816), .ZN(n18221) );
  NAND2_X1 U12805 ( .A1(n16109), .A2(n16108), .ZN(n18506) );
  INV_X1 U12806 ( .A(n18474), .ZN(n18329) );
  OR3_X1 U12807 ( .A1(n14737), .A2(n14725), .A3(n18489), .ZN(n18494) );
  INV_X1 U12808 ( .A(n18500), .ZN(n18476) );
  NAND2_X1 U12809 ( .A1(n14243), .A2(n14246), .ZN(n19239) );
  NOR2_X1 U12810 ( .A1(n19634), .A2(n19633), .ZN(n19378) );
  AND2_X1 U12811 ( .A1(n13589), .A2(n18619), .ZN(n19531) );
  INV_X1 U12812 ( .A(n17241), .ZN(n17267) );
  INV_X1 U12813 ( .A(n17163), .ZN(n17198) );
  INV_X1 U12814 ( .A(n18244), .ZN(n18511) );
  NAND2_X1 U12815 ( .A1(n14150), .A2(n14525), .ZN(n16767) );
  INV_X1 U12816 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19255) );
  AOI21_X1 U12817 ( .B1(n19311), .B2(n19310), .A(n19639), .ZN(n19754) );
  INV_X1 U12818 ( .A(n19750), .ZN(n19741) );
  NAND2_X1 U12819 ( .A1(n19258), .A2(n19254), .ZN(n19733) );
  NAND2_X1 U12820 ( .A1(n19258), .A2(n19240), .ZN(n19721) );
  NAND2_X1 U12821 ( .A1(n19225), .A2(n19254), .ZN(n19708) );
  NAND2_X1 U12822 ( .A1(n19240), .A2(n19225), .ZN(n19695) );
  NAND2_X1 U12823 ( .A1(n19178), .A2(n19221), .ZN(n19688) );
  NAND2_X1 U12824 ( .A1(n19240), .A2(n19178), .ZN(n19676) );
  AND2_X1 U12825 ( .A1(n19138), .A2(n19137), .ZN(n19435) );
  OR2_X1 U12826 ( .A1(n19143), .A2(n19283), .ZN(n19657) );
  OR2_X1 U12827 ( .A1(n19143), .A2(n19147), .ZN(n19537) );
  AND2_X1 U12828 ( .A1(n14550), .A2(n14549), .ZN(n18617) );
  NAND2_X1 U12829 ( .A1(n21266), .A2(n21236), .ZN(n21270) );
  AND2_X1 U12830 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17595), .ZN(n17611) );
  AND2_X1 U12831 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17317), .ZN(n17431) );
  AND2_X1 U12832 ( .A1(n17438), .A2(n20693), .ZN(n17685) );
  NOR2_X1 U12833 ( .A1(n12524), .A2(n12523), .ZN(n20631) );
  NOR2_X1 U12834 ( .A1(n21253), .A2(n18145), .ZN(n18159) );
  NAND2_X1 U12835 ( .A1(n17688), .A2(n16824), .ZN(n18144) );
  INV_X1 U12836 ( .A(n20151), .ZN(n20145) );
  INV_X1 U12837 ( .A(n18004), .ZN(n17967) );
  INV_X1 U12838 ( .A(n18081), .ZN(n18090) );
  INV_X1 U12839 ( .A(n21194), .ZN(n21150) );
  NAND2_X1 U12840 ( .A1(n10961), .A2(n21068), .ZN(n21086) );
  INV_X1 U12841 ( .A(n20560), .ZN(n21247) );
  INV_X1 U12842 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21252) );
  INV_X1 U12843 ( .A(n21682), .ZN(n21724) );
  INV_X1 U12844 ( .A(n18194), .ZN(n18207) );
  INV_X1 U12845 ( .A(n21682), .ZN(n18214) );
  NAND3_X1 U12846 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .ZN(n21461) );
  INV_X1 U12847 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21460) );
  NOR2_X1 U12848 ( .A1(n21461), .A2(n21460), .ZN(n21467) );
  NAND2_X1 U12849 ( .A1(n21467), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n21479) );
  INV_X1 U12850 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n19852) );
  NOR2_X1 U12851 ( .A1(n21479), .A2(n19852), .ZN(n21494) );
  NAND2_X1 U12852 ( .A1(n21494), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n14746) );
  INV_X1 U12853 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n19855) );
  NOR2_X1 U12854 ( .A1(n14746), .A2(n19855), .ZN(n14816) );
  NAND2_X1 U12855 ( .A1(n14816), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14955) );
  INV_X1 U12856 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n19857) );
  NOR2_X1 U12857 ( .A1(n14955), .A2(n19857), .ZN(n15652) );
  INV_X1 U12858 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11411) );
  INV_X1 U12859 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11412) );
  AND2_X4 U12860 ( .A1(n11420), .A2(n11417), .ZN(n11521) );
  AOI22_X1 U12861 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11416) );
  NOR2_X4 U12862 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U12863 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11460), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11415) );
  AND2_X4 U12864 ( .A1(n11418), .A2(n11422), .ZN(n11736) );
  AOI22_X1 U12865 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11722), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11414) );
  AND2_X2 U12866 ( .A1(n14270), .A2(n16085), .ZN(n11447) );
  AOI22_X1 U12867 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11413) );
  AND2_X4 U12868 ( .A1(n11417), .A2(n11422), .ZN(n12150) );
  AOI22_X1 U12869 ( .A1(n11841), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U12870 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11426) );
  AND2_X2 U12871 ( .A1(n11420), .A2(n11421), .ZN(n11871) );
  AOI22_X1 U12872 ( .A1(n11871), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11503), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11425) );
  AND2_X2 U12873 ( .A1(n16085), .A2(n11422), .ZN(n11516) );
  NOR2_X1 U12874 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11423) );
  AND2_X2 U12875 ( .A1(n14269), .A2(n11423), .ZN(n11741) );
  AOI22_X1 U12876 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11424) );
  NAND2_X1 U12877 ( .A1(n11407), .A2(n11410), .ZN(n11573) );
  AOI22_X1 U12878 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U12879 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U12880 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11722), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U12881 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11503), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11429) );
  NAND4_X1 U12882 ( .A1(n11432), .A2(n11431), .A3(n11430), .A4(n11429), .ZN(
        n11438) );
  AOI22_X1 U12883 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U12884 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11871), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U12885 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U12886 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11433) );
  NAND4_X1 U12887 ( .A1(n11436), .A2(n11435), .A3(n11434), .A4(n11433), .ZN(
        n11437) );
  NAND2_X1 U12889 ( .A1(n11841), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11442) );
  NAND2_X1 U12890 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11441) );
  NAND2_X1 U12891 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11440) );
  NAND2_X1 U12892 ( .A1(n11722), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11439) );
  NAND2_X1 U12893 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11446) );
  NAND2_X1 U12894 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11445) );
  NAND2_X1 U12895 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11444) );
  NAND2_X1 U12896 ( .A1(n11503), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11443) );
  NAND2_X1 U12897 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11451) );
  NAND2_X1 U12898 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11450) );
  NAND2_X1 U12899 ( .A1(n12340), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11449) );
  NAND2_X1 U12900 ( .A1(n11447), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11448) );
  NAND2_X1 U12901 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11455) );
  NAND2_X1 U12902 ( .A1(n11871), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11454) );
  NAND2_X1 U12903 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11453) );
  NAND2_X1 U12904 ( .A1(n11741), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11452) );
  AOI22_X1 U12905 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U12906 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U12907 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11722), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U12908 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11503), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11461) );
  NAND4_X1 U12909 ( .A1(n11464), .A2(n11463), .A3(n11462), .A4(n11461), .ZN(
        n11470) );
  AOI22_X1 U12910 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U12911 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11871), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11467) );
  AOI22_X1 U12912 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U12913 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11465) );
  NAND4_X1 U12914 ( .A1(n11468), .A2(n11467), .A3(n11466), .A4(n11465), .ZN(
        n11469) );
  OR2_X4 U12915 ( .A1(n11470), .A2(n11469), .ZN(n11680) );
  AOI22_X1 U12916 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U12917 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U12918 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11722), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U12919 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11503), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U12920 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U12921 ( .A1(n11475), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U12922 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11871), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11476) );
  NAND2_X1 U12923 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11485) );
  NAND2_X1 U12924 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11484) );
  NAND2_X1 U12925 ( .A1(n11871), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11483) );
  NAND2_X1 U12926 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11482) );
  NAND2_X1 U12927 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11489) );
  NAND2_X1 U12928 ( .A1(n11447), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11488) );
  NAND2_X1 U12929 ( .A1(n11503), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11487) );
  NAND2_X1 U12930 ( .A1(n11741), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11486) );
  NAND2_X1 U12931 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11495) );
  NAND2_X1 U12932 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11494) );
  NAND2_X1 U12933 ( .A1(n11722), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11493) );
  NAND2_X1 U12934 ( .A1(n12340), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11492) );
  NAND2_X1 U12935 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11499) );
  NAND2_X1 U12936 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11498) );
  NAND2_X1 U12937 ( .A1(n11841), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11497) );
  NAND2_X1 U12938 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11496) );
  AND3_X4 U12939 ( .A1(n11502), .A2(n11501), .A3(n11500), .ZN(n11682) );
  NAND3_X1 U12940 ( .A1(n11700), .A2(n11709), .A3(n11682), .ZN(n12395) );
  NOR2_X2 U12941 ( .A1(n11012), .A2(n12395), .ZN(n15566) );
  AOI22_X1 U12942 ( .A1(n11460), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U12943 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U12944 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11722), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U12945 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11503), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11504) );
  NAND4_X1 U12946 ( .A1(n11507), .A2(n11506), .A3(n11505), .A4(n11504), .ZN(
        n11513) );
  AOI22_X1 U12947 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U12948 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11871), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U12949 ( .A1(n11515), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U12950 ( .A1(n11516), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11508) );
  NAND4_X1 U12951 ( .A1(n11511), .A2(n11510), .A3(n11509), .A4(n11508), .ZN(
        n11512) );
  NAND2_X1 U12953 ( .A1(n11686), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11749) );
  INV_X1 U12954 ( .A(n11941), .ZN(n11526) );
  NAND2_X1 U12955 ( .A1(n21892), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11544) );
  INV_X1 U12956 ( .A(n11544), .ZN(n11514) );
  AOI21_X1 U12957 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n13961), .A(
        n11514), .ZN(n11527) );
  INV_X1 U12958 ( .A(n11527), .ZN(n11525) );
  AOI22_X1 U12959 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11515), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U12960 ( .A1(n12366), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11871), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U12961 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11518) );
  AOI22_X1 U12962 ( .A1(n11722), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U12963 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U12964 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11741), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11522) );
  OAI21_X1 U12965 ( .B1(n11526), .B2(n11525), .A(n11568), .ZN(n11536) );
  INV_X1 U12966 ( .A(n11538), .ZN(n11530) );
  NAND2_X1 U12967 ( .A1(n11530), .A2(n14410), .ZN(n11533) );
  XNOR2_X1 U12968 ( .A(n11531), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11532) );
  XNOR2_X1 U12969 ( .A(n11532), .B(n11544), .ZN(n11580) );
  NAND3_X1 U12970 ( .A1(n11536), .A2(n11535), .A3(n11534), .ZN(n11542) );
  NAND3_X1 U12971 ( .A1(n11941), .A2(n11685), .A3(n11580), .ZN(n11541) );
  NOR2_X1 U12972 ( .A1(n11944), .A2(n11580), .ZN(n11539) );
  OAI22_X1 U12973 ( .A1(n11539), .A2(n11538), .B1(n11537), .B2(n11580), .ZN(
        n11540) );
  NAND3_X1 U12974 ( .A1(n11542), .A2(n11541), .A3(n11540), .ZN(n11550) );
  MUX2_X1 U12975 ( .A(n16851), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11551) );
  NAND2_X1 U12976 ( .A1(n21880), .A2(n11531), .ZN(n11543) );
  AOI22_X1 U12977 ( .A1(n11544), .A2(n11543), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n11718), .ZN(n11552) );
  XOR2_X1 U12978 ( .A(n11551), .B(n11552), .Z(n11578) );
  NAND2_X1 U12979 ( .A1(n11941), .A2(n11578), .ZN(n11545) );
  OAI211_X1 U12980 ( .C1(n11578), .C2(n11944), .A(n11546), .B(n11545), .ZN(
        n11549) );
  INV_X1 U12981 ( .A(n11545), .ZN(n11548) );
  INV_X1 U12982 ( .A(n11546), .ZN(n11547) );
  AOI22_X1 U12983 ( .A1(n11550), .A2(n11549), .B1(n11548), .B2(n11547), .ZN(
        n11563) );
  NAND2_X1 U12984 ( .A1(n11552), .A2(n11551), .ZN(n11554) );
  NAND2_X1 U12985 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n16851), .ZN(
        n11553) );
  NAND2_X1 U12986 ( .A1(n11554), .A2(n11553), .ZN(n11559) );
  NAND2_X1 U12987 ( .A1(n11559), .A2(n11555), .ZN(n11557) );
  INV_X1 U12988 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11834) );
  NAND2_X1 U12989 ( .A1(n11834), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11556) );
  NAND2_X1 U12990 ( .A1(n11557), .A2(n11556), .ZN(n11565) );
  INV_X1 U12991 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16815) );
  NAND2_X1 U12992 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16815), .ZN(
        n11566) );
  MUX2_X1 U12993 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n11834), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11558) );
  XNOR2_X1 U12994 ( .A(n11559), .B(n11558), .ZN(n11560) );
  OAI21_X1 U12995 ( .B1(n11565), .B2(n11566), .A(n11560), .ZN(n11561) );
  INV_X1 U12996 ( .A(n11561), .ZN(n11579) );
  NOR2_X1 U12997 ( .A1(n11853), .A2(n11579), .ZN(n11562) );
  OAI22_X1 U12998 ( .A1(n11563), .A2(n11562), .B1(n11579), .B2(n11568), .ZN(
        n11570) );
  AND2_X1 U12999 ( .A1(n21655), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11569) );
  INV_X1 U13000 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16888) );
  AND2_X1 U13001 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16888), .ZN(
        n11564) );
  INV_X1 U13002 ( .A(n11582), .ZN(n11571) );
  NAND2_X1 U13003 ( .A1(n14568), .A2(n11680), .ZN(n11572) );
  MUX2_X1 U13004 ( .A(n11572), .B(n12400), .S(n11709), .Z(n11575) );
  INV_X1 U13005 ( .A(n12777), .ZN(n14392) );
  OR2_X2 U13006 ( .A1(n11683), .A2(n14392), .ZN(n11711) );
  AOI21_X2 U13007 ( .B1(n11689), .B2(n14056), .A(n12394), .ZN(n11574) );
  NOR2_X2 U13008 ( .A1(n11697), .A2(n11576), .ZN(n11705) );
  NAND3_X1 U13009 ( .A1(n11580), .A2(n11579), .A3(n11578), .ZN(n11581) );
  AND2_X1 U13010 ( .A1(n11582), .A2(n11581), .ZN(n15571) );
  NAND2_X1 U13011 ( .A1(n11577), .A2(n15571), .ZN(n13822) );
  NAND2_X1 U13012 ( .A1(n16813), .A2(n21655), .ZN(n12768) );
  NOR2_X1 U13013 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11583) );
  NAND2_X1 U13014 ( .A1(n12378), .A2(n21655), .ZN(n16884) );
  NOR2_X1 U13015 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21659) );
  NAND2_X1 U13016 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21659), .ZN(n16882) );
  OAI22_X1 U13017 ( .A1(n16886), .A2(n16884), .B1(n21655), .B2(n16882), .ZN(
        n11584) );
  INV_X1 U13018 ( .A(n21483), .ZN(n14660) );
  INV_X2 U13019 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21922) );
  NAND2_X1 U13020 ( .A1(n11585), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n11586) );
  OR2_X1 U13021 ( .A1(n11699), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n21692) );
  NAND2_X1 U13022 ( .A1(n14410), .A2(n21692), .ZN(n14050) );
  NAND2_X1 U13023 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21683) );
  AND2_X1 U13024 ( .A1(n21683), .A2(n14439), .ZN(n11672) );
  NAND2_X1 U13025 ( .A1(n15652), .A2(n21493), .ZN(n21510) );
  INV_X1 U13026 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n19969) );
  INV_X1 U13027 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n19861) );
  INV_X1 U13028 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n19866) );
  NAND2_X1 U13029 ( .A1(n15236), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n21540) );
  INV_X1 U13030 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21539) );
  INV_X1 U13031 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n19870) );
  INV_X1 U13032 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21592) );
  NAND2_X1 U13033 ( .A1(n21588), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n21599) );
  INV_X1 U13034 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21600) );
  INV_X1 U13035 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n19877) );
  INV_X1 U13036 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n19884) );
  NAND2_X1 U13037 ( .A1(n15612), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15597) );
  INV_X1 U13038 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n19888) );
  INV_X1 U13039 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n15807) );
  INV_X1 U13040 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n19891) );
  OR2_X4 U13041 ( .A1(n12777), .A2(n11686), .ZN(n11656) );
  OR2_X1 U13042 ( .A1(n15578), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n11587) );
  OAI21_X1 U13043 ( .B1(n11696), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11587), .ZN(n15587) );
  INV_X4 U13044 ( .A(n11663), .ZN(n13950) );
  INV_X1 U13045 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14616) );
  NAND2_X1 U13046 ( .A1(n11653), .A2(n14616), .ZN(n11588) );
  NAND2_X1 U13047 ( .A1(n11589), .A2(n11588), .ZN(n11591) );
  INV_X1 U13048 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11590) );
  OAI22_X1 U13049 ( .A1(n11656), .A2(n11590), .B1(n13950), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13986) );
  XNOR2_X1 U13050 ( .A(n11591), .B(n13986), .ZN(n14173) );
  AOI21_X1 U13051 ( .B1(n14173), .B2(n11023), .A(n11591), .ZN(n14416) );
  MUX2_X1 U13052 ( .A(n11659), .B(n13950), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n11593) );
  INV_X1 U13053 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21300) );
  NAND2_X1 U13054 ( .A1(n11653), .A2(n21300), .ZN(n11592) );
  AND2_X1 U13055 ( .A1(n11593), .A2(n11592), .ZN(n14415) );
  INV_X1 U13056 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11594) );
  NAND2_X1 U13057 ( .A1(n11656), .A2(n11594), .ZN(n11595) );
  OAI211_X1 U13058 ( .C1(n15578), .C2(P1_EBX_REG_3__SCAN_IN), .A(n13950), .B(
        n11595), .ZN(n11596) );
  OAI21_X1 U13059 ( .B1(n11662), .B2(P1_EBX_REG_3__SCAN_IN), .A(n11596), .ZN(
        n14427) );
  NAND2_X1 U13060 ( .A1(n14428), .A2(n14427), .ZN(n14426) );
  MUX2_X1 U13061 ( .A(n11659), .B(n13950), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n11598) );
  INV_X1 U13062 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12812) );
  NAND2_X1 U13063 ( .A1(n11653), .A2(n12812), .ZN(n11597) );
  NAND2_X1 U13064 ( .A1(n11598), .A2(n11597), .ZN(n14649) );
  NAND2_X1 U13065 ( .A1(n13950), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11599) );
  NAND2_X1 U13066 ( .A1(n11656), .A2(n11599), .ZN(n11600) );
  OAI21_X1 U13067 ( .B1(n15578), .B2(P1_EBX_REG_5__SCAN_IN), .A(n11600), .ZN(
        n11601) );
  OAI21_X1 U13068 ( .B1(n11662), .B2(P1_EBX_REG_5__SCAN_IN), .A(n11601), .ZN(
        n14653) );
  MUX2_X1 U13069 ( .A(n11659), .B(n13950), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n11602) );
  NAND2_X1 U13070 ( .A1(n11602), .A2(n11392), .ZN(n14799) );
  MUX2_X1 U13071 ( .A(n11659), .B(n13950), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n11603) );
  AND2_X1 U13072 ( .A1(n11603), .A2(n11399), .ZN(n14751) );
  INV_X1 U13073 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21334) );
  NAND2_X1 U13074 ( .A1(n11656), .A2(n21334), .ZN(n11604) );
  OAI211_X1 U13075 ( .C1(n15578), .C2(P1_EBX_REG_7__SCAN_IN), .A(n13950), .B(
        n11604), .ZN(n11605) );
  OAI21_X1 U13076 ( .B1(n11662), .B2(P1_EBX_REG_7__SCAN_IN), .A(n11605), .ZN(
        n19939) );
  NAND2_X1 U13077 ( .A1(n14751), .A2(n19939), .ZN(n11606) );
  INV_X1 U13078 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n11607) );
  NAND2_X1 U13079 ( .A1(n11642), .A2(n11607), .ZN(n11610) );
  INV_X1 U13080 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15933) );
  NAND2_X1 U13081 ( .A1(n11656), .A2(n15933), .ZN(n11608) );
  OAI211_X1 U13082 ( .C1(n15578), .C2(P1_EBX_REG_9__SCAN_IN), .A(n13950), .B(
        n11608), .ZN(n11609) );
  MUX2_X1 U13083 ( .A(n11659), .B(n13950), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n11612) );
  INV_X1 U13084 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15932) );
  NAND2_X1 U13085 ( .A1(n11653), .A2(n15932), .ZN(n11611) );
  NAND2_X1 U13086 ( .A1(n11612), .A2(n11611), .ZN(n14943) );
  NOR2_X1 U13087 ( .A1(n14940), .A2(n14943), .ZN(n11613) );
  INV_X1 U13088 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n21506) );
  NAND2_X1 U13089 ( .A1(n11642), .A2(n21506), .ZN(n11617) );
  INV_X1 U13090 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11614) );
  NAND2_X1 U13091 ( .A1(n11656), .A2(n11614), .ZN(n11615) );
  OAI211_X1 U13092 ( .C1(n15578), .C2(P1_EBX_REG_11__SCAN_IN), .A(n13950), .B(
        n11615), .ZN(n11616) );
  NAND2_X1 U13093 ( .A1(n13950), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11618) );
  OAI211_X1 U13094 ( .C1(n15578), .C2(P1_EBX_REG_12__SCAN_IN), .A(n11656), .B(
        n11618), .ZN(n11619) );
  OAI21_X1 U13095 ( .B1(n11659), .B2(P1_EBX_REG_12__SCAN_IN), .A(n11619), .ZN(
        n19920) );
  INV_X1 U13096 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15656) );
  NAND2_X1 U13097 ( .A1(n11642), .A2(n15656), .ZN(n11622) );
  INV_X1 U13098 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21282) );
  NAND2_X1 U13099 ( .A1(n11656), .A2(n21282), .ZN(n11620) );
  OAI211_X1 U13100 ( .C1(n15578), .C2(P1_EBX_REG_13__SCAN_IN), .A(n10954), .B(
        n11620), .ZN(n11621) );
  INV_X1 U13101 ( .A(n11659), .ZN(n11646) );
  MUX2_X1 U13102 ( .A(n11646), .B(n11663), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n11624) );
  NOR2_X1 U13103 ( .A1(n11696), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11623) );
  NOR2_X1 U13104 ( .A1(n11624), .A2(n11623), .ZN(n15203) );
  INV_X1 U13105 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16058) );
  NAND2_X1 U13106 ( .A1(n11656), .A2(n16058), .ZN(n11625) );
  OAI211_X1 U13107 ( .C1(n15578), .C2(P1_EBX_REG_15__SCAN_IN), .A(n10954), .B(
        n11625), .ZN(n11626) );
  OAI21_X1 U13108 ( .B1(n11662), .B2(P1_EBX_REG_15__SCAN_IN), .A(n11626), .ZN(
        n15237) );
  MUX2_X1 U13109 ( .A(n11659), .B(n13950), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n11627) );
  OAI21_X1 U13110 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n11696), .A(
        n11627), .ZN(n15645) );
  INV_X1 U13111 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n21534) );
  NAND2_X1 U13112 ( .A1(n11642), .A2(n21534), .ZN(n11630) );
  INV_X1 U13113 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15896) );
  NAND2_X1 U13114 ( .A1(n11656), .A2(n15896), .ZN(n11628) );
  OAI211_X1 U13115 ( .C1(n15578), .C2(P1_EBX_REG_17__SCAN_IN), .A(n10954), .B(
        n11628), .ZN(n11629) );
  MUX2_X1 U13116 ( .A(n11659), .B(n13950), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n11631) );
  NAND2_X1 U13117 ( .A1(n11631), .A2(n11405), .ZN(n15714) );
  INV_X1 U13118 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15876) );
  NAND2_X1 U13119 ( .A1(n11656), .A2(n15876), .ZN(n11632) );
  OAI211_X1 U13120 ( .C1(n15578), .C2(P1_EBX_REG_19__SCAN_IN), .A(n13950), .B(
        n11632), .ZN(n11633) );
  OAI21_X1 U13121 ( .B1(n11662), .B2(P1_EBX_REG_19__SCAN_IN), .A(n11633), .ZN(
        n15706) );
  INV_X1 U13122 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n21565) );
  NAND2_X1 U13123 ( .A1(n11646), .A2(n21565), .ZN(n11636) );
  NAND2_X1 U13124 ( .A1(n13950), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11634) );
  OAI211_X1 U13125 ( .C1(n15578), .C2(P1_EBX_REG_20__SCAN_IN), .A(n11656), .B(
        n11634), .ZN(n11635) );
  AND2_X1 U13126 ( .A1(n11636), .A2(n11635), .ZN(n19934) );
  INV_X1 U13127 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12869) );
  NAND2_X1 U13128 ( .A1(n11656), .A2(n12869), .ZN(n11637) );
  OAI211_X1 U13129 ( .C1(n15578), .C2(P1_EBX_REG_21__SCAN_IN), .A(n10954), .B(
        n11637), .ZN(n11638) );
  OAI21_X1 U13130 ( .B1(n11662), .B2(P1_EBX_REG_21__SCAN_IN), .A(n11638), .ZN(
        n15696) );
  MUX2_X1 U13131 ( .A(n11659), .B(n13950), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11640) );
  INV_X1 U13132 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21406) );
  NAND2_X1 U13133 ( .A1(n11653), .A2(n21406), .ZN(n11639) );
  NAND2_X1 U13134 ( .A1(n11640), .A2(n11639), .ZN(n15691) );
  INV_X1 U13135 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n11641) );
  NAND2_X1 U13136 ( .A1(n11642), .A2(n11641), .ZN(n11645) );
  INV_X1 U13137 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15939) );
  NAND2_X1 U13138 ( .A1(n11656), .A2(n15939), .ZN(n11643) );
  OAI211_X1 U13139 ( .C1(n15578), .C2(P1_EBX_REG_23__SCAN_IN), .A(n10954), .B(
        n11643), .ZN(n11644) );
  AND2_X1 U13140 ( .A1(n11645), .A2(n11644), .ZN(n15678) );
  INV_X1 U13141 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n21611) );
  NAND2_X1 U13142 ( .A1(n11646), .A2(n21611), .ZN(n11649) );
  NAND2_X1 U13143 ( .A1(n13950), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11647) );
  OAI211_X1 U13144 ( .C1(n15578), .C2(P1_EBX_REG_24__SCAN_IN), .A(n11656), .B(
        n11647), .ZN(n11648) );
  AND2_X1 U13145 ( .A1(n11649), .A2(n11648), .ZN(n19928) );
  NAND2_X1 U13146 ( .A1(n13950), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11650) );
  NAND2_X1 U13147 ( .A1(n11656), .A2(n11650), .ZN(n11651) );
  OAI21_X1 U13148 ( .B1(n15578), .B2(P1_EBX_REG_25__SCAN_IN), .A(n11651), .ZN(
        n11652) );
  OAI21_X1 U13149 ( .B1(n11662), .B2(P1_EBX_REG_25__SCAN_IN), .A(n11652), .ZN(
        n15672) );
  MUX2_X1 U13150 ( .A(n11659), .B(n13950), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n11655) );
  INV_X1 U13151 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15998) );
  NAND2_X1 U13152 ( .A1(n11653), .A2(n15998), .ZN(n11654) );
  NAND2_X1 U13153 ( .A1(n11655), .A2(n11654), .ZN(n15632) );
  INV_X1 U13154 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15990) );
  NAND2_X1 U13155 ( .A1(n11656), .A2(n15990), .ZN(n11657) );
  OAI211_X1 U13156 ( .C1(n15578), .C2(P1_EBX_REG_27__SCAN_IN), .A(n10954), .B(
        n11657), .ZN(n11658) );
  OAI21_X1 U13157 ( .B1(n11662), .B2(P1_EBX_REG_27__SCAN_IN), .A(n11658), .ZN(
        n15607) );
  INV_X1 U13158 ( .A(n15607), .ZN(n15622) );
  MUX2_X1 U13159 ( .A(n11659), .B(n13950), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n11660) );
  OAI21_X1 U13160 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n11696), .A(
        n11660), .ZN(n15610) );
  OR2_X1 U13161 ( .A1(n15578), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n11661) );
  OAI21_X1 U13162 ( .B1(n11696), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11661), .ZN(n15585) );
  OAI22_X1 U13163 ( .A1(n15585), .A2(n11663), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n11662), .ZN(n15599) );
  NAND2_X1 U13164 ( .A1(n10978), .A2(n15599), .ZN(n15598) );
  NAND2_X1 U13165 ( .A1(n11696), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n11665) );
  NAND2_X1 U13166 ( .A1(n15578), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11664) );
  NAND2_X1 U13167 ( .A1(n11665), .A2(n11664), .ZN(n11667) );
  NAND2_X1 U13168 ( .A1(n11666), .A2(n11667), .ZN(n11671) );
  NOR2_X1 U13169 ( .A1(n15598), .A2(n15587), .ZN(n11669) );
  INV_X1 U13170 ( .A(n11667), .ZN(n11668) );
  NAND2_X1 U13171 ( .A1(n11669), .A2(n11668), .ZN(n11670) );
  NAND2_X1 U13172 ( .A1(n11685), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n11674) );
  NOR2_X1 U13173 ( .A1(n11674), .A2(n11672), .ZN(n11673) );
  NAND2_X1 U13174 ( .A1(n11045), .A2(n11674), .ZN(n11675) );
  AOI22_X1 U13175 ( .A1(n21615), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n21597), .ZN(n11677) );
  NAND2_X1 U13176 ( .A1(n21483), .A2(n21484), .ZN(n21627) );
  OR2_X1 U13177 ( .A1(n15590), .A2(n19891), .ZN(n11679) );
  INV_X1 U13178 ( .A(n15576), .ZN(n11681) );
  NAND2_X1 U13179 ( .A1(n12766), .A2(n11682), .ZN(n11687) );
  INV_X1 U13180 ( .A(n11687), .ZN(n11684) );
  NAND2_X1 U13181 ( .A1(n11684), .A2(n12758), .ZN(n13933) );
  NAND2_X1 U13182 ( .A1(n13933), .A2(n13956), .ZN(n11694) );
  NAND2_X1 U13183 ( .A1(n11688), .A2(n14056), .ZN(n13946) );
  NOR2_X2 U13184 ( .A1(n14056), .A2(n12777), .ZN(n14268) );
  NAND2_X1 U13185 ( .A1(n11686), .A2(n11685), .ZN(n14598) );
  NAND2_X1 U13186 ( .A1(n11697), .A2(n11686), .ZN(n11714) );
  AOI21_X1 U13187 ( .B1(n11704), .B2(n11703), .A(n14070), .ZN(n11706) );
  NAND2_X1 U13188 ( .A1(n11705), .A2(n14410), .ZN(n13954) );
  AND2_X2 U13189 ( .A1(n11706), .A2(n13954), .ZN(n11719) );
  NAND2_X2 U13190 ( .A1(n11707), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11785) );
  MUX2_X1 U13191 ( .A(n21649), .B(n12768), .S(n21892), .Z(n11708) );
  OAI21_X2 U13192 ( .B1(n11785), .B2(n13961), .A(n11708), .ZN(n11758) );
  INV_X1 U13193 ( .A(n11702), .ZN(n15579) );
  NAND2_X1 U13194 ( .A1(n14268), .A2(n14404), .ZN(n14074) );
  NAND4_X1 U13195 ( .A1(n14074), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n16813), 
        .A4(n14598), .ZN(n11710) );
  AOI21_X1 U13196 ( .B1(n13861), .B2(n11711), .A(n11710), .ZN(n11715) );
  NAND3_X1 U13197 ( .A1(n13933), .A2(n11685), .A3(n13956), .ZN(n11712) );
  NAND4_X1 U13198 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n11756) );
  XNOR2_X1 U13199 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21830) );
  OR2_X1 U13200 ( .A1(n21649), .A2(n21880), .ZN(n11780) );
  OAI21_X1 U13201 ( .B1(n12768), .B2(n21830), .A(n11780), .ZN(n11716) );
  INV_X1 U13202 ( .A(n11716), .ZN(n11717) );
  INV_X1 U13203 ( .A(n11719), .ZN(n11720) );
  NAND2_X1 U13204 ( .A1(n14382), .A2(n11721), .ZN(n14438) );
  INV_X1 U13205 ( .A(n11777), .ZN(n11769) );
  AOI22_X1 U13206 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U13207 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U13208 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U13209 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11723) );
  NAND4_X1 U13210 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(
        n11732) );
  AOI22_X1 U13211 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U13212 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U13213 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11728) );
  AOI22_X1 U13214 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11727) );
  NAND4_X1 U13215 ( .A1(n11730), .A2(n11729), .A3(n11728), .A4(n11727), .ZN(
        n11731) );
  NAND2_X1 U13216 ( .A1(n11769), .A2(n12789), .ZN(n11733) );
  INV_X1 U13217 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11734) );
  OR2_X1 U13218 ( .A1(n11944), .A2(n11734), .ZN(n11752) );
  INV_X1 U13219 ( .A(n12789), .ZN(n11748) );
  AOI22_X1 U13220 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U13221 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11739) );
  BUF_X1 U13222 ( .A(n11841), .Z(n11735) );
  AOI22_X1 U13223 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U13224 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11737) );
  NAND4_X1 U13225 ( .A1(n11740), .A2(n11739), .A3(n11738), .A4(n11737), .ZN(
        n11747) );
  AOI22_X1 U13226 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U13227 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11744) );
  AOI22_X1 U13228 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U13229 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11742) );
  NAND4_X1 U13230 ( .A1(n11745), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n11746) );
  OAI22_X1 U13231 ( .A1(n11749), .A2(n11748), .B1(n11777), .B2(n12846), .ZN(
        n11750) );
  INV_X1 U13232 ( .A(n11750), .ZN(n11751) );
  NAND2_X1 U13233 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  NAND2_X1 U13234 ( .A1(n11754), .A2(n11753), .ZN(n11755) );
  OR2_X2 U13235 ( .A1(n11754), .A2(n11753), .ZN(n11779) );
  INV_X1 U13236 ( .A(n11756), .ZN(n11757) );
  AOI22_X1 U13237 ( .A1(n12320), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U13238 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12321), .B1(
        n10971), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U13239 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n10977), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U13240 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11759) );
  NAND4_X1 U13241 ( .A1(n11762), .A2(n11761), .A3(n11760), .A4(n11759), .ZN(
        n11768) );
  AOI22_X1 U13242 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U13243 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U13244 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U13245 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11763) );
  NAND4_X1 U13246 ( .A1(n11766), .A2(n11765), .A3(n11764), .A4(n11763), .ZN(
        n11767) );
  XNOR2_X1 U13247 ( .A(n11778), .B(n12790), .ZN(n11770) );
  NAND2_X1 U13248 ( .A1(n11770), .A2(n11769), .ZN(n11771) );
  INV_X1 U13249 ( .A(n12790), .ZN(n11776) );
  INV_X1 U13250 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11773) );
  OR2_X1 U13251 ( .A1(n11944), .A2(n11773), .ZN(n11775) );
  AOI21_X1 U13252 ( .B1(n11682), .B2(n12846), .A(n21655), .ZN(n11774) );
  OAI211_X1 U13253 ( .C1(n11776), .C2(n11688), .A(n11775), .B(n11774), .ZN(
        n11821) );
  NOR2_X1 U13254 ( .A1(n11778), .A2(n11777), .ZN(n12842) );
  INV_X1 U13255 ( .A(n11780), .ZN(n11782) );
  INV_X1 U13256 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13979) );
  INV_X1 U13257 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16851) );
  NAND2_X1 U13258 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11786) );
  NAND2_X1 U13259 ( .A1(n16851), .A2(n11786), .ZN(n11788) );
  NAND2_X1 U13260 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21921) );
  INV_X1 U13261 ( .A(n21921), .ZN(n11787) );
  NAND2_X1 U13262 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11787), .ZN(
        n21919) );
  NAND2_X1 U13263 ( .A1(n11788), .A2(n21919), .ZN(n14766) );
  OAI22_X1 U13264 ( .A1(n12768), .A2(n14766), .B1(n21649), .B2(n16851), .ZN(
        n11789) );
  INV_X1 U13265 ( .A(n11789), .ZN(n11790) );
  NAND2_X2 U13266 ( .A1(n11793), .A2(n11792), .ZN(n14286) );
  AOI22_X1 U13267 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U13268 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U13269 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12340), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U13270 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11795) );
  NAND4_X1 U13271 ( .A1(n11798), .A2(n11797), .A3(n11796), .A4(n11795), .ZN(
        n11804) );
  AOI22_X1 U13272 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U13273 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U13274 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U13275 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11799) );
  NAND4_X1 U13276 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11803) );
  AOI22_X1 U13277 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11941), .B2(n12791), .ZN(n11805) );
  NAND2_X1 U13278 ( .A1(n12788), .A2(n12069), .ZN(n11811) );
  NAND2_X1 U13279 ( .A1(n12418), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11861) );
  XNOR2_X1 U13280 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21441) );
  AOI21_X1 U13281 ( .B1(n12378), .B2(n21441), .A(n12385), .ZN(n11808) );
  NAND2_X1 U13282 ( .A1(n12386), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11807) );
  OAI211_X1 U13283 ( .C1(n11861), .C2(n13979), .A(n11808), .B(n11807), .ZN(
        n11809) );
  INV_X1 U13284 ( .A(n11809), .ZN(n11810) );
  NAND2_X1 U13285 ( .A1(n11811), .A2(n11810), .ZN(n11812) );
  NAND2_X1 U13286 ( .A1(n12385), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11830) );
  NAND2_X1 U13287 ( .A1(n11812), .A2(n11830), .ZN(n14307) );
  INV_X1 U13288 ( .A(n11813), .ZN(n11814) );
  NAND2_X1 U13289 ( .A1(n11027), .A2(n11814), .ZN(n11815) );
  NAND2_X1 U13290 ( .A1(n11816), .A2(n11815), .ZN(n14298) );
  NAND2_X1 U13291 ( .A1(n14298), .A2(n12069), .ZN(n11820) );
  AOI22_X1 U13292 ( .A1(n12386), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21922), .ZN(n11818) );
  INV_X1 U13293 ( .A(n11861), .ZN(n11881) );
  NAND2_X1 U13294 ( .A1(n11881), .A2(n11531), .ZN(n11817) );
  AND2_X1 U13295 ( .A1(n11818), .A2(n11817), .ZN(n11819) );
  NAND2_X1 U13296 ( .A1(n11820), .A2(n11819), .ZN(n14175) );
  XNOR2_X2 U13297 ( .A(n11822), .B(n11821), .ZN(n12775) );
  NAND2_X1 U13298 ( .A1(n12775), .A2(n14404), .ZN(n11823) );
  NAND2_X1 U13299 ( .A1(n11823), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13992) );
  NAND2_X1 U13300 ( .A1(n21922), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11826) );
  NAND2_X1 U13301 ( .A1(n11824), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11825) );
  OAI211_X1 U13302 ( .C1(n11861), .C2(n13961), .A(n11826), .B(n11825), .ZN(
        n11827) );
  OR2_X1 U13303 ( .A1(n13992), .A2(n11828), .ZN(n13993) );
  OR2_X1 U13304 ( .A1(n11369), .A2(n12384), .ZN(n11829) );
  NAND2_X1 U13305 ( .A1(n13993), .A2(n11829), .ZN(n14174) );
  NAND2_X1 U13306 ( .A1(n14175), .A2(n14174), .ZN(n14308) );
  OAI21_X2 U13307 ( .B1(n14307), .B2(n14308), .A(n11830), .ZN(n14423) );
  INV_X1 U13308 ( .A(n11831), .ZN(n11833) );
  NAND2_X1 U13309 ( .A1(n11833), .A2(n11832), .ZN(n11865) );
  INV_X1 U13310 ( .A(n12768), .ZN(n11837) );
  INV_X1 U13311 ( .A(n21919), .ZN(n11835) );
  NAND2_X1 U13312 ( .A1(n11835), .A2(n11834), .ZN(n14572) );
  NAND2_X1 U13313 ( .A1(n21919), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11836) );
  NAND2_X1 U13314 ( .A1(n14572), .A2(n11836), .ZN(n21831) );
  INV_X1 U13315 ( .A(n21649), .ZN(n16876) );
  AOI22_X1 U13316 ( .A1(n11837), .A2(n21831), .B1(n16876), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11838) );
  XNOR2_X2 U13317 ( .A(n14286), .B(n14381), .ZN(n21829) );
  AOI22_X1 U13318 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U13319 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U13320 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U13321 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11842) );
  NAND4_X1 U13322 ( .A1(n11845), .A2(n11844), .A3(n11843), .A4(n11842), .ZN(
        n11852) );
  AOI22_X1 U13323 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11850) );
  BUF_X1 U13324 ( .A(n11846), .Z(n12321) );
  AOI22_X1 U13325 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U13326 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U13327 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11847) );
  NAND4_X1 U13328 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11851) );
  AOI22_X1 U13329 ( .A1(n11853), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11941), .B2(n12803), .ZN(n11854) );
  NAND2_X2 U13330 ( .A1(n11855), .A2(n11854), .ZN(n14368) );
  NAND2_X1 U13331 ( .A1(n12799), .A2(n12069), .ZN(n11864) );
  NAND2_X1 U13332 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11856) );
  INV_X1 U13333 ( .A(n11856), .ZN(n11858) );
  INV_X1 U13334 ( .A(n11908), .ZN(n11857) );
  OAI21_X1 U13335 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11858), .A(
        n11857), .ZN(n14624) );
  AOI22_X1 U13336 ( .A1(n12378), .A2(n14624), .B1(n12385), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11860) );
  NAND2_X1 U13337 ( .A1(n12386), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11859) );
  OAI211_X1 U13338 ( .C1(n11861), .C2(n11376), .A(n11860), .B(n11859), .ZN(
        n11862) );
  INV_X1 U13339 ( .A(n11862), .ZN(n11863) );
  NAND2_X1 U13340 ( .A1(n14423), .A2(n14425), .ZN(n14424) );
  INV_X1 U13341 ( .A(n11865), .ZN(n11889) );
  NAND2_X1 U13342 ( .A1(n11889), .A2(n14368), .ZN(n11880) );
  INV_X1 U13343 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11866) );
  OR2_X1 U13344 ( .A1(n11944), .A2(n11866), .ZN(n11879) );
  AOI22_X1 U13345 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U13346 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U13347 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U13348 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11867) );
  NAND4_X1 U13349 ( .A1(n11870), .A2(n11869), .A3(n11868), .A4(n11867), .ZN(
        n11877) );
  AOI22_X1 U13350 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U13352 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U13353 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U13354 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11872) );
  NAND4_X1 U13355 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11876) );
  NAND2_X1 U13356 ( .A1(n11941), .A2(n12815), .ZN(n11878) );
  NAND2_X1 U13357 ( .A1(n11879), .A2(n11878), .ZN(n11888) );
  NAND2_X1 U13358 ( .A1(n11881), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11886) );
  INV_X1 U13359 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11882) );
  AOI21_X1 U13360 ( .B1(n11882), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11883) );
  AOI21_X1 U13361 ( .B1(n12386), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11883), .ZN(
        n11885) );
  XNOR2_X1 U13362 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B(n11908), .ZN(
        n21466) );
  INV_X1 U13363 ( .A(n21466), .ZN(n11884) );
  AOI22_X1 U13364 ( .A1(n11886), .A2(n11885), .B1(n12378), .B2(n11884), .ZN(
        n11887) );
  NOR2_X2 U13365 ( .A1(n14424), .A2(n14647), .ZN(n14656) );
  INV_X1 U13366 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11890) );
  OR2_X1 U13367 ( .A1(n11944), .A2(n11890), .ZN(n11902) );
  AOI22_X1 U13368 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U13369 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U13370 ( .A1(n12268), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U13371 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11891) );
  NAND4_X1 U13372 ( .A1(n11894), .A2(n11893), .A3(n11892), .A4(n11891), .ZN(
        n11900) );
  AOI22_X1 U13373 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U13374 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U13375 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12340), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U13376 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11895) );
  NAND4_X1 U13377 ( .A1(n11898), .A2(n11897), .A3(n11896), .A4(n11895), .ZN(
        n11899) );
  NAND2_X1 U13378 ( .A1(n11941), .A2(n12826), .ZN(n11901) );
  NAND2_X1 U13379 ( .A1(n11906), .A2(n11905), .ZN(n11907) );
  NAND2_X1 U13380 ( .A1(n11938), .A2(n11907), .ZN(n12820) );
  INV_X1 U13381 ( .A(n11928), .ZN(n11930) );
  INV_X1 U13382 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11910) );
  NAND2_X1 U13383 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11908), .ZN(
        n11909) );
  NAND2_X1 U13384 ( .A1(n11910), .A2(n11909), .ZN(n11911) );
  NAND2_X1 U13385 ( .A1(n11930), .A2(n11911), .ZN(n21478) );
  AOI22_X1 U13386 ( .A1(n21478), .A2(n12378), .B1(n12385), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11912) );
  INV_X1 U13387 ( .A(n11912), .ZN(n11913) );
  INV_X1 U13388 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11915) );
  OR2_X1 U13389 ( .A1(n11944), .A2(n11915), .ZN(n11927) );
  AOI22_X1 U13390 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U13391 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U13392 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11917) );
  AOI22_X1 U13393 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11916) );
  NAND4_X1 U13394 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11925) );
  AOI22_X1 U13395 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U13396 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11922) );
  AOI22_X1 U13397 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11921) );
  AOI22_X1 U13398 ( .A1(n12340), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11920) );
  NAND4_X1 U13399 ( .A1(n11923), .A2(n11922), .A3(n11921), .A4(n11920), .ZN(
        n11924) );
  NAND2_X1 U13400 ( .A1(n11941), .A2(n12835), .ZN(n11926) );
  NAND2_X1 U13401 ( .A1(n12824), .A2(n12069), .ZN(n11937) );
  INV_X1 U13402 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11934) );
  INV_X1 U13403 ( .A(n11946), .ZN(n11932) );
  INV_X1 U13404 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11929) );
  NAND2_X1 U13405 ( .A1(n11930), .A2(n11929), .ZN(n11931) );
  NAND2_X1 U13406 ( .A1(n11932), .A2(n11931), .ZN(n21492) );
  AOI22_X1 U13407 ( .A1(n21492), .A2(n12378), .B1(n12385), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11933) );
  OAI21_X1 U13408 ( .B1(n12330), .B2(n11934), .A(n11933), .ZN(n11935) );
  NAND3_X1 U13409 ( .A1(n14656), .A2(n14657), .A3(n14800), .ZN(n14698) );
  INV_X1 U13410 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11943) );
  NAND2_X1 U13411 ( .A1(n11941), .A2(n12846), .ZN(n11942) );
  OAI21_X1 U13412 ( .B1(n11944), .B2(n11943), .A(n11942), .ZN(n11945) );
  INV_X1 U13413 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11948) );
  OAI21_X1 U13414 ( .B1(n11946), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n11966), .ZN(n21505) );
  AOI22_X1 U13415 ( .A1(n21505), .A2(n12378), .B1(n12385), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11947) );
  OAI21_X1 U13416 ( .B1(n12330), .B2(n11948), .A(n11947), .ZN(n11949) );
  AOI21_X1 U13417 ( .B1(n12833), .B2(n12069), .A(n11949), .ZN(n14697) );
  INV_X1 U13418 ( .A(n14697), .ZN(n11950) );
  AOI22_X1 U13419 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U13420 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n10977), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U13421 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U13422 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n12150), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11952) );
  NAND4_X1 U13423 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(
        n11961) );
  AOI22_X1 U13424 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U13425 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n11736), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U13426 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n10971), .B1(
        n12340), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U13427 ( .A1(n12320), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11956) );
  NAND4_X1 U13428 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11960) );
  OAI21_X1 U13429 ( .B1(n11961), .B2(n11960), .A(n12069), .ZN(n11965) );
  NAND2_X1 U13430 ( .A1(n12386), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11964) );
  INV_X1 U13431 ( .A(n11966), .ZN(n11962) );
  XNOR2_X1 U13432 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11962), .ZN(
        n15090) );
  AOI22_X1 U13433 ( .A1(n12378), .A2(n15090), .B1(n12385), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11963) );
  XOR2_X1 U13434 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11992), .Z(n15228) );
  INV_X1 U13435 ( .A(n15228), .ZN(n14813) );
  AOI22_X1 U13436 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U13437 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12340), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11969) );
  AOI22_X1 U13438 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U13439 ( .A1(n12320), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11967) );
  NAND4_X1 U13440 ( .A1(n11970), .A2(n11969), .A3(n11968), .A4(n11967), .ZN(
        n11976) );
  AOI22_X1 U13441 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U13442 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U13443 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U13444 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11971) );
  NAND4_X1 U13445 ( .A1(n11974), .A2(n11973), .A3(n11972), .A4(n11971), .ZN(
        n11975) );
  OAI21_X1 U13446 ( .B1(n11976), .B2(n11975), .A(n12069), .ZN(n11979) );
  NAND2_X1 U13447 ( .A1(n12386), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11978) );
  NAND2_X1 U13448 ( .A1(n12385), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11977) );
  NAND3_X1 U13449 ( .A1(n11979), .A2(n11978), .A3(n11977), .ZN(n11980) );
  AOI21_X1 U13450 ( .B1(n14813), .B2(n11583), .A(n11980), .ZN(n14810) );
  AOI22_X1 U13451 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11871), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U13452 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U13453 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U13454 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11982) );
  NAND4_X1 U13455 ( .A1(n11985), .A2(n11984), .A3(n11983), .A4(n11982), .ZN(
        n11991) );
  AOI22_X1 U13456 ( .A1(n11841), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U13457 ( .A1(n12340), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U13458 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U13459 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11986) );
  NAND4_X1 U13460 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n11990) );
  NOR2_X1 U13461 ( .A1(n11991), .A2(n11990), .ZN(n11995) );
  XNOR2_X1 U13462 ( .A(n11997), .B(n11996), .ZN(n15926) );
  NAND2_X1 U13463 ( .A1(n15926), .A2(n11583), .ZN(n11994) );
  AOI22_X1 U13464 ( .A1(n12386), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12385), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11993) );
  OAI211_X1 U13465 ( .C1(n11995), .C2(n11371), .A(n11994), .B(n11993), .ZN(
        n14936) );
  NAND2_X1 U13466 ( .A1(n14808), .A2(n14936), .ZN(n14935) );
  OR2_X1 U13467 ( .A1(n11998), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11999) );
  NAND2_X1 U13468 ( .A1(n11999), .A2(n12038), .ZN(n21515) );
  INV_X1 U13469 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15168) );
  INV_X1 U13470 ( .A(n12385), .ZN(n12106) );
  INV_X1 U13471 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12000) );
  OAI22_X1 U13472 ( .A1(n12330), .A2(n15168), .B1(n12106), .B2(n12000), .ZN(
        n12001) );
  AOI21_X1 U13473 ( .B1(n21515), .B2(n11583), .A(n12001), .ZN(n15161) );
  AOI22_X1 U13474 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U13475 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U13476 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U13477 ( .A1(n12320), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12002) );
  NAND4_X1 U13478 ( .A1(n12005), .A2(n12004), .A3(n12003), .A4(n12002), .ZN(
        n12011) );
  AOI22_X1 U13479 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U13480 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U13481 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12007) );
  AOI22_X1 U13482 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12006) );
  NAND4_X1 U13483 ( .A1(n12009), .A2(n12008), .A3(n12007), .A4(n12006), .ZN(
        n12010) );
  OR2_X1 U13484 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  NAND2_X1 U13485 ( .A1(n12069), .A2(n12012), .ZN(n15169) );
  AOI22_X1 U13486 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U13487 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U13488 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U13489 ( .A1(n12320), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12014) );
  NAND4_X1 U13490 ( .A1(n12017), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12023) );
  AOI22_X1 U13491 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U13492 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U13493 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U13494 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12018) );
  NAND4_X1 U13495 ( .A1(n12021), .A2(n12020), .A3(n12019), .A4(n12018), .ZN(
        n12022) );
  NOR2_X1 U13496 ( .A1(n12023), .A2(n12022), .ZN(n12027) );
  INV_X1 U13497 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12024) );
  XNOR2_X1 U13498 ( .A(n12044), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15917) );
  NAND2_X1 U13499 ( .A1(n15917), .A2(n11583), .ZN(n12026) );
  AOI22_X1 U13500 ( .A1(n12386), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n12385), 
        .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12025) );
  OAI211_X1 U13501 ( .C1(n12027), .C2(n11371), .A(n12026), .B(n12025), .ZN(
        n15216) );
  AOI22_X1 U13502 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U13503 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U13504 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U13505 ( .A1(n11447), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12028) );
  NAND4_X1 U13506 ( .A1(n12031), .A2(n12030), .A3(n12029), .A4(n12028), .ZN(
        n12037) );
  AOI22_X1 U13507 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U13508 ( .A1(n12320), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U13509 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U13510 ( .A1(n12340), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11516), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12032) );
  NAND4_X1 U13511 ( .A1(n12035), .A2(n12034), .A3(n12033), .A4(n12032), .ZN(
        n12036) );
  NOR2_X1 U13512 ( .A1(n12037), .A2(n12036), .ZN(n12042) );
  XNOR2_X1 U13513 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12038), .ZN(
        n21521) );
  INV_X1 U13514 ( .A(n21521), .ZN(n12039) );
  AOI22_X1 U13515 ( .A1(n12039), .A2(n11583), .B1(n12385), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12041) );
  NAND2_X1 U13516 ( .A1(n12386), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12040) );
  OAI211_X1 U13517 ( .C1(n11371), .C2(n12042), .A(n12041), .B(n12040), .ZN(
        n15171) );
  NAND2_X1 U13518 ( .A1(n15216), .A2(n15171), .ZN(n12043) );
  XOR2_X1 U13519 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n12059), .Z(
        n21527) );
  AOI22_X1 U13520 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U13521 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U13522 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U13523 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12045) );
  NAND4_X1 U13524 ( .A1(n12048), .A2(n12047), .A3(n12046), .A4(n12045), .ZN(
        n12055) );
  AOI22_X1 U13525 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U13526 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U13527 ( .A1(n11871), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U13528 ( .A1(n12340), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12050) );
  NAND4_X1 U13529 ( .A1(n12053), .A2(n12052), .A3(n12051), .A4(n12050), .ZN(
        n12054) );
  OR2_X1 U13530 ( .A1(n12055), .A2(n12054), .ZN(n12056) );
  AOI22_X1 U13531 ( .A1(n12069), .A2(n12056), .B1(n12385), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12058) );
  NAND2_X1 U13532 ( .A1(n12386), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12057) );
  OAI211_X1 U13533 ( .C1(n21527), .C2(n12384), .A(n12058), .B(n12057), .ZN(
        n15201) );
  INV_X1 U13534 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12060) );
  XNOR2_X1 U13535 ( .A(n12078), .B(n12060), .ZN(n15905) );
  AOI22_X1 U13536 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U13537 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U13538 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U13539 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12061) );
  NAND4_X1 U13540 ( .A1(n12064), .A2(n12063), .A3(n12062), .A4(n12061), .ZN(
        n12071) );
  AOI22_X1 U13541 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U13542 ( .A1(n12340), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U13543 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U13544 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12065) );
  NAND4_X1 U13545 ( .A1(n12068), .A2(n12067), .A3(n12066), .A4(n12065), .ZN(
        n12070) );
  OAI21_X1 U13546 ( .B1(n12071), .B2(n12070), .A(n12069), .ZN(n12074) );
  NAND2_X1 U13547 ( .A1(n12386), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12073) );
  NAND2_X1 U13548 ( .A1(n12385), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12072) );
  NAND3_X1 U13549 ( .A1(n12074), .A2(n12073), .A3(n12072), .ZN(n12075) );
  AOI21_X1 U13550 ( .B1(n15905), .B2(n12378), .A(n12075), .ZN(n15234) );
  OR2_X1 U13551 ( .A1(n12079), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12080) );
  NAND2_X1 U13552 ( .A1(n12080), .A2(n12124), .ZN(n20000) );
  AOI22_X1 U13553 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n10971), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U13554 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U13555 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n10977), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U13556 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12081) );
  NAND4_X1 U13557 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12090) );
  AOI22_X1 U13558 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n11736), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U13559 ( .A1(n11871), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U13560 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U13561 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12085) );
  NAND4_X1 U13562 ( .A1(n12088), .A2(n12087), .A3(n12086), .A4(n12085), .ZN(
        n12089) );
  NOR2_X1 U13563 ( .A1(n12090), .A2(n12089), .ZN(n12091) );
  NOR2_X1 U13564 ( .A1(n12381), .A2(n12091), .ZN(n12094) );
  INV_X1 U13565 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15785) );
  NAND2_X1 U13566 ( .A1(n21922), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12092) );
  OAI211_X1 U13567 ( .C1(n12330), .C2(n15785), .A(n12384), .B(n12092), .ZN(
        n12093) );
  OAI22_X1 U13568 ( .A1(n20000), .A2(n12384), .B1(n12094), .B2(n12093), .ZN(
        n15642) );
  AOI22_X1 U13569 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10977), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U13570 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U13571 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U13572 ( .A1(n12320), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U13573 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12104) );
  AOI22_X1 U13574 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U13575 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U13576 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U13577 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12099) );
  NAND4_X1 U13578 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12103) );
  OR2_X1 U13579 ( .A1(n12104), .A2(n12103), .ZN(n12105) );
  NAND2_X1 U13580 ( .A1(n12353), .A2(n12105), .ZN(n12109) );
  XNOR2_X1 U13581 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12124), .ZN(
        n21537) );
  OAI22_X1 U13582 ( .A1(n12384), .A2(n21537), .B1(n12106), .B2(n21535), .ZN(
        n12107) );
  AOI21_X1 U13583 ( .B1(n12386), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12107), .ZN(
        n12108) );
  NAND2_X1 U13584 ( .A1(n12109), .A2(n12108), .ZN(n15716) );
  AOI22_X1 U13585 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U13586 ( .A1(n11841), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U13587 ( .A1(n11871), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U13588 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12110) );
  NAND4_X1 U13589 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12119) );
  AOI22_X1 U13590 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U13591 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U13592 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U13593 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12114) );
  NAND4_X1 U13594 ( .A1(n12117), .A2(n12116), .A3(n12115), .A4(n12114), .ZN(
        n12118) );
  NOR2_X1 U13595 ( .A1(n12119), .A2(n12118), .ZN(n12123) );
  OAI21_X1 U13596 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n14439), .A(
        n21922), .ZN(n12120) );
  INV_X1 U13597 ( .A(n12120), .ZN(n12121) );
  AOI21_X1 U13598 ( .B1(n12386), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12121), .ZN(
        n12122) );
  OAI21_X1 U13599 ( .B1(n12381), .B2(n12123), .A(n12122), .ZN(n12127) );
  INV_X1 U13600 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n21535) );
  OAI21_X1 U13601 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12125), .A(
        n12147), .ZN(n15884) );
  INV_X1 U13602 ( .A(n15884), .ZN(n21546) );
  NAND2_X1 U13603 ( .A1(n21546), .A2(n11583), .ZN(n12126) );
  AOI22_X1 U13604 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U13605 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U13606 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U13607 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12128) );
  NAND4_X1 U13608 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12137) );
  AOI22_X1 U13609 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U13610 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U13611 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U13612 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12132) );
  NAND4_X1 U13613 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12136) );
  NOR2_X1 U13614 ( .A1(n12137), .A2(n12136), .ZN(n12141) );
  NAND2_X1 U13615 ( .A1(n21922), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12138) );
  NAND2_X1 U13616 ( .A1(n12384), .A2(n12138), .ZN(n12139) );
  AOI21_X1 U13617 ( .B1(n12386), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12139), .ZN(
        n12140) );
  OAI21_X1 U13618 ( .B1(n12381), .B2(n12141), .A(n12140), .ZN(n12145) );
  INV_X1 U13619 ( .A(n12147), .ZN(n12142) );
  XNOR2_X1 U13620 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12142), .ZN(
        n21564) );
  INV_X1 U13621 ( .A(n21564), .ZN(n12143) );
  NAND2_X1 U13622 ( .A1(n12143), .A2(n11583), .ZN(n12144) );
  INV_X1 U13623 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12146) );
  OR2_X1 U13624 ( .A1(n12148), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12149) );
  NAND2_X1 U13625 ( .A1(n12149), .A2(n12196), .ZN(n21566) );
  AOI22_X1 U13626 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U13627 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U13628 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U13629 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12151) );
  NAND4_X1 U13630 ( .A1(n12154), .A2(n12153), .A3(n12152), .A4(n12151), .ZN(
        n12160) );
  AOI22_X1 U13631 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U13632 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U13633 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U13634 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12155) );
  NAND4_X1 U13635 ( .A1(n12158), .A2(n12157), .A3(n12156), .A4(n12155), .ZN(
        n12159) );
  NOR2_X1 U13636 ( .A1(n12160), .A2(n12159), .ZN(n12163) );
  OAI21_X1 U13637 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n14439), .A(
        n21922), .ZN(n12162) );
  NAND2_X1 U13638 ( .A1(n12386), .A2(P1_EAX_REG_20__SCAN_IN), .ZN(n12161) );
  OAI211_X1 U13639 ( .C1(n12381), .C2(n12163), .A(n12162), .B(n12161), .ZN(
        n12164) );
  OAI21_X1 U13640 ( .B1(n21566), .B2(n12384), .A(n12164), .ZN(n15765) );
  INV_X1 U13641 ( .A(n15765), .ZN(n12165) );
  NAND2_X1 U13642 ( .A1(n15702), .A2(n12165), .ZN(n15693) );
  AOI22_X1 U13643 ( .A1(n11871), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U13644 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U13645 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U13646 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12166) );
  NAND4_X1 U13647 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n12175) );
  AOI22_X1 U13648 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U13649 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U13650 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U13651 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12170) );
  NAND4_X1 U13652 ( .A1(n12173), .A2(n12172), .A3(n12171), .A4(n12170), .ZN(
        n12174) );
  NOR2_X1 U13653 ( .A1(n12175), .A2(n12174), .ZN(n12179) );
  NAND2_X1 U13654 ( .A1(n21922), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12176) );
  NAND2_X1 U13655 ( .A1(n12384), .A2(n12176), .ZN(n12177) );
  AOI21_X1 U13656 ( .B1(n12386), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12177), .ZN(
        n12178) );
  OAI21_X1 U13657 ( .B1(n12381), .B2(n12179), .A(n12178), .ZN(n12181) );
  XNOR2_X1 U13658 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12196), .ZN(
        n21580) );
  NAND2_X1 U13659 ( .A1(n12378), .A2(n21580), .ZN(n12180) );
  NAND2_X1 U13660 ( .A1(n12181), .A2(n12180), .ZN(n15695) );
  NOR2_X2 U13661 ( .A1(n15693), .A2(n15695), .ZN(n15684) );
  AOI22_X1 U13662 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10971), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U13663 ( .A1(n11871), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U13664 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U13665 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12182) );
  NAND4_X1 U13666 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        n12191) );
  AOI22_X1 U13667 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U13668 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U13669 ( .A1(n12340), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U13670 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12186) );
  NAND4_X1 U13671 ( .A1(n12189), .A2(n12188), .A3(n12187), .A4(n12186), .ZN(
        n12190) );
  NOR2_X1 U13672 ( .A1(n12191), .A2(n12190), .ZN(n12195) );
  NAND2_X1 U13673 ( .A1(n21922), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12192) );
  NAND2_X1 U13674 ( .A1(n12384), .A2(n12192), .ZN(n12193) );
  AOI21_X1 U13675 ( .B1(n12386), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12193), .ZN(
        n12194) );
  OAI21_X1 U13676 ( .B1(n12381), .B2(n12195), .A(n12194), .ZN(n12199) );
  INV_X1 U13677 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21577) );
  OAI21_X1 U13678 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12197), .A(
        n12227), .ZN(n20013) );
  INV_X1 U13679 ( .A(n20013), .ZN(n21586) );
  NAND2_X1 U13680 ( .A1(n21586), .A2(n11583), .ZN(n12198) );
  NAND2_X1 U13681 ( .A1(n15684), .A2(n15683), .ZN(n15674) );
  AOI22_X1 U13682 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n10977), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U13683 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12360), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U13684 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U13685 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12200) );
  NAND4_X1 U13686 ( .A1(n12203), .A2(n12202), .A3(n12201), .A4(n12200), .ZN(
        n12209) );
  AOI22_X1 U13687 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n11735), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U13688 ( .A1(n12320), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U13689 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U13690 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12204) );
  NAND4_X1 U13691 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n12204), .ZN(
        n12208) );
  NOR2_X1 U13692 ( .A1(n12209), .A2(n12208), .ZN(n12231) );
  AOI22_X1 U13693 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10971), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U13694 ( .A1(n11735), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11736), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U13695 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U13696 ( .A1(n12320), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12210) );
  NAND4_X1 U13697 ( .A1(n12213), .A2(n12212), .A3(n12211), .A4(n12210), .ZN(
        n12219) );
  AOI22_X1 U13698 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U13699 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U13700 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U13701 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12214) );
  NAND4_X1 U13702 ( .A1(n12217), .A2(n12216), .A3(n12215), .A4(n12214), .ZN(
        n12218) );
  NOR2_X1 U13703 ( .A1(n12219), .A2(n12218), .ZN(n12230) );
  XOR2_X1 U13704 ( .A(n12231), .B(n12230), .Z(n12220) );
  NAND2_X1 U13705 ( .A1(n12220), .A2(n12353), .ZN(n12224) );
  NAND2_X1 U13706 ( .A1(n21922), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12221) );
  NAND2_X1 U13707 ( .A1(n12384), .A2(n12221), .ZN(n12222) );
  AOI21_X1 U13708 ( .B1(n12386), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12222), .ZN(
        n12223) );
  NAND2_X1 U13709 ( .A1(n12224), .A2(n12223), .ZN(n12226) );
  XNOR2_X1 U13710 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12227), .ZN(
        n21598) );
  NAND2_X1 U13711 ( .A1(n12378), .A2(n21598), .ZN(n12225) );
  NAND2_X1 U13712 ( .A1(n12226), .A2(n12225), .ZN(n15675) );
  NOR2_X2 U13713 ( .A1(n15674), .A2(n15675), .ZN(n15676) );
  INV_X1 U13714 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21609) );
  OR2_X1 U13715 ( .A1(n12228), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12229) );
  NAND2_X1 U13716 ( .A1(n12229), .A2(n12283), .ZN(n21612) );
  NOR2_X1 U13717 ( .A1(n12231), .A2(n12230), .ZN(n12259) );
  AOI22_X1 U13718 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U13719 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U13720 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U13721 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12232) );
  NAND4_X1 U13722 ( .A1(n12235), .A2(n12234), .A3(n12233), .A4(n12232), .ZN(
        n12241) );
  AOI22_X1 U13723 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U13724 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U13725 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U13726 ( .A1(n12340), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12236) );
  NAND4_X1 U13727 ( .A1(n12239), .A2(n12238), .A3(n12237), .A4(n12236), .ZN(
        n12240) );
  OR2_X1 U13728 ( .A1(n12241), .A2(n12240), .ZN(n12258) );
  XNOR2_X1 U13729 ( .A(n12259), .B(n12258), .ZN(n12245) );
  NAND2_X1 U13730 ( .A1(n21922), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12242) );
  NAND2_X1 U13731 ( .A1(n12384), .A2(n12242), .ZN(n12243) );
  AOI21_X1 U13732 ( .B1(n12386), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12243), .ZN(
        n12244) );
  OAI21_X1 U13733 ( .B1(n12245), .B2(n12381), .A(n12244), .ZN(n12246) );
  OAI21_X1 U13734 ( .B1(n21612), .B2(n12384), .A(n12246), .ZN(n15746) );
  AOI22_X1 U13735 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U13736 ( .A1(n12320), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U13737 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U13738 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12248) );
  NAND4_X1 U13739 ( .A1(n12251), .A2(n12250), .A3(n12249), .A4(n12248), .ZN(
        n12257) );
  AOI22_X1 U13740 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U13741 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U13742 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12340), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U13743 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12252) );
  NAND4_X1 U13744 ( .A1(n12255), .A2(n12254), .A3(n12253), .A4(n12252), .ZN(
        n12256) );
  NOR2_X1 U13745 ( .A1(n12257), .A2(n12256), .ZN(n12267) );
  NAND2_X1 U13746 ( .A1(n12259), .A2(n12258), .ZN(n12266) );
  XOR2_X1 U13747 ( .A(n12267), .B(n12266), .Z(n12260) );
  NAND2_X1 U13748 ( .A1(n12260), .A2(n12353), .ZN(n12265) );
  NAND2_X1 U13749 ( .A1(n21922), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12261) );
  NAND2_X1 U13750 ( .A1(n12384), .A2(n12261), .ZN(n12262) );
  AOI21_X1 U13751 ( .B1(n12386), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12262), .ZN(
        n12264) );
  XNOR2_X1 U13752 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n12283), .ZN(
        n21635) );
  AOI21_X1 U13753 ( .B1(n12265), .B2(n12264), .A(n12263), .ZN(n15670) );
  NOR2_X1 U13754 ( .A1(n12267), .A2(n12266), .ZN(n12304) );
  AOI22_X1 U13755 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U13756 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U13757 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U13758 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12269) );
  NAND4_X1 U13759 ( .A1(n12272), .A2(n12271), .A3(n12270), .A4(n12269), .ZN(
        n12278) );
  AOI22_X1 U13760 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U13761 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U13762 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U13763 ( .A1(n12365), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12273) );
  NAND4_X1 U13764 ( .A1(n12276), .A2(n12275), .A3(n12274), .A4(n12273), .ZN(
        n12277) );
  OR2_X1 U13765 ( .A1(n12278), .A2(n12277), .ZN(n12303) );
  INV_X1 U13766 ( .A(n12303), .ZN(n12279) );
  XNOR2_X1 U13767 ( .A(n12304), .B(n12279), .ZN(n12280) );
  NAND2_X1 U13768 ( .A1(n12280), .A2(n12353), .ZN(n12291) );
  NAND2_X1 U13769 ( .A1(n21922), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12281) );
  NAND2_X1 U13770 ( .A1(n12384), .A2(n12281), .ZN(n12282) );
  AOI21_X1 U13771 ( .B1(n12386), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12282), .ZN(
        n12290) );
  INV_X1 U13772 ( .A(n12283), .ZN(n12284) );
  INV_X1 U13773 ( .A(n12285), .ZN(n12287) );
  INV_X1 U13774 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12286) );
  NAND2_X1 U13775 ( .A1(n12287), .A2(n12286), .ZN(n12288) );
  NAND2_X1 U13776 ( .A1(n12333), .A2(n12288), .ZN(n15846) );
  NOR2_X1 U13777 ( .A1(n12384), .A2(n15846), .ZN(n12289) );
  AOI21_X1 U13778 ( .B1(n12291), .B2(n12290), .A(n12289), .ZN(n15630) );
  AOI22_X1 U13779 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U13780 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12340), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U13781 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U13782 ( .A1(n11871), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12292) );
  NAND4_X1 U13783 ( .A1(n12295), .A2(n12294), .A3(n12293), .A4(n12292), .ZN(
        n12302) );
  AOI22_X1 U13784 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U13785 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U13786 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U13787 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12297) );
  NAND4_X1 U13788 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n12301) );
  NOR2_X1 U13789 ( .A1(n12302), .A2(n12301), .ZN(n12314) );
  NAND2_X1 U13790 ( .A1(n12304), .A2(n12303), .ZN(n12313) );
  XOR2_X1 U13791 ( .A(n12314), .B(n12313), .Z(n12305) );
  NAND2_X1 U13792 ( .A1(n12305), .A2(n12353), .ZN(n12308) );
  INV_X1 U13793 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15841) );
  AOI21_X1 U13794 ( .B1(n15841), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12306) );
  AOI21_X1 U13795 ( .B1(n12386), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12306), .ZN(
        n12307) );
  NAND2_X1 U13796 ( .A1(n12308), .A2(n12307), .ZN(n12310) );
  XNOR2_X1 U13797 ( .A(n12333), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15839) );
  NAND2_X1 U13798 ( .A1(n15839), .A2(n11583), .ZN(n12309) );
  NAND2_X1 U13799 ( .A1(n12310), .A2(n12309), .ZN(n15621) );
  NOR2_X1 U13800 ( .A1(n12314), .A2(n12313), .ZN(n12352) );
  AOI22_X1 U13801 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U13802 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U13803 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U13804 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12316) );
  NAND4_X1 U13805 ( .A1(n12319), .A2(n12318), .A3(n12317), .A4(n12316), .ZN(
        n12327) );
  AOI22_X1 U13806 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U13807 ( .A1(n12321), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U13808 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U13809 ( .A1(n12340), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12367), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12322) );
  NAND4_X1 U13810 ( .A1(n12325), .A2(n12324), .A3(n12323), .A4(n12322), .ZN(
        n12326) );
  OR2_X1 U13811 ( .A1(n12327), .A2(n12326), .ZN(n12351) );
  INV_X1 U13812 ( .A(n12351), .ZN(n12328) );
  XNOR2_X1 U13813 ( .A(n12352), .B(n12328), .ZN(n12332) );
  INV_X1 U13814 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n15730) );
  NAND2_X1 U13815 ( .A1(n21922), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12329) );
  OAI211_X1 U13816 ( .C1(n12330), .C2(n15730), .A(n12384), .B(n12329), .ZN(
        n12331) );
  AOI21_X1 U13817 ( .B1(n12332), .B2(n12353), .A(n12331), .ZN(n12339) );
  NAND2_X1 U13818 ( .A1(n12334), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12358) );
  INV_X1 U13819 ( .A(n12334), .ZN(n12336) );
  INV_X1 U13820 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12335) );
  NAND2_X1 U13821 ( .A1(n12336), .A2(n12335), .ZN(n12337) );
  NAND2_X1 U13822 ( .A1(n12358), .A2(n12337), .ZN(n15833) );
  NOR2_X1 U13823 ( .A1(n15833), .A2(n12384), .ZN(n12338) );
  AOI22_X1 U13824 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U13825 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11735), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U13826 ( .A1(n11871), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12340), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U13827 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12341) );
  NAND4_X1 U13828 ( .A1(n12344), .A2(n12343), .A3(n12342), .A4(n12341), .ZN(
        n12350) );
  AOI22_X1 U13829 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12150), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12348) );
  AOI22_X1 U13830 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U13831 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U13832 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12345) );
  NAND4_X1 U13833 ( .A1(n12348), .A2(n12347), .A3(n12346), .A4(n12345), .ZN(
        n12349) );
  NOR2_X1 U13834 ( .A1(n12350), .A2(n12349), .ZN(n12375) );
  NAND2_X1 U13835 ( .A1(n12352), .A2(n12351), .ZN(n12374) );
  XOR2_X1 U13836 ( .A(n12375), .B(n12374), .Z(n12354) );
  NAND2_X1 U13837 ( .A1(n12354), .A2(n12353), .ZN(n12357) );
  INV_X1 U13838 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15813) );
  NOR2_X1 U13839 ( .A1(n15813), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12355) );
  AOI211_X1 U13840 ( .C1(n12386), .C2(P1_EAX_REG_29__SCAN_IN), .A(n12378), .B(
        n12355), .ZN(n12356) );
  XNOR2_X1 U13841 ( .A(n12358), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15815) );
  AOI22_X1 U13842 ( .A1(n12357), .A2(n12356), .B1(n12378), .B2(n15815), .ZN(
        n15596) );
  INV_X1 U13843 ( .A(n12358), .ZN(n12359) );
  XNOR2_X1 U13844 ( .A(n12388), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15809) );
  AOI22_X1 U13845 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11841), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U13846 ( .A1(n11736), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12315), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U13847 ( .A1(n12150), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12268), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U13848 ( .A1(n11846), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11981), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12361) );
  NAND4_X1 U13849 ( .A1(n12364), .A2(n12363), .A3(n12362), .A4(n12361), .ZN(
        n12373) );
  AOI22_X1 U13850 ( .A1(n10977), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11521), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U13851 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12320), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U13852 ( .A1(n10971), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12365), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U13853 ( .A1(n12367), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12368) );
  NAND4_X1 U13854 ( .A1(n12371), .A2(n12370), .A3(n12369), .A4(n12368), .ZN(
        n12372) );
  NOR2_X1 U13855 ( .A1(n12373), .A2(n12372), .ZN(n12377) );
  NOR2_X1 U13856 ( .A1(n12375), .A2(n12374), .ZN(n12376) );
  XOR2_X1 U13857 ( .A(n12377), .B(n12376), .Z(n12382) );
  AOI21_X1 U13858 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21922), .A(
        n12378), .ZN(n12380) );
  NAND2_X1 U13859 ( .A1(n12386), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n12379) );
  OAI211_X1 U13860 ( .C1(n12382), .C2(n12381), .A(n12380), .B(n12379), .ZN(
        n12383) );
  OAI21_X1 U13861 ( .B1(n12384), .B2(n15809), .A(n12383), .ZN(n12757) );
  AOI22_X1 U13862 ( .A1(n12386), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12385), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12387) );
  NAND2_X1 U13863 ( .A1(n12388), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12390) );
  INV_X1 U13864 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12389) );
  XNOR2_X1 U13865 ( .A(n12390), .B(n12389), .ZN(n14595) );
  NOR2_X1 U13866 ( .A1(n14595), .A2(n16886), .ZN(n12391) );
  NAND2_X1 U13867 ( .A1(n12774), .A2(n21618), .ZN(n12392) );
  NOR2_X1 U13868 ( .A1(n11695), .A2(n11681), .ZN(n12397) );
  INV_X1 U13869 ( .A(n12395), .ZN(n12396) );
  NAND2_X1 U13870 ( .A1(n12397), .A2(n12396), .ZN(n14069) );
  OR2_X1 U13871 ( .A1(n14069), .A2(n15578), .ZN(n14063) );
  INV_X1 U13872 ( .A(n21683), .ZN(n21691) );
  INV_X1 U13873 ( .A(n11695), .ZN(n13935) );
  AND2_X1 U13874 ( .A1(n13935), .A2(n11702), .ZN(n12398) );
  NAND2_X1 U13875 ( .A1(n12398), .A2(n16079), .ZN(n15567) );
  OAI21_X1 U13876 ( .B1(n14063), .B2(n21691), .A(n15567), .ZN(n13927) );
  NAND2_X1 U13877 ( .A1(n12393), .A2(n13927), .ZN(n12405) );
  NAND2_X1 U13878 ( .A1(n14410), .A2(n21683), .ZN(n12399) );
  OR2_X1 U13879 ( .A1(n13822), .A2(n12399), .ZN(n13938) );
  NOR2_X1 U13880 ( .A1(n12400), .A2(n21664), .ZN(n12402) );
  NOR2_X1 U13881 ( .A1(n11680), .A2(n15576), .ZN(n12401) );
  NAND4_X1 U13882 ( .A1(n14268), .A2(n12402), .A3(n12401), .A4(n11806), .ZN(
        n13989) );
  OAI22_X1 U13883 ( .A1(n13938), .A2(n21664), .B1(n15579), .B2(n13989), .ZN(
        n12403) );
  INV_X1 U13884 ( .A(n12403), .ZN(n12404) );
  AND2_X1 U13885 ( .A1(n15794), .A2(n11681), .ZN(n12406) );
  NOR4_X1 U13886 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12410) );
  NOR4_X1 U13887 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12409) );
  NOR4_X1 U13888 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12408) );
  NOR4_X1 U13889 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12407) );
  AND4_X1 U13890 ( .A1(n12410), .A2(n12409), .A3(n12408), .A4(n12407), .ZN(
        n12415) );
  NOR4_X1 U13891 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12413) );
  NOR4_X1 U13892 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12412) );
  NOR4_X1 U13893 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12411) );
  INV_X1 U13894 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n19845) );
  AND4_X1 U13895 ( .A1(n12413), .A2(n12412), .A3(n12411), .A4(n19845), .ZN(
        n12414) );
  NAND2_X1 U13896 ( .A1(n12415), .A2(n12414), .ZN(n12416) );
  AND2_X1 U13897 ( .A1(n12418), .A2(n15727), .ZN(n12417) );
  NAND2_X1 U13898 ( .A1(n15794), .A2(n12417), .ZN(n15786) );
  INV_X1 U13899 ( .A(DATAI_31_), .ZN(n14396) );
  NOR2_X1 U13900 ( .A1(n15786), .A2(n14396), .ZN(n12421) );
  INV_X1 U13901 ( .A(n12418), .ZN(n14051) );
  NOR3_X4 U13902 ( .A1(n15798), .A2(n14051), .A3(n15727), .ZN(n15788) );
  AOI22_X1 U13903 ( .A1(n15788), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n15798), .ZN(n12419) );
  NOR2_X1 U13904 ( .A1(n12421), .A2(n12420), .ZN(n12422) );
  NAND2_X1 U13905 ( .A1(n12423), .A2(n12422), .ZN(P1_U2873) );
  INV_X1 U13906 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12545) );
  BUF_X4 U13907 ( .A(n17640), .Z(n17667) );
  NOR2_X2 U13908 ( .A1(n12431), .A2(n12432), .ZN(n12474) );
  AOI22_X1 U13909 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12429) );
  INV_X2 U13910 ( .A(n17598), .ZN(n17641) );
  AOI22_X1 U13911 ( .A1(n17641), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12428) );
  AOI22_X1 U13912 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12427) );
  NOR3_X1 U13913 ( .A1(n20784), .A2(n12698), .A3(n20821), .ZN(n12424) );
  INV_X1 U13914 ( .A(n12424), .ZN(n12463) );
  INV_X2 U13915 ( .A(n12463), .ZN(n17353) );
  AOI22_X1 U13916 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12426) );
  NAND4_X1 U13917 ( .A1(n12429), .A2(n12428), .A3(n12427), .A4(n12426), .ZN(
        n12440) );
  BUF_X4 U13918 ( .A(n12475), .Z(n17668) );
  BUF_X4 U13919 ( .A(n12481), .Z(n17664) );
  AOI22_X1 U13920 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U13921 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12465), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12437) );
  NOR2_X2 U13922 ( .A1(n12434), .A2(n20821), .ZN(n17658) );
  AOI22_X1 U13923 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U13924 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12435) );
  NAND4_X1 U13925 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        n12439) );
  AOI22_X1 U13926 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10960), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17658), .ZN(n12444) );
  AOI22_X1 U13927 ( .A1(n12512), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12474), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U13928 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12517), .B1(
        n12529), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12442) );
  INV_X2 U13929 ( .A(n12463), .ZN(n17627) );
  AOI22_X1 U13930 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12425), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12424), .ZN(n12441) );
  NAND4_X1 U13931 ( .A1(n12444), .A2(n12443), .A3(n12442), .A4(n12441), .ZN(
        n12450) );
  AOI22_X1 U13932 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12452), .B1(
        n12557), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U13933 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12451), .B1(
        n12482), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U13934 ( .A1(n12475), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17641), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U13935 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12465), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n12481), .ZN(n12445) );
  NAND4_X1 U13936 ( .A1(n12448), .A2(n12447), .A3(n12446), .A4(n12445), .ZN(
        n12449) );
  INV_X2 U13937 ( .A(n12572), .ZN(n17666) );
  AOI22_X1 U13938 ( .A1(n17641), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17666), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U13939 ( .A1(n12475), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12452), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U13940 ( .A1(n12424), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12481), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U13941 ( .A1(n12529), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12425), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12453) );
  NAND4_X1 U13942 ( .A1(n12456), .A2(n12455), .A3(n12454), .A4(n12453), .ZN(
        n12462) );
  AOI22_X1 U13943 ( .A1(n12512), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12482), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12460) );
  AOI22_X1 U13944 ( .A1(n12465), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12474), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U13945 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10980), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U13946 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17658), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12457) );
  NAND4_X1 U13947 ( .A1(n12460), .A2(n12459), .A3(n12458), .A4(n12457), .ZN(
        n12461) );
  OR2_X2 U13948 ( .A1(n12462), .A2(n12461), .ZN(n20647) );
  INV_X1 U13949 ( .A(n12672), .ZN(n12473) );
  AOI22_X1 U13950 ( .A1(n10980), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U13951 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12471) );
  INV_X1 U13952 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17509) );
  AOI22_X1 U13953 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12464) );
  OAI21_X1 U13954 ( .B1(n20196), .B2(n17509), .A(n12464), .ZN(n12470) );
  AOI22_X1 U13955 ( .A1(n17641), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17658), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U13956 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12468) );
  AOI22_X1 U13957 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17536), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12467) );
  AOI22_X1 U13958 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12466) );
  XOR2_X1 U13959 ( .A(n20639), .B(n12508), .Z(n12496) );
  INV_X1 U13960 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20871) );
  XNOR2_X1 U13961 ( .A(n20774), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18077) );
  AOI22_X1 U13962 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17658), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U13963 ( .A1(n12529), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12465), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U13964 ( .A1(n12475), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12474), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U13965 ( .A1(n12512), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17641), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U13966 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17640), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12488) );
  INV_X1 U13967 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17326) );
  OAI21_X1 U13968 ( .B1(n12463), .B2(n17326), .A(n12480), .ZN(n12486) );
  AOI22_X1 U13969 ( .A1(n12451), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12481), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12484) );
  NAND2_X1 U13970 ( .A1(n12484), .A2(n12483), .ZN(n12485) );
  NAND3_X1 U13971 ( .A1(n11401), .A2(n12488), .A3(n12487), .ZN(n20775) );
  INV_X1 U13972 ( .A(n20774), .ZN(n12490) );
  NOR2_X1 U13973 ( .A1(n20871), .A2(n12492), .ZN(n12493) );
  NOR2_X2 U13974 ( .A1(n18067), .A2(n12493), .ZN(n12494) );
  INV_X1 U13975 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20878) );
  NOR2_X1 U13976 ( .A1(n12494), .A2(n20878), .ZN(n12495) );
  XNOR2_X1 U13977 ( .A(n12494), .B(n20878), .ZN(n18057) );
  XOR2_X1 U13978 ( .A(n20644), .B(n12672), .Z(n18056) );
  NOR2_X1 U13979 ( .A1(n18057), .A2(n18056), .ZN(n18055) );
  NOR2_X1 U13980 ( .A1(n12495), .A2(n18055), .ZN(n18045) );
  XNOR2_X1 U13981 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12496), .ZN(
        n18044) );
  NOR2_X1 U13982 ( .A1(n18045), .A2(n18044), .ZN(n18043) );
  NOR2_X2 U13983 ( .A1(n12497), .A2(n18043), .ZN(n12509) );
  AOI22_X1 U13984 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12507) );
  AOI22_X1 U13985 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17656), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12506) );
  INV_X1 U13986 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17522) );
  AOI22_X1 U13987 ( .A1(n17659), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12498) );
  OAI21_X1 U13988 ( .B1(n20196), .B2(n17522), .A(n12498), .ZN(n12504) );
  AOI22_X1 U13989 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12465), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U13990 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17666), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12501) );
  INV_X2 U13991 ( .A(n17598), .ZN(n17657) );
  AOI22_X1 U13992 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17657), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U13993 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12499) );
  NAND4_X1 U13994 ( .A1(n12502), .A2(n12501), .A3(n12500), .A4(n12499), .ZN(
        n12503) );
  AOI211_X1 U13995 ( .C1(n10960), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n12504), .B(n12503), .ZN(n12505) );
  NAND3_X1 U13996 ( .A1(n12507), .A2(n12506), .A3(n12505), .ZN(n12666) );
  XNOR2_X1 U13997 ( .A(n12666), .B(n12525), .ZN(n12510) );
  NOR2_X1 U13998 ( .A1(n12509), .A2(n12510), .ZN(n12511) );
  INV_X1 U13999 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20903) );
  XNOR2_X1 U14000 ( .A(n12510), .B(n12509), .ZN(n18035) );
  AOI22_X1 U14001 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17640), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12516) );
  AOI22_X1 U14002 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12515) );
  AOI22_X1 U14003 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12514) );
  AOI22_X1 U14004 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12513) );
  NAND4_X1 U14005 ( .A1(n12516), .A2(n12515), .A3(n12514), .A4(n12513), .ZN(
        n12524) );
  AOI22_X1 U14006 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17666), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12522) );
  AOI22_X1 U14007 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12521) );
  AOI22_X1 U14008 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12520) );
  AOI22_X1 U14009 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12519) );
  NAND4_X1 U14010 ( .A1(n12522), .A2(n12521), .A3(n12520), .A4(n12519), .ZN(
        n12523) );
  NAND2_X1 U14011 ( .A1(n12525), .A2(n12666), .ZN(n12527) );
  XOR2_X1 U14012 ( .A(n20631), .B(n12527), .Z(n12526) );
  XNOR2_X1 U14013 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12526), .ZN(
        n18025) );
  AOI22_X1 U14014 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12538) );
  AOI22_X1 U14015 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10980), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12537) );
  INV_X1 U14016 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17315) );
  AOI22_X1 U14017 ( .A1(n17659), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12528) );
  OAI21_X1 U14018 ( .B1(n20196), .B2(n17315), .A(n12528), .ZN(n12535) );
  AOI22_X1 U14019 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12533) );
  AOI22_X1 U14020 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U14021 ( .A1(n17641), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17666), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U14022 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12530) );
  NAND4_X1 U14023 ( .A1(n12533), .A2(n12532), .A3(n12531), .A4(n12530), .ZN(
        n12534) );
  AOI211_X1 U14024 ( .C1(n17640), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n12535), .B(n12534), .ZN(n12536) );
  NAND3_X1 U14025 ( .A1(n12538), .A2(n12537), .A3(n12536), .ZN(n12663) );
  OAI21_X1 U14026 ( .B1(n12539), .B2(n12663), .A(n17869), .ZN(n12540) );
  NOR2_X1 U14027 ( .A1(n17718), .A2(n12540), .ZN(n12541) );
  INV_X1 U14028 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20927) );
  NOR2_X2 U14029 ( .A1(n20927), .A2(n18018), .ZN(n18017) );
  INV_X1 U14030 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20943) );
  AOI22_X1 U14031 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17971), .B1(
        n17869), .B2(n20943), .ZN(n17998) );
  NOR2_X1 U14032 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17976) );
  INV_X1 U14033 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20956) );
  INV_X1 U14034 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21166) );
  NAND2_X1 U14035 ( .A1(n17756), .A2(n21166), .ZN(n17720) );
  INV_X1 U14036 ( .A(n17720), .ZN(n12544) );
  NAND3_X1 U14037 ( .A1(n12545), .A2(n17950), .A3(n12544), .ZN(n12546) );
  NAND2_X1 U14038 ( .A1(n12546), .A2(n17869), .ZN(n12549) );
  NAND2_X1 U14039 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n20946) );
  INV_X1 U14040 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n20968) );
  NOR3_X1 U14041 ( .A1(n20946), .A2(n20968), .A3(n20956), .ZN(n20957) );
  NAND2_X1 U14042 ( .A1(n20957), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17719) );
  INV_X1 U14043 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17950) );
  NOR2_X1 U14044 ( .A1(n17719), .A2(n17950), .ZN(n20995) );
  NAND2_X1 U14045 ( .A1(n20995), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21139) );
  INV_X1 U14046 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21155) );
  OAI22_X2 U14047 ( .A1(n12550), .A2(n21155), .B1(n17869), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U14048 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21132) );
  INV_X1 U14049 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17790) );
  INV_X1 U14050 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21120) );
  NOR2_X1 U14051 ( .A1(n17790), .A2(n21120), .ZN(n20841) );
  NAND2_X1 U14052 ( .A1(n20841), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21019) );
  INV_X1 U14053 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17703) );
  NAND2_X1 U14054 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17827) );
  NOR2_X1 U14055 ( .A1(n21132), .A2(n17703), .ZN(n17704) );
  INV_X1 U14056 ( .A(n21019), .ZN(n12743) );
  NAND2_X1 U14057 ( .A1(n17704), .A2(n12743), .ZN(n17765) );
  NOR2_X1 U14058 ( .A1(n17971), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17788) );
  NOR2_X1 U14059 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17780) );
  INV_X1 U14060 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21007) );
  NAND3_X1 U14061 ( .A1(n17788), .A2(n17780), .A3(n21007), .ZN(n17763) );
  NOR2_X1 U14062 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17763), .ZN(
        n17808) );
  INV_X1 U14063 ( .A(n17808), .ZN(n12551) );
  OAI22_X1 U14064 ( .A1(n11398), .A2(n17732), .B1(n12551), .B2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12552) );
  INV_X1 U14065 ( .A(n12552), .ZN(n12553) );
  INV_X1 U14066 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21101) );
  INV_X1 U14067 ( .A(n17827), .ZN(n12554) );
  INV_X1 U14068 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21057) );
  INV_X1 U14069 ( .A(n12751), .ZN(n12890) );
  NOR2_X2 U14070 ( .A1(n12556), .A2(n21057), .ZN(n12662) );
  NOR2_X1 U14071 ( .A1(n12890), .A2(n12662), .ZN(n17853) );
  NAND2_X1 U14072 ( .A1(n17853), .A2(n17971), .ZN(n17852) );
  NAND2_X1 U14073 ( .A1(n17852), .A2(n12751), .ZN(n17846) );
  NOR2_X1 U14074 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17971), .ZN(
        n12889) );
  AOI21_X1 U14075 ( .B1(n17971), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12889), .ZN(n17847) );
  AOI22_X1 U14076 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U14077 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12560) );
  AOI22_X1 U14078 ( .A1(n17664), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17658), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U14079 ( .A1(n17353), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12558) );
  NAND4_X1 U14080 ( .A1(n12561), .A2(n12560), .A3(n12559), .A4(n12558), .ZN(
        n12567) );
  AOI22_X1 U14081 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17657), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U14082 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17668), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U14083 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10980), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U14084 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12562) );
  NAND4_X1 U14085 ( .A1(n12565), .A2(n12564), .A3(n12563), .A4(n12562), .ZN(
        n12566) );
  NOR2_X4 U14086 ( .A1(n12567), .A2(n12566), .ZN(n20158) );
  INV_X1 U14087 ( .A(n20158), .ZN(n12661) );
  AOI22_X1 U14088 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12571) );
  AOI22_X1 U14089 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17536), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U14090 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U14091 ( .A1(n17353), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12568) );
  NAND4_X1 U14092 ( .A1(n12571), .A2(n12570), .A3(n12569), .A4(n12568), .ZN(
        n12578) );
  AOI22_X1 U14093 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17658), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U14094 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U14095 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17640), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U14096 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12474), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12573) );
  NAND4_X1 U14097 ( .A1(n12576), .A2(n12575), .A3(n12574), .A4(n12573), .ZN(
        n12577) );
  AOI22_X1 U14098 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17668), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U14099 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12588) );
  INV_X1 U14100 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17597) );
  AOI22_X1 U14101 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17658), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12580) );
  OAI21_X1 U14102 ( .B1(n12579), .B2(n17597), .A(n12580), .ZN(n12586) );
  AOI22_X1 U14103 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10980), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U14104 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12474), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U14105 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U14106 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17627), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12581) );
  NAND4_X1 U14107 ( .A1(n12584), .A2(n12583), .A3(n12582), .A4(n12581), .ZN(
        n12585) );
  AOI211_X1 U14108 ( .C1(n17656), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n12586), .B(n12585), .ZN(n12587) );
  NAND3_X1 U14109 ( .A1(n12589), .A2(n12588), .A3(n12587), .ZN(n12621) );
  NAND2_X1 U14110 ( .A1(n18772), .A2(n12621), .ZN(n12720) );
  AOI22_X1 U14111 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17657), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U14112 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17666), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U14113 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U14114 ( .A1(n17353), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12590) );
  NAND4_X1 U14115 ( .A1(n12593), .A2(n12592), .A3(n12591), .A4(n12590), .ZN(
        n12599) );
  AOI22_X1 U14116 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17658), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U14117 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U14118 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U14119 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12594) );
  NAND4_X1 U14120 ( .A1(n12597), .A2(n12596), .A3(n12595), .A4(n12594), .ZN(
        n12598) );
  AOI22_X1 U14121 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U14122 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10980), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12608) );
  INV_X1 U14123 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17405) );
  AOI22_X1 U14124 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12600) );
  OAI21_X1 U14125 ( .B1(n12579), .B2(n17405), .A(n12600), .ZN(n12606) );
  AOI22_X1 U14126 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12474), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U14127 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12603) );
  AOI22_X1 U14128 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17658), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U14129 ( .A1(n17353), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12601) );
  NAND4_X1 U14130 ( .A1(n12604), .A2(n12603), .A3(n12602), .A4(n12601), .ZN(
        n12605) );
  AOI211_X1 U14131 ( .C1(n17668), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n12606), .B(n12605), .ZN(n12607) );
  NAND3_X1 U14132 ( .A1(n12609), .A2(n12608), .A3(n12607), .ZN(n12650) );
  INV_X2 U14133 ( .A(n12650), .ZN(n18891) );
  NOR2_X2 U14134 ( .A1(n18772), .A2(n12621), .ZN(n20602) );
  INV_X1 U14135 ( .A(n12621), .ZN(n20656) );
  AOI22_X1 U14136 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17658), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U14137 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12618) );
  INV_X1 U14138 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17295) );
  AOI22_X1 U14139 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12474), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12610) );
  OAI21_X1 U14140 ( .B1(n12579), .B2(n17295), .A(n12610), .ZN(n12616) );
  AOI22_X1 U14141 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U14142 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U14143 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U14144 ( .A1(n17353), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12611) );
  NAND4_X1 U14145 ( .A1(n12614), .A2(n12613), .A3(n12612), .A4(n12611), .ZN(
        n12615) );
  AOI211_X1 U14146 ( .C1(n17599), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n12616), .B(n12615), .ZN(n12617) );
  NAND3_X1 U14147 ( .A1(n12619), .A2(n12618), .A3(n12617), .ZN(n12730) );
  NAND2_X1 U14148 ( .A1(n20656), .A2(n12730), .ZN(n20796) );
  INV_X1 U14149 ( .A(n20796), .ZN(n12620) );
  NAND2_X1 U14150 ( .A1(n12621), .A2(n20655), .ZN(n12734) );
  AOI22_X1 U14151 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U14152 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U14153 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12622) );
  OAI21_X1 U14154 ( .B1(n12579), .B2(n17315), .A(n12622), .ZN(n12628) );
  AOI22_X1 U14155 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12626) );
  AOI22_X1 U14156 ( .A1(n17659), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17658), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U14157 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U14158 ( .A1(n17353), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12623) );
  NAND4_X1 U14159 ( .A1(n12626), .A2(n12625), .A3(n12624), .A4(n12623), .ZN(
        n12627) );
  NOR2_X1 U14160 ( .A1(n20156), .A2(n12661), .ZN(n12659) );
  INV_X1 U14161 ( .A(n20602), .ZN(n20782) );
  NAND2_X1 U14162 ( .A1(n20693), .A2(n20782), .ZN(n20600) );
  NAND2_X1 U14163 ( .A1(n12659), .A2(n20600), .ZN(n12726) );
  OAI211_X1 U14164 ( .C1(n12734), .C2(n18811), .A(n20693), .B(n12726), .ZN(
        n12648) );
  AOI22_X1 U14165 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U14166 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U14167 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17640), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U14168 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12632) );
  NAND4_X1 U14169 ( .A1(n12635), .A2(n12634), .A3(n12633), .A4(n12632), .ZN(
        n12641) );
  AOI22_X1 U14170 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12639) );
  AOI22_X1 U14171 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12638) );
  AOI22_X1 U14172 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12637) );
  AOI22_X1 U14173 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12636) );
  NAND4_X1 U14174 ( .A1(n12639), .A2(n12638), .A3(n12637), .A4(n12636), .ZN(
        n12640) );
  NAND2_X1 U14175 ( .A1(n18891), .A2(n18811), .ZN(n12727) );
  INV_X1 U14176 ( .A(n12727), .ZN(n12642) );
  NOR2_X1 U14177 ( .A1(n18772), .A2(n12650), .ZN(n12719) );
  OAI21_X1 U14178 ( .B1(n12642), .B2(n12719), .A(n12720), .ZN(n12643) );
  INV_X1 U14179 ( .A(n12643), .ZN(n12651) );
  NOR2_X1 U14180 ( .A1(n20592), .A2(n20158), .ZN(n12658) );
  INV_X1 U14181 ( .A(n12658), .ZN(n12654) );
  NAND2_X1 U14182 ( .A1(n18891), .A2(n12654), .ZN(n12724) );
  NAND2_X1 U14183 ( .A1(n12734), .A2(n12724), .ZN(n12644) );
  OAI21_X1 U14184 ( .B1(n12651), .B2(n18851), .A(n12644), .ZN(n12645) );
  AOI21_X1 U14185 ( .B1(n18851), .B2(n12657), .A(n12645), .ZN(n12646) );
  INV_X1 U14186 ( .A(n12646), .ZN(n12647) );
  AOI211_X2 U14187 ( .C1(n12720), .C2(n12652), .A(n12648), .B(n12647), .ZN(
        n12693) );
  INV_X1 U14188 ( .A(n12693), .ZN(n20798) );
  NAND2_X1 U14189 ( .A1(n18891), .A2(n18851), .ZN(n20795) );
  NOR2_X1 U14190 ( .A1(n12720), .A2(n20795), .ZN(n17291) );
  NAND2_X1 U14191 ( .A1(n20158), .A2(n17291), .ZN(n12656) );
  INV_X1 U14192 ( .A(n18851), .ZN(n12649) );
  NAND2_X1 U14193 ( .A1(n10972), .A2(n12650), .ZN(n12722) );
  INV_X1 U14194 ( .A(n12722), .ZN(n12653) );
  NOR2_X2 U14195 ( .A1(n12653), .A2(n12655), .ZN(n21198) );
  NAND2_X1 U14196 ( .A1(n20158), .A2(n12655), .ZN(n21239) );
  NOR2_X1 U14197 ( .A1(n12659), .A2(n12658), .ZN(n20102) );
  INV_X1 U14198 ( .A(n17697), .ZN(n21209) );
  INV_X1 U14199 ( .A(n12663), .ZN(n20626) );
  NAND3_X1 U14200 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17971), .A3(
        n12662), .ZN(n17910) );
  NAND2_X1 U14201 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12900) );
  INV_X1 U14202 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21016) );
  NAND2_X1 U14203 ( .A1(n17869), .A2(n17999), .ZN(n17955) );
  INV_X2 U14204 ( .A(n21130), .ZN(n20958) );
  INV_X1 U14205 ( .A(n17719), .ZN(n20969) );
  NAND2_X1 U14206 ( .A1(n20958), .A2(n20969), .ZN(n17948) );
  NAND2_X1 U14207 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21084), .ZN(
        n17822) );
  NOR2_X1 U14208 ( .A1(n21016), .A2(n17822), .ZN(n17821) );
  NAND2_X1 U14209 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17821), .ZN(
        n21034) );
  NOR2_X1 U14210 ( .A1(n12900), .A2(n21034), .ZN(n21058) );
  INV_X1 U14211 ( .A(n21131), .ZN(n21063) );
  INV_X1 U14212 ( .A(n20775), .ZN(n12674) );
  NOR2_X1 U14213 ( .A1(n20774), .A2(n12674), .ZN(n12676) );
  NAND2_X1 U14214 ( .A1(n20644), .A2(n12671), .ZN(n12669) );
  NOR2_X1 U14215 ( .A1(n12669), .A2(n20639), .ZN(n12667) );
  NAND2_X1 U14216 ( .A1(n12666), .A2(n12667), .ZN(n12665) );
  NOR2_X1 U14217 ( .A1(n12665), .A2(n20631), .ZN(n12664) );
  AND2_X1 U14218 ( .A1(n12663), .A2(n12664), .ZN(n12689) );
  XNOR2_X1 U14219 ( .A(n20626), .B(n12664), .ZN(n18011) );
  XOR2_X1 U14220 ( .A(n20631), .B(n12665), .Z(n12683) );
  INV_X1 U14221 ( .A(n12666), .ZN(n20634) );
  XNOR2_X1 U14222 ( .A(n20634), .B(n12667), .ZN(n12668) );
  NAND2_X1 U14223 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12668), .ZN(
        n12682) );
  XNOR2_X1 U14224 ( .A(n20903), .B(n12668), .ZN(n18033) );
  XOR2_X1 U14225 ( .A(n20639), .B(n12669), .Z(n12679) );
  NAND2_X1 U14226 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12670), .ZN(
        n12678) );
  XNOR2_X1 U14227 ( .A(n20878), .B(n12670), .ZN(n18054) );
  OAI21_X1 U14228 ( .B1(n12674), .B2(n12672), .A(n12671), .ZN(n12673) );
  NAND2_X1 U14229 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12673), .ZN(
        n12677) );
  XOR2_X1 U14230 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12673), .Z(
        n18073) );
  NOR2_X1 U14231 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12490), .ZN(
        n12675) );
  INV_X1 U14232 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20860) );
  NAND2_X1 U14233 ( .A1(n12674), .A2(n20860), .ZN(n18085) );
  INV_X1 U14234 ( .A(n18077), .ZN(n18079) );
  NOR2_X1 U14235 ( .A1(n18085), .A2(n18079), .ZN(n18078) );
  NOR3_X1 U14236 ( .A1(n12676), .A2(n12675), .A3(n18078), .ZN(n18072) );
  NAND2_X1 U14237 ( .A1(n18073), .A2(n18072), .ZN(n18071) );
  NAND2_X1 U14238 ( .A1(n12677), .A2(n18071), .ZN(n18053) );
  NAND2_X1 U14239 ( .A1(n18054), .A2(n18053), .ZN(n18052) );
  NAND2_X1 U14240 ( .A1(n12678), .A2(n18052), .ZN(n12680) );
  NAND2_X1 U14241 ( .A1(n12679), .A2(n12680), .ZN(n12681) );
  XOR2_X1 U14242 ( .A(n12680), .B(n12679), .Z(n18042) );
  NAND2_X1 U14243 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18042), .ZN(
        n18041) );
  NAND2_X1 U14244 ( .A1(n12683), .A2(n12684), .ZN(n12685) );
  NAND2_X1 U14245 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18023), .ZN(
        n18022) );
  NAND2_X1 U14246 ( .A1(n12689), .A2(n12686), .ZN(n12690) );
  NAND2_X1 U14247 ( .A1(n18011), .A2(n18012), .ZN(n18010) );
  NAND2_X1 U14248 ( .A1(n12689), .A2(n12688), .ZN(n12687) );
  OAI211_X1 U14249 ( .C1(n12689), .C2(n12688), .A(n18010), .B(n12687), .ZN(
        n18001) );
  NAND2_X1 U14250 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18001), .ZN(
        n18000) );
  NAND2_X1 U14251 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21087), .ZN(
        n17824) );
  NOR2_X1 U14252 ( .A1(n12900), .A2(n21032), .ZN(n21061) );
  OAI22_X1 U14253 ( .A1(n21058), .A2(n21063), .B1(n21061), .B2(n21202), .ZN(
        n12691) );
  INV_X1 U14254 ( .A(n21203), .ZN(n21133) );
  INV_X1 U14255 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21038) );
  NAND4_X1 U14256 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21031) );
  NOR2_X1 U14257 ( .A1(n21038), .A2(n21031), .ZN(n17904) );
  INV_X1 U14258 ( .A(n17904), .ZN(n21044) );
  INV_X1 U14259 ( .A(n21139), .ZN(n20832) );
  NAND2_X1 U14260 ( .A1(n20832), .A2(n17704), .ZN(n12742) );
  OAI21_X1 U14261 ( .B1(n12489), .B2(n20860), .A(n20871), .ZN(n20873) );
  INV_X1 U14262 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12692) );
  NOR3_X1 U14263 ( .A1(n20903), .A2(n20878), .A3(n12692), .ZN(n20906) );
  AND2_X1 U14264 ( .A1(n20873), .A2(n20906), .ZN(n20897) );
  NAND4_X1 U14265 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n20897), .ZN(n20936) );
  NOR2_X1 U14266 ( .A1(n12742), .A2(n20936), .ZN(n20836) );
  NAND2_X1 U14267 ( .A1(n20836), .A2(n12743), .ZN(n21015) );
  OAI21_X1 U14268 ( .B1(n21044), .B2(n21015), .A(n21133), .ZN(n12898) );
  NAND2_X1 U14269 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n12898), .ZN(
        n21045) );
  OAI21_X1 U14270 ( .B1(n20786), .B2(n20795), .A(n12693), .ZN(n20954) );
  INV_X1 U14271 ( .A(n20954), .ZN(n21004) );
  NAND2_X1 U14272 ( .A1(n17904), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12744) );
  INV_X1 U14273 ( .A(n12744), .ZN(n17844) );
  NAND3_X1 U14274 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12694) );
  NAND3_X1 U14275 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n20906), .ZN(n20895) );
  NOR2_X1 U14276 ( .A1(n12694), .A2(n20895), .ZN(n21184) );
  NAND2_X1 U14277 ( .A1(n20832), .A2(n21184), .ZN(n21134) );
  NOR2_X1 U14278 ( .A1(n21134), .A2(n17765), .ZN(n21013) );
  NAND2_X1 U14279 ( .A1(n20860), .A2(n20954), .ZN(n21049) );
  OAI221_X1 U14280 ( .B1(n21004), .B2(n17844), .C1(n21004), .C2(n21013), .A(
        n21049), .ZN(n12896) );
  AOI21_X1 U14281 ( .B1(n21133), .B2(n21045), .A(n12896), .ZN(n21067) );
  NAND2_X1 U14282 ( .A1(n17904), .A2(n21013), .ZN(n21047) );
  INV_X1 U14283 ( .A(n20786), .ZN(n12697) );
  NAND2_X1 U14284 ( .A1(n10972), .A2(n12695), .ZN(n21204) );
  NAND2_X1 U14285 ( .A1(n12697), .A2(n21204), .ZN(n20955) );
  OAI21_X1 U14286 ( .B1(n21045), .B2(n21047), .A(n20955), .ZN(n12739) );
  NOR2_X1 U14287 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21255) );
  NAND2_X1 U14288 ( .A1(n21255), .A2(n21252), .ZN(n17691) );
  INV_X1 U14289 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18652) );
  AOI22_X1 U14290 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18652), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20808), .ZN(n12704) );
  AOI22_X1 U14291 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21217), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n20794), .ZN(n12717) );
  INV_X1 U14292 ( .A(n12717), .ZN(n12703) );
  NAND2_X1 U14293 ( .A1(n21216), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12716) );
  NAND2_X1 U14294 ( .A1(n12704), .A2(n12705), .ZN(n12700) );
  OAI21_X1 U14295 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20808), .A(
        n12700), .ZN(n12701) );
  OAI22_X1 U14296 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16822), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12701), .ZN(n12706) );
  NOR2_X1 U14297 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16822), .ZN(
        n12702) );
  NAND2_X1 U14298 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12701), .ZN(
        n12707) );
  AOI22_X1 U14299 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12706), .B1(
        n12702), .B2(n12707), .ZN(n12712) );
  OAI21_X1 U14300 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21216), .A(
        n12716), .ZN(n12732) );
  NOR2_X1 U14301 ( .A1(n12703), .A2(n12732), .ZN(n12711) );
  XNOR2_X1 U14302 ( .A(n12705), .B(n12704), .ZN(n12710) );
  INV_X1 U14303 ( .A(n12712), .ZN(n12709) );
  AOI21_X1 U14304 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12707), .A(
        n12706), .ZN(n12708) );
  AOI21_X1 U14305 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n16822), .A(
        n12708), .ZN(n12714) );
  OAI21_X1 U14306 ( .B1(n12710), .B2(n12709), .A(n12714), .ZN(n12713) );
  AOI21_X1 U14307 ( .B1(n12712), .B2(n12711), .A(n12713), .ZN(n17696) );
  INV_X1 U14308 ( .A(n12713), .ZN(n12731) );
  OAI21_X1 U14309 ( .B1(n12717), .B2(n12716), .A(n12714), .ZN(n12715) );
  AOI21_X1 U14310 ( .B1(n12717), .B2(n12716), .A(n12715), .ZN(n12733) );
  XOR2_X1 U14311 ( .A(n20158), .B(n18891), .Z(n12718) );
  NAND2_X1 U14312 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n21678), .ZN(n21721) );
  INV_X1 U14313 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21726) );
  AOI21_X1 U14314 ( .B1(n21724), .B2(n21721), .A(n18205), .ZN(n20155) );
  NAND2_X1 U14315 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n21723) );
  OAI21_X1 U14316 ( .B1(n12718), .B2(n20155), .A(n21723), .ZN(n21201) );
  NOR3_X1 U14317 ( .A1(n12719), .A2(n21207), .A3(n21201), .ZN(n12729) );
  OAI211_X1 U14318 ( .C1(n20602), .C2(n18811), .A(n12721), .B(n12720), .ZN(
        n12723) );
  OAI21_X1 U14319 ( .B1(n12724), .B2(n12723), .A(n12722), .ZN(n12725) );
  OAI211_X1 U14320 ( .C1(n12728), .C2(n12727), .A(n12726), .B(n12725), .ZN(
        n16806) );
  AOI211_X1 U14321 ( .C1(n17696), .C2(n12730), .A(n12729), .B(n16806), .ZN(
        n12738) );
  AOI21_X1 U14322 ( .B1(n12733), .B2(n12732), .A(n12731), .ZN(n21210) );
  NOR2_X1 U14323 ( .A1(n20158), .A2(n21210), .ZN(n12736) );
  INV_X1 U14324 ( .A(n12734), .ZN(n12735) );
  OAI211_X1 U14325 ( .C1(n12736), .C2(n17696), .A(n12735), .B(n18891), .ZN(
        n12737) );
  INV_X1 U14326 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n17690) );
  NOR2_X1 U14327 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17690), .ZN(n21243) );
  NAND2_X1 U14328 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21243), .ZN(n21263) );
  AOI21_X2 U14329 ( .B1(n12738), .B2(n12737), .A(n21263), .ZN(n21078) );
  NAND4_X1 U14330 ( .A1(n12740), .A2(n21067), .A3(n12739), .A4(n21086), .ZN(
        n12750) );
  AOI22_X1 U14331 ( .A1(n21111), .A2(n17957), .B1(n21131), .B2(n20958), .ZN(
        n20944) );
  NOR2_X1 U14332 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20955), .ZN(
        n20852) );
  NOR2_X1 U14333 ( .A1(n20874), .A2(n20852), .ZN(n20872) );
  INV_X1 U14334 ( .A(n17704), .ZN(n20833) );
  NOR2_X1 U14335 ( .A1(n20833), .A2(n21134), .ZN(n12741) );
  AOI22_X1 U14336 ( .A1(n21133), .A2(n20836), .B1(n20872), .B2(n12741), .ZN(
        n21020) );
  OAI21_X1 U14337 ( .B1(n20944), .B2(n12742), .A(n21020), .ZN(n20829) );
  NAND2_X1 U14338 ( .A1(n12743), .A2(n20829), .ZN(n21093) );
  OAI22_X1 U14339 ( .A1(n17869), .A2(n12745), .B1(n21093), .B2(n12744), .ZN(
        n12746) );
  NAND2_X1 U14340 ( .A1(n12746), .A2(n21078), .ZN(n12748) );
  NAND2_X1 U14341 ( .A1(n12748), .A2(n12747), .ZN(n12749) );
  NAND3_X1 U14342 ( .A1(n12750), .A2(n12749), .A3(n10961), .ZN(n12754) );
  NAND2_X1 U14343 ( .A1(n21078), .A2(n21209), .ZN(n20923) );
  NAND2_X1 U14344 ( .A1(n21189), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17841) );
  INV_X1 U14345 ( .A(n17841), .ZN(n12752) );
  NAND2_X1 U14346 ( .A1(n12754), .A2(n12753), .ZN(P3_U2834) );
  AOI21_X1 U14347 ( .B1(n12757), .B2(n12755), .A(n12756), .ZN(n15811) );
  INV_X1 U14348 ( .A(n15811), .ZN(n15663) );
  NAND2_X1 U14349 ( .A1(n12758), .A2(n15576), .ZN(n14218) );
  NOR3_X4 U14350 ( .A1(n15798), .A2(n12394), .A3(n11680), .ZN(n15790) );
  MUX2_X1 U14351 ( .A(BUF1_REG_14__SCAN_IN), .B(DATAI_14_), .S(n15727), .Z(
        n21770) );
  AOI22_X1 U14352 ( .A1(n15790), .A2(n21770), .B1(n15788), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12759) );
  INV_X1 U14353 ( .A(n12759), .ZN(n12762) );
  INV_X1 U14354 ( .A(DATAI_30_), .ZN(n16909) );
  INV_X1 U14355 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12760) );
  OAI22_X1 U14356 ( .A1(n15786), .A2(n16909), .B1(n12760), .B2(n15794), .ZN(
        n12761) );
  NOR2_X1 U14357 ( .A1(n12762), .A2(n12761), .ZN(n12763) );
  OAI21_X1 U14358 ( .B1(n15663), .B2(n15801), .A(n12763), .ZN(P1_U2874) );
  NAND3_X1 U14359 ( .A1(n21655), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n21652) );
  INV_X1 U14360 ( .A(n21652), .ZN(n12764) );
  NAND2_X1 U14361 ( .A1(n11683), .A2(n11682), .ZN(n12765) );
  AND2_X1 U14362 ( .A1(n12766), .A2(n12765), .ZN(n13951) );
  NOR2_X1 U14363 ( .A1(n11695), .A2(n11689), .ZN(n12767) );
  NAND2_X1 U14364 ( .A1(n13956), .A2(n11686), .ZN(n13934) );
  INV_X1 U14365 ( .A(n21900), .ZN(n21924) );
  NAND2_X1 U14366 ( .A1(n21924), .A2(n12768), .ZN(n21277) );
  NAND2_X1 U14367 ( .A1(n21277), .A2(n21655), .ZN(n12769) );
  NAND2_X1 U14368 ( .A1(n21655), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16877) );
  NAND2_X1 U14369 ( .A1(n14439), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12770) );
  AND2_X1 U14370 ( .A1(n16877), .A2(n12770), .ZN(n14177) );
  INV_X1 U14371 ( .A(n14177), .ZN(n12771) );
  INV_X2 U14372 ( .A(n15898), .ZN(n20014) );
  NOR2_X1 U14373 ( .A1(n21419), .A2(n19891), .ZN(n15954) );
  AOI21_X1 U14374 ( .B1(n20014), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15954), .ZN(n12772) );
  OAI21_X1 U14375 ( .B1(n20024), .B2(n14595), .A(n12772), .ZN(n12773) );
  AOI21_X1 U14376 ( .B1(n12774), .B2(n20021), .A(n12773), .ZN(n12888) );
  INV_X1 U14377 ( .A(n12775), .ZN(n14379) );
  AND2_X1 U14378 ( .A1(n11680), .A2(n11685), .ZN(n13930) );
  NAND2_X1 U14379 ( .A1(n14379), .A2(n13930), .ZN(n12780) );
  INV_X1 U14380 ( .A(n21274), .ZN(n14068) );
  NAND2_X1 U14381 ( .A1(n11686), .A2(n12777), .ZN(n12792) );
  OAI21_X1 U14382 ( .B1(n14068), .B2(n12790), .A(n12792), .ZN(n12778) );
  INV_X1 U14383 ( .A(n12778), .ZN(n12779) );
  NAND2_X1 U14384 ( .A1(n12780), .A2(n12779), .ZN(n14047) );
  INV_X1 U14385 ( .A(n13930), .ZN(n12843) );
  OR2_X1 U14386 ( .A1(n11754), .A2(n12843), .ZN(n12784) );
  XNOR2_X1 U14387 ( .A(n12790), .B(n12789), .ZN(n12781) );
  OAI211_X1 U14388 ( .C1(n12781), .C2(n14068), .A(n13935), .B(n11680), .ZN(
        n12782) );
  INV_X1 U14389 ( .A(n12782), .ZN(n12783) );
  NAND2_X1 U14390 ( .A1(n12784), .A2(n12783), .ZN(n12785) );
  INV_X1 U14391 ( .A(n12785), .ZN(n12786) );
  OR2_X1 U14392 ( .A1(n14049), .A2(n12786), .ZN(n12787) );
  XNOR2_X1 U14393 ( .A(n12797), .B(n21300), .ZN(n14306) );
  NAND2_X1 U14394 ( .A1(n10975), .A2(n13930), .ZN(n12796) );
  NAND2_X1 U14395 ( .A1(n12790), .A2(n12789), .ZN(n12801) );
  INV_X1 U14396 ( .A(n12791), .ZN(n12800) );
  XNOR2_X1 U14397 ( .A(n12801), .B(n12800), .ZN(n12794) );
  INV_X1 U14398 ( .A(n12792), .ZN(n12793) );
  AOI21_X1 U14399 ( .B1(n12794), .B2(n21274), .A(n12793), .ZN(n12795) );
  NAND2_X1 U14400 ( .A1(n12796), .A2(n12795), .ZN(n14305) );
  NAND2_X1 U14401 ( .A1(n12797), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12798) );
  NAND2_X1 U14402 ( .A1(n12799), .A2(n13930), .ZN(n12805) );
  NAND2_X1 U14403 ( .A1(n12801), .A2(n12800), .ZN(n12802) );
  NAND2_X1 U14404 ( .A1(n12802), .A2(n12803), .ZN(n12817) );
  OAI211_X1 U14405 ( .C1(n12803), .C2(n12802), .A(n12817), .B(n21274), .ZN(
        n12804) );
  NAND2_X1 U14406 ( .A1(n12805), .A2(n12804), .ZN(n14613) );
  NAND2_X1 U14407 ( .A1(n12806), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14610) );
  NAND2_X1 U14408 ( .A1(n12807), .A2(n14610), .ZN(n19949) );
  NAND2_X1 U14409 ( .A1(n12808), .A2(n13930), .ZN(n12811) );
  XNOR2_X1 U14410 ( .A(n12817), .B(n12815), .ZN(n12809) );
  NAND2_X1 U14411 ( .A1(n12809), .A2(n21274), .ZN(n12810) );
  NAND2_X1 U14412 ( .A1(n12811), .A2(n12810), .ZN(n12813) );
  XNOR2_X1 U14413 ( .A(n12813), .B(n12812), .ZN(n19948) );
  NAND2_X1 U14414 ( .A1(n19949), .A2(n19948), .ZN(n19947) );
  NAND2_X1 U14415 ( .A1(n12813), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12814) );
  INV_X1 U14416 ( .A(n12815), .ZN(n12816) );
  OR2_X1 U14417 ( .A1(n12817), .A2(n12816), .ZN(n12825) );
  XNOR2_X1 U14418 ( .A(n12825), .B(n12826), .ZN(n12818) );
  NAND2_X1 U14419 ( .A1(n12818), .A2(n21274), .ZN(n12819) );
  OAI21_X1 U14420 ( .B1(n12820), .B2(n12843), .A(n12819), .ZN(n12821) );
  XNOR2_X1 U14421 ( .A(n12821), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14684) );
  OR2_X1 U14422 ( .A1(n12821), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12822) );
  NAND3_X1 U14423 ( .A1(n12823), .A2(n13930), .A3(n12824), .ZN(n12830) );
  INV_X1 U14424 ( .A(n12825), .ZN(n12827) );
  NAND2_X1 U14425 ( .A1(n12827), .A2(n12826), .ZN(n12834) );
  XNOR2_X1 U14426 ( .A(n12834), .B(n12835), .ZN(n12828) );
  NAND2_X1 U14427 ( .A1(n12828), .A2(n21274), .ZN(n12829) );
  NAND2_X1 U14428 ( .A1(n12830), .A2(n12829), .ZN(n12831) );
  XNOR2_X1 U14429 ( .A(n12831), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19960) );
  NAND2_X1 U14430 ( .A1(n12831), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12832) );
  NAND2_X1 U14431 ( .A1(n19957), .A2(n12832), .ZN(n19965) );
  NAND2_X1 U14432 ( .A1(n12833), .A2(n13930), .ZN(n12839) );
  INV_X1 U14433 ( .A(n12834), .ZN(n12836) );
  NAND2_X1 U14434 ( .A1(n12836), .A2(n12835), .ZN(n12848) );
  XNOR2_X1 U14435 ( .A(n12848), .B(n12846), .ZN(n12837) );
  NAND2_X1 U14436 ( .A1(n12837), .A2(n21274), .ZN(n12838) );
  NAND2_X1 U14437 ( .A1(n12839), .A2(n12838), .ZN(n12840) );
  XNOR2_X1 U14438 ( .A(n12840), .B(n21334), .ZN(n19964) );
  NAND2_X1 U14439 ( .A1(n19965), .A2(n19964), .ZN(n19963) );
  NAND2_X1 U14440 ( .A1(n12840), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12841) );
  INV_X1 U14441 ( .A(n12842), .ZN(n12844) );
  NOR2_X1 U14442 ( .A1(n12844), .A2(n12843), .ZN(n12845) );
  NAND2_X2 U14443 ( .A1(n12823), .A2(n12845), .ZN(n12852) );
  NAND2_X1 U14444 ( .A1(n21274), .A2(n12846), .ZN(n12847) );
  OR2_X1 U14445 ( .A1(n12848), .A2(n12847), .ZN(n12849) );
  NAND2_X1 U14446 ( .A1(n12852), .A2(n12849), .ZN(n12850) );
  INV_X1 U14447 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21340) );
  XNOR2_X1 U14448 ( .A(n12850), .B(n21340), .ZN(n15089) );
  OR2_X1 U14449 ( .A1(n12850), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12851) );
  XNOR2_X1 U14450 ( .A(n19971), .B(n15933), .ZN(n15225) );
  NAND2_X1 U14451 ( .A1(n19971), .A2(n21282), .ZN(n12855) );
  NAND2_X1 U14452 ( .A1(n19983), .A2(n12855), .ZN(n15914) );
  INV_X1 U14453 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12861) );
  NAND2_X1 U14454 ( .A1(n19971), .A2(n12861), .ZN(n15913) );
  NAND2_X1 U14455 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12856) );
  NAND2_X1 U14456 ( .A1(n19971), .A2(n12856), .ZN(n15911) );
  NAND2_X1 U14457 ( .A1(n15913), .A2(n15911), .ZN(n12857) );
  INV_X1 U14458 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21287) );
  AND2_X1 U14459 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16046) );
  NAND2_X1 U14460 ( .A1(n16046), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16040) );
  NAND2_X1 U14461 ( .A1(n19971), .A2(n16040), .ZN(n12859) );
  NOR2_X1 U14462 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12860) );
  NAND2_X1 U14463 ( .A1(n15909), .A2(n15912), .ZN(n15888) );
  NOR2_X1 U14464 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12862) );
  NOR2_X1 U14465 ( .A1(n19971), .A2(n12862), .ZN(n12863) );
  NOR2_X1 U14466 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21392) );
  AND2_X1 U14467 ( .A1(n21392), .A2(n15896), .ZN(n12864) );
  NOR2_X1 U14468 ( .A1(n19971), .A2(n12864), .ZN(n12865) );
  NOR2_X1 U14469 ( .A1(n15902), .A2(n12865), .ZN(n12866) );
  AND2_X1 U14470 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21405) );
  NAND2_X1 U14471 ( .A1(n21405), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21408) );
  INV_X1 U14472 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16041) );
  NOR2_X1 U14473 ( .A1(n21408), .A2(n16041), .ZN(n12867) );
  NAND2_X1 U14474 ( .A1(n12868), .A2(n19971), .ZN(n20008) );
  NAND2_X1 U14475 ( .A1(n20008), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12871) );
  NOR2_X1 U14476 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21398) );
  NAND3_X1 U14477 ( .A1(n21398), .A2(n12869), .A3(n16041), .ZN(n12870) );
  OAI21_X1 U14478 ( .B1(n15868), .B2(n12870), .A(n19993), .ZN(n20009) );
  INV_X1 U14479 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21429) );
  INV_X1 U14480 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16011) );
  NAND3_X1 U14481 ( .A1(n21429), .A2(n15939), .A3(n16011), .ZN(n15827) );
  NAND2_X1 U14482 ( .A1(n12871), .A2(n19971), .ZN(n15854) );
  NOR2_X1 U14483 ( .A1(n21429), .A2(n15939), .ZN(n15951) );
  AND2_X1 U14484 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n15951), .ZN(
        n15943) );
  INV_X1 U14485 ( .A(n15943), .ZN(n12872) );
  NAND2_X1 U14486 ( .A1(n19971), .A2(n12872), .ZN(n15848) );
  NAND3_X1 U14487 ( .A1(n15854), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15848), .ZN(n12873) );
  NOR2_X1 U14488 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15981) );
  NOR2_X1 U14489 ( .A1(n20015), .A2(n15981), .ZN(n12874) );
  AND2_X1 U14490 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15980) );
  INV_X1 U14491 ( .A(n15980), .ZN(n12875) );
  INV_X1 U14492 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15969) );
  NAND2_X1 U14493 ( .A1(n19971), .A2(n15969), .ZN(n15816) );
  INV_X1 U14494 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15946) );
  XNOR2_X1 U14495 ( .A(n20015), .B(n15946), .ZN(n12879) );
  INV_X1 U14496 ( .A(n12879), .ZN(n12877) );
  INV_X1 U14497 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15952) );
  NAND2_X1 U14498 ( .A1(n19971), .A2(n15952), .ZN(n12881) );
  NAND2_X1 U14499 ( .A1(n12877), .A2(n12881), .ZN(n12885) );
  NAND2_X1 U14500 ( .A1(n19993), .A2(n11404), .ZN(n12878) );
  AND2_X1 U14501 ( .A1(n12879), .A2(n12878), .ZN(n12880) );
  OR2_X1 U14502 ( .A1(n20015), .A2(n15969), .ZN(n15820) );
  OAI211_X1 U14503 ( .C1(n20015), .C2(n15952), .A(n15820), .B(n12881), .ZN(
        n12882) );
  NAND2_X1 U14504 ( .A1(n12882), .A2(n15946), .ZN(n12883) );
  OAI211_X1 U14505 ( .C1(n15817), .C2(n12885), .A(n12884), .B(n12883), .ZN(
        n15958) );
  INV_X1 U14506 ( .A(n15958), .ZN(n12886) );
  NAND2_X1 U14507 ( .A1(n12888), .A2(n12887), .ZN(P1_U2968) );
  NAND2_X1 U14508 ( .A1(n12890), .A2(n12889), .ZN(n17911) );
  INV_X1 U14509 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21074) );
  INV_X1 U14510 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21075) );
  OAI33_X1 U14511 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n17911), .B1(n21074), .B2(
        n17910), .B3(n21075), .ZN(n12892) );
  XNOR2_X1 U14512 ( .A(n12892), .B(n12891), .ZN(n17891) );
  NAND2_X1 U14513 ( .A1(n17891), .A2(n21194), .ZN(n12908) );
  NOR2_X1 U14514 ( .A1(n12900), .A2(n21075), .ZN(n17903) );
  INV_X1 U14515 ( .A(n17903), .ZN(n12897) );
  NAND2_X1 U14516 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n21062), .ZN(
        n12893) );
  XOR2_X1 U14517 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12893), .Z(
        n17888) );
  NAND2_X1 U14518 ( .A1(n21078), .A2(n21111), .ZN(n20921) );
  NOR2_X1 U14519 ( .A1(n21034), .A2(n12897), .ZN(n21064) );
  NAND2_X1 U14520 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n21064), .ZN(
        n12894) );
  XOR2_X1 U14521 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12894), .Z(
        n17894) );
  NOR2_X1 U14522 ( .A1(n21044), .A2(n12900), .ZN(n12895) );
  AOI21_X1 U14523 ( .B1(n21013), .B2(n12895), .A(n21162), .ZN(n21065) );
  AOI211_X1 U14524 ( .C1(n21153), .C2(n12897), .A(n21065), .B(n12896), .ZN(
        n12899) );
  NAND3_X1 U14525 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n12899), .A3(
        n12898), .ZN(n21080) );
  NAND3_X1 U14526 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21153), .A3(
        n21080), .ZN(n12902) );
  NOR4_X1 U14527 ( .A1(n21020), .A2(n21019), .A3(n21044), .A4(n12900), .ZN(
        n21060) );
  NAND4_X1 U14528 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n21060), .A4(n12891), .ZN(
        n12901) );
  OAI211_X1 U14529 ( .C1(n17894), .C2(n21063), .A(n12902), .B(n12901), .ZN(
        n12903) );
  INV_X1 U14530 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18208) );
  NOR2_X1 U14531 ( .A1(n10961), .A2(n18208), .ZN(n17887) );
  AOI21_X1 U14532 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21092), .A(
        n17887), .ZN(n12904) );
  INV_X1 U14533 ( .A(n12906), .ZN(n12907) );
  NAND2_X1 U14534 ( .A1(n12908), .A2(n12907), .ZN(P3_U2831) );
  AOI22_X1 U14535 ( .A1(n13396), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12913) );
  AOI22_X1 U14536 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12912) );
  AOI22_X1 U14537 ( .A1(n13134), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12911) );
  AND2_X2 U14538 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13125) );
  AND2_X4 U14539 ( .A1(n13125), .A2(n14481), .ZN(n13135) );
  AND2_X4 U14540 ( .A1(n13125), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13136) );
  NAND4_X1 U14541 ( .A1(n12913), .A2(n12912), .A3(n12911), .A4(n12910), .ZN(
        n12914) );
  AOI22_X1 U14542 ( .A1(n13476), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U14543 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U14544 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12915) );
  NAND4_X1 U14545 ( .A1(n12918), .A2(n12917), .A3(n12916), .A4(n12915), .ZN(
        n12919) );
  INV_X2 U14546 ( .A(n13462), .ZN(n13339) );
  AOI22_X1 U14547 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12923) );
  AOI22_X1 U14548 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12922) );
  AOI22_X1 U14549 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U14550 ( .A1(n13476), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U14551 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12926) );
  AOI22_X1 U14552 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12925) );
  AOI22_X1 U14553 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12924) );
  XNOR2_X1 U14554 ( .A(n13799), .B(n13579), .ZN(n13905) );
  AOI22_X1 U14555 ( .A1(n13396), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U14556 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12930) );
  AOI22_X1 U14557 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12929) );
  AOI22_X1 U14558 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U14559 ( .A1(n13396), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12936) );
  AOI22_X1 U14560 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U14561 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12934) );
  AOI22_X1 U14562 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12933) );
  NAND2_X2 U14563 ( .A1(n12939), .A2(n12938), .ZN(n12992) );
  AOI22_X1 U14564 ( .A1(n13476), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U14565 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13142), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U14566 ( .A1(n13134), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12941) );
  AOI22_X1 U14567 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12940) );
  NAND4_X1 U14568 ( .A1(n12943), .A2(n12942), .A3(n12941), .A4(n12940), .ZN(
        n12944) );
  NAND2_X1 U14569 ( .A1(n12944), .A2(n13511), .ZN(n12951) );
  AOI22_X1 U14570 ( .A1(n13396), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U14571 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U14572 ( .A1(n13134), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U14573 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12945) );
  NAND4_X1 U14574 ( .A1(n12948), .A2(n12947), .A3(n12946), .A4(n12945), .ZN(
        n12949) );
  NAND2_X1 U14575 ( .A1(n12949), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12950) );
  INV_X1 U14576 ( .A(n13011), .ZN(n13597) );
  AOI22_X1 U14577 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U14578 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12956) );
  AOI22_X1 U14579 ( .A1(n13396), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12955) );
  AOI22_X1 U14580 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12954) );
  NAND4_X1 U14581 ( .A1(n12957), .A2(n12956), .A3(n12955), .A4(n12954), .ZN(
        n12963) );
  AOI22_X1 U14582 ( .A1(n13396), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12960) );
  AOI22_X1 U14583 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U14584 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12958) );
  NAND4_X1 U14585 ( .A1(n12961), .A2(n12960), .A3(n12959), .A4(n12958), .ZN(
        n12962) );
  AND2_X2 U14586 ( .A1(n12965), .A2(n11393), .ZN(n13041) );
  AOI22_X1 U14587 ( .A1(n13476), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U14588 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U14589 ( .A1(n13134), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U14590 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12967) );
  NAND4_X1 U14591 ( .A1(n12970), .A2(n12969), .A3(n12968), .A4(n12967), .ZN(
        n12971) );
  NAND2_X1 U14592 ( .A1(n12971), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12978) );
  AOI22_X1 U14593 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12975) );
  AOI22_X1 U14594 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12974) );
  AOI22_X1 U14595 ( .A1(n13396), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12973) );
  NAND4_X1 U14596 ( .A1(n12975), .A2(n12974), .A3(n12973), .A4(n12972), .ZN(
        n12976) );
  NAND2_X1 U14597 ( .A1(n12976), .A2(n13511), .ZN(n12977) );
  AOI22_X1 U14598 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12982) );
  AOI22_X1 U14599 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12981) );
  AOI22_X1 U14600 ( .A1(n13476), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12980) );
  AOI22_X1 U14601 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12979) );
  NAND4_X1 U14602 ( .A1(n12982), .A2(n12981), .A3(n12980), .A4(n12979), .ZN(
        n12983) );
  AOI22_X1 U14603 ( .A1(n13134), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U14604 ( .A1(n13476), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U14605 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U14606 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12984) );
  NAND4_X1 U14607 ( .A1(n12987), .A2(n12986), .A3(n12985), .A4(n12984), .ZN(
        n12988) );
  NAND2_X2 U14608 ( .A1(n12990), .A2(n12989), .ZN(n14727) );
  NOR2_X2 U14609 ( .A1(n13783), .A2(n12992), .ZN(n13901) );
  NAND2_X1 U14610 ( .A1(n12992), .A2(n12991), .ZN(n13014) );
  INV_X1 U14611 ( .A(n13014), .ZN(n13005) );
  AOI22_X1 U14612 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U14613 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12995) );
  AOI22_X1 U14614 ( .A1(n13476), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U14615 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U14616 ( .A1(n13339), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13128), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U14617 ( .A1(n13142), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U14618 ( .A1(n13396), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13141), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U14619 ( .A1(n13135), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13136), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12998) );
  NAND2_X1 U14620 ( .A1(n13002), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13003) );
  OR2_X2 U14621 ( .A1(n13008), .A2(n13006), .ZN(n13583) );
  NAND2_X1 U14622 ( .A1(n13799), .A2(n13579), .ZN(n13016) );
  NAND2_X1 U14623 ( .A1(n13016), .A2(n19534), .ZN(n13007) );
  OAI21_X1 U14624 ( .B1(n13008), .B2(n13007), .A(n19642), .ZN(n13009) );
  INV_X1 U14625 ( .A(n13009), .ZN(n13010) );
  INV_X1 U14626 ( .A(n13041), .ZN(n13013) );
  AND2_X1 U14627 ( .A1(n13011), .A2(n10967), .ZN(n13012) );
  NAND2_X1 U14628 ( .A1(n13013), .A2(n13012), .ZN(n13054) );
  NAND2_X1 U14629 ( .A1(n19534), .A2(n14142), .ZN(n13018) );
  NAND2_X1 U14630 ( .A1(n13020), .A2(n13019), .ZN(n13030) );
  NAND2_X1 U14631 ( .A1(n14714), .A2(n15263), .ZN(n18595) );
  NAND2_X1 U14632 ( .A1(n19642), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13029) );
  AND2_X1 U14633 ( .A1(n19642), .A2(n13799), .ZN(n13026) );
  NAND3_X1 U14634 ( .A1(n13026), .A2(n14136), .A3(n13025), .ZN(n14114) );
  INV_X1 U14635 ( .A(n14114), .ZN(n13027) );
  NAND2_X1 U14636 ( .A1(n13027), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13028) );
  INV_X1 U14637 ( .A(n13038), .ZN(n13033) );
  INV_X1 U14638 ( .A(n13030), .ZN(n13032) );
  OAI211_X1 U14639 ( .C1(n18595), .C2(n19260), .A(n13033), .B(n13812), .ZN(
        n13034) );
  NAND2_X1 U14640 ( .A1(n13036), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13061) );
  OR2_X4 U14641 ( .A1(n13812), .A2(n19585), .ZN(n15300) );
  INV_X1 U14642 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n13869) );
  INV_X1 U14643 ( .A(n13837), .ZN(n13040) );
  NAND2_X1 U14644 ( .A1(n13108), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n13043) );
  NAND2_X1 U14645 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13042) );
  NOR2_X1 U14646 ( .A1(n13045), .A2(n13044), .ZN(n13046) );
  OR2_X2 U14647 ( .A1(n13047), .A2(n13046), .ZN(n13097) );
  NAND2_X1 U14648 ( .A1(n13047), .A2(n13046), .ZN(n13099) );
  INV_X1 U14649 ( .A(n13090), .ZN(n13065) );
  INV_X1 U14650 ( .A(n13048), .ZN(n14320) );
  NAND2_X1 U14651 ( .A1(n10965), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13059) );
  INV_X1 U14652 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18240) );
  NAND2_X1 U14653 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13049) );
  NAND2_X1 U14654 ( .A1(n18595), .A2(n13049), .ZN(n13050) );
  AOI21_X1 U14655 ( .B1(n13108), .B2(P2_EBX_REG_0__SCAN_IN), .A(n13050), .ZN(
        n13052) );
  OAI211_X1 U14656 ( .C1(n15300), .C2(n18240), .A(n13052), .B(n13051), .ZN(
        n13053) );
  INV_X1 U14657 ( .A(n13053), .ZN(n13058) );
  NAND2_X1 U14658 ( .A1(n11024), .A2(n13054), .ZN(n14125) );
  NAND3_X1 U14659 ( .A1(n13059), .A2(n13058), .A3(n13057), .ZN(n13085) );
  NAND2_X1 U14660 ( .A1(n15264), .A2(n14490), .ZN(n13060) );
  INV_X1 U14661 ( .A(n18595), .ZN(n13105) );
  NAND2_X1 U14662 ( .A1(n13105), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13062) );
  NAND2_X1 U14663 ( .A1(n13064), .A2(n13063), .ZN(n13086) );
  NAND2_X1 U14664 ( .A1(n13085), .A2(n13086), .ZN(n13098) );
  NAND2_X1 U14665 ( .A1(n13065), .A2(n13098), .ZN(n14979) );
  NAND2_X1 U14666 ( .A1(n14979), .A2(n13099), .ZN(n13077) );
  OAI21_X1 U14667 ( .B1(n19256), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15263), 
        .ZN(n13066) );
  INV_X1 U14668 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n18577) );
  NAND2_X1 U14669 ( .A1(n15285), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n13068) );
  NAND2_X1 U14670 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13067) );
  NAND2_X1 U14671 ( .A1(n13073), .A2(n13072), .ZN(n13102) );
  INV_X1 U14672 ( .A(n13073), .ZN(n13074) );
  XNOR2_X2 U14673 ( .A(n13077), .B(n13076), .ZN(n14995) );
  NAND2_X1 U14674 ( .A1(n14714), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14557) );
  INV_X1 U14675 ( .A(n14557), .ZN(n13087) );
  NAND2_X1 U14676 ( .A1(n15005), .A2(n13087), .ZN(n13081) );
  NAND2_X1 U14677 ( .A1(n13799), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13078) );
  NAND2_X1 U14678 ( .A1(n13078), .A2(n17222), .ZN(n13114) );
  AND2_X1 U14679 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19192) );
  NAND2_X1 U14680 ( .A1(n19192), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13111) );
  INV_X1 U14681 ( .A(n19192), .ZN(n19257) );
  NAND2_X1 U14682 ( .A1(n19257), .A2(n19256), .ZN(n13079) );
  AND2_X1 U14683 ( .A1(n13111), .A2(n13079), .ZN(n19148) );
  AOI22_X1 U14684 ( .A1(n13114), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19304), .B2(n19148), .ZN(n13080) );
  NAND2_X1 U14685 ( .A1(n13081), .A2(n13080), .ZN(n13084) );
  NAND2_X1 U14686 ( .A1(n13082), .A2(n13035), .ZN(n13387) );
  INV_X1 U14687 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19574) );
  NOR2_X1 U14688 ( .A1(n13387), .A2(n19574), .ZN(n13083) );
  AOI22_X1 U14689 ( .A1(n13114), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19304), .B2(n19288), .ZN(n13088) );
  NAND2_X1 U14690 ( .A1(n13445), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13093) );
  NAND2_X1 U14691 ( .A1(n19288), .A2(n19260), .ZN(n19303) );
  NAND2_X1 U14692 ( .A1(n19257), .A2(n19303), .ZN(n19217) );
  NOR2_X1 U14693 ( .A1(n19217), .A2(n19290), .ZN(n19272) );
  AOI21_X1 U14694 ( .B1(n13114), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19272), .ZN(n13091) );
  NAND2_X1 U14695 ( .A1(n14169), .A2(n14168), .ZN(n13096) );
  INV_X1 U14696 ( .A(n13964), .ZN(n13094) );
  NAND2_X1 U14697 ( .A1(n13094), .A2(n13093), .ZN(n13095) );
  NAND3_X1 U14698 ( .A1(n13098), .A2(n13100), .A3(n13097), .ZN(n13104) );
  INV_X1 U14699 ( .A(n13099), .ZN(n13101) );
  NAND2_X1 U14700 ( .A1(n13101), .A2(n13100), .ZN(n13103) );
  NAND2_X1 U14701 ( .A1(n13105), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13106) );
  INV_X1 U14702 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13662) );
  NAND2_X1 U14703 ( .A1(n10965), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13110) );
  AOI22_X1 U14704 ( .A1(n15556), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13109) );
  OAI211_X1 U14705 ( .C1(n15300), .C2(n13662), .A(n13110), .B(n13109), .ZN(
        n14326) );
  AOI21_X1 U14706 ( .B1(n13111), .B2(n19255), .A(n19290), .ZN(n13113) );
  INV_X1 U14707 ( .A(n13111), .ZN(n13112) );
  NAND2_X1 U14708 ( .A1(n13112), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19111) );
  AOI22_X1 U14709 ( .A1(n13114), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13113), .B2(n19111), .ZN(n13115) );
  NAND2_X1 U14710 ( .A1(n13445), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13117) );
  NAND2_X1 U14711 ( .A1(n13118), .A2(n13117), .ZN(n13119) );
  NAND2_X1 U14712 ( .A1(n13799), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13120) );
  INV_X1 U14713 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19469) );
  NOR2_X1 U14714 ( .A1(n13387), .A2(n19469), .ZN(n14338) );
  INV_X1 U14715 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19369) );
  INV_X1 U14716 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19320) );
  AND2_X1 U14717 ( .A1(n14487), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13124) );
  AOI22_X1 U14718 ( .A1(n13599), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13155), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13132) );
  AND2_X1 U14719 ( .A1(n14490), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13126) );
  AOI22_X1 U14720 ( .A1(n13600), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13131) );
  NAND2_X1 U14721 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13130) );
  NAND2_X1 U14722 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13129) );
  AND4_X1 U14723 ( .A1(n13132), .A2(n13131), .A3(n13130), .A4(n13129), .ZN(
        n13140) );
  INV_X1 U14724 ( .A(n13457), .ZN(n13133) );
  AND2_X2 U14725 ( .A1(n10979), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13606) );
  AOI22_X1 U14726 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13605), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13139) );
  INV_X1 U14727 ( .A(n13136), .ZN(n14505) );
  INV_X1 U14728 ( .A(n14505), .ZN(n13137) );
  AOI22_X1 U14729 ( .A1(n13301), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13138) );
  NAND3_X1 U14730 ( .A1(n13140), .A2(n13139), .A3(n13138), .ZN(n13151) );
  AND2_X2 U14731 ( .A1(n13495), .A2(n13511), .ZN(n13705) );
  AOI22_X1 U14732 ( .A1(n10957), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13149) );
  INV_X1 U14733 ( .A(n13142), .ZN(n13340) );
  AND2_X1 U14734 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13145) );
  AOI22_X1 U14735 ( .A1(n13525), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13706), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13148) );
  AND2_X2 U14736 ( .A1(n13492), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13834) );
  AOI22_X1 U14737 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13147) );
  NAND3_X1 U14738 ( .A1(n13149), .A2(n13148), .A3(n13147), .ZN(n13150) );
  NAND2_X1 U14739 ( .A1(n14681), .A2(n14680), .ZN(n14679) );
  AOI22_X1 U14740 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10958), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13154) );
  AOI22_X1 U14741 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n13706), .ZN(n13153) );
  AOI22_X1 U14742 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n13525), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13152) );
  AND3_X1 U14743 ( .A1(n13154), .A2(n13153), .A3(n13152), .ZN(n13168) );
  AOI22_X1 U14744 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13155), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13160) );
  AOI22_X1 U14745 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13600), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13159) );
  NAND2_X1 U14746 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13158) );
  NAND2_X1 U14747 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13157) );
  NAND4_X1 U14748 ( .A1(n13160), .A2(n13159), .A3(n13158), .A4(n13157), .ZN(
        n13166) );
  NAND2_X1 U14749 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13164) );
  NAND2_X1 U14750 ( .A1(n13605), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13163) );
  NAND2_X1 U14751 ( .A1(n13301), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13162) );
  NAND2_X1 U14752 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13161) );
  NAND4_X1 U14753 ( .A1(n13164), .A2(n13163), .A3(n13162), .A4(n13161), .ZN(
        n13165) );
  NOR2_X1 U14754 ( .A1(n13166), .A2(n13165), .ZN(n13167) );
  AOI22_X1 U14755 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n13705), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13172) );
  AOI22_X1 U14756 ( .A1(n13707), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n13706), .ZN(n13171) );
  AOI22_X1 U14757 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n13525), .B1(
        n13834), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13170) );
  AND3_X1 U14758 ( .A1(n13172), .A2(n13171), .A3(n13170), .ZN(n13184) );
  AOI22_X1 U14759 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13155), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13176) );
  AOI22_X1 U14760 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n13600), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13175) );
  NAND2_X1 U14761 ( .A1(n13605), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13174) );
  NAND2_X1 U14762 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13173) );
  NAND4_X1 U14763 ( .A1(n13176), .A2(n13175), .A3(n13174), .A4(n13173), .ZN(
        n13182) );
  NAND2_X1 U14764 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13180) );
  NAND2_X1 U14765 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13179) );
  NAND2_X1 U14766 ( .A1(n10957), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13178) );
  NAND2_X1 U14767 ( .A1(n13301), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13177) );
  NAND4_X1 U14768 ( .A1(n13180), .A2(n13179), .A3(n13178), .A4(n13177), .ZN(
        n13181) );
  NOR2_X1 U14769 ( .A1(n13182), .A2(n13181), .ZN(n13183) );
  AOI22_X1 U14770 ( .A1(n13600), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13188) );
  NAND2_X1 U14771 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n13187) );
  NAND2_X1 U14772 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n13186) );
  AOI22_X1 U14773 ( .A1(n13598), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13706), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13185) );
  AND4_X1 U14774 ( .A1(n13188), .A2(n13187), .A3(n13186), .A4(n13185), .ZN(
        n13191) );
  AOI22_X1 U14775 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13605), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U14776 ( .A1(n13301), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13189) );
  NAND3_X1 U14777 ( .A1(n13191), .A2(n13190), .A3(n13189), .ZN(n13196) );
  AOI22_X1 U14778 ( .A1(n10958), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U14779 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13155), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13193) );
  AOI22_X1 U14780 ( .A1(n13525), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13192) );
  NAND3_X1 U14781 ( .A1(n13194), .A2(n13193), .A3(n13192), .ZN(n13195) );
  OR2_X1 U14782 ( .A1(n13196), .A2(n13195), .ZN(n14921) );
  AOI22_X1 U14783 ( .A1(n13598), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13155), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13200) );
  AOI22_X1 U14784 ( .A1(n13600), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13199) );
  NAND2_X1 U14785 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13198) );
  NAND2_X1 U14786 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13197) );
  AND4_X1 U14787 ( .A1(n13200), .A2(n13199), .A3(n13198), .A4(n13197), .ZN(
        n13203) );
  AOI22_X1 U14788 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13605), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13202) );
  AOI22_X1 U14789 ( .A1(n13301), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13201) );
  NAND3_X1 U14790 ( .A1(n13203), .A2(n13202), .A3(n13201), .ZN(n13208) );
  AOI22_X1 U14791 ( .A1(n10957), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13206) );
  AOI22_X1 U14792 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13706), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U14793 ( .A1(n13525), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13204) );
  NAND3_X1 U14794 ( .A1(n13206), .A2(n13205), .A3(n13204), .ZN(n13207) );
  OR2_X1 U14795 ( .A1(n13208), .A2(n13207), .ZN(n14896) );
  AOI22_X1 U14796 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13155), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13212) );
  AOI22_X1 U14797 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13600), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13211) );
  NAND2_X1 U14798 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n13210) );
  NAND2_X1 U14799 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n13209) );
  AND4_X1 U14800 ( .A1(n13212), .A2(n13211), .A3(n13210), .A4(n13209), .ZN(
        n13215) );
  AOI22_X1 U14801 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n13606), .B1(
        n13605), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U14802 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n13301), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13213) );
  NAND3_X1 U14803 ( .A1(n13215), .A2(n13214), .A3(n13213), .ZN(n13220) );
  AOI22_X1 U14804 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10958), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13218) );
  AOI22_X1 U14805 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n13706), .ZN(n13217) );
  AOI22_X1 U14806 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n13525), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13216) );
  NAND3_X1 U14807 ( .A1(n13218), .A2(n13217), .A3(n13216), .ZN(n13219) );
  OR2_X1 U14808 ( .A1(n13220), .A2(n13219), .ZN(n14948) );
  AOI22_X1 U14809 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13155), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13224) );
  AOI22_X1 U14810 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13600), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13223) );
  NAND2_X1 U14811 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13222) );
  NAND2_X1 U14812 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13221) );
  AND4_X1 U14813 ( .A1(n13224), .A2(n13223), .A3(n13222), .A4(n13221), .ZN(
        n13227) );
  AOI22_X1 U14814 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13271), .B1(
        n13605), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13226) );
  AOI22_X1 U14815 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n13301), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13225) );
  NAND3_X1 U14816 ( .A1(n13227), .A2(n13226), .A3(n13225), .ZN(n13232) );
  AOI22_X1 U14817 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10958), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13230) );
  AOI22_X1 U14818 ( .A1(n13525), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n13706), .ZN(n13229) );
  AOI22_X1 U14819 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13707), .B1(
        n13834), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13228) );
  NAND3_X1 U14820 ( .A1(n13230), .A2(n13229), .A3(n13228), .ZN(n13231) );
  OR2_X1 U14821 ( .A1(n13232), .A2(n13231), .ZN(n14947) );
  AND2_X1 U14822 ( .A1(n14948), .A2(n14947), .ZN(n14894) );
  AND2_X1 U14823 ( .A1(n14896), .A2(n14894), .ZN(n14895) );
  AND2_X1 U14824 ( .A1(n14921), .A2(n14895), .ZN(n13233) );
  AOI22_X1 U14825 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13155), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13237) );
  AOI22_X1 U14826 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13600), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13236) );
  NAND2_X1 U14827 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13235) );
  NAND2_X1 U14828 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n13234) );
  AND4_X1 U14829 ( .A1(n13237), .A2(n13236), .A3(n13235), .A4(n13234), .ZN(
        n13240) );
  AOI22_X1 U14830 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n13606), .B1(
        n13605), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13239) );
  AOI22_X1 U14831 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n13301), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13238) );
  NAND3_X1 U14832 ( .A1(n13240), .A2(n13239), .A3(n13238), .ZN(n13245) );
  AOI22_X1 U14833 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10958), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U14834 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n13706), .ZN(n13242) );
  AOI22_X1 U14835 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n13525), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13241) );
  NAND3_X1 U14836 ( .A1(n13243), .A2(n13242), .A3(n13241), .ZN(n13244) );
  OR2_X1 U14837 ( .A1(n13245), .A2(n13244), .ZN(n14965) );
  AOI22_X1 U14838 ( .A1(n13598), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13155), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13249) );
  AOI22_X1 U14839 ( .A1(n13600), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13248) );
  NAND2_X1 U14840 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13247) );
  NAND2_X1 U14841 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13246) );
  AND4_X1 U14842 ( .A1(n13249), .A2(n13248), .A3(n13247), .A4(n13246), .ZN(
        n13252) );
  AOI22_X1 U14843 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13605), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13251) );
  AOI22_X1 U14844 ( .A1(n13301), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13250) );
  NAND3_X1 U14845 ( .A1(n13252), .A2(n13251), .A3(n13250), .ZN(n13257) );
  AOI22_X1 U14846 ( .A1(n10958), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13255) );
  AOI22_X1 U14847 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13706), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13254) );
  AOI22_X1 U14848 ( .A1(n13525), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13253) );
  NAND3_X1 U14849 ( .A1(n13255), .A2(n13254), .A3(n13253), .ZN(n13256) );
  NOR2_X1 U14850 ( .A1(n13257), .A2(n13256), .ZN(n15182) );
  INV_X1 U14851 ( .A(n15182), .ZN(n13258) );
  AOI22_X1 U14852 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13155), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13262) );
  AOI22_X1 U14853 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13600), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13261) );
  NAND2_X1 U14854 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13260) );
  NAND2_X1 U14855 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13259) );
  AND4_X1 U14856 ( .A1(n13262), .A2(n13261), .A3(n13260), .A4(n13259), .ZN(
        n13265) );
  AOI22_X1 U14857 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n13605), .B1(
        n13606), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13264) );
  AOI22_X1 U14858 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n13301), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13263) );
  NAND3_X1 U14859 ( .A1(n13265), .A2(n13264), .A3(n13263), .ZN(n13270) );
  AOI22_X1 U14860 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10958), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13268) );
  AOI22_X1 U14861 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n13706), .ZN(n13267) );
  AOI22_X1 U14862 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n13525), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13266) );
  NAND3_X1 U14863 ( .A1(n13268), .A2(n13267), .A3(n13266), .ZN(n13269) );
  OR2_X1 U14864 ( .A1(n13270), .A2(n13269), .ZN(n15208) );
  AOI22_X1 U14865 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n13155), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13275) );
  AOI22_X1 U14866 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n13600), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13274) );
  NAND2_X1 U14867 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13273) );
  NAND2_X1 U14868 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13272) );
  AND4_X1 U14869 ( .A1(n13275), .A2(n13274), .A3(n13273), .A4(n13272), .ZN(
        n13278) );
  AOI22_X1 U14870 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n13605), .B1(
        n13606), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13277) );
  AOI22_X1 U14871 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n13301), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13276) );
  NAND3_X1 U14872 ( .A1(n13278), .A2(n13277), .A3(n13276), .ZN(n13283) );
  AOI22_X1 U14873 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10958), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U14874 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n13706), .ZN(n13280) );
  AOI22_X1 U14875 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n13525), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13279) );
  NAND3_X1 U14876 ( .A1(n13281), .A2(n13280), .A3(n13279), .ZN(n13282) );
  NOR2_X1 U14877 ( .A1(n13283), .A2(n13282), .ZN(n16265) );
  AOI22_X1 U14878 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13155), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13287) );
  AOI22_X1 U14879 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n13600), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13286) );
  NAND2_X1 U14880 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13285) );
  NAND2_X1 U14881 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13284) );
  AND4_X1 U14882 ( .A1(n13287), .A2(n13286), .A3(n13285), .A4(n13284), .ZN(
        n13290) );
  AOI22_X1 U14883 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n13605), .B1(
        n13606), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13289) );
  AOI22_X1 U14884 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n13301), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13288) );
  NAND3_X1 U14885 ( .A1(n13290), .A2(n13289), .A3(n13288), .ZN(n13295) );
  AOI22_X1 U14886 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10957), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13293) );
  AOI22_X1 U14887 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n13706), .ZN(n13292) );
  AOI22_X1 U14888 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n13525), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13291) );
  NAND3_X1 U14889 ( .A1(n13293), .A2(n13292), .A3(n13291), .ZN(n13294) );
  NOR2_X1 U14890 ( .A1(n13295), .A2(n13294), .ZN(n16256) );
  INV_X1 U14891 ( .A(n16256), .ZN(n13296) );
  AOI22_X1 U14892 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13155), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U14893 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13600), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13299) );
  NAND2_X1 U14894 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13298) );
  NAND2_X1 U14895 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13297) );
  AND4_X1 U14896 ( .A1(n13300), .A2(n13299), .A3(n13298), .A4(n13297), .ZN(
        n13304) );
  AOI22_X1 U14897 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n13605), .B1(
        n13606), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13303) );
  AOI22_X1 U14898 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n13301), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13302) );
  NAND3_X1 U14899 ( .A1(n13304), .A2(n13303), .A3(n13302), .ZN(n13310) );
  AOI22_X1 U14900 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10957), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13308) );
  AOI22_X1 U14901 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n13706), .ZN(n13307) );
  AOI22_X1 U14902 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n13525), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13306) );
  NAND3_X1 U14903 ( .A1(n13308), .A2(n13307), .A3(n13306), .ZN(n13309) );
  OR2_X1 U14904 ( .A1(n13310), .A2(n13309), .ZN(n16244) );
  INV_X1 U14905 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15101) );
  NOR2_X1 U14906 ( .A1(n13692), .A2(n15101), .ZN(n13313) );
  INV_X1 U14907 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15105) );
  INV_X1 U14908 ( .A(n14512), .ZN(n13538) );
  INV_X1 U14909 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13311) );
  OAI22_X1 U14910 ( .A1(n11395), .A2(n15105), .B1(n13538), .B2(n13311), .ZN(
        n13312) );
  AOI211_X1 U14911 ( .C1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .C2(n13606), .A(
        n13313), .B(n13312), .ZN(n13317) );
  AOI22_X1 U14912 ( .A1(n13600), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13316) );
  AOI22_X1 U14913 ( .A1(n13598), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13155), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13315) );
  AOI22_X1 U14914 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13271), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13314) );
  AND4_X1 U14915 ( .A1(n13317), .A2(n13316), .A3(n13315), .A4(n13314), .ZN(
        n13321) );
  AOI22_X1 U14916 ( .A1(n10957), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13320) );
  INV_X1 U14917 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19419) );
  AOI22_X1 U14918 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13706), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13319) );
  AOI22_X1 U14919 ( .A1(n13525), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13318) );
  NAND4_X1 U14920 ( .A1(n13321), .A2(n13320), .A3(n13319), .A4(n13318), .ZN(
        n16239) );
  AOI22_X1 U14921 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13271), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U14922 ( .A1(n13600), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U14923 ( .A1(n13598), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13155), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13322) );
  NAND3_X1 U14924 ( .A1(n13324), .A2(n13323), .A3(n13322), .ZN(n13333) );
  INV_X1 U14925 ( .A(n13606), .ZN(n13536) );
  INV_X1 U14926 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13325) );
  INV_X1 U14927 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15325) );
  OAI22_X1 U14928 ( .A1(n13536), .A2(n13325), .B1(n13692), .B2(n15325), .ZN(
        n13332) );
  INV_X1 U14929 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15327) );
  INV_X1 U14930 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13326) );
  OAI22_X1 U14931 ( .A1(n11395), .A2(n15327), .B1(n13538), .B2(n13326), .ZN(
        n13331) );
  AOI22_X1 U14932 ( .A1(n10957), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13329) );
  AOI22_X1 U14933 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13706), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13328) );
  AOI22_X1 U14934 ( .A1(n13525), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13327) );
  NAND3_X1 U14935 ( .A1(n13329), .A2(n13328), .A3(n13327), .ZN(n13330) );
  NOR4_X1 U14936 ( .A1(n13333), .A2(n13332), .A3(n13331), .A4(n13330), .ZN(
        n16235) );
  INV_X1 U14937 ( .A(n13334), .ZN(n13491) );
  AOI22_X1 U14938 ( .A1(n13491), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13344) );
  AND2_X1 U14939 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13336) );
  OR2_X1 U14940 ( .A1(n13336), .A2(n13335), .ZN(n13496) );
  INV_X1 U14941 ( .A(n13496), .ZN(n13432) );
  NAND2_X1 U14942 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13338) );
  NAND2_X1 U14943 ( .A1(n13492), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13337) );
  AND3_X1 U14944 ( .A1(n13432), .A2(n13338), .A3(n13337), .ZN(n13343) );
  AOI22_X1 U14945 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U14946 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13341) );
  NAND4_X1 U14947 ( .A1(n13344), .A2(n13343), .A3(n13342), .A4(n13341), .ZN(
        n13352) );
  AOI22_X1 U14948 ( .A1(n13491), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13350) );
  AOI22_X1 U14949 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13349) );
  AOI22_X1 U14950 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13348) );
  NAND2_X1 U14951 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13346) );
  NAND2_X1 U14952 ( .A1(n13492), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13345) );
  AND3_X1 U14953 ( .A1(n13346), .A2(n13496), .A3(n13345), .ZN(n13347) );
  NAND4_X1 U14954 ( .A1(n13350), .A2(n13349), .A3(n13348), .A4(n13347), .ZN(
        n13351) );
  NAND2_X1 U14955 ( .A1(n13352), .A2(n13351), .ZN(n13366) );
  AOI22_X1 U14956 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13598), .B1(
        n13155), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13356) );
  AOI22_X1 U14957 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n13600), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13355) );
  NAND2_X1 U14958 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n13354) );
  NAND2_X1 U14959 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13353) );
  AND4_X1 U14960 ( .A1(n13356), .A2(n13355), .A3(n13354), .A4(n13353), .ZN(
        n13359) );
  AOI22_X1 U14961 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n13605), .B1(
        n13606), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13358) );
  AOI22_X1 U14962 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n13301), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13357) );
  NAND3_X1 U14963 ( .A1(n13359), .A2(n13358), .A3(n13357), .ZN(n13364) );
  AOI22_X1 U14964 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10957), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13362) );
  AOI22_X1 U14965 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n13706), .ZN(n13361) );
  AOI22_X1 U14966 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n13525), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13360) );
  NAND3_X1 U14967 ( .A1(n13362), .A2(n13361), .A3(n13360), .ZN(n13363) );
  NOR2_X1 U14968 ( .A1(n13364), .A2(n13363), .ZN(n13365) );
  XOR2_X1 U14969 ( .A(n13366), .B(n13365), .Z(n16224) );
  INV_X1 U14970 ( .A(n13365), .ZN(n13368) );
  INV_X1 U14971 ( .A(n13366), .ZN(n13367) );
  AND2_X1 U14972 ( .A1(n13368), .A2(n13367), .ZN(n13384) );
  AOI22_X1 U14973 ( .A1(n13491), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13374) );
  NAND2_X1 U14974 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13370) );
  NAND2_X1 U14975 ( .A1(n13492), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13369) );
  AND3_X1 U14976 ( .A1(n13432), .A2(n13370), .A3(n13369), .ZN(n13373) );
  AOI22_X1 U14977 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13372) );
  AOI22_X1 U14978 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13371) );
  NAND4_X1 U14979 ( .A1(n13374), .A2(n13373), .A3(n13372), .A4(n13371), .ZN(
        n13382) );
  AOI22_X1 U14980 ( .A1(n13491), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13380) );
  AOI22_X1 U14981 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13379) );
  AOI22_X1 U14982 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13378) );
  NAND2_X1 U14983 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13376) );
  NAND2_X1 U14984 ( .A1(n13492), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13375) );
  AND3_X1 U14985 ( .A1(n13376), .A2(n13496), .A3(n13375), .ZN(n13377) );
  NAND4_X1 U14986 ( .A1(n13380), .A2(n13379), .A3(n13378), .A4(n13377), .ZN(
        n13381) );
  NAND2_X1 U14987 ( .A1(n13382), .A2(n13381), .ZN(n13385) );
  INV_X1 U14988 ( .A(n13385), .ZN(n13383) );
  NAND2_X1 U14989 ( .A1(n13384), .A2(n13383), .ZN(n13389) );
  INV_X1 U14990 ( .A(n13384), .ZN(n13386) );
  OAI21_X1 U14991 ( .B1(n13387), .B2(n13386), .A(n13385), .ZN(n13388) );
  OAI21_X1 U14992 ( .B1(n19585), .B2(n13389), .A(n13388), .ZN(n16219) );
  INV_X1 U14993 ( .A(n13389), .ZN(n13405) );
  AOI22_X1 U14994 ( .A1(n13491), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13395) );
  NAND2_X1 U14995 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13391) );
  NAND2_X1 U14996 ( .A1(n13492), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13390) );
  AND3_X1 U14997 ( .A1(n13432), .A2(n13391), .A3(n13390), .ZN(n13394) );
  AOI22_X1 U14998 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13393) );
  AOI22_X1 U14999 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13392) );
  NAND4_X1 U15000 ( .A1(n13395), .A2(n13394), .A3(n13393), .A4(n13392), .ZN(
        n13404) );
  AOI22_X1 U15001 ( .A1(n13396), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U15002 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13401) );
  AOI22_X1 U15003 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13400) );
  NAND2_X1 U15004 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n13398) );
  NAND2_X1 U15005 ( .A1(n13492), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13397) );
  AND3_X1 U15006 ( .A1(n13398), .A2(n13496), .A3(n13397), .ZN(n13399) );
  NAND4_X1 U15007 ( .A1(n13402), .A2(n13401), .A3(n13400), .A4(n13399), .ZN(
        n13403) );
  AND2_X1 U15008 ( .A1(n13404), .A2(n13403), .ZN(n13406) );
  NAND2_X1 U15009 ( .A1(n13405), .A2(n13406), .ZN(n13429) );
  OAI211_X1 U15010 ( .C1(n13405), .C2(n13406), .A(n13445), .B(n13429), .ZN(
        n13408) );
  INV_X1 U15011 ( .A(n13406), .ZN(n13407) );
  NOR2_X1 U15012 ( .A1(n14142), .A2(n13407), .ZN(n16207) );
  AOI22_X1 U15013 ( .A1(n13491), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13415) );
  NAND2_X1 U15014 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13411) );
  NAND2_X1 U15015 ( .A1(n13492), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n13410) );
  AND3_X1 U15016 ( .A1(n13432), .A2(n13411), .A3(n13410), .ZN(n13414) );
  AOI22_X1 U15017 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U15018 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13412) );
  NAND4_X1 U15019 ( .A1(n13415), .A2(n13414), .A3(n13413), .A4(n13412), .ZN(
        n13423) );
  AOI22_X1 U15020 ( .A1(n13491), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13421) );
  AOI22_X1 U15021 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13420) );
  AOI22_X1 U15022 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13419) );
  NAND2_X1 U15023 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n13417) );
  NAND2_X1 U15024 ( .A1(n13492), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13416) );
  AND3_X1 U15025 ( .A1(n13417), .A2(n13496), .A3(n13416), .ZN(n13418) );
  NAND4_X1 U15026 ( .A1(n13421), .A2(n13420), .A3(n13419), .A4(n13418), .ZN(
        n13422) );
  AND2_X1 U15027 ( .A1(n13423), .A2(n13422), .ZN(n13427) );
  XNOR2_X1 U15028 ( .A(n13429), .B(n13427), .ZN(n13424) );
  XNOR2_X1 U15029 ( .A(n13425), .B(n11394), .ZN(n16203) );
  NAND2_X1 U15030 ( .A1(n19585), .A2(n13427), .ZN(n16202) );
  INV_X1 U15031 ( .A(n13427), .ZN(n13428) );
  NOR2_X1 U15032 ( .A1(n13429), .A2(n13428), .ZN(n13446) );
  AOI22_X1 U15033 ( .A1(n13491), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13436) );
  NAND2_X1 U15034 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13431) );
  NAND2_X1 U15035 ( .A1(n13492), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n13430) );
  AND3_X1 U15036 ( .A1(n13432), .A2(n13431), .A3(n13430), .ZN(n13435) );
  AOI22_X1 U15037 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13434) );
  AOI22_X1 U15038 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13433) );
  NAND4_X1 U15039 ( .A1(n13436), .A2(n13435), .A3(n13434), .A4(n13433), .ZN(
        n13444) );
  AOI22_X1 U15040 ( .A1(n13491), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13442) );
  AOI22_X1 U15041 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13441) );
  AOI22_X1 U15042 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13440) );
  NAND2_X1 U15043 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n13438) );
  NAND2_X1 U15044 ( .A1(n13492), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13437) );
  AND3_X1 U15045 ( .A1(n13438), .A2(n13496), .A3(n13437), .ZN(n13439) );
  NAND4_X1 U15046 ( .A1(n13442), .A2(n13441), .A3(n13440), .A4(n13439), .ZN(
        n13443) );
  AND2_X1 U15047 ( .A1(n13444), .A2(n13443), .ZN(n13447) );
  NAND2_X1 U15048 ( .A1(n13446), .A2(n13447), .ZN(n13470) );
  OAI211_X1 U15049 ( .C1(n13446), .C2(n13447), .A(n13445), .B(n13470), .ZN(
        n13468) );
  INV_X1 U15050 ( .A(n13447), .ZN(n13448) );
  NOR2_X1 U15051 ( .A1(n14142), .A2(n13448), .ZN(n16191) );
  INV_X1 U15052 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13451) );
  AOI21_X1 U15053 ( .B1(n13492), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n13496), .ZN(n13450) );
  AOI22_X1 U15054 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13449) );
  OAI211_X1 U15055 ( .C1(n14505), .C2(n13451), .A(n13450), .B(n13449), .ZN(
        n13456) );
  INV_X1 U15056 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13452) );
  OAI22_X1 U15057 ( .A1(n13334), .A2(n15101), .B1(n13457), .B2(n13452), .ZN(
        n13455) );
  INV_X1 U15058 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13453) );
  OAI22_X1 U15059 ( .A1(n13462), .A2(n13453), .B1(n13340), .B2(n15105), .ZN(
        n13454) );
  NOR3_X1 U15060 ( .A1(n13456), .A2(n13455), .A3(n13454), .ZN(n13467) );
  INV_X1 U15061 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15106) );
  OAI22_X1 U15062 ( .A1(n13334), .A2(n15106), .B1(n13457), .B2(n19419), .ZN(
        n13465) );
  AOI22_X1 U15063 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13460) );
  NAND2_X1 U15064 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n13459) );
  NAND2_X1 U15065 ( .A1(n13492), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13458) );
  NAND4_X1 U15066 ( .A1(n13460), .A2(n13496), .A3(n13459), .A4(n13458), .ZN(
        n13464) );
  INV_X1 U15067 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13461) );
  INV_X1 U15068 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15102) );
  OAI22_X1 U15069 ( .A1(n13462), .A2(n13461), .B1(n13340), .B2(n15102), .ZN(
        n13463) );
  NOR3_X1 U15070 ( .A1(n13465), .A2(n13464), .A3(n13463), .ZN(n13466) );
  NOR2_X1 U15071 ( .A1(n13467), .A2(n13466), .ZN(n16182) );
  NAND2_X1 U15072 ( .A1(n13469), .A2(n13468), .ZN(n16188) );
  INV_X1 U15073 ( .A(n13470), .ZN(n16181) );
  NAND3_X1 U15074 ( .A1(n16181), .A2(n16182), .A3(n14142), .ZN(n16176) );
  AOI22_X1 U15075 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13472) );
  AOI22_X1 U15076 ( .A1(n13491), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13471) );
  NAND2_X1 U15077 ( .A1(n13472), .A2(n13471), .ZN(n13485) );
  INV_X1 U15078 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13475) );
  AOI21_X1 U15079 ( .B1(n13492), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n13496), .ZN(n13474) );
  AOI22_X1 U15080 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13473) );
  OAI211_X1 U15081 ( .C1(n14505), .C2(n13475), .A(n13474), .B(n13473), .ZN(
        n13484) );
  AOI22_X1 U15082 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13476), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13478) );
  AOI22_X1 U15083 ( .A1(n13133), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13492), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13477) );
  NAND2_X1 U15084 ( .A1(n13478), .A2(n13477), .ZN(n13483) );
  AOI22_X1 U15085 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13481) );
  NAND2_X1 U15086 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n13480) );
  NAND2_X1 U15087 ( .A1(n13143), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n13479) );
  NAND4_X1 U15088 ( .A1(n13481), .A2(n13496), .A3(n13480), .A4(n13479), .ZN(
        n13482) );
  OAI22_X1 U15089 ( .A1(n13485), .A2(n13484), .B1(n13483), .B2(n13482), .ZN(
        n16175) );
  AOI21_X1 U15090 ( .B1(n16174), .B2(n16176), .A(n16175), .ZN(n13506) );
  AOI22_X1 U15091 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13491), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13487) );
  AOI22_X1 U15092 ( .A1(n13133), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13143), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13486) );
  NAND2_X1 U15093 ( .A1(n13487), .A2(n13486), .ZN(n13503) );
  INV_X1 U15094 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13490) );
  AOI21_X1 U15095 ( .B1(n13492), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n13496), .ZN(n13489) );
  AOI22_X1 U15096 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13488) );
  OAI211_X1 U15097 ( .C1(n14505), .C2(n13490), .A(n13489), .B(n13488), .ZN(
        n13502) );
  AOI22_X1 U15098 ( .A1(n13491), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13494) );
  AOI22_X1 U15099 ( .A1(n10959), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13492), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13493) );
  NAND2_X1 U15100 ( .A1(n13494), .A2(n13493), .ZN(n13501) );
  AOI22_X1 U15101 ( .A1(n13495), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13135), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13499) );
  NAND2_X1 U15102 ( .A1(n13143), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13498) );
  NAND2_X1 U15103 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n13497) );
  NAND4_X1 U15104 ( .A1(n13499), .A2(n13498), .A3(n13497), .A4(n13496), .ZN(
        n13500) );
  OAI22_X1 U15105 ( .A1(n13503), .A2(n13502), .B1(n13501), .B2(n13500), .ZN(
        n13504) );
  INV_X1 U15106 ( .A(n13504), .ZN(n13505) );
  XNOR2_X1 U15107 ( .A(n13506), .B(n13505), .ZN(n15303) );
  XNOR2_X1 U15108 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13841) );
  NAND2_X1 U15109 ( .A1(n13841), .A2(n13563), .ZN(n13508) );
  NAND2_X1 U15110 ( .A1(n19260), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13507) );
  NAND2_X1 U15111 ( .A1(n13508), .A2(n13507), .ZN(n13561) );
  XNOR2_X1 U15112 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13559) );
  NAND2_X1 U15113 ( .A1(n13561), .A2(n13559), .ZN(n13510) );
  NAND2_X1 U15114 ( .A1(n19256), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13509) );
  XNOR2_X1 U15115 ( .A(n13511), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13557) );
  INV_X1 U15116 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16838) );
  NOR2_X1 U15117 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16838), .ZN(
        n13514) );
  NAND3_X1 U15118 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13515), .A3(
        n13917), .ZN(n13830) );
  NOR2_X1 U15119 ( .A1(n13830), .A2(n13837), .ZN(n13516) );
  OR2_X1 U15120 ( .A1(n13844), .A2(n13516), .ZN(n13575) );
  AOI22_X1 U15121 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13155), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13520) );
  AOI22_X1 U15122 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n13599), .B1(
        n13600), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13519) );
  NAND2_X1 U15123 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n13518) );
  NAND2_X1 U15124 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n13517) );
  AND4_X1 U15125 ( .A1(n13520), .A2(n13519), .A3(n13518), .A4(n13517), .ZN(
        n13534) );
  NAND2_X1 U15126 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13524) );
  NAND2_X1 U15127 ( .A1(n13605), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13523) );
  NAND2_X1 U15128 ( .A1(n13301), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n13522) );
  NAND2_X1 U15129 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n13521) );
  AOI22_X1 U15130 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13705), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13532) );
  INV_X1 U15131 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13527) );
  INV_X1 U15132 ( .A(n13525), .ZN(n13547) );
  INV_X1 U15133 ( .A(n13707), .ZN(n13546) );
  INV_X1 U15134 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13526) );
  OAI22_X1 U15135 ( .A1(n13527), .A2(n13547), .B1(n13546), .B2(n13526), .ZN(
        n13530) );
  INV_X1 U15136 ( .A(n13834), .ZN(n13550) );
  INV_X1 U15137 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13528) );
  INV_X1 U15138 ( .A(n13706), .ZN(n13549) );
  OAI22_X1 U15139 ( .A1(n13550), .A2(n13528), .B1(n19469), .B2(n13549), .ZN(
        n13529) );
  NOR2_X1 U15140 ( .A1(n13530), .A2(n13529), .ZN(n13531) );
  NAND4_X1 U15141 ( .A1(n13534), .A2(n13533), .A3(n13532), .A4(n13531), .ZN(
        n15052) );
  MUX2_X1 U15142 ( .A(n13830), .B(n15052), .S(n11085), .Z(n14840) );
  INV_X1 U15143 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13537) );
  INV_X1 U15144 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13535) );
  OAI22_X1 U15145 ( .A1(n13537), .A2(n13536), .B1(n13692), .B2(n13535), .ZN(
        n13541) );
  INV_X1 U15146 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13539) );
  INV_X1 U15147 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14996) );
  OAI22_X1 U15148 ( .A1(n13539), .A2(n13538), .B1(n11395), .B2(n14996), .ZN(
        n13540) );
  NOR2_X1 U15149 ( .A1(n13541), .A2(n13540), .ZN(n13556) );
  AOI22_X1 U15150 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13155), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13545) );
  AOI22_X1 U15151 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n13599), .B1(
        n13600), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13544) );
  NAND2_X1 U15152 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n13543) );
  NAND2_X1 U15153 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n13542) );
  AND4_X1 U15154 ( .A1(n13545), .A2(n13544), .A3(n13543), .A4(n13542), .ZN(
        n13555) );
  AOI22_X1 U15155 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13705), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13554) );
  INV_X1 U15156 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13548) );
  INV_X1 U15157 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15002) );
  OAI22_X1 U15158 ( .A1(n13548), .A2(n13547), .B1(n13546), .B2(n15002), .ZN(
        n13552) );
  INV_X1 U15159 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14997) );
  INV_X1 U15160 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19517) );
  OAI22_X1 U15161 ( .A1(n13550), .A2(n14997), .B1(n19517), .B2(n13549), .ZN(
        n13551) );
  NOR2_X1 U15162 ( .A1(n13552), .A2(n13551), .ZN(n13553) );
  NAND4_X1 U15163 ( .A1(n13556), .A2(n13555), .A3(n13554), .A4(n13553), .ZN(
        n15014) );
  XNOR2_X1 U15164 ( .A(n13558), .B(n13557), .ZN(n13829) );
  MUX2_X1 U15165 ( .A(n15014), .B(n13829), .S(n13837), .Z(n14722) );
  NAND2_X1 U15166 ( .A1(n14840), .A2(n14722), .ZN(n13843) );
  INV_X1 U15167 ( .A(n13559), .ZN(n13560) );
  XNOR2_X1 U15168 ( .A(n13561), .B(n13560), .ZN(n13828) );
  NAND2_X1 U15169 ( .A1(n13837), .A2(n13828), .ZN(n13839) );
  INV_X1 U15170 ( .A(n13839), .ZN(n13572) );
  AOI21_X1 U15171 ( .B1(n18227), .B2(n14142), .A(n13828), .ZN(n13571) );
  INV_X1 U15172 ( .A(n13828), .ZN(n13569) );
  INV_X1 U15173 ( .A(n13563), .ZN(n13566) );
  NAND2_X1 U15174 ( .A1(n14490), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13564) );
  AND2_X1 U15175 ( .A1(n13566), .A2(n13564), .ZN(n13838) );
  NAND2_X1 U15176 ( .A1(n13838), .A2(n13841), .ZN(n13565) );
  NAND2_X1 U15177 ( .A1(n11085), .A2(n13565), .ZN(n13568) );
  XNOR2_X1 U15178 ( .A(n13841), .B(n13566), .ZN(n13581) );
  OAI211_X1 U15179 ( .C1(n14142), .C2(n13838), .A(n19642), .B(n13581), .ZN(
        n13567) );
  OAI211_X1 U15180 ( .C1(n13562), .C2(n13569), .A(n13568), .B(n13567), .ZN(
        n13570) );
  OAI21_X1 U15181 ( .B1(n13572), .B2(n13571), .A(n13570), .ZN(n13573) );
  AOI22_X1 U15182 ( .A1(n13843), .A2(n13837), .B1(n13829), .B2(n13573), .ZN(
        n13574) );
  NOR2_X1 U15183 ( .A1(n13575), .A2(n13574), .ZN(n13576) );
  MUX2_X1 U15184 ( .A(n13917), .B(n13576), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n14098) );
  AND2_X1 U15185 ( .A1(n13844), .A2(n13031), .ZN(n13577) );
  AND3_X1 U15186 ( .A1(n19585), .A2(n19534), .A3(n15490), .ZN(n13580) );
  AND2_X1 U15187 ( .A1(n13578), .A2(n13580), .ZN(n14523) );
  AND4_X1 U15188 ( .A1(n13830), .A2(n13828), .A3(n13829), .A4(n13581), .ZN(
        n13582) );
  OR2_X1 U15189 ( .A1(n13844), .A2(n13582), .ZN(n14538) );
  INV_X1 U15190 ( .A(n13583), .ZN(n13584) );
  NAND2_X1 U15191 ( .A1(n13584), .A2(n19642), .ZN(n14115) );
  OR2_X1 U15192 ( .A1(n14555), .A2(n19642), .ZN(n14116) );
  NAND2_X1 U15193 ( .A1(n14115), .A2(n14116), .ZN(n14536) );
  NAND2_X1 U15194 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n18222) );
  AND2_X1 U15195 ( .A1(n13585), .A2(n18222), .ZN(n14534) );
  NAND2_X1 U15196 ( .A1(n14536), .A2(n14534), .ZN(n13586) );
  NOR2_X1 U15197 ( .A1(n14538), .A2(n13586), .ZN(n13587) );
  AOI21_X1 U15198 ( .B1(n14561), .B2(n14523), .A(n13587), .ZN(n13910) );
  INV_X1 U15199 ( .A(n13562), .ZN(n14122) );
  NAND3_X1 U15200 ( .A1(n13041), .A2(n14122), .A3(n14136), .ZN(n13588) );
  NAND2_X1 U15201 ( .A1(n13910), .A2(n13588), .ZN(n13589) );
  AND2_X1 U15202 ( .A1(n15263), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14551) );
  NAND2_X1 U15203 ( .A1(n19531), .A2(n13597), .ZN(n19579) );
  AND2_X1 U15204 ( .A1(n13968), .A2(n17222), .ZN(n13590) );
  NAND2_X1 U15205 ( .A1(n13591), .A2(n13590), .ZN(n13727) );
  OR2_X1 U15206 ( .A1(n13727), .A2(n18240), .ZN(n13596) );
  INV_X1 U15207 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13593) );
  INV_X1 U15208 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16783) );
  NAND2_X1 U15209 ( .A1(n14142), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13592) );
  OAI211_X1 U15210 ( .C1(n13968), .C2(n13593), .A(n13592), .B(n17222), .ZN(
        n13594) );
  INV_X1 U15211 ( .A(n13594), .ZN(n13595) );
  NAND2_X1 U15212 ( .A1(n13596), .A2(n13595), .ZN(n14160) );
  AND2_X2 U15213 ( .A1(n13024), .A2(n17222), .ZN(n13655) );
  NAND2_X1 U15214 ( .A1(n13597), .A2(n13655), .ZN(n13650) );
  MUX2_X1 U15215 ( .A(n13968), .B(n19288), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13616) );
  AOI22_X1 U15216 ( .A1(n13598), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13155), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13604) );
  AOI22_X1 U15217 ( .A1(n13600), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13603) );
  NAND2_X1 U15218 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13602) );
  NAND2_X1 U15219 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13601) );
  AND4_X1 U15220 ( .A1(n13604), .A2(n13603), .A3(n13602), .A4(n13601), .ZN(
        n13609) );
  AOI22_X1 U15221 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13605), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13608) );
  AOI22_X1 U15222 ( .A1(n13301), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14512), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13607) );
  NAND3_X1 U15223 ( .A1(n13609), .A2(n13608), .A3(n13607), .ZN(n13614) );
  AOI22_X1 U15224 ( .A1(n10958), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13612) );
  INV_X1 U15225 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U15226 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13706), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13611) );
  AOI22_X1 U15227 ( .A1(n13525), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13610) );
  NAND3_X1 U15228 ( .A1(n13612), .A2(n13611), .A3(n13610), .ZN(n13613) );
  NAND2_X1 U15229 ( .A1(n13748), .A2(n13867), .ZN(n13615) );
  NAND3_X1 U15230 ( .A1(n13650), .A2(n13616), .A3(n13615), .ZN(n14159) );
  OR2_X1 U15231 ( .A1(n13727), .A2(n13869), .ZN(n13618) );
  NOR2_X1 U15232 ( .A1(n13968), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13654) );
  INV_X1 U15233 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16789) );
  AOI22_X1 U15234 ( .A1(n13654), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13655), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13617) );
  NAND2_X1 U15235 ( .A1(n13618), .A2(n13617), .ZN(n13636) );
  INV_X1 U15236 ( .A(n13636), .ZN(n13619) );
  NAND2_X1 U15237 ( .A1(n12952), .A2(n13968), .ZN(n13620) );
  MUX2_X1 U15238 ( .A(n13620), .B(n19260), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13634) );
  AOI22_X1 U15239 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13155), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13624) );
  AOI22_X1 U15240 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13599), .B1(
        n13600), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13623) );
  NAND2_X1 U15241 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13622) );
  NAND2_X1 U15242 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13621) );
  AND4_X1 U15243 ( .A1(n13624), .A2(n13623), .A3(n13622), .A4(n13621), .ZN(
        n13627) );
  AOI22_X1 U15244 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n13606), .B1(
        n13605), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13626) );
  AOI22_X1 U15245 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14512), .B1(
        n13301), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13625) );
  NAND3_X1 U15246 ( .A1(n13627), .A2(n13626), .A3(n13625), .ZN(n13632) );
  AOI22_X1 U15247 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13705), .B1(
        n10957), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13630) );
  AOI22_X1 U15248 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n13706), .ZN(n13629) );
  AOI22_X1 U15249 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n13525), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13628) );
  NAND3_X1 U15250 ( .A1(n13630), .A2(n13629), .A3(n13628), .ZN(n13631) );
  NAND2_X1 U15251 ( .A1(n10955), .A2(n13884), .ZN(n13633) );
  NAND2_X1 U15252 ( .A1(n13634), .A2(n13633), .ZN(n14146) );
  INV_X1 U15253 ( .A(n14146), .ZN(n13635) );
  NAND2_X1 U15254 ( .A1(n14145), .A2(n13635), .ZN(n14149) );
  AOI22_X1 U15255 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n13155), .B1(
        n13598), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13640) );
  AOI22_X1 U15256 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n13599), .B1(
        n13600), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13639) );
  NAND2_X1 U15257 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n13638) );
  NAND2_X1 U15258 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13637) );
  AND4_X1 U15259 ( .A1(n13640), .A2(n13639), .A3(n13638), .A4(n13637), .ZN(
        n13643) );
  AOI22_X1 U15260 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n13606), .B1(
        n13605), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13642) );
  AOI22_X1 U15261 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n14512), .B1(
        n13301), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13641) );
  NAND3_X1 U15262 ( .A1(n13643), .A2(n13642), .A3(n13641), .ZN(n13648) );
  AOI22_X1 U15263 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13705), .B1(
        n13305), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13646) );
  AOI22_X1 U15264 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n13706), .ZN(n13645) );
  AOI22_X1 U15265 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n13525), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13644) );
  NAND3_X1 U15266 ( .A1(n13646), .A2(n13645), .A3(n13644), .ZN(n13647) );
  OR2_X2 U15267 ( .A1(n13648), .A2(n13647), .ZN(n15034) );
  NAND2_X1 U15268 ( .A1(n10955), .A2(n15034), .ZN(n13649) );
  OAI211_X1 U15269 ( .C1(n17222), .C2(n19256), .A(n13650), .B(n13649), .ZN(
        n13651) );
  AND3_X1 U15270 ( .A1(n14149), .A2(n13652), .A3(n13651), .ZN(n13653) );
  OR2_X1 U15271 ( .A1(n13775), .A2(n18577), .ZN(n13657) );
  AOI22_X1 U15272 ( .A1(n15550), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13655), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13656) );
  NAND2_X1 U15273 ( .A1(n13657), .A2(n13656), .ZN(n14926) );
  NOR2_X1 U15274 ( .A1(n14927), .A2(n14926), .ZN(n13658) );
  NOR2_X1 U15275 ( .A1(n13659), .A2(n13658), .ZN(n14718) );
  AOI22_X1 U15276 ( .A1(n10955), .A2(n15014), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13655), .ZN(n13661) );
  AOI22_X1 U15277 ( .A1(n15550), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13660) );
  OAI211_X1 U15278 ( .C1(n13775), .C2(n13662), .A(n13661), .B(n13660), .ZN(
        n14717) );
  NAND2_X1 U15279 ( .A1(n14718), .A2(n14717), .ZN(n14846) );
  INV_X1 U15280 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n13663) );
  OR2_X1 U15281 ( .A1(n13775), .A2(n13663), .ZN(n13666) );
  AOI22_X1 U15282 ( .A1(n15550), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13655), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13665) );
  NAND2_X1 U15283 ( .A1(n10955), .A2(n15052), .ZN(n13664) );
  AOI22_X1 U15284 ( .A1(n10958), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13669) );
  AOI22_X1 U15285 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13706), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13668) );
  AOI22_X1 U15286 ( .A1(n13525), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13667) );
  AND3_X1 U15287 ( .A1(n13669), .A2(n13668), .A3(n13667), .ZN(n13681) );
  AOI22_X1 U15288 ( .A1(n13598), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13155), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13673) );
  AOI22_X1 U15289 ( .A1(n13600), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13672) );
  NAND2_X1 U15290 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13671) );
  NAND2_X1 U15291 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n13670) );
  NAND4_X1 U15292 ( .A1(n13673), .A2(n13672), .A3(n13671), .A4(n13670), .ZN(
        n13679) );
  NAND2_X1 U15293 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13677) );
  NAND2_X1 U15294 ( .A1(n13605), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13676) );
  NAND2_X1 U15295 ( .A1(n13301), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n13675) );
  NAND2_X1 U15296 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n13674) );
  NAND4_X1 U15297 ( .A1(n13677), .A2(n13676), .A3(n13675), .A4(n13674), .ZN(
        n13678) );
  NOR2_X1 U15298 ( .A1(n13679), .A2(n13678), .ZN(n13680) );
  AOI22_X1 U15299 ( .A1(n13682), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n10955), 
        .B2(n14871), .ZN(n13684) );
  AOI22_X1 U15300 ( .A1(n15550), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n13655), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13683) );
  NAND2_X1 U15301 ( .A1(n13684), .A2(n13683), .ZN(n15147) );
  AOI22_X1 U15302 ( .A1(n10958), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13705), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13687) );
  AOI22_X1 U15303 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13706), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13686) );
  AOI22_X1 U15304 ( .A1(n13525), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13685) );
  AND3_X1 U15305 ( .A1(n13687), .A2(n13686), .A3(n13685), .ZN(n13700) );
  AOI22_X1 U15306 ( .A1(n13598), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13155), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13691) );
  AOI22_X1 U15307 ( .A1(n13600), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13599), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13690) );
  NAND2_X1 U15308 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n13689) );
  NAND2_X1 U15309 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n13688) );
  NAND4_X1 U15310 ( .A1(n13691), .A2(n13690), .A3(n13689), .A4(n13688), .ZN(
        n13698) );
  NAND2_X1 U15311 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13696) );
  NAND2_X1 U15312 ( .A1(n13605), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n13695) );
  NAND2_X1 U15313 ( .A1(n13301), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n13694) );
  NAND2_X1 U15314 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n13693) );
  NAND4_X1 U15315 ( .A1(n13696), .A2(n13695), .A3(n13694), .A4(n13693), .ZN(
        n13697) );
  NOR2_X1 U15316 ( .A1(n13698), .A2(n13697), .ZN(n13699) );
  INV_X1 U15317 ( .A(n15336), .ZN(n13701) );
  NAND2_X1 U15318 ( .A1(n10955), .A2(n13701), .ZN(n13702) );
  INV_X1 U15319 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n17272) );
  OR2_X1 U15320 ( .A1(n13775), .A2(n17272), .ZN(n13704) );
  AOI22_X1 U15321 ( .A1(n15550), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n13655), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13703) );
  NAND2_X1 U15322 ( .A1(n13704), .A2(n13703), .ZN(n14880) );
  AOI22_X1 U15323 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13705), .B1(
        n10958), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13710) );
  AOI22_X1 U15324 ( .A1(n13834), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n13706), .ZN(n13709) );
  AOI22_X1 U15325 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n13525), .B1(
        n13707), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13708) );
  AND3_X1 U15326 ( .A1(n13710), .A2(n13709), .A3(n13708), .ZN(n13722) );
  AOI22_X1 U15327 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n13598), .B1(
        n13155), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13714) );
  AOI22_X1 U15328 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n13599), .B1(
        n13600), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13713) );
  NAND2_X1 U15329 ( .A1(n13156), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n13712) );
  NAND2_X1 U15330 ( .A1(n13271), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n13711) );
  NAND4_X1 U15331 ( .A1(n13714), .A2(n13713), .A3(n13712), .A4(n13711), .ZN(
        n13720) );
  NAND2_X1 U15332 ( .A1(n13606), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13718) );
  NAND2_X1 U15333 ( .A1(n13605), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n13717) );
  NAND2_X1 U15334 ( .A1(n13301), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n13716) );
  NAND2_X1 U15335 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n13715) );
  NAND4_X1 U15336 ( .A1(n13718), .A2(n13717), .A3(n13716), .A4(n13715), .ZN(
        n13719) );
  NOR2_X1 U15337 ( .A1(n13720), .A2(n13719), .ZN(n13721) );
  NAND2_X1 U15338 ( .A1(n10955), .A2(n11050), .ZN(n13723) );
  INV_X1 U15339 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n18265) );
  OR2_X1 U15340 ( .A1(n13775), .A2(n18265), .ZN(n13726) );
  AOI22_X1 U15341 ( .A1(n15550), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n13655), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13725) );
  NAND2_X1 U15342 ( .A1(n13726), .A2(n13725), .ZN(n16737) );
  INV_X1 U15343 ( .A(n10955), .ZN(n13742) );
  INV_X1 U15344 ( .A(n14680), .ZN(n13729) );
  AOI22_X1 U15345 ( .A1(n15550), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n13655), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13728) );
  OAI21_X1 U15346 ( .B1(n13742), .B2(n13729), .A(n13728), .ZN(n13730) );
  AOI21_X1 U15347 ( .B1(n13682), .B2(P2_REIP_REG_8__SCAN_IN), .A(n13730), .ZN(
        n14869) );
  NOR2_X2 U15348 ( .A1(n16739), .A2(n14869), .ZN(n16723) );
  INV_X1 U15349 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n14704) );
  AOI22_X1 U15350 ( .A1(n15550), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n13655), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13732) );
  NAND2_X1 U15351 ( .A1(n10955), .A2(n11406), .ZN(n13731) );
  OAI211_X1 U15352 ( .C1(n13775), .C2(n14704), .A(n13732), .B(n13731), .ZN(
        n16724) );
  INV_X1 U15353 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n13733) );
  OR2_X1 U15354 ( .A1(n13775), .A2(n13733), .ZN(n13737) );
  AOI22_X1 U15355 ( .A1(n15550), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13736) );
  INV_X1 U15356 ( .A(n13734), .ZN(n14858) );
  NAND2_X1 U15357 ( .A1(n10955), .A2(n14858), .ZN(n13735) );
  AOI22_X1 U15358 ( .A1(n13682), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n15550), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13739) );
  AOI22_X1 U15359 ( .A1(n10955), .A2(n14948), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n13655), .ZN(n13738) );
  NAND2_X1 U15360 ( .A1(n13739), .A2(n13738), .ZN(n16690) );
  INV_X1 U15361 ( .A(n14947), .ZN(n13741) );
  AOI22_X1 U15362 ( .A1(n15550), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13740) );
  OAI21_X1 U15363 ( .B1(n13742), .B2(n13741), .A(n13740), .ZN(n13743) );
  AOI21_X1 U15364 ( .B1(n13682), .B2(P2_REIP_REG_12__SCAN_IN), .A(n13743), 
        .ZN(n16136) );
  INV_X1 U15365 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n16453) );
  AOI22_X1 U15366 ( .A1(n15550), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13745) );
  NAND2_X1 U15367 ( .A1(n10955), .A2(n14896), .ZN(n13744) );
  OAI211_X1 U15368 ( .C1(n13775), .C2(n16453), .A(n13745), .B(n13744), .ZN(
        n16126) );
  INV_X1 U15369 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n17274) );
  AOI22_X1 U15370 ( .A1(n15550), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13747) );
  NAND2_X1 U15371 ( .A1(n10955), .A2(n14921), .ZN(n13746) );
  OAI211_X1 U15372 ( .C1(n13775), .C2(n17274), .A(n13747), .B(n13746), .ZN(
        n15079) );
  INV_X1 U15373 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n14969) );
  AOI22_X1 U15374 ( .A1(n15550), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13750) );
  NAND2_X1 U15375 ( .A1(n10955), .A2(n14965), .ZN(n13749) );
  OAI211_X1 U15376 ( .C1(n13775), .C2(n14969), .A(n13750), .B(n13749), .ZN(
        n16650) );
  NAND2_X2 U15377 ( .A1(n16651), .A2(n16650), .ZN(n16652) );
  INV_X1 U15378 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15174) );
  OR2_X1 U15379 ( .A1(n13775), .A2(n15174), .ZN(n13752) );
  AOI22_X1 U15380 ( .A1(n15550), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13751) );
  INV_X1 U15381 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n17275) );
  OR2_X1 U15382 ( .A1(n13775), .A2(n17275), .ZN(n13754) );
  AOI22_X1 U15383 ( .A1(n15550), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13753) );
  NAND2_X1 U15384 ( .A1(n13754), .A2(n13753), .ZN(n16334) );
  AOI222_X1 U15385 ( .A1(n13682), .A2(P2_REIP_REG_18__SCAN_IN), .B1(n15550), 
        .B2(P2_EAX_REG_18__SCAN_IN), .C1(n13655), .C2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18351) );
  INV_X1 U15386 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n17276) );
  OR2_X1 U15387 ( .A1(n13775), .A2(n17276), .ZN(n13756) );
  AOI22_X1 U15388 ( .A1(n15550), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13755) );
  NAND2_X1 U15389 ( .A1(n13756), .A2(n13755), .ZN(n16328) );
  INV_X1 U15390 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15260) );
  OR2_X1 U15391 ( .A1(n13775), .A2(n15260), .ZN(n13758) );
  AOI22_X1 U15392 ( .A1(n15550), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13757) );
  INV_X1 U15393 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n17277) );
  OR2_X1 U15394 ( .A1(n13775), .A2(n17277), .ZN(n13760) );
  AOI22_X1 U15395 ( .A1(n15550), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13759) );
  NAND2_X1 U15396 ( .A1(n13760), .A2(n13759), .ZN(n16321) );
  AOI222_X1 U15397 ( .A1(n13682), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n13655), .C1(n15550), .C2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16577) );
  INV_X1 U15398 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n17278) );
  OR2_X1 U15399 ( .A1(n13775), .A2(n17278), .ZN(n13762) );
  AOI22_X1 U15400 ( .A1(n15550), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13761) );
  NAND2_X1 U15401 ( .A1(n13762), .A2(n13761), .ZN(n16315) );
  INV_X1 U15402 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n15277) );
  OR2_X1 U15403 ( .A1(n13775), .A2(n15277), .ZN(n13764) );
  AOI22_X1 U15404 ( .A1(n15550), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13763) );
  NAND2_X1 U15405 ( .A1(n13764), .A2(n13763), .ZN(n16308) );
  INV_X1 U15406 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n17279) );
  OR2_X1 U15407 ( .A1(n13775), .A2(n17279), .ZN(n13766) );
  AOI22_X1 U15408 ( .A1(n15550), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13765) );
  AND2_X1 U15409 ( .A1(n13766), .A2(n13765), .ZN(n16301) );
  INV_X1 U15410 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n17280) );
  OR2_X1 U15411 ( .A1(n13775), .A2(n17280), .ZN(n13768) );
  AOI22_X1 U15412 ( .A1(n15550), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13767) );
  NAND2_X1 U15413 ( .A1(n13768), .A2(n13767), .ZN(n16294) );
  INV_X1 U15414 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n18448) );
  OR2_X1 U15415 ( .A1(n13775), .A2(n18448), .ZN(n13770) );
  AOI22_X1 U15416 ( .A1(n15550), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13769) );
  AND2_X1 U15417 ( .A1(n13770), .A2(n13769), .ZN(n16283) );
  INV_X1 U15418 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n15291) );
  OR2_X1 U15419 ( .A1(n13775), .A2(n15291), .ZN(n13772) );
  AOI22_X1 U15420 ( .A1(n15550), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13771) );
  AND2_X1 U15421 ( .A1(n13772), .A2(n13771), .ZN(n16276) );
  INV_X1 U15422 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n17282) );
  OR2_X1 U15423 ( .A1(n13775), .A2(n17282), .ZN(n13774) );
  AOI22_X1 U15424 ( .A1(n15550), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13773) );
  INV_X1 U15425 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n17283) );
  OR2_X1 U15426 ( .A1(n13775), .A2(n17283), .ZN(n13777) );
  AOI22_X1 U15427 ( .A1(n15550), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n13655), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13776) );
  NAND2_X1 U15428 ( .A1(n13777), .A2(n13776), .ZN(n13779) );
  INV_X1 U15429 ( .A(n13778), .ZN(n13781) );
  INV_X1 U15430 ( .A(n13779), .ZN(n13780) );
  NAND2_X1 U15431 ( .A1(n13781), .A2(n13780), .ZN(n13782) );
  AND2_X1 U15432 ( .A1(n19381), .A2(n13968), .ZN(n13784) );
  NAND2_X1 U15433 ( .A1(n19531), .A2(n13784), .ZN(n16337) );
  NOR4_X1 U15434 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13788) );
  NOR4_X1 U15435 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13787) );
  NOR4_X1 U15436 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13786) );
  NOR4_X1 U15437 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13785) );
  NAND4_X1 U15438 ( .A1(n13788), .A2(n13787), .A3(n13786), .A4(n13785), .ZN(
        n13793) );
  NOR4_X1 U15439 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13791) );
  NOR4_X1 U15440 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13790) );
  NOR4_X1 U15441 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13789) );
  INV_X1 U15442 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19757) );
  NAND4_X1 U15443 ( .A1(n13791), .A2(n13790), .A3(n13789), .A4(n19757), .ZN(
        n13792) );
  NAND2_X1 U15444 ( .A1(n19108), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13795) );
  INV_X1 U15445 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20057) );
  OR2_X1 U15446 ( .A1(n14088), .A2(n20057), .ZN(n13794) );
  NAND2_X1 U15447 ( .A1(n13795), .A2(n13794), .ZN(n19083) );
  INV_X1 U15448 ( .A(n19083), .ZN(n13797) );
  INV_X1 U15449 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13796) );
  OAI22_X1 U15450 ( .A1(n16337), .A2(n13797), .B1(n19531), .B2(n13796), .ZN(
        n13798) );
  AOI21_X1 U15451 ( .B1(n16113), .B2(n19633), .A(n13798), .ZN(n13802) );
  AND2_X1 U15452 ( .A1(n13799), .A2(n13968), .ZN(n13800) );
  NAND2_X1 U15453 ( .A1(n19531), .A2(n13800), .ZN(n14157) );
  NOR2_X2 U15454 ( .A1(n14157), .A2(n19109), .ZN(n19630) );
  NOR2_X2 U15455 ( .A1(n14157), .A2(n19108), .ZN(n19631) );
  AOI22_X1 U15456 ( .A1(n19630), .A2(BUF2_REG_30__SCAN_IN), .B1(n19631), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n13801) );
  AND2_X1 U15457 ( .A1(n13802), .A2(n13801), .ZN(n13803) );
  OAI21_X1 U15458 ( .B1(n15303), .B2(n19579), .A(n13803), .ZN(P2_U2889) );
  INV_X1 U15459 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20095) );
  INV_X1 U15460 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22277) );
  NOR4_X1 U15461 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20095), .A4(n22277), .ZN(n13805) );
  NOR4_X1 U15462 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13804) );
  NAND3_X1 U15463 ( .A1(n14377), .A2(n13805), .A3(n13804), .ZN(U214) );
  NOR2_X1 U15464 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n13807) );
  NOR4_X1 U15465 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13806) );
  NAND4_X1 U15466 ( .A1(n13807), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n13806), .ZN(n13808) );
  NOR2_X1 U15467 ( .A1(n14088), .A2(n13808), .ZN(n20027) );
  NAND2_X1 U15468 ( .A1(n20027), .A2(U214), .ZN(U212) );
  NOR2_X1 U15469 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13808), .ZN(n18649)
         );
  INV_X1 U15470 ( .A(n18619), .ZN(n18616) );
  OR2_X1 U15471 ( .A1(n14538), .A2(n18616), .ZN(n13817) );
  INV_X1 U15472 ( .A(n13817), .ZN(n13810) );
  INV_X1 U15473 ( .A(n14115), .ZN(n13809) );
  NAND2_X1 U15474 ( .A1(n13810), .A2(n13809), .ZN(n18241) );
  INV_X1 U15475 ( .A(n18241), .ZN(n13815) );
  INV_X1 U15476 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n17237) );
  NAND2_X1 U15477 ( .A1(n19304), .A2(n15263), .ZN(n13819) );
  INV_X1 U15478 ( .A(n14551), .ZN(n13811) );
  OR2_X1 U15479 ( .A1(n13812), .A2(n13811), .ZN(n13813) );
  NOR2_X1 U15480 ( .A1(n14538), .A2(n13813), .ZN(n13981) );
  INV_X1 U15481 ( .A(n13981), .ZN(n13814) );
  OAI211_X1 U15482 ( .C1(n13815), .C2(n17237), .A(n13819), .B(n13814), .ZN(
        P2_U2814) );
  INV_X1 U15483 ( .A(n14536), .ZN(n13816) );
  NOR2_X1 U15484 ( .A1(n18221), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13820)
         );
  INV_X1 U15485 ( .A(n13585), .ZN(n13818) );
  AOI22_X1 U15486 ( .A1(n13820), .A2(n13819), .B1(n13818), .B2(n18221), .ZN(
        P2_U3612) );
  AND2_X1 U15487 ( .A1(n13822), .A2(n11134), .ZN(n13823) );
  AOI21_X1 U15488 ( .B1(n13821), .B2(n15579), .A(n13823), .ZN(n15581) );
  INV_X1 U15489 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n16996) );
  AOI21_X1 U15490 ( .B1(n15581), .B2(n15582), .A(n16996), .ZN(n13825) );
  INV_X1 U15491 ( .A(n16813), .ZN(n21645) );
  NOR3_X1 U15492 ( .A1(n21645), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n21655), 
        .ZN(n13824) );
  OR2_X1 U15493 ( .A1(n13825), .A2(n13824), .ZN(P1_U2803) );
  AND2_X1 U15494 ( .A1(n21900), .A2(n16886), .ZN(n14745) );
  AOI21_X1 U15495 ( .B1(n13826), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14745), 
        .ZN(n13827) );
  NAND2_X1 U15496 ( .A1(n14259), .A2(n13827), .ZN(P1_U2801) );
  NAND4_X1 U15497 ( .A1(n13830), .A2(n13829), .A3(n13828), .A4(n13838), .ZN(
        n13831) );
  NAND2_X1 U15498 ( .A1(n13831), .A2(n15263), .ZN(n13832) );
  OR2_X1 U15499 ( .A1(n14538), .A2(n13832), .ZN(n13836) );
  NAND2_X1 U15500 ( .A1(n14502), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13833) );
  NAND2_X1 U15501 ( .A1(n13833), .A2(n13917), .ZN(n13915) );
  INV_X1 U15502 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18624) );
  OAI21_X1 U15503 ( .B1(n13834), .B2(n13915), .A(n18624), .ZN(n13835) );
  NAND2_X1 U15504 ( .A1(n13835), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17209) );
  NAND2_X1 U15505 ( .A1(n13836), .A2(n17209), .ZN(n16836) );
  AND2_X1 U15506 ( .A1(n14101), .A2(n11085), .ZN(n14525) );
  NAND2_X1 U15507 ( .A1(n16836), .A2(n14525), .ZN(n13847) );
  MUX2_X1 U15508 ( .A(n13867), .B(n13838), .S(n13837), .Z(n13849) );
  NAND2_X1 U15509 ( .A1(n11085), .A2(n15034), .ZN(n13840) );
  NAND2_X1 U15510 ( .A1(n13840), .A2(n13839), .ZN(n13880) );
  AOI21_X1 U15511 ( .B1(n13849), .B2(n13841), .A(n13880), .ZN(n13842) );
  NOR2_X1 U15512 ( .A1(n13843), .A2(n13842), .ZN(n13845) );
  OR2_X1 U15513 ( .A1(n13845), .A2(n13844), .ZN(n14526) );
  INV_X1 U15514 ( .A(n14526), .ZN(n13846) );
  AND2_X1 U15515 ( .A1(n19585), .A2(n14727), .ZN(n14553) );
  AND2_X1 U15516 ( .A1(n14101), .A2(n14553), .ZN(n14527) );
  NAND2_X1 U15517 ( .A1(n13846), .A2(n14527), .ZN(n14106) );
  NAND2_X1 U15518 ( .A1(n13847), .A2(n14106), .ZN(n14543) );
  NAND2_X1 U15519 ( .A1(n14543), .A2(n18619), .ZN(n18623) );
  NAND2_X1 U15520 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n16835) );
  NAND3_X1 U15521 ( .A1(n14714), .A2(n17222), .A3(n16835), .ZN(n13848) );
  AND2_X1 U15522 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n16832) );
  OR2_X1 U15523 ( .A1(n18623), .A2(n19585), .ZN(n17156) );
  MUX2_X1 U15524 ( .A(n13849), .B(P2_EBX_REG_0__SCAN_IN), .S(n19381), .Z(
        n18237) );
  XNOR2_X1 U15525 ( .A(n18237), .B(n16783), .ZN(n18507) );
  OR2_X1 U15526 ( .A1(n19290), .A2(n18595), .ZN(n14141) );
  NAND2_X1 U15527 ( .A1(n18559), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n18510) );
  INV_X1 U15528 ( .A(n18510), .ZN(n13853) );
  OR2_X1 U15529 ( .A1(n18623), .A2(n14142), .ZN(n17152) );
  AND2_X1 U15530 ( .A1(n19585), .A2(n13867), .ZN(n13885) );
  INV_X1 U15531 ( .A(n13885), .ZN(n13850) );
  NAND2_X1 U15532 ( .A1(n13850), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13886) );
  NAND2_X1 U15533 ( .A1(n13885), .A2(n16783), .ZN(n13851) );
  NAND2_X1 U15534 ( .A1(n13886), .A2(n13851), .ZN(n18509) );
  NOR2_X1 U15535 ( .A1(n17152), .A2(n18509), .ZN(n13852) );
  AOI211_X1 U15536 ( .C1(n17202), .C2(n18507), .A(n13853), .B(n13852), .ZN(
        n13857) );
  INV_X1 U15537 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n13854) );
  NAND2_X1 U15538 ( .A1(n13854), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13855) );
  NAND2_X1 U15539 ( .A1(n14557), .A2(n13855), .ZN(n13870) );
  OAI21_X1 U15540 ( .B1(n17200), .B2(n13870), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13856) );
  OAI211_X1 U15541 ( .C1(n17207), .C2(n18511), .A(n13857), .B(n13856), .ZN(
        P2_U3014) );
  INV_X1 U15542 ( .A(n13858), .ZN(n13860) );
  OAI21_X1 U15543 ( .B1(n14745), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13860), 
        .ZN(n13859) );
  OAI21_X1 U15544 ( .B1(n13861), .B2(n13860), .A(n13859), .ZN(P1_U3487) );
  INV_X1 U15545 ( .A(n18237), .ZN(n13862) );
  NOR2_X1 U15546 ( .A1(n13862), .A2(n16783), .ZN(n13865) );
  NOR2_X1 U15547 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n13863) );
  MUX2_X1 U15548 ( .A(n13863), .B(n13884), .S(n15490), .Z(n13881) );
  AND3_X1 U15549 ( .A1(n19381), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n13864) );
  NOR2_X1 U15550 ( .A1(n13881), .A2(n13864), .ZN(n16165) );
  AND2_X1 U15551 ( .A1(n13865), .A2(n16165), .ZN(n13876) );
  NOR2_X1 U15552 ( .A1(n13865), .A2(n16165), .ZN(n13878) );
  NOR2_X1 U15553 ( .A1(n13876), .A2(n13878), .ZN(n13866) );
  XNOR2_X1 U15554 ( .A(n13866), .B(n16789), .ZN(n14140) );
  INV_X1 U15555 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13873) );
  XNOR2_X1 U15556 ( .A(n13884), .B(n13867), .ZN(n13887) );
  XNOR2_X1 U15557 ( .A(n13887), .B(n13886), .ZN(n13868) );
  NOR2_X1 U15558 ( .A1(n16789), .A2(n13868), .ZN(n13888) );
  AOI21_X1 U15559 ( .B1(n16789), .B2(n13868), .A(n13888), .ZN(n14151) );
  NOR2_X1 U15560 ( .A1(n14141), .A2(n13869), .ZN(n14139) );
  AOI21_X1 U15561 ( .B1(n17203), .B2(n14151), .A(n14139), .ZN(n13872) );
  NAND2_X1 U15562 ( .A1(n17163), .A2(n13873), .ZN(n13871) );
  OAI211_X1 U15563 ( .C1(n17151), .C2(n13873), .A(n13872), .B(n13871), .ZN(
        n13874) );
  AOI21_X1 U15564 ( .B1(n17202), .B2(n14140), .A(n13874), .ZN(n13875) );
  OAI21_X1 U15565 ( .B1(n10973), .B2(n17207), .A(n13875), .ZN(P2_U3013) );
  INV_X1 U15566 ( .A(n14995), .ZN(n14986) );
  NOR2_X1 U15567 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13876), .ZN(
        n13877) );
  NOR2_X1 U15568 ( .A1(n13878), .A2(n13877), .ZN(n15040) );
  INV_X1 U15569 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13879) );
  MUX2_X1 U15570 ( .A(n13880), .B(n13879), .S(n19381), .Z(n13882) );
  NAND2_X1 U15571 ( .A1(n13882), .A2(n13881), .ZN(n14721) );
  OAI21_X1 U15572 ( .B1(n13882), .B2(n13881), .A(n14721), .ZN(n16156) );
  XNOR2_X1 U15573 ( .A(n16156), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15039) );
  INV_X1 U15574 ( .A(n15039), .ZN(n13883) );
  XNOR2_X1 U15575 ( .A(n15040), .B(n13883), .ZN(n18583) );
  OAI21_X1 U15576 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n14712), .ZN(n16150) );
  AND2_X1 U15577 ( .A1(n13885), .A2(n13884), .ZN(n15035) );
  XOR2_X1 U15578 ( .A(n15034), .B(n15035), .Z(n13891) );
  INV_X1 U15579 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18593) );
  NOR2_X1 U15580 ( .A1(n13887), .A2(n13886), .ZN(n13889) );
  NOR2_X1 U15581 ( .A1(n13889), .A2(n13888), .ZN(n15047) );
  XNOR2_X1 U15582 ( .A(n18593), .B(n15047), .ZN(n13890) );
  NOR2_X1 U15583 ( .A1(n13891), .A2(n13890), .ZN(n15049) );
  AOI21_X1 U15584 ( .B1(n13891), .B2(n13890), .A(n15049), .ZN(n18569) );
  INV_X1 U15585 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16152) );
  OAI22_X1 U15586 ( .A1(n17151), .A2(n16152), .B1(n18577), .B2(n14141), .ZN(
        n13892) );
  AOI21_X1 U15587 ( .B1(n18569), .B2(n17203), .A(n13892), .ZN(n13893) );
  OAI21_X1 U15588 ( .B1(n16150), .B2(n17198), .A(n13893), .ZN(n13894) );
  AOI21_X1 U15589 ( .B1(n18583), .B2(n17202), .A(n13894), .ZN(n13895) );
  OAI21_X1 U15590 ( .B1(n16157), .B2(n17207), .A(n13895), .ZN(P2_U3012) );
  INV_X1 U15591 ( .A(n14561), .ZN(n14524) );
  INV_X1 U15592 ( .A(n13896), .ZN(n13897) );
  NAND2_X1 U15593 ( .A1(n13897), .A2(n13578), .ZN(n14474) );
  INV_X1 U15594 ( .A(n14474), .ZN(n14531) );
  NAND2_X1 U15595 ( .A1(n14524), .A2(n14531), .ZN(n13966) );
  INV_X1 U15596 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n17269) );
  NAND2_X1 U15597 ( .A1(n17269), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21702) );
  INV_X1 U15598 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21713) );
  NAND2_X2 U15599 ( .A1(n17281), .A2(n21713), .ZN(n17284) );
  NOR2_X1 U15600 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n16829) );
  NAND2_X1 U15601 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n16829), .ZN(n17268) );
  NAND2_X1 U15602 ( .A1(n17284), .A2(n17268), .ZN(n18228) );
  NAND2_X1 U15603 ( .A1(n18222), .A2(n18228), .ZN(n14552) );
  OR2_X1 U15604 ( .A1(n14555), .A2(n14552), .ZN(n13898) );
  OR2_X1 U15605 ( .A1(n14538), .A2(n13898), .ZN(n13909) );
  NAND2_X1 U15606 ( .A1(n13899), .A2(n19534), .ZN(n13907) );
  NAND2_X1 U15607 ( .A1(n13905), .A2(n13968), .ZN(n13900) );
  AND2_X1 U15608 ( .A1(n13900), .A2(n14553), .ZN(n14127) );
  NAND2_X1 U15609 ( .A1(n13901), .A2(n19585), .ZN(n13902) );
  OAI211_X1 U15610 ( .C1(n19642), .C2(n11083), .A(n13902), .B(n19534), .ZN(
        n13904) );
  OAI211_X1 U15611 ( .C1(n12953), .C2(n13905), .A(n13904), .B(n13903), .ZN(
        n13906) );
  AOI211_X1 U15612 ( .C1(n14115), .C2(n13907), .A(n14127), .B(n13906), .ZN(
        n13908) );
  AND2_X1 U15613 ( .A1(n13909), .A2(n13908), .ZN(n14107) );
  NAND3_X1 U15614 ( .A1(n13910), .A2(n13966), .A3(n14107), .ZN(n13913) );
  NAND2_X1 U15615 ( .A1(n14561), .A2(n14142), .ZN(n14112) );
  OR2_X1 U15616 ( .A1(n14115), .A2(n14552), .ZN(n13911) );
  NOR2_X1 U15617 ( .A1(n14112), .A2(n13911), .ZN(n13912) );
  NOR2_X1 U15618 ( .A1(n13913), .A2(n13912), .ZN(n14522) );
  INV_X1 U15619 ( .A(n16835), .ZN(n17208) );
  NAND2_X1 U15620 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17208), .ZN(n16837) );
  INV_X1 U15621 ( .A(n16837), .ZN(n16833) );
  NOR2_X1 U15622 ( .A1(n17222), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14559) );
  AOI21_X1 U15623 ( .B1(n16833), .B2(P2_FLUSH_REG_SCAN_IN), .A(n14559), .ZN(
        n13914) );
  OAI21_X1 U15624 ( .B1(n14522), .B2(n18616), .A(n13914), .ZN(n16792) );
  INV_X1 U15625 ( .A(n16792), .ZN(n16799) );
  INV_X1 U15626 ( .A(n13915), .ZN(n14540) );
  NAND2_X1 U15627 ( .A1(n15263), .A2(n17222), .ZN(n18596) );
  OR2_X1 U15628 ( .A1(n14115), .A2(n14142), .ZN(n14539) );
  OR4_X1 U15629 ( .A1(n16799), .A2(n14540), .A3(n18596), .A4(n14539), .ZN(
        n13916) );
  OAI21_X1 U15630 ( .B1(n13917), .B2(n16792), .A(n13916), .ZN(P2_U3595) );
  INV_X1 U15631 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13921) );
  OR2_X1 U15632 ( .A1(n14115), .A2(n18616), .ZN(n13918) );
  NAND2_X1 U15633 ( .A1(n13981), .A2(n19585), .ZN(n14095) );
  OAI21_X1 U15634 ( .B1(n14112), .B2(n13918), .A(n14095), .ZN(n13919) );
  AND2_X1 U15635 ( .A1(n13919), .A2(n18228), .ZN(n17241) );
  NAND2_X1 U15636 ( .A1(n17241), .A2(n13031), .ZN(n14208) );
  NOR2_X1 U15637 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16835), .ZN(n17256) );
  AOI22_X1 U15638 ( .A1(n17256), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17254), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13920) );
  OAI21_X1 U15639 ( .B1(n13921), .B2(n14208), .A(n13920), .ZN(P2_U2933) );
  INV_X1 U15640 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13923) );
  AOI22_X1 U15641 ( .A1(n17256), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17254), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13922) );
  OAI21_X1 U15642 ( .B1(n13923), .B2(n14208), .A(n13922), .ZN(P2_U2934) );
  INV_X1 U15643 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21837) );
  INV_X1 U15644 ( .A(n13821), .ZN(n13925) );
  NOR2_X1 U15645 ( .A1(n21692), .A2(n21691), .ZN(n13924) );
  NAND2_X1 U15646 ( .A1(n13925), .A2(n13924), .ZN(n16875) );
  NAND2_X1 U15647 ( .A1(n11577), .A2(n11685), .ZN(n16081) );
  AND2_X1 U15648 ( .A1(n16081), .A2(n14069), .ZN(n13926) );
  OR2_X1 U15649 ( .A1(n16875), .A2(n13926), .ZN(n13945) );
  INV_X1 U15650 ( .A(n13927), .ZN(n13942) );
  NOR2_X1 U15651 ( .A1(n15578), .A2(n11695), .ZN(n13928) );
  NAND2_X1 U15652 ( .A1(n13928), .A2(n16079), .ZN(n15575) );
  INV_X1 U15653 ( .A(n15575), .ZN(n13929) );
  NAND2_X1 U15654 ( .A1(n13821), .A2(n13929), .ZN(n13941) );
  INV_X1 U15655 ( .A(n11577), .ZN(n13937) );
  AND2_X1 U15656 ( .A1(n13930), .A2(n14404), .ZN(n14054) );
  INV_X1 U15657 ( .A(n14054), .ZN(n13931) );
  AND2_X1 U15658 ( .A1(n13931), .A2(n11688), .ZN(n13932) );
  NAND2_X1 U15659 ( .A1(n13933), .A2(n13932), .ZN(n13949) );
  NAND4_X1 U15660 ( .A1(n13949), .A2(n13935), .A3(n13951), .A4(n13934), .ZN(
        n13936) );
  NAND2_X1 U15661 ( .A1(n13937), .A2(n13936), .ZN(n14058) );
  OAI211_X1 U15662 ( .C1(n14598), .C2(n14056), .A(n13938), .B(n14058), .ZN(
        n13939) );
  INV_X1 U15663 ( .A(n13939), .ZN(n13940) );
  OAI211_X1 U15664 ( .C1(n13821), .C2(n13942), .A(n13941), .B(n13940), .ZN(
        n13943) );
  INV_X1 U15665 ( .A(n13943), .ZN(n13944) );
  NAND2_X1 U15666 ( .A1(n13945), .A2(n13944), .ZN(n14285) );
  NAND2_X1 U15667 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n21654) );
  NOR2_X1 U15668 ( .A1(n21655), .A2(n21654), .ZN(n14295) );
  AOI22_X1 U15669 ( .A1(n15582), .A2(n14285), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n14295), .ZN(n16817) );
  OAI21_X1 U15670 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21837), .A(n16817), 
        .ZN(n21647) );
  NAND2_X1 U15671 ( .A1(n11693), .A2(n11689), .ZN(n13947) );
  AND2_X1 U15672 ( .A1(n13947), .A2(n13946), .ZN(n13948) );
  OAI211_X1 U15673 ( .C1(n13951), .C2(n13950), .A(n13949), .B(n13948), .ZN(
        n13952) );
  INV_X1 U15674 ( .A(n13952), .ZN(n13953) );
  NAND2_X1 U15675 ( .A1(n13953), .A2(n11047), .ZN(n14076) );
  NAND2_X1 U15676 ( .A1(n13954), .A2(n11680), .ZN(n13955) );
  OR2_X1 U15677 ( .A1(n14076), .A2(n13955), .ZN(n16083) );
  NOR2_X1 U15678 ( .A1(n13956), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13957) );
  INV_X1 U15679 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U15680 ( .A1(n13961), .A2(n21658), .B1(n14078), .B2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n13958) );
  OAI21_X1 U15681 ( .B1(n16854), .B2(n21645), .A(n13958), .ZN(n13959) );
  NOR2_X1 U15682 ( .A1(n16081), .A2(n13961), .ZN(n16852) );
  AOI22_X1 U15683 ( .A1(n21647), .A2(n13959), .B1(n16813), .B2(n16852), .ZN(
        n13960) );
  OAI21_X1 U15684 ( .B1(n21647), .B2(n13961), .A(n13960), .ZN(P1_U3474) );
  NAND2_X1 U15685 ( .A1(n14142), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13962) );
  AND4_X1 U15686 ( .A1(n13035), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13962), 
        .A4(n17222), .ZN(n13963) );
  INV_X1 U15687 ( .A(n13965), .ZN(n14470) );
  NAND2_X1 U15688 ( .A1(n13966), .A2(n14470), .ZN(n13967) );
  NAND2_X1 U15689 ( .A1(n11059), .A2(n13968), .ZN(n16253) );
  INV_X1 U15690 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13969) );
  MUX2_X1 U15691 ( .A(n18511), .B(n13969), .S(n10963), .Z(n13970) );
  OAI21_X1 U15692 ( .B1(n19141), .B2(n16253), .A(n13970), .ZN(P2_U2887) );
  INV_X1 U15693 ( .A(n16083), .ZN(n13974) );
  OR2_X1 U15694 ( .A1(n21877), .A2(n13974), .ZN(n13976) );
  XNOR2_X1 U15695 ( .A(n16085), .B(n13979), .ZN(n13977) );
  AND2_X1 U15696 ( .A1(n14268), .A2(n13977), .ZN(n13973) );
  XNOR2_X1 U15697 ( .A(n11531), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13971) );
  AND2_X1 U15698 ( .A1(n15567), .A2(n15575), .ZN(n14275) );
  OAI22_X1 U15699 ( .A1(n16081), .A2(n13971), .B1(n14275), .B2(n13977), .ZN(
        n13972) );
  AOI21_X1 U15700 ( .B1(n13974), .B2(n13973), .A(n13972), .ZN(n13975) );
  NAND2_X1 U15701 ( .A1(n13976), .A2(n13975), .ZN(n14265) );
  NOR2_X1 U15702 ( .A1(n16886), .A2(n14078), .ZN(n16087) );
  AOI22_X1 U15703 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n15946), .B2(n14616), .ZN(
        n16084) );
  AOI222_X1 U15704 ( .A1(n14265), .A2(n16813), .B1(n16087), .B2(n16084), .C1(
        n13977), .C2(n21658), .ZN(n13978) );
  MUX2_X1 U15705 ( .A(n13979), .B(n13978), .S(n21647), .Z(n13980) );
  INV_X1 U15706 ( .A(n13980), .ZN(P1_U3472) );
  AND2_X1 U15707 ( .A1(n13981), .A2(n18222), .ZN(n13983) );
  INV_X1 U15708 ( .A(n13983), .ZN(n13982) );
  INV_X1 U15709 ( .A(n14091), .ZN(n13985) );
  AOI22_X1 U15710 ( .A1(n19109), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19108), .ZN(n19079) );
  INV_X2 U15711 ( .A(n14095), .ZN(n14044) );
  OR2_X1 U15712 ( .A1(n14044), .A2(n13983), .ZN(n13997) );
  INV_X1 U15713 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13984) );
  INV_X1 U15714 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19080) );
  OAI222_X1 U15715 ( .A1(n13985), .A2(n19079), .B1(n13997), .B2(n13984), .C1(
        n14095), .C2(n19080), .ZN(P2_U2982) );
  NOR2_X1 U15716 ( .A1(n11696), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13987) );
  NOR2_X1 U15717 ( .A1(n13987), .A2(n13986), .ZN(n21434) );
  NOR2_X1 U15718 ( .A1(n15575), .A2(n21664), .ZN(n13988) );
  NAND2_X1 U15719 ( .A1(n13821), .A2(n13988), .ZN(n13991) );
  OR2_X1 U15720 ( .A1(n13989), .A2(n15578), .ZN(n13990) );
  INV_X1 U15721 ( .A(n13992), .ZN(n13994) );
  OAI21_X1 U15722 ( .B1(n13994), .B2(n11369), .A(n13993), .ZN(n21438) );
  OAI222_X1 U15723 ( .A1(n11375), .A2(n19942), .B1(n19946), .B2(n11590), .C1(
        n21438), .C2(n15726), .ZN(P1_U2872) );
  INV_X2 U15724 ( .A(n13997), .ZN(n14085) );
  AOI22_X1 U15725 ( .A1(n14085), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n14044), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13996) );
  AOI22_X1 U15726 ( .A1(n19109), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n14088), .ZN(n19093) );
  INV_X1 U15727 ( .A(n19093), .ZN(n13995) );
  NAND2_X1 U15728 ( .A1(n14091), .A2(n13995), .ZN(n14030) );
  NAND2_X1 U15729 ( .A1(n13996), .A2(n14030), .ZN(P2_U2978) );
  AOI22_X1 U15730 ( .A1(n14085), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n14044), .ZN(n13998) );
  OAI22_X1 U15731 ( .A1(n14088), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19109), .ZN(n19329) );
  INV_X1 U15732 ( .A(n19329), .ZN(n19321) );
  NAND2_X1 U15733 ( .A1(n14091), .A2(n19321), .ZN(n14045) );
  NAND2_X1 U15734 ( .A1(n13998), .A2(n14045), .ZN(P2_U2958) );
  AOI22_X1 U15735 ( .A1(n14085), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n14044), .ZN(n13999) );
  INV_X1 U15736 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20029) );
  INV_X1 U15737 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n20747) );
  AOI22_X1 U15738 ( .A1(n19109), .A2(n20029), .B1(n20747), .B2(n19108), .ZN(
        n19628) );
  NAND2_X1 U15739 ( .A1(n14091), .A2(n19628), .ZN(n14038) );
  NAND2_X1 U15740 ( .A1(n13999), .A2(n14038), .ZN(P2_U2952) );
  AOI22_X1 U15741 ( .A1(n14085), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n14044), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n14000) );
  INV_X1 U15742 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20033) );
  INV_X1 U15743 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n20130) );
  AOI22_X1 U15744 ( .A1(n19109), .A2(n20033), .B1(n20130), .B2(n19108), .ZN(
        n19532) );
  NAND2_X1 U15745 ( .A1(n14091), .A2(n19532), .ZN(n14028) );
  NAND2_X1 U15746 ( .A1(n14000), .A2(n14028), .ZN(P2_U2969) );
  AOI22_X1 U15747 ( .A1(n14085), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n14044), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n14002) );
  AOI22_X1 U15748 ( .A1(n19109), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14088), .ZN(n19477) );
  INV_X1 U15749 ( .A(n19477), .ZN(n14001) );
  NAND2_X1 U15750 ( .A1(n14091), .A2(n14001), .ZN(n14014) );
  NAND2_X1 U15751 ( .A1(n14002), .A2(n14014), .ZN(P2_U2955) );
  AOI22_X1 U15752 ( .A1(n14085), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n14044), .ZN(n14003) );
  INV_X1 U15753 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20037) );
  INV_X1 U15754 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n20643) );
  AOI22_X1 U15755 ( .A1(n19109), .A2(n20037), .B1(n20643), .B2(n19108), .ZN(
        n19428) );
  NAND2_X1 U15756 ( .A1(n14091), .A2(n19428), .ZN(n14016) );
  NAND2_X1 U15757 ( .A1(n14003), .A2(n14016), .ZN(P2_U2956) );
  AOI22_X1 U15758 ( .A1(n14085), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(n14044), .ZN(n14007) );
  OR2_X1 U15759 ( .A1(n14088), .A2(n20049), .ZN(n14005) );
  NAND2_X1 U15760 ( .A1(n19108), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14004) );
  AND2_X1 U15761 ( .A1(n14005), .A2(n14004), .ZN(n19096) );
  INV_X1 U15762 ( .A(n19096), .ZN(n14006) );
  NAND2_X1 U15763 ( .A1(n14091), .A2(n14006), .ZN(n14020) );
  NAND2_X1 U15764 ( .A1(n14007), .A2(n14020), .ZN(P2_U2977) );
  AOI22_X1 U15765 ( .A1(n14085), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n14044), .ZN(n14009) );
  AOI22_X1 U15766 ( .A1(n19109), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n14088), .ZN(n19103) );
  INV_X1 U15767 ( .A(n19103), .ZN(n14008) );
  NAND2_X1 U15768 ( .A1(n14091), .A2(n14008), .ZN(n14010) );
  NAND2_X1 U15769 ( .A1(n14009), .A2(n14010), .ZN(P2_U2975) );
  AOI22_X1 U15770 ( .A1(n14085), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n14044), .ZN(n14011) );
  NAND2_X1 U15771 ( .A1(n14011), .A2(n14010), .ZN(P2_U2960) );
  AOI22_X1 U15772 ( .A1(n14085), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n14044), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n14013) );
  AOI22_X1 U15773 ( .A1(n19109), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n19108), .ZN(n19099) );
  INV_X1 U15774 ( .A(n19099), .ZN(n14012) );
  NAND2_X1 U15775 ( .A1(n14091), .A2(n14012), .ZN(n14042) );
  NAND2_X1 U15776 ( .A1(n14013), .A2(n14042), .ZN(P2_U2961) );
  AOI22_X1 U15777 ( .A1(n14085), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n14044), .ZN(n14015) );
  NAND2_X1 U15778 ( .A1(n14015), .A2(n14014), .ZN(P2_U2970) );
  AOI22_X1 U15779 ( .A1(n14085), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n14044), .ZN(n14017) );
  NAND2_X1 U15780 ( .A1(n14017), .A2(n14016), .ZN(P2_U2971) );
  AOI22_X1 U15781 ( .A1(n14085), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n14044), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n14019) );
  AOI22_X1 U15782 ( .A1(n19109), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14088), .ZN(n19584) );
  INV_X1 U15783 ( .A(n19584), .ZN(n14018) );
  NAND2_X1 U15784 ( .A1(n14091), .A2(n14018), .ZN(n14026) );
  NAND2_X1 U15785 ( .A1(n14019), .A2(n14026), .ZN(P2_U2953) );
  AOI22_X1 U15786 ( .A1(n14085), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_26__SCAN_IN), .B2(n14044), .ZN(n14021) );
  NAND2_X1 U15787 ( .A1(n14021), .A2(n14020), .ZN(P2_U2962) );
  AOI22_X1 U15788 ( .A1(n14085), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n14044), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n14023) );
  AOI22_X1 U15789 ( .A1(n19109), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14088), .ZN(n19113) );
  INV_X1 U15790 ( .A(n19113), .ZN(n14022) );
  NAND2_X1 U15791 ( .A1(n14091), .A2(n14022), .ZN(n14024) );
  NAND2_X1 U15792 ( .A1(n14023), .A2(n14024), .ZN(P2_U2974) );
  AOI22_X1 U15793 ( .A1(n14085), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n14044), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n14025) );
  NAND2_X1 U15794 ( .A1(n14025), .A2(n14024), .ZN(P2_U2959) );
  AOI22_X1 U15795 ( .A1(n14085), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n14044), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n14027) );
  NAND2_X1 U15796 ( .A1(n14027), .A2(n14026), .ZN(P2_U2968) );
  AOI22_X1 U15797 ( .A1(n14085), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n14044), .ZN(n14029) );
  NAND2_X1 U15798 ( .A1(n14029), .A2(n14028), .ZN(P2_U2954) );
  AOI22_X1 U15799 ( .A1(n14085), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n14044), .ZN(n14031) );
  NAND2_X1 U15800 ( .A1(n14031), .A2(n14030), .ZN(P2_U2963) );
  AOI22_X1 U15801 ( .A1(n14085), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n14044), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n14033) );
  AOI22_X1 U15802 ( .A1(n19109), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19108), .ZN(n19379) );
  INV_X1 U15803 ( .A(n19379), .ZN(n14032) );
  NAND2_X1 U15804 ( .A1(n14091), .A2(n14032), .ZN(n14040) );
  NAND2_X1 U15805 ( .A1(n14033), .A2(n14040), .ZN(P2_U2972) );
  AOI22_X1 U15806 ( .A1(n14085), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n14044), .ZN(n14035) );
  AOI22_X1 U15807 ( .A1(n19109), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19108), .ZN(n19087) );
  INV_X1 U15808 ( .A(n19087), .ZN(n14034) );
  NAND2_X1 U15809 ( .A1(n14091), .A2(n14034), .ZN(n14036) );
  NAND2_X1 U15810 ( .A1(n14035), .A2(n14036), .ZN(P2_U2980) );
  AOI22_X1 U15811 ( .A1(n14085), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n14044), .ZN(n14037) );
  NAND2_X1 U15812 ( .A1(n14037), .A2(n14036), .ZN(P2_U2965) );
  AOI22_X1 U15813 ( .A1(n14085), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n14044), .ZN(n14039) );
  NAND2_X1 U15814 ( .A1(n14039), .A2(n14038), .ZN(P2_U2967) );
  AOI22_X1 U15815 ( .A1(n14085), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n14044), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n14041) );
  NAND2_X1 U15816 ( .A1(n14041), .A2(n14040), .ZN(P2_U2957) );
  AOI22_X1 U15817 ( .A1(n14085), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n14044), .ZN(n14043) );
  NAND2_X1 U15818 ( .A1(n14043), .A2(n14042), .ZN(P2_U2976) );
  AOI22_X1 U15819 ( .A1(n14085), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n14044), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n14046) );
  NAND2_X1 U15820 ( .A1(n14046), .A2(n14045), .ZN(P2_U2973) );
  OR2_X1 U15821 ( .A1(n14047), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14048) );
  NAND2_X1 U15822 ( .A1(n14049), .A2(n14048), .ZN(n14178) );
  NAND2_X1 U15823 ( .A1(n14050), .A2(n21683), .ZN(n14052) );
  OAI211_X1 U15824 ( .C1(n14069), .C2(n14052), .A(n11688), .B(n14051), .ZN(
        n14053) );
  NAND3_X1 U15825 ( .A1(n12393), .A2(n14568), .A3(n14053), .ZN(n14062) );
  NAND2_X1 U15826 ( .A1(n13821), .A2(n14054), .ZN(n14059) );
  NAND2_X1 U15827 ( .A1(n11685), .A2(n21692), .ZN(n14055) );
  NAND4_X1 U15828 ( .A1(n15571), .A2(n14056), .A3(n21683), .A4(n14055), .ZN(
        n14057) );
  NAND3_X1 U15829 ( .A1(n14059), .A2(n14058), .A3(n14057), .ZN(n14060) );
  NAND2_X1 U15830 ( .A1(n14060), .A2(n15582), .ZN(n14061) );
  OAI211_X1 U15831 ( .C1(n11682), .C2(n14064), .A(n14063), .B(n15567), .ZN(
        n14065) );
  NOR2_X1 U15832 ( .A1(n14065), .A2(n16868), .ZN(n14066) );
  AND2_X1 U15833 ( .A1(n13954), .A2(n14066), .ZN(n14067) );
  NAND2_X1 U15834 ( .A1(n14070), .A2(n11682), .ZN(n14071) );
  AND2_X1 U15835 ( .A1(n16880), .A2(n14071), .ZN(n14072) );
  AND2_X1 U15836 ( .A1(n14073), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14180) );
  INV_X1 U15837 ( .A(n14074), .ZN(n14075) );
  NOR2_X1 U15838 ( .A1(n14076), .A2(n14075), .ZN(n14077) );
  NAND2_X1 U15839 ( .A1(n21368), .A2(n15942), .ZN(n15945) );
  NAND2_X1 U15840 ( .A1(n14078), .A2(n15945), .ZN(n14211) );
  INV_X1 U15841 ( .A(n14211), .ZN(n14079) );
  AOI211_X1 U15842 ( .C1(n21421), .C2(n21434), .A(n14180), .B(n14079), .ZN(
        n14083) );
  NAND2_X1 U15843 ( .A1(n14080), .A2(n21419), .ZN(n14615) );
  INV_X1 U15844 ( .A(n14615), .ZN(n14081) );
  OAI21_X1 U15845 ( .B1(n14614), .B2(n14081), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14082) );
  OAI211_X1 U15846 ( .C1(n14178), .C2(n21382), .A(n14083), .B(n14082), .ZN(
        P1_U3031) );
  INV_X1 U15847 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n17263) );
  NAND2_X1 U15848 ( .A1(n14085), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n14084) );
  NAND2_X1 U15849 ( .A1(n14091), .A2(n19083), .ZN(n14086) );
  OAI211_X1 U15850 ( .C1(n17263), .C2(n14095), .A(n14084), .B(n14086), .ZN(
        P2_U2981) );
  NAND2_X1 U15851 ( .A1(n14085), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14087) );
  OAI211_X1 U15852 ( .C1(n13796), .C2(n14095), .A(n14087), .B(n14086), .ZN(
        P2_U2966) );
  INV_X1 U15853 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14188) );
  NAND2_X1 U15854 ( .A1(n14085), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14092) );
  NAND2_X1 U15855 ( .A1(n19108), .A2(BUF2_REG_12__SCAN_IN), .ZN(n14090) );
  INV_X1 U15856 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20053) );
  OR2_X1 U15857 ( .A1(n14088), .A2(n20053), .ZN(n14089) );
  NAND2_X1 U15858 ( .A1(n14090), .A2(n14089), .ZN(n19090) );
  NAND2_X1 U15859 ( .A1(n14091), .A2(n19090), .ZN(n14093) );
  OAI211_X1 U15860 ( .C1(n14188), .C2(n14095), .A(n14092), .B(n14093), .ZN(
        P2_U2964) );
  INV_X1 U15861 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n17260) );
  NAND2_X1 U15862 ( .A1(n14085), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n14094) );
  OAI211_X1 U15863 ( .C1(n17260), .C2(n14095), .A(n14094), .B(n14093), .ZN(
        P2_U2979) );
  INV_X1 U15864 ( .A(n14552), .ZN(n14096) );
  NAND2_X1 U15865 ( .A1(n14097), .A2(n14096), .ZN(n14111) );
  OAI21_X1 U15866 ( .B1(n14098), .B2(n14727), .A(n12953), .ZN(n14099) );
  INV_X1 U15867 ( .A(n14099), .ZN(n14100) );
  NAND2_X1 U15868 ( .A1(n14100), .A2(n14112), .ZN(n14110) );
  NAND3_X1 U15869 ( .A1(n16836), .A2(n14101), .A3(n14142), .ZN(n14108) );
  MUX2_X1 U15870 ( .A(n19534), .B(n14555), .S(n14142), .Z(n14102) );
  INV_X1 U15871 ( .A(n14102), .ZN(n14103) );
  NAND2_X1 U15872 ( .A1(n14103), .A2(n18222), .ZN(n14104) );
  OR2_X1 U15873 ( .A1(n14538), .A2(n14104), .ZN(n14105) );
  AND4_X1 U15874 ( .A1(n14108), .A2(n14107), .A3(n14106), .A4(n14105), .ZN(
        n14109) );
  OAI211_X1 U15875 ( .C1(n14112), .C2(n14111), .A(n14110), .B(n14109), .ZN(
        n14113) );
  NAND2_X1 U15876 ( .A1(n14115), .A2(n14114), .ZN(n14118) );
  INV_X1 U15877 ( .A(n14116), .ZN(n14117) );
  OR2_X1 U15878 ( .A1(n14118), .A2(n14117), .ZN(n14504) );
  NAND2_X1 U15879 ( .A1(n14504), .A2(n19585), .ZN(n14120) );
  NAND2_X1 U15880 ( .A1(n14120), .A2(n14119), .ZN(n14121) );
  NAND2_X1 U15881 ( .A1(n14150), .A2(n14121), .ZN(n18512) );
  NAND2_X1 U15882 ( .A1(n13041), .A2(n14122), .ZN(n14123) );
  AND2_X1 U15883 ( .A1(n14123), .A2(n13585), .ZN(n14124) );
  NAND2_X1 U15884 ( .A1(n14125), .A2(n14124), .ZN(n14137) );
  NAND2_X1 U15885 ( .A1(n14126), .A2(n14142), .ZN(n14484) );
  INV_X1 U15886 ( .A(n14127), .ZN(n14128) );
  NAND2_X1 U15887 ( .A1(n14484), .A2(n14128), .ZN(n14130) );
  NAND2_X1 U15888 ( .A1(n14130), .A2(n14129), .ZN(n14134) );
  OAI22_X1 U15889 ( .A1(n13585), .A2(n12992), .B1(n19642), .B2(n19534), .ZN(
        n14131) );
  INV_X1 U15890 ( .A(n14131), .ZN(n14133) );
  NAND3_X1 U15891 ( .A1(n14134), .A2(n14133), .A3(n14132), .ZN(n14135) );
  AOI21_X1 U15892 ( .B1(n14137), .B2(n14136), .A(n14135), .ZN(n14498) );
  NAND2_X1 U15893 ( .A1(n14498), .A2(n14470), .ZN(n14138) );
  NOR2_X1 U15894 ( .A1(n18573), .A2(n18568), .ZN(n18517) );
  INV_X1 U15895 ( .A(n18517), .ZN(n18519) );
  NAND2_X1 U15896 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18567) );
  OAI211_X1 U15897 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n18519), .B(n18567), .ZN(n14155) );
  AOI21_X1 U15898 ( .B1(n18582), .B2(n14140), .A(n14139), .ZN(n14154) );
  NOR2_X1 U15900 ( .A1(n14150), .A2(n18559), .ZN(n18566) );
  NAND2_X1 U15901 ( .A1(n14536), .A2(n14142), .ZN(n14143) );
  NAND2_X1 U15902 ( .A1(n14474), .A2(n14143), .ZN(n14144) );
  NAND2_X1 U15903 ( .A1(n14150), .A2(n14144), .ZN(n18579) );
  INV_X1 U15904 ( .A(n14145), .ZN(n14147) );
  NAND2_X1 U15905 ( .A1(n14147), .A2(n14146), .ZN(n14148) );
  NAND2_X1 U15906 ( .A1(n14149), .A2(n14148), .ZN(n19575) );
  AOI22_X1 U15907 ( .A1(n18566), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n18553), .B2(n19575), .ZN(n14153) );
  NAND2_X1 U15908 ( .A1(n14150), .A2(n14527), .ZN(n18576) );
  NAND2_X1 U15909 ( .A1(n18556), .A2(n14151), .ZN(n14152) );
  AND4_X1 U15910 ( .A1(n14155), .A2(n14154), .A3(n14153), .A4(n14152), .ZN(
        n14156) );
  OAI21_X1 U15911 ( .B1(n10973), .B2(n18512), .A(n14156), .ZN(P2_U3045) );
  NAND2_X1 U15912 ( .A1(n16337), .A2(n14157), .ZN(n19524) );
  INV_X1 U15913 ( .A(n19628), .ZN(n19640) );
  INV_X1 U15914 ( .A(n14158), .ZN(n14164) );
  INV_X1 U15915 ( .A(n14159), .ZN(n14162) );
  INV_X1 U15916 ( .A(n14160), .ZN(n14161) );
  NAND2_X1 U15917 ( .A1(n14162), .A2(n14161), .ZN(n14163) );
  NAND2_X1 U15918 ( .A1(n14164), .A2(n14163), .ZN(n18508) );
  INV_X1 U15919 ( .A(n18508), .ZN(n18236) );
  NOR2_X1 U15920 ( .A1(n19141), .A2(n18508), .ZN(n19577) );
  INV_X1 U15921 ( .A(n19577), .ZN(n14165) );
  OAI211_X1 U15922 ( .C1(n19123), .C2(n18236), .A(n14165), .B(n19634), .ZN(
        n14167) );
  AOI22_X1 U15923 ( .A1(n19633), .A2(n18236), .B1(n19627), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n14166) );
  OAI211_X1 U15924 ( .C1(n19583), .C2(n19640), .A(n14167), .B(n14166), .ZN(
        P2_U2919) );
  NOR2_X1 U15925 ( .A1(n10973), .A2(n10963), .ZN(n14171) );
  AOI21_X1 U15926 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n10963), .A(n14171), .ZN(
        n14172) );
  OAI21_X1 U15927 ( .B1(n19142), .B2(n16253), .A(n14172), .ZN(P2_U2886) );
  XNOR2_X1 U15928 ( .A(n14173), .B(n15578), .ZN(n14665) );
  INV_X1 U15929 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14176) );
  OAI21_X1 U15930 ( .B1(n14175), .B2(n14174), .A(n14308), .ZN(n14670) );
  OAI222_X1 U15931 ( .A1(n14665), .A2(n19942), .B1(n14176), .B2(n19946), .C1(
        n14670), .C2(n15726), .ZN(P1_U2871) );
  NAND2_X1 U15932 ( .A1(n14177), .A2(n15898), .ZN(n14181) );
  NOR2_X1 U15933 ( .A1(n14178), .A2(n21639), .ZN(n14179) );
  AOI211_X1 U15934 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n14181), .A(
        n14180), .B(n14179), .ZN(n14182) );
  OAI21_X1 U15935 ( .B1(n19975), .B2(n21438), .A(n14182), .ZN(P1_U2999) );
  INV_X1 U15936 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14184) );
  AOI22_X1 U15937 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n17265), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17264), .ZN(n14183) );
  OAI21_X1 U15938 ( .B1(n14184), .B2(n14208), .A(n14183), .ZN(P2_U2935) );
  INV_X1 U15939 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14186) );
  AOI22_X1 U15940 ( .A1(n17265), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14185) );
  OAI21_X1 U15941 ( .B1(n14186), .B2(n14208), .A(n14185), .ZN(P2_U2924) );
  AOI22_X1 U15942 ( .A1(n17265), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14187) );
  OAI21_X1 U15943 ( .B1(n14188), .B2(n14208), .A(n14187), .ZN(P2_U2923) );
  INV_X1 U15944 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14190) );
  AOI22_X1 U15945 ( .A1(n17265), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14189) );
  OAI21_X1 U15946 ( .B1(n14190), .B2(n14208), .A(n14189), .ZN(P2_U2927) );
  INV_X1 U15947 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14192) );
  AOI22_X1 U15948 ( .A1(n17265), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14191) );
  OAI21_X1 U15949 ( .B1(n14192), .B2(n14208), .A(n14191), .ZN(P2_U2926) );
  INV_X1 U15950 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14194) );
  AOI22_X1 U15951 ( .A1(n17265), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14193) );
  OAI21_X1 U15952 ( .B1(n14194), .B2(n14208), .A(n14193), .ZN(P2_U2925) );
  INV_X1 U15953 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14196) );
  AOI22_X1 U15954 ( .A1(n17265), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14195) );
  OAI21_X1 U15955 ( .B1(n14196), .B2(n14208), .A(n14195), .ZN(P2_U2930) );
  INV_X1 U15956 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14198) );
  AOI22_X1 U15957 ( .A1(n17265), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14197) );
  OAI21_X1 U15958 ( .B1(n14198), .B2(n14208), .A(n14197), .ZN(P2_U2922) );
  INV_X1 U15959 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14200) );
  AOI22_X1 U15960 ( .A1(n17265), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14199) );
  OAI21_X1 U15961 ( .B1(n14200), .B2(n14208), .A(n14199), .ZN(P2_U2928) );
  INV_X1 U15962 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14202) );
  AOI22_X1 U15963 ( .A1(n17265), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14201) );
  OAI21_X1 U15964 ( .B1(n14202), .B2(n14208), .A(n14201), .ZN(P2_U2931) );
  INV_X1 U15965 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14204) );
  AOI22_X1 U15966 ( .A1(n17265), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14203) );
  OAI21_X1 U15967 ( .B1(n14204), .B2(n14208), .A(n14203), .ZN(P2_U2929) );
  INV_X1 U15968 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14206) );
  AOI22_X1 U15969 ( .A1(n17256), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14205) );
  OAI21_X1 U15970 ( .B1(n14206), .B2(n14208), .A(n14205), .ZN(P2_U2932) );
  AOI22_X1 U15971 ( .A1(n17256), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14207) );
  OAI21_X1 U15972 ( .B1(n13796), .B2(n14208), .A(n14207), .ZN(P2_U2921) );
  INV_X1 U15973 ( .A(n15945), .ZN(n14209) );
  AND2_X1 U15974 ( .A1(n16062), .A2(n14209), .ZN(n16032) );
  NOR2_X1 U15975 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14614), .ZN(
        n14618) );
  NOR3_X1 U15976 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16032), .A3(
        n14618), .ZN(n14214) );
  NOR2_X1 U15977 ( .A1(n21414), .A2(n14665), .ZN(n14213) );
  INV_X1 U15978 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n14210) );
  NOR2_X1 U15979 ( .A1(n21419), .A2(n14210), .ZN(n14249) );
  AOI21_X1 U15980 ( .B1(n14615), .B2(n14211), .A(n14616), .ZN(n14212) );
  NOR4_X1 U15981 ( .A1(n14214), .A2(n14213), .A3(n14249), .A4(n14212), .ZN(
        n14217) );
  OR2_X1 U15982 ( .A1(n14215), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14251) );
  NAND3_X1 U15983 ( .A1(n14251), .A2(n14250), .A3(n21422), .ZN(n14216) );
  NAND2_X1 U15984 ( .A1(n14217), .A2(n14216), .ZN(P1_U3030) );
  INV_X1 U15985 ( .A(DATAI_0_), .ZN(n16950) );
  NOR2_X1 U15986 ( .A1(n15727), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14219) );
  AOI21_X1 U15987 ( .B1(n16950), .B2(n15727), .A(n14219), .ZN(n15789) );
  INV_X1 U15988 ( .A(n15789), .ZN(n14220) );
  INV_X1 U15989 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19822) );
  OAI222_X1 U15990 ( .A1(n15796), .A2(n14220), .B1(n15794), .B2(n19822), .C1(
        n15801), .C2(n21438), .ZN(P1_U2904) );
  INV_X1 U15991 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20031) );
  NOR2_X1 U15992 ( .A1(n14377), .A2(DATAI_1_), .ZN(n14221) );
  AOI21_X1 U15993 ( .B1(n14377), .B2(n20031), .A(n14221), .ZN(n15782) );
  INV_X1 U15994 ( .A(n15782), .ZN(n14222) );
  INV_X1 U15995 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19824) );
  OAI222_X1 U15996 ( .A1(n15796), .A2(n14222), .B1(n15794), .B2(n19824), .C1(
        n15801), .C2(n14670), .ZN(P1_U2903) );
  INV_X1 U15997 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21749) );
  INV_X1 U15998 ( .A(n16880), .ZN(n14223) );
  INV_X1 U15999 ( .A(n16081), .ZN(n14224) );
  NAND2_X1 U16000 ( .A1(n12393), .A2(n14224), .ZN(n14225) );
  NAND2_X1 U16001 ( .A1(n21777), .A2(n14225), .ZN(n14227) );
  INV_X1 U16002 ( .A(n21692), .ZN(n14226) );
  NAND2_X1 U16003 ( .A1(n19820), .A2(n11688), .ZN(n14637) );
  NOR2_X1 U16004 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21654), .ZN(n14630) );
  AOI22_X1 U16005 ( .A1(n14630), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n14629), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14228) );
  OAI21_X1 U16006 ( .B1(n21749), .B2(n14637), .A(n14228), .ZN(P1_U2910) );
  INV_X1 U16007 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n21736) );
  AOI22_X1 U16008 ( .A1(n14630), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n14629), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14229) );
  OAI21_X1 U16009 ( .B1(n21736), .B2(n14637), .A(n14229), .ZN(P1_U2912) );
  INV_X1 U16010 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14231) );
  AOI22_X1 U16011 ( .A1(n14630), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n14629), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14230) );
  OAI21_X1 U16012 ( .B1(n14231), .B2(n14637), .A(n14230), .ZN(P1_U2917) );
  INV_X1 U16013 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14233) );
  AOI22_X1 U16014 ( .A1(n14630), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n14629), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14232) );
  OAI21_X1 U16015 ( .B1(n14233), .B2(n14637), .A(n14232), .ZN(P1_U2914) );
  INV_X1 U16016 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n21754) );
  AOI22_X1 U16017 ( .A1(n14630), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n14629), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14234) );
  OAI21_X1 U16018 ( .B1(n21754), .B2(n14637), .A(n14234), .ZN(P1_U2909) );
  INV_X1 U16019 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14236) );
  AOI22_X1 U16020 ( .A1(n14630), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n14629), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14235) );
  OAI21_X1 U16021 ( .B1(n14236), .B2(n14637), .A(n14235), .ZN(P1_U2915) );
  INV_X1 U16022 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21743) );
  AOI22_X1 U16023 ( .A1(n14630), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n14629), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14237) );
  OAI21_X1 U16024 ( .B1(n21743), .B2(n14637), .A(n14237), .ZN(P1_U2911) );
  INV_X1 U16025 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14239) );
  AOI22_X1 U16026 ( .A1(n14630), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n14629), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14238) );
  OAI21_X1 U16027 ( .B1(n14239), .B2(n14637), .A(n14238), .ZN(P1_U2919) );
  INV_X1 U16028 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n15768) );
  AOI22_X1 U16029 ( .A1(n14630), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n14629), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14240) );
  OAI21_X1 U16030 ( .B1(n15768), .B2(n14637), .A(n14240), .ZN(P1_U2916) );
  AOI22_X1 U16031 ( .A1(n21278), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n14629), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14241) );
  OAI21_X1 U16032 ( .B1(n15785), .B2(n14637), .A(n14241), .ZN(P1_U2920) );
  AOI22_X1 U16033 ( .A1(n21278), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n14629), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14242) );
  OAI21_X1 U16034 ( .B1(n12760), .B2(n14637), .A(n14242), .ZN(P1_U2906) );
  INV_X1 U16035 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n14732) );
  MUX2_X1 U16036 ( .A(n14732), .B(n17101), .S(n11059), .Z(n14247) );
  OAI21_X1 U16037 ( .B1(n19239), .B2(n16253), .A(n14247), .ZN(P2_U2884) );
  NOR2_X1 U16038 ( .A1(n20024), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14248) );
  AOI211_X1 U16039 ( .C1(n20014), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14249), .B(n14248), .ZN(n14253) );
  NAND3_X1 U16040 ( .A1(n14251), .A2(n14250), .A3(n20020), .ZN(n14252) );
  OAI211_X1 U16041 ( .C1(n19975), .C2(n14670), .A(n14253), .B(n14252), .ZN(
        P1_U2998) );
  MUX2_X1 U16042 ( .A(n13879), .B(n16157), .S(n11059), .Z(n14257) );
  OAI21_X1 U16043 ( .B1(n19238), .B2(n16253), .A(n14257), .ZN(P2_U2885) );
  INV_X1 U16044 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19844) );
  NOR2_X1 U16045 ( .A1(n21274), .A2(n21683), .ZN(n14258) );
  INV_X1 U16046 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14260) );
  OR2_X1 U16047 ( .A1(n15727), .A2(n14260), .ZN(n14262) );
  NAND2_X1 U16048 ( .A1(n15727), .A2(DATAI_15_), .ZN(n14261) );
  AND2_X1 U16049 ( .A1(n14262), .A2(n14261), .ZN(n15795) );
  INV_X1 U16050 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14263) );
  OAI222_X1 U16051 ( .A1(n21777), .A2(n19844), .B1(n21772), .B2(n15795), .C1(
        n14264), .C2(n14263), .ZN(P1_U2967) );
  MUX2_X1 U16052 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14265), .S(
        n14285), .Z(n16860) );
  INV_X1 U16053 ( .A(n14285), .ZN(n16856) );
  NAND2_X1 U16054 ( .A1(n16856), .A2(n11376), .ZN(n14282) );
  NAND2_X1 U16055 ( .A1(n16085), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14266) );
  NAND2_X1 U16056 ( .A1(n14266), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14267) );
  NAND2_X1 U16057 ( .A1(n11428), .A2(n14267), .ZN(n21642) );
  NAND2_X1 U16058 ( .A1(n14268), .A2(n21642), .ZN(n14279) );
  XNOR2_X1 U16059 ( .A(n14269), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14276) );
  INV_X1 U16060 ( .A(n14270), .ZN(n14271) );
  MUX2_X1 U16061 ( .A(n14271), .B(n11376), .S(n16085), .Z(n14273) );
  INV_X1 U16062 ( .A(n11422), .ZN(n14272) );
  NAND2_X1 U16063 ( .A1(n14273), .A2(n14272), .ZN(n14274) );
  OAI22_X1 U16064 ( .A1(n16081), .A2(n14276), .B1(n14275), .B2(n14274), .ZN(
        n14277) );
  INV_X1 U16065 ( .A(n14277), .ZN(n14278) );
  OAI21_X1 U16066 ( .B1(n16083), .B2(n14279), .A(n14278), .ZN(n14280) );
  AOI21_X1 U16067 ( .B1(n21829), .B2(n16083), .A(n14280), .ZN(n21646) );
  NAND2_X1 U16068 ( .A1(n21646), .A2(n14285), .ZN(n14281) );
  AND2_X1 U16069 ( .A1(n14282), .A2(n14281), .ZN(n16865) );
  NAND2_X1 U16070 ( .A1(n16860), .A2(n16865), .ZN(n14284) );
  NAND2_X1 U16071 ( .A1(n11422), .A2(n21640), .ZN(n14283) );
  MUX2_X1 U16072 ( .A(n14284), .B(n14283), .S(P1_STATE2_REG_1__SCAN_IN), .Z(
        n14292) );
  NAND2_X1 U16073 ( .A1(n14285), .A2(n16886), .ZN(n14291) );
  INV_X1 U16074 ( .A(n14381), .ZN(n21876) );
  OR2_X1 U16075 ( .A1(n14286), .A2(n21876), .ZN(n14287) );
  XNOR2_X1 U16076 ( .A(n14287), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n21457) );
  INV_X1 U16077 ( .A(n13954), .ZN(n14288) );
  AND2_X1 U16078 ( .A1(n21457), .A2(n14288), .ZN(n16814) );
  AND2_X1 U16079 ( .A1(n14291), .A2(n16815), .ZN(n14289) );
  AOI21_X1 U16080 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(P1_FLUSH_REG_SCAN_IN), 
        .A(n14289), .ZN(n14290) );
  OAI21_X1 U16081 ( .B1(n14291), .B2(n16814), .A(n14290), .ZN(n14293) );
  NAND2_X1 U16082 ( .A1(n14292), .A2(n14293), .ZN(n16874) );
  NAND2_X1 U16083 ( .A1(n14293), .A2(n11421), .ZN(n14294) );
  NAND2_X1 U16084 ( .A1(n16874), .A2(n14294), .ZN(n14314) );
  INV_X1 U16085 ( .A(n14314), .ZN(n14296) );
  OAI21_X1 U16086 ( .B1(n14296), .B2(P1_FLUSH_REG_SCAN_IN), .A(n14295), .ZN(
        n14297) );
  INV_X1 U16087 ( .A(n21659), .ZN(n21275) );
  NAND2_X1 U16088 ( .A1(n14297), .A2(n21783), .ZN(n16887) );
  AND2_X1 U16089 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21837), .ZN(n16075) );
  AND2_X1 U16090 ( .A1(n21900), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14299) );
  NAND2_X1 U16091 ( .A1(n16073), .A2(n14299), .ZN(n14372) );
  NAND2_X1 U16092 ( .A1(n16073), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14300) );
  INV_X1 U16093 ( .A(n21862), .ZN(n14369) );
  MUX2_X1 U16094 ( .A(n14372), .B(n14369), .S(n10975), .Z(n14301) );
  OAI21_X1 U16095 ( .B1(n16075), .B2(n21877), .A(n14301), .ZN(n14302) );
  NAND2_X1 U16096 ( .A1(n16887), .A2(n14302), .ZN(n14303) );
  OAI21_X1 U16097 ( .B1(n16887), .B2(n16851), .A(n14303), .ZN(P1_U3476) );
  OAI21_X1 U16098 ( .B1(n14306), .B2(n14305), .A(n14304), .ZN(n21297) );
  INV_X1 U16099 ( .A(n14308), .ZN(n14309) );
  XNOR2_X1 U16100 ( .A(n14307), .B(n14309), .ZN(n21451) );
  INV_X1 U16101 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21443) );
  NOR2_X1 U16102 ( .A1(n21419), .A2(n21443), .ZN(n21294) );
  AOI21_X1 U16103 ( .B1(n20014), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n21294), .ZN(n14310) );
  OAI21_X1 U16104 ( .B1(n20024), .B2(n21441), .A(n14310), .ZN(n14311) );
  AOI21_X1 U16105 ( .B1(n21451), .B2(n20021), .A(n14311), .ZN(n14312) );
  OAI21_X1 U16106 ( .B1(n21639), .B2(n21297), .A(n14312), .ZN(P1_U2997) );
  INV_X1 U16107 ( .A(n21654), .ZN(n14313) );
  AND2_X1 U16108 ( .A1(n14314), .A2(n14313), .ZN(n21662) );
  OAI22_X1 U16109 ( .A1(n12775), .A2(n21924), .B1(n14315), .B2(n16075), .ZN(
        n14316) );
  OAI21_X1 U16110 ( .B1(n21662), .B2(n14316), .A(n16887), .ZN(n14317) );
  OAI21_X1 U16111 ( .B1(n16887), .B2(n21892), .A(n14317), .ZN(P1_U3478) );
  INV_X1 U16112 ( .A(n21451), .ZN(n14417) );
  MUX2_X1 U16113 ( .A(BUF1_REG_2__SCAN_IN), .B(DATAI_2_), .S(n15727), .Z(
        n15777) );
  INV_X1 U16114 ( .A(n15777), .ZN(n14318) );
  INV_X1 U16115 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19826) );
  OAI222_X1 U16116 ( .A1(n14417), .A2(n15801), .B1(n15796), .B2(n14318), .C1(
        n15794), .C2(n19826), .ZN(P1_U2902) );
  XOR2_X1 U16117 ( .A(n14319), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14337)
         );
  INV_X1 U16118 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18248) );
  INV_X1 U16119 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15501) );
  OAI22_X1 U16120 ( .A1(n15264), .A2(n18248), .B1(n15263), .B2(n18249), .ZN(
        n14321) );
  AOI21_X1 U16121 ( .B1(n15294), .B2(P2_REIP_REG_5__SCAN_IN), .A(n14321), .ZN(
        n14322) );
  OAI21_X1 U16122 ( .B1(n15297), .B2(n15501), .A(n14322), .ZN(n14323) );
  INV_X1 U16123 ( .A(n14323), .ZN(n14335) );
  NAND2_X1 U16124 ( .A1(n14325), .A2(n14324), .ZN(n14329) );
  OR2_X1 U16125 ( .A1(n14327), .A2(n14326), .ZN(n14328) );
  NAND2_X1 U16126 ( .A1(n14329), .A2(n14328), .ZN(n14341) );
  INV_X1 U16127 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15502) );
  INV_X1 U16128 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14839) );
  INV_X1 U16129 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14844) );
  OAI22_X1 U16130 ( .A1(n15264), .A2(n14839), .B1(n15263), .B2(n14844), .ZN(
        n14330) );
  AOI21_X1 U16131 ( .B1(n15294), .B2(P2_REIP_REG_4__SCAN_IN), .A(n14330), .ZN(
        n14331) );
  OAI21_X1 U16132 ( .B1(n15297), .B2(n15502), .A(n14331), .ZN(n14332) );
  INV_X1 U16133 ( .A(n14332), .ZN(n14340) );
  INV_X1 U16134 ( .A(n14588), .ZN(n14334) );
  AOI21_X1 U16135 ( .B1(n14335), .B2(n14333), .A(n14334), .ZN(n18256) );
  INV_X1 U16136 ( .A(n18256), .ZN(n15154) );
  MUX2_X1 U16137 ( .A(n18248), .B(n15154), .S(n11059), .Z(n14336) );
  OAI21_X1 U16138 ( .B1(n14337), .B2(n16253), .A(n14336), .ZN(P2_U2882) );
  OAI21_X1 U16139 ( .B1(n14339), .B2(n14338), .A(n14319), .ZN(n19372) );
  NAND2_X1 U16140 ( .A1(n14341), .A2(n14340), .ZN(n14342) );
  AND2_X1 U16141 ( .A1(n14333), .A2(n14342), .ZN(n17108) );
  NOR2_X1 U16142 ( .A1(n11059), .A2(n14839), .ZN(n14343) );
  AOI21_X1 U16143 ( .B1(n17108), .B2(n11059), .A(n14343), .ZN(n14344) );
  OAI21_X1 U16144 ( .B1(n19372), .B2(n16253), .A(n14344), .ZN(P2_U2883) );
  INV_X1 U16145 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20035) );
  NOR2_X1 U16146 ( .A1(n14377), .A2(DATAI_3_), .ZN(n14345) );
  AOI21_X1 U16147 ( .B1(n14377), .B2(n20035), .A(n14345), .ZN(n15773) );
  NAND2_X1 U16148 ( .A1(n21740), .A2(n15773), .ZN(n14360) );
  AOI22_X1 U16149 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_19__SCAN_IN), .ZN(n14346) );
  NAND2_X1 U16150 ( .A1(n14360), .A2(n14346), .ZN(P1_U2940) );
  NOR2_X1 U16151 ( .A1(n14377), .A2(DATAI_4_), .ZN(n14347) );
  AOI21_X1 U16152 ( .B1(n14377), .B2(n20037), .A(n14347), .ZN(n15770) );
  NAND2_X1 U16153 ( .A1(n21740), .A2(n15770), .ZN(n14352) );
  AOI22_X1 U16154 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_20__SCAN_IN), .ZN(n14348) );
  NAND2_X1 U16155 ( .A1(n14352), .A2(n14348), .ZN(P1_U2941) );
  INV_X1 U16156 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20041) );
  NOR2_X1 U16157 ( .A1(n14377), .A2(DATAI_6_), .ZN(n14349) );
  AOI21_X1 U16158 ( .B1(n14377), .B2(n20041), .A(n14349), .ZN(n15758) );
  NAND2_X1 U16159 ( .A1(n21740), .A2(n15758), .ZN(n14354) );
  AOI22_X1 U16160 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_22__SCAN_IN), .ZN(n14350) );
  NAND2_X1 U16161 ( .A1(n14354), .A2(n14350), .ZN(P1_U2943) );
  AOI22_X1 U16162 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_4__SCAN_IN), .ZN(n14351) );
  NAND2_X1 U16163 ( .A1(n14352), .A2(n14351), .ZN(P1_U2956) );
  AOI22_X1 U16164 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_6__SCAN_IN), .ZN(n14353) );
  NAND2_X1 U16165 ( .A1(n14354), .A2(n14353), .ZN(P1_U2958) );
  INV_X1 U16166 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20039) );
  NOR2_X1 U16167 ( .A1(n14377), .A2(DATAI_5_), .ZN(n14355) );
  AOI21_X1 U16168 ( .B1(n14377), .B2(n20039), .A(n14355), .ZN(n15762) );
  NAND2_X1 U16169 ( .A1(n21740), .A2(n15762), .ZN(n14358) );
  AOI22_X1 U16170 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_5__SCAN_IN), .ZN(n14356) );
  NAND2_X1 U16171 ( .A1(n14358), .A2(n14356), .ZN(P1_U2957) );
  AOI22_X1 U16172 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_21__SCAN_IN), .ZN(n14357) );
  NAND2_X1 U16173 ( .A1(n14358), .A2(n14357), .ZN(P1_U2942) );
  AOI22_X1 U16174 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_3__SCAN_IN), .ZN(n14359) );
  NAND2_X1 U16175 ( .A1(n14360), .A2(n14359), .ZN(P1_U2955) );
  INV_X1 U16176 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20043) );
  NOR2_X1 U16177 ( .A1(n14377), .A2(DATAI_7_), .ZN(n14361) );
  AOI21_X1 U16178 ( .B1(n14377), .B2(n20043), .A(n14361), .ZN(n15755) );
  NAND2_X1 U16179 ( .A1(n21740), .A2(n15755), .ZN(n14364) );
  AOI22_X1 U16180 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_7__SCAN_IN), .ZN(n14362) );
  NAND2_X1 U16181 ( .A1(n14364), .A2(n14362), .ZN(P1_U2959) );
  AOI22_X1 U16182 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_23__SCAN_IN), .ZN(n14363) );
  NAND2_X1 U16183 ( .A1(n14364), .A2(n14363), .ZN(P1_U2944) );
  NAND2_X1 U16184 ( .A1(n21740), .A2(n15789), .ZN(n14432) );
  AOI22_X1 U16185 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_0__SCAN_IN), .ZN(n14365) );
  NAND2_X1 U16186 ( .A1(n14432), .A2(n14365), .ZN(P1_U2952) );
  NAND2_X1 U16187 ( .A1(n21740), .A2(n15777), .ZN(n14434) );
  AOI22_X1 U16188 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_2__SCAN_IN), .ZN(n14366) );
  NAND2_X1 U16189 ( .A1(n14434), .A2(n14366), .ZN(P1_U2954) );
  NAND2_X1 U16190 ( .A1(n21740), .A2(n15782), .ZN(n14436) );
  AOI22_X1 U16191 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_1__SCAN_IN), .ZN(n14367) );
  NAND2_X1 U16192 ( .A1(n14436), .A2(n14367), .ZN(P1_U2953) );
  INV_X1 U16193 ( .A(n16887), .ZN(n14376) );
  OAI21_X1 U16194 ( .B1(n21905), .B2(n21924), .A(n14369), .ZN(n21929) );
  INV_X1 U16195 ( .A(n21829), .ZN(n14370) );
  NOR2_X1 U16196 ( .A1(n14370), .A2(n16075), .ZN(n14373) );
  NAND2_X1 U16197 ( .A1(n10975), .A2(n14371), .ZN(n14441) );
  NOR2_X1 U16198 ( .A1(n14441), .A2(n14372), .ZN(n14378) );
  NAND2_X1 U16199 ( .A1(n14376), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14374) );
  OAI21_X1 U16200 ( .B1(n14376), .B2(n14375), .A(n14374), .ZN(P1_U3475) );
  INV_X1 U16201 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20085) );
  INV_X1 U16202 ( .A(DATAI_28_), .ZN(n15731) );
  OAI22_X1 U16203 ( .A1(n20085), .A2(n14567), .B1(n15731), .B2(n14566), .ZN(
        n22088) );
  INV_X1 U16204 ( .A(n22088), .ZN(n22098) );
  NOR2_X1 U16205 ( .A1(n21921), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14384) );
  OAI21_X1 U16206 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n21837), .A(
        n14570), .ZN(n21928) );
  INV_X1 U16207 ( .A(n21928), .ZN(n21898) );
  OAI21_X1 U16208 ( .B1(n14378), .B2(n14384), .A(n21898), .ZN(n14565) );
  NAND2_X1 U16209 ( .A1(n14565), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14390) );
  OR2_X1 U16210 ( .A1(n14441), .A2(n21868), .ZN(n14422) );
  INV_X1 U16211 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20068) );
  INV_X1 U16212 ( .A(DATAI_20_), .ZN(n17021) );
  OAI22_X1 U16213 ( .A1(n20068), .A2(n14567), .B1(n17021), .B2(n14566), .ZN(
        n22082) );
  NOR2_X1 U16214 ( .A1(n14569), .A2(n11682), .ZN(n22091) );
  INV_X1 U16215 ( .A(n22091), .ZN(n22076) );
  NOR2_X1 U16216 ( .A1(n21877), .A2(n14381), .ZN(n21817) );
  INV_X1 U16217 ( .A(n14572), .ZN(n14383) );
  AOI21_X1 U16218 ( .B1(n21817), .B2(n10998), .A(n14383), .ZN(n14386) );
  INV_X1 U16219 ( .A(n14384), .ZN(n14385) );
  OAI22_X1 U16220 ( .A1(n14386), .A2(n21924), .B1(n14385), .B2(n21922), .ZN(
        n14387) );
  INV_X1 U16221 ( .A(n14387), .ZN(n14571) );
  NAND2_X1 U16222 ( .A1(n14570), .A2(n15770), .ZN(n22085) );
  OAI22_X1 U16223 ( .A1(n22076), .A2(n14572), .B1(n14571), .B2(n22085), .ZN(
        n14388) );
  AOI21_X1 U16224 ( .B1(n22217), .B2(n22082), .A(n14388), .ZN(n14389) );
  OAI211_X1 U16225 ( .C1(n22067), .C2(n22098), .A(n14390), .B(n14389), .ZN(
        P1_U3093) );
  INV_X1 U16226 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20083) );
  INV_X1 U16227 ( .A(DATAI_27_), .ZN(n14391) );
  OAI22_X1 U16228 ( .A1(n20083), .A2(n14567), .B1(n14391), .B2(n14566), .ZN(
        n22046) );
  INV_X1 U16229 ( .A(n22046), .ZN(n22056) );
  NAND2_X1 U16230 ( .A1(n14565), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14395) );
  INV_X1 U16231 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20066) );
  INV_X1 U16232 ( .A(DATAI_19_), .ZN(n17001) );
  NOR2_X1 U16233 ( .A1(n14569), .A2(n14392), .ZN(n22049) );
  INV_X1 U16234 ( .A(n22049), .ZN(n22034) );
  NAND2_X1 U16235 ( .A1(n14570), .A2(n15773), .ZN(n22043) );
  OAI22_X1 U16236 ( .A1(n22034), .A2(n14572), .B1(n14571), .B2(n22043), .ZN(
        n14393) );
  AOI21_X1 U16237 ( .B1(n22217), .B2(n22040), .A(n14393), .ZN(n14394) );
  OAI211_X1 U16238 ( .C1(n22067), .C2(n22056), .A(n14395), .B(n14394), .ZN(
        P1_U3092) );
  INV_X1 U16239 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20093) );
  OAI22_X1 U16240 ( .A1(n14396), .A2(n14566), .B1(n20093), .B2(n14567), .ZN(
        n22258) );
  INV_X1 U16241 ( .A(n22258), .ZN(n22275) );
  NAND2_X1 U16242 ( .A1(n14565), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14400) );
  INV_X1 U16243 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20075) );
  INV_X1 U16244 ( .A(DATAI_23_), .ZN(n14397) );
  OAI22_X1 U16245 ( .A1(n20075), .A2(n14567), .B1(n14397), .B2(n14566), .ZN(
        n22242) );
  NOR2_X1 U16246 ( .A1(n14569), .A2(n11681), .ZN(n22264) );
  INV_X1 U16247 ( .A(n22264), .ZN(n22228) );
  NAND2_X1 U16248 ( .A1(n14570), .A2(n15755), .ZN(n22247) );
  OAI22_X1 U16249 ( .A1(n22228), .A2(n14572), .B1(n14571), .B2(n22247), .ZN(
        n14398) );
  AOI21_X1 U16250 ( .B1(n22217), .B2(n22242), .A(n14398), .ZN(n14399) );
  OAI211_X1 U16251 ( .C1(n22067), .C2(n22275), .A(n14400), .B(n14399), .ZN(
        P1_U3096) );
  INV_X1 U16252 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20087) );
  INV_X1 U16253 ( .A(DATAI_29_), .ZN(n16910) );
  OAI22_X1 U16254 ( .A1(n20087), .A2(n14567), .B1(n16910), .B2(n14566), .ZN(
        n22127) );
  INV_X1 U16255 ( .A(n22127), .ZN(n22137) );
  NAND2_X1 U16256 ( .A1(n14565), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14403) );
  INV_X1 U16257 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20070) );
  INV_X1 U16258 ( .A(DATAI_21_), .ZN(n17017) );
  NOR2_X1 U16259 ( .A1(n14569), .A2(n11700), .ZN(n22130) );
  INV_X1 U16260 ( .A(n22130), .ZN(n22115) );
  NAND2_X1 U16261 ( .A1(n14570), .A2(n15762), .ZN(n22124) );
  OAI22_X1 U16262 ( .A1(n22115), .A2(n14572), .B1(n14571), .B2(n22124), .ZN(
        n14401) );
  AOI21_X1 U16263 ( .B1(n22217), .B2(n22121), .A(n14401), .ZN(n14402) );
  OAI211_X1 U16264 ( .C1(n22067), .C2(n22137), .A(n14403), .B(n14402), .ZN(
        P1_U3094) );
  INV_X1 U16265 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20091) );
  OAI22_X1 U16266 ( .A1(n20091), .A2(n14567), .B1(n16909), .B2(n14566), .ZN(
        n22170) );
  INV_X1 U16267 ( .A(n22170), .ZN(n22180) );
  NAND2_X1 U16268 ( .A1(n14565), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14407) );
  INV_X1 U16269 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20072) );
  INV_X1 U16270 ( .A(DATAI_22_), .ZN(n16916) );
  NOR2_X1 U16271 ( .A1(n14569), .A2(n14404), .ZN(n22173) );
  INV_X1 U16272 ( .A(n22173), .ZN(n22156) );
  NAND2_X1 U16273 ( .A1(n14570), .A2(n15758), .ZN(n22167) );
  OAI22_X1 U16274 ( .A1(n22156), .A2(n14572), .B1(n14571), .B2(n22167), .ZN(
        n14405) );
  AOI21_X1 U16275 ( .B1(n22217), .B2(n22164), .A(n14405), .ZN(n14406) );
  OAI211_X1 U16276 ( .C1(n22067), .C2(n22180), .A(n14407), .B(n14406), .ZN(
        P1_U3095) );
  INV_X1 U16277 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20079) );
  INV_X1 U16278 ( .A(DATAI_25_), .ZN(n14408) );
  OAI22_X1 U16279 ( .A1(n20079), .A2(n14567), .B1(n14408), .B2(n14566), .ZN(
        n21968) );
  INV_X1 U16280 ( .A(n21968), .ZN(n21978) );
  NAND2_X1 U16281 ( .A1(n14565), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14413) );
  INV_X1 U16282 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20062) );
  INV_X1 U16283 ( .A(DATAI_17_), .ZN(n14409) );
  OAI22_X1 U16284 ( .A1(n20062), .A2(n14567), .B1(n14409), .B2(n14566), .ZN(
        n21962) );
  NOR2_X1 U16285 ( .A1(n14569), .A2(n14410), .ZN(n21971) );
  INV_X1 U16286 ( .A(n21971), .ZN(n21956) );
  NAND2_X1 U16287 ( .A1(n14570), .A2(n15782), .ZN(n21965) );
  OAI22_X1 U16288 ( .A1(n21956), .A2(n14572), .B1(n14571), .B2(n21965), .ZN(
        n14411) );
  AOI21_X1 U16289 ( .B1(n22217), .B2(n21962), .A(n14411), .ZN(n14412) );
  OAI211_X1 U16290 ( .C1(n22067), .C2(n21978), .A(n14413), .B(n14412), .ZN(
        P1_U3090) );
  INV_X1 U16291 ( .A(n14428), .ZN(n14414) );
  OAI21_X1 U16292 ( .B1(n14416), .B2(n14415), .A(n14414), .ZN(n21293) );
  INV_X1 U16293 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14418) );
  OAI222_X1 U16294 ( .A1(n21293), .A2(n19942), .B1(n14418), .B2(n19946), .C1(
        n15726), .C2(n14417), .ZN(P1_U2870) );
  INV_X1 U16295 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20060) );
  INV_X1 U16296 ( .A(DATAI_16_), .ZN(n17026) );
  OAI22_X1 U16297 ( .A1(n20060), .A2(n14567), .B1(n17026), .B2(n14566), .ZN(
        n21881) );
  INV_X1 U16298 ( .A(n21881), .ZN(n21934) );
  NAND2_X1 U16299 ( .A1(n14565), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14421) );
  INV_X1 U16300 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20077) );
  INV_X1 U16301 ( .A(DATAI_24_), .ZN(n17010) );
  OAI22_X1 U16302 ( .A1(n20077), .A2(n14567), .B1(n17010), .B2(n14566), .ZN(
        n21916) );
  NOR2_X1 U16303 ( .A1(n14569), .A2(n11686), .ZN(n21925) );
  INV_X1 U16304 ( .A(n21925), .ZN(n21852) );
  NAND2_X1 U16305 ( .A1(n14570), .A2(n15789), .ZN(n21889) );
  OAI22_X1 U16306 ( .A1(n21852), .A2(n14572), .B1(n14571), .B2(n21889), .ZN(
        n14419) );
  AOI21_X1 U16307 ( .B1(n22210), .B2(n21916), .A(n14419), .ZN(n14420) );
  OAI211_X1 U16308 ( .C1(n14422), .C2(n21934), .A(n14421), .B(n14420), .ZN(
        P1_U3089) );
  OAI21_X1 U16309 ( .B1(n14423), .B2(n14425), .A(n14648), .ZN(n14622) );
  OAI21_X1 U16310 ( .B1(n14428), .B2(n14427), .A(n14426), .ZN(n14617) );
  INV_X1 U16311 ( .A(n14617), .ZN(n14429) );
  INV_X1 U16312 ( .A(n19946), .ZN(n15724) );
  AOI22_X1 U16313 ( .A1(n19925), .A2(n14429), .B1(n15724), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n14430) );
  OAI21_X1 U16314 ( .B1(n14622), .B2(n15726), .A(n14430), .ZN(P1_U2869) );
  NAND2_X1 U16315 ( .A1(n21775), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14431) );
  OAI211_X1 U16316 ( .C1(n21777), .C2(n15785), .A(n14432), .B(n14431), .ZN(
        P1_U2937) );
  INV_X1 U16317 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14632) );
  NAND2_X1 U16318 ( .A1(n21775), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14433) );
  OAI211_X1 U16319 ( .C1(n21777), .C2(n14632), .A(n14434), .B(n14433), .ZN(
        P1_U2939) );
  NAND2_X1 U16320 ( .A1(n21775), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14435) );
  OAI211_X1 U16321 ( .C1(n21777), .C2(n14239), .A(n14436), .B(n14435), .ZN(
        P1_U2938) );
  INV_X1 U16322 ( .A(n16073), .ZN(n14437) );
  INV_X1 U16323 ( .A(n21916), .ZN(n21938) );
  NAND3_X1 U16324 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n11834), .A3(
        n21880), .ZN(n14762) );
  INV_X1 U16325 ( .A(n14762), .ZN(n14445) );
  INV_X1 U16326 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n14439) );
  INV_X1 U16327 ( .A(n14438), .ZN(n21893) );
  NOR2_X1 U16328 ( .A1(n21892), .A2(n14762), .ZN(n14442) );
  AOI21_X1 U16329 ( .B1(n21817), .B2(n21893), .A(n14442), .ZN(n14443) );
  OAI211_X1 U16330 ( .C1(n14441), .C2(n14439), .A(n21900), .B(n14443), .ZN(
        n14440) );
  OAI211_X1 U16331 ( .C1(n21900), .C2(n14445), .A(n14440), .B(n21898), .ZN(
        n14576) );
  NAND2_X1 U16332 ( .A1(n14576), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n14450) );
  INV_X1 U16333 ( .A(n21890), .ZN(n21844) );
  INV_X1 U16334 ( .A(n14442), .ZN(n14578) );
  INV_X1 U16335 ( .A(n14443), .ZN(n14444) );
  NAND2_X1 U16336 ( .A1(n14444), .A2(n21900), .ZN(n14447) );
  NAND2_X1 U16337 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14445), .ZN(n14446) );
  AND2_X1 U16338 ( .A1(n14447), .A2(n14446), .ZN(n14577) );
  OAI22_X1 U16339 ( .A1(n21852), .A2(n14578), .B1(n21889), .B2(n14577), .ZN(
        n14448) );
  AOI21_X1 U16340 ( .B1(n22069), .B2(n21881), .A(n14448), .ZN(n14449) );
  OAI211_X1 U16341 ( .C1(n14582), .C2(n21938), .A(n14450), .B(n14449), .ZN(
        P1_U3073) );
  NAND2_X1 U16342 ( .A1(n14576), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n14453) );
  OAI22_X1 U16343 ( .A1(n21956), .A2(n14578), .B1(n21965), .B2(n14577), .ZN(
        n14451) );
  AOI21_X1 U16344 ( .B1(n22069), .B2(n21962), .A(n14451), .ZN(n14452) );
  OAI211_X1 U16345 ( .C1(n14582), .C2(n21978), .A(n14453), .B(n14452), .ZN(
        P1_U3074) );
  NAND2_X1 U16346 ( .A1(n14576), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n14456) );
  OAI22_X1 U16347 ( .A1(n22034), .A2(n14578), .B1(n22043), .B2(n14577), .ZN(
        n14454) );
  AOI21_X1 U16348 ( .B1(n22069), .B2(n22040), .A(n14454), .ZN(n14455) );
  OAI211_X1 U16349 ( .C1(n14582), .C2(n22056), .A(n14456), .B(n14455), .ZN(
        P1_U3076) );
  NAND2_X1 U16350 ( .A1(n14576), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n14459) );
  OAI22_X1 U16351 ( .A1(n22156), .A2(n14578), .B1(n22167), .B2(n14577), .ZN(
        n14457) );
  AOI21_X1 U16352 ( .B1(n22069), .B2(n22164), .A(n14457), .ZN(n14458) );
  OAI211_X1 U16353 ( .C1(n14582), .C2(n22180), .A(n14459), .B(n14458), .ZN(
        P1_U3079) );
  NAND2_X1 U16354 ( .A1(n14576), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n14462) );
  OAI22_X1 U16355 ( .A1(n22228), .A2(n14578), .B1(n22247), .B2(n14577), .ZN(
        n14460) );
  AOI21_X1 U16356 ( .B1(n22069), .B2(n22242), .A(n14460), .ZN(n14461) );
  OAI211_X1 U16357 ( .C1(n14582), .C2(n22275), .A(n14462), .B(n14461), .ZN(
        P1_U3080) );
  NAND2_X1 U16358 ( .A1(n14576), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14465) );
  OAI22_X1 U16359 ( .A1(n22115), .A2(n14578), .B1(n22124), .B2(n14577), .ZN(
        n14463) );
  AOI21_X1 U16360 ( .B1(n22069), .B2(n22121), .A(n14463), .ZN(n14464) );
  OAI211_X1 U16361 ( .C1(n14582), .C2(n22137), .A(n14465), .B(n14464), .ZN(
        P1_U3078) );
  NAND2_X1 U16362 ( .A1(n14576), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n14468) );
  OAI22_X1 U16363 ( .A1(n22076), .A2(n14578), .B1(n22085), .B2(n14577), .ZN(
        n14466) );
  AOI21_X1 U16364 ( .B1(n22069), .B2(n22082), .A(n14466), .ZN(n14467) );
  OAI211_X1 U16365 ( .C1(n14582), .C2(n22098), .A(n14468), .B(n14467), .ZN(
        P1_U3077) );
  INV_X1 U16366 ( .A(n14498), .ZN(n14493) );
  NAND2_X1 U16367 ( .A1(n15005), .A2(n14493), .ZN(n14480) );
  NOR2_X1 U16368 ( .A1(n14469), .A2(n14502), .ZN(n14472) );
  NAND2_X1 U16369 ( .A1(n14119), .A2(n14470), .ZN(n14506) );
  INV_X1 U16370 ( .A(n13125), .ZN(n14471) );
  NAND2_X1 U16371 ( .A1(n14471), .A2(n14481), .ZN(n14508) );
  AND2_X1 U16372 ( .A1(n14505), .A2(n14508), .ZN(n14475) );
  AOI22_X1 U16373 ( .A1(n14504), .A2(n14472), .B1(n14506), .B2(n14475), .ZN(
        n14478) );
  INV_X1 U16374 ( .A(n14523), .ZN(n14473) );
  NAND2_X1 U16375 ( .A1(n14474), .A2(n14473), .ZN(n14499) );
  INV_X1 U16376 ( .A(n14475), .ZN(n14476) );
  NAND2_X1 U16377 ( .A1(n14499), .A2(n14476), .ZN(n14477) );
  AND2_X1 U16378 ( .A1(n14478), .A2(n14477), .ZN(n14479) );
  NAND2_X1 U16379 ( .A1(n14480), .A2(n14479), .ZN(n16797) );
  OR2_X1 U16380 ( .A1(n16797), .A2(n14522), .ZN(n14483) );
  NAND2_X1 U16381 ( .A1(n14522), .A2(n14481), .ZN(n14482) );
  NAND2_X1 U16382 ( .A1(n14483), .A2(n14482), .ZN(n14521) );
  OR2_X1 U16383 ( .A1(n10973), .A2(n14498), .ZN(n14489) );
  INV_X1 U16384 ( .A(n13578), .ZN(n14485) );
  NAND2_X1 U16385 ( .A1(n14485), .A2(n14484), .ZN(n14491) );
  NOR2_X1 U16386 ( .A1(n13127), .A2(n13125), .ZN(n14486) );
  AOI22_X1 U16387 ( .A1(n14504), .A2(n14487), .B1(n14491), .B2(n14486), .ZN(
        n14488) );
  AND2_X1 U16388 ( .A1(n14489), .A2(n14488), .ZN(n16791) );
  MUX2_X1 U16389 ( .A(n14504), .B(n14491), .S(n14490), .Z(n14492) );
  AOI21_X1 U16390 ( .B1(n18244), .B2(n14493), .A(n14492), .ZN(n16784) );
  OAI211_X1 U16391 ( .C1(n16791), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16784), .ZN(n14495) );
  AOI21_X1 U16392 ( .B1(n16791), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n14522), .ZN(n14494) );
  NAND2_X1 U16393 ( .A1(n14495), .A2(n14494), .ZN(n14496) );
  OAI21_X1 U16394 ( .B1(n14521), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n14496), .ZN(n14497) );
  OAI21_X1 U16395 ( .B1(n16797), .B2(n19256), .A(n14497), .ZN(n14517) );
  OR2_X1 U16396 ( .A1(n17101), .A2(n14498), .ZN(n14515) );
  NAND2_X1 U16397 ( .A1(n14499), .A2(n14508), .ZN(n14501) );
  NAND2_X1 U16398 ( .A1(n14504), .A2(n14502), .ZN(n14500) );
  NAND2_X1 U16399 ( .A1(n14501), .A2(n14500), .ZN(n14511) );
  INV_X1 U16400 ( .A(n14502), .ZN(n14503) );
  NAND2_X1 U16401 ( .A1(n14504), .A2(n14503), .ZN(n14509) );
  NAND2_X1 U16402 ( .A1(n14506), .A2(n14505), .ZN(n14507) );
  NAND3_X1 U16403 ( .A1(n14509), .A2(n14508), .A3(n14507), .ZN(n14510) );
  MUX2_X1 U16404 ( .A(n14511), .B(n14510), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14513) );
  NOR2_X1 U16405 ( .A1(n14513), .A2(n14512), .ZN(n14514) );
  NAND2_X1 U16406 ( .A1(n14515), .A2(n14514), .ZN(n14562) );
  MUX2_X1 U16407 ( .A(n14562), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14522), .Z(n14547) );
  INV_X1 U16408 ( .A(n14547), .ZN(n14518) );
  OR2_X1 U16409 ( .A1(n14518), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14516) );
  NAND2_X1 U16410 ( .A1(n14517), .A2(n14516), .ZN(n14520) );
  AOI21_X1 U16411 ( .B1(n14518), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n14519) );
  NAND2_X1 U16412 ( .A1(n14520), .A2(n14519), .ZN(n14550) );
  INV_X1 U16413 ( .A(n14521), .ZN(n14548) );
  NAND2_X1 U16414 ( .A1(n14522), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14545) );
  NAND2_X1 U16415 ( .A1(n14524), .A2(n14523), .ZN(n14533) );
  INV_X1 U16416 ( .A(n14525), .ZN(n14529) );
  AOI22_X1 U16417 ( .A1(n14527), .A2(n14526), .B1(n14538), .B2(n14536), .ZN(
        n14528) );
  OAI21_X1 U16418 ( .B1(n16836), .B2(n14529), .A(n14528), .ZN(n14530) );
  AOI21_X1 U16419 ( .B1(n14561), .B2(n14531), .A(n14530), .ZN(n14532) );
  AND2_X1 U16420 ( .A1(n14533), .A2(n14532), .ZN(n18621) );
  INV_X1 U16421 ( .A(n14534), .ZN(n14535) );
  NAND3_X1 U16422 ( .A1(n14536), .A2(n14552), .A3(n14535), .ZN(n14537) );
  OR2_X1 U16423 ( .A1(n14538), .A2(n14537), .ZN(n18618) );
  NOR2_X1 U16424 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n14541) );
  OAI22_X1 U16425 ( .A1(n18618), .A2(n14541), .B1(n14540), .B2(n14539), .ZN(
        n14542) );
  NOR2_X1 U16426 ( .A1(n14543), .A2(n14542), .ZN(n14544) );
  NAND3_X1 U16427 ( .A1(n14545), .A2(n18621), .A3(n14544), .ZN(n14546) );
  AOI21_X1 U16428 ( .B1(n14548), .B2(n14547), .A(n14546), .ZN(n14549) );
  NAND2_X1 U16429 ( .A1(n18617), .A2(n14551), .ZN(n14558) );
  NOR2_X1 U16430 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14552), .ZN(n14726) );
  AND2_X1 U16431 ( .A1(n14553), .A2(n14726), .ZN(n14720) );
  INV_X1 U16432 ( .A(n14720), .ZN(n14554) );
  NOR2_X1 U16433 ( .A1(n14555), .A2(n14554), .ZN(n14556) );
  AOI21_X1 U16434 ( .B1(n14558), .B2(n14557), .A(n14556), .ZN(n18613) );
  AOI211_X1 U16435 ( .C1(n18613), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n16833), 
        .B(n14559), .ZN(n14560) );
  INV_X1 U16436 ( .A(n14560), .ZN(P2_U3593) );
  INV_X1 U16437 ( .A(n18606), .ZN(n16794) );
  INV_X1 U16438 ( .A(n18596), .ZN(n17213) );
  AOI22_X1 U16439 ( .A1(n19110), .A2(n16794), .B1(n17213), .B2(n14562), .ZN(
        n14563) );
  MUX2_X1 U16440 ( .A(n13511), .B(n14563), .S(n16792), .Z(n14564) );
  INV_X1 U16441 ( .A(n14564), .ZN(P2_U3596) );
  INV_X1 U16442 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20081) );
  INV_X1 U16443 ( .A(DATAI_26_), .ZN(n16906) );
  OAI22_X1 U16444 ( .A1(n20081), .A2(n14567), .B1(n16906), .B2(n14566), .ZN(
        n22007) );
  INV_X1 U16445 ( .A(n22007), .ZN(n22017) );
  NAND2_X1 U16446 ( .A1(n14565), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14575) );
  INV_X1 U16447 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20064) );
  INV_X1 U16448 ( .A(DATAI_18_), .ZN(n17002) );
  NOR2_X1 U16449 ( .A1(n14569), .A2(n14568), .ZN(n22010) );
  INV_X1 U16450 ( .A(n22010), .ZN(n21995) );
  NAND2_X1 U16451 ( .A1(n14570), .A2(n15777), .ZN(n22004) );
  OAI22_X1 U16452 ( .A1(n21995), .A2(n14572), .B1(n14571), .B2(n22004), .ZN(
        n14573) );
  AOI21_X1 U16453 ( .B1(n22217), .B2(n22001), .A(n14573), .ZN(n14574) );
  OAI211_X1 U16454 ( .C1(n22067), .C2(n22017), .A(n14575), .B(n14574), .ZN(
        P1_U3091) );
  NAND2_X1 U16455 ( .A1(n14576), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n14581) );
  OAI22_X1 U16456 ( .A1(n21995), .A2(n14578), .B1(n22004), .B2(n14577), .ZN(
        n14579) );
  AOI21_X1 U16457 ( .B1(n22069), .B2(n22001), .A(n14579), .ZN(n14580) );
  OAI211_X1 U16458 ( .C1(n14582), .C2(n22017), .A(n14581), .B(n14580), .ZN(
        P1_U3075) );
  INV_X1 U16459 ( .A(n15773), .ZN(n14583) );
  INV_X1 U16460 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19828) );
  OAI222_X1 U16461 ( .A1(n15796), .A2(n14583), .B1(n15794), .B2(n19828), .C1(
        n15801), .C2(n14622), .ZN(P1_U2901) );
  NAND2_X1 U16462 ( .A1(n15285), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n14585) );
  NAND2_X1 U16463 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n14584) );
  OAI211_X1 U16464 ( .C1(n15300), .C2(n17272), .A(n14585), .B(n14584), .ZN(
        n14586) );
  AOI21_X1 U16465 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14586), .ZN(n14587) );
  AND2_X1 U16466 ( .A1(n14588), .A2(n14587), .ZN(n14589) );
  OR2_X1 U16467 ( .A1(n14589), .A2(n14642), .ZN(n17114) );
  NOR2_X1 U16468 ( .A1(n14319), .A2(n19419), .ZN(n14590) );
  OAI211_X1 U16469 ( .C1(n14590), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n16266), .B(n14638), .ZN(n14592) );
  NAND2_X1 U16470 ( .A1(n10963), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n14591) );
  OAI211_X1 U16471 ( .C1(n17114), .C2(n10963), .A(n14592), .B(n14591), .ZN(
        P2_U2881) );
  AND2_X1 U16472 ( .A1(n11702), .A2(n14593), .ZN(n14594) );
  NOR2_X1 U16473 ( .A1(n21618), .A2(n14594), .ZN(n21440) );
  INV_X1 U16474 ( .A(n14624), .ZN(n14608) );
  AND2_X1 U16475 ( .A1(n14595), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14596) );
  NOR2_X1 U16476 ( .A1(n14598), .A2(n14597), .ZN(n21456) );
  NOR2_X1 U16477 ( .A1(n14617), .A2(n21638), .ZN(n14604) );
  INV_X1 U16478 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14602) );
  INV_X1 U16479 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n19847) );
  NAND4_X1 U16480 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(n21493), .A4(n19847), .ZN(n14601) );
  OAI221_X1 U16481 ( .B1(n21484), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n21484), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n21483), .ZN(n14599) );
  NAND2_X1 U16482 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n14599), .ZN(n14600) );
  OAI211_X1 U16483 ( .C1(n21623), .C2(n14602), .A(n14601), .B(n14600), .ZN(
        n14603) );
  AOI211_X1 U16484 ( .C1(n21829), .C2(n21456), .A(n14604), .B(n14603), .ZN(
        n14605) );
  OAI21_X1 U16485 ( .B1(n21626), .B2(n14606), .A(n14605), .ZN(n14607) );
  AOI21_X1 U16486 ( .B1(n14608), .B2(n21634), .A(n14607), .ZN(n14609) );
  OAI21_X1 U16487 ( .B1(n14622), .B2(n21440), .A(n14609), .ZN(P1_U2837) );
  NAND2_X1 U16488 ( .A1(n14611), .A2(n14610), .ZN(n14612) );
  XOR2_X1 U16489 ( .A(n14613), .B(n14612), .Z(n14628) );
  INV_X1 U16490 ( .A(n15941), .ZN(n21366) );
  OAI21_X1 U16491 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15942), .A(
        n14615), .ZN(n21401) );
  AOI21_X1 U16492 ( .B1(n14616), .B2(n21366), .A(n21401), .ZN(n21295) );
  INV_X1 U16493 ( .A(n21368), .ZN(n16033) );
  AOI21_X1 U16494 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14688) );
  NAND2_X1 U16495 ( .A1(n16033), .A2(n14688), .ZN(n21303) );
  OAI211_X1 U16496 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n15941), .A(
        n21295), .B(n21303), .ZN(n21306) );
  OAI22_X1 U16497 ( .A1(n21414), .A2(n14617), .B1(n19847), .B2(n21419), .ZN(
        n14620) );
  NAND3_X1 U16498 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21301), .ZN(n21316) );
  OAI21_X1 U16499 ( .B1(n14688), .B2(n21368), .A(n21316), .ZN(n21312) );
  INV_X1 U16500 ( .A(n21312), .ZN(n14691) );
  NOR2_X1 U16501 ( .A1(n14691), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14619) );
  AOI211_X1 U16502 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n21306), .A(
        n14620), .B(n14619), .ZN(n14621) );
  OAI21_X1 U16503 ( .B1(n14628), .B2(n21382), .A(n14621), .ZN(P1_U3028) );
  INV_X1 U16504 ( .A(n14622), .ZN(n14626) );
  AOI22_X1 U16505 ( .A1(n20014), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n14073), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n14623) );
  OAI21_X1 U16506 ( .B1(n20024), .B2(n14624), .A(n14623), .ZN(n14625) );
  AOI21_X1 U16507 ( .B1(n14626), .B2(n20021), .A(n14625), .ZN(n14627) );
  OAI21_X1 U16508 ( .B1(n14628), .B2(n21639), .A(n14627), .ZN(P1_U2996) );
  AOI22_X1 U16509 ( .A1(n14630), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14631) );
  OAI21_X1 U16510 ( .B1(n14632), .B2(n14637), .A(n14631), .ZN(P1_U2918) );
  INV_X1 U16511 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14634) );
  AOI22_X1 U16512 ( .A1(n21278), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14633) );
  OAI21_X1 U16513 ( .B1(n14634), .B2(n14637), .A(n14633), .ZN(P1_U2913) );
  AOI22_X1 U16514 ( .A1(n21278), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14635) );
  OAI21_X1 U16515 ( .B1(n15730), .B2(n14637), .A(n14635), .ZN(P1_U2908) );
  INV_X1 U16516 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n21766) );
  AOI22_X1 U16517 ( .A1(n21278), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14636) );
  OAI21_X1 U16518 ( .B1(n21766), .B2(n14637), .A(n14636), .ZN(P1_U2907) );
  XOR2_X1 U16519 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n14638), .Z(n14646)
         );
  INV_X1 U16520 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16745) );
  AOI22_X1 U16521 ( .A1(n15556), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14640) );
  NAND2_X1 U16522 ( .A1(n15294), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n14639) );
  OAI211_X1 U16523 ( .C1(n15297), .C2(n16745), .A(n14640), .B(n14639), .ZN(
        n14641) );
  NAND2_X1 U16524 ( .A1(n14642), .A2(n14641), .ZN(n14677) );
  OR2_X1 U16525 ( .A1(n14642), .A2(n14641), .ZN(n14643) );
  NAND2_X1 U16526 ( .A1(n14677), .A2(n14643), .ZN(n18269) );
  INV_X1 U16527 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n14644) );
  MUX2_X1 U16528 ( .A(n18269), .B(n14644), .S(n10963), .Z(n14645) );
  OAI21_X1 U16529 ( .B1(n14646), .B2(n16253), .A(n14645), .ZN(P2_U2880) );
  XOR2_X1 U16530 ( .A(n14648), .B(n14647), .Z(n21463) );
  INV_X1 U16531 ( .A(n21463), .ZN(n14651) );
  AOI21_X1 U16532 ( .B1(n14649), .B2(n14426), .A(n14654), .ZN(n21455) );
  AOI22_X1 U16533 ( .A1(n19925), .A2(n21455), .B1(n15724), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n14650) );
  OAI21_X1 U16534 ( .B1(n14651), .B2(n15726), .A(n14650), .ZN(P1_U2868) );
  INV_X1 U16535 ( .A(n15770), .ZN(n14652) );
  INV_X1 U16536 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19830) );
  OAI222_X1 U16537 ( .A1(n15796), .A2(n14652), .B1(n15801), .B2(n14651), .C1(
        n19830), .C2(n15794), .ZN(P1_U2900) );
  OR2_X1 U16538 ( .A1(n14654), .A2(n14653), .ZN(n14655) );
  NAND2_X1 U16539 ( .A1(n14798), .A2(n14655), .ZN(n21471) );
  INV_X1 U16540 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14659) );
  AND2_X1 U16541 ( .A1(n14656), .A2(n14657), .ZN(n14801) );
  NOR2_X1 U16542 ( .A1(n14656), .A2(n14657), .ZN(n14658) );
  OAI222_X1 U16543 ( .A1(n21471), .A2(n19942), .B1(n14659), .B2(n19946), .C1(
        n19953), .C2(n15726), .ZN(P1_U2867) );
  INV_X1 U16544 ( .A(n14662), .ZN(n21906) );
  NAND2_X1 U16545 ( .A1(n21906), .A2(n21456), .ZN(n14664) );
  AOI22_X1 U16546 ( .A1(n21597), .A2(P1_EBX_REG_1__SCAN_IN), .B1(n21493), .B2(
        n14210), .ZN(n14663) );
  OAI211_X1 U16547 ( .C1(n14665), .C2(n21638), .A(n14664), .B(n14663), .ZN(
        n14666) );
  AOI21_X1 U16548 ( .B1(n14660), .B2(P1_REIP_REG_1__SCAN_IN), .A(n14666), .ZN(
        n14667) );
  OAI21_X1 U16549 ( .B1(n21613), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14667), .ZN(n14668) );
  AOI21_X1 U16550 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21615), .A(
        n14668), .ZN(n14669) );
  OAI21_X1 U16551 ( .B1(n21440), .B2(n14670), .A(n14669), .ZN(P1_U2839) );
  INV_X1 U16552 ( .A(n15762), .ZN(n14671) );
  INV_X1 U16553 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n19832) );
  OAI222_X1 U16554 ( .A1(n15796), .A2(n14671), .B1(n15794), .B2(n19832), .C1(
        n15801), .C2(n19953), .ZN(P1_U2899) );
  INV_X1 U16555 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15348) );
  INV_X1 U16556 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n14872) );
  INV_X1 U16557 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14672) );
  OAI22_X1 U16558 ( .A1(n15264), .A2(n14872), .B1(n15263), .B2(n14672), .ZN(
        n14673) );
  AOI21_X1 U16559 ( .B1(n15294), .B2(P2_REIP_REG_8__SCAN_IN), .A(n14673), .ZN(
        n14674) );
  OAI21_X1 U16560 ( .B1(n15297), .B2(n15348), .A(n14674), .ZN(n14675) );
  INV_X1 U16561 ( .A(n14675), .ZN(n14678) );
  AOI21_X1 U16562 ( .B1(n14678), .B2(n14677), .A(n11210), .ZN(n18557) );
  INV_X1 U16563 ( .A(n18557), .ZN(n14879) );
  OAI211_X1 U16564 ( .C1(n14681), .C2(n14680), .A(n14679), .B(n16266), .ZN(
        n14683) );
  NAND2_X1 U16565 ( .A1(n10963), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14682) );
  OAI211_X1 U16566 ( .C1(n14879), .C2(n10963), .A(n14683), .B(n14682), .ZN(
        P2_U2879) );
  NAND2_X1 U16567 ( .A1(n14685), .A2(n14684), .ZN(n14686) );
  NAND2_X1 U16568 ( .A1(n14687), .A2(n14686), .ZN(n19954) );
  NAND2_X1 U16569 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21308) );
  INV_X1 U16570 ( .A(n21308), .ZN(n21313) );
  INV_X1 U16571 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14690) );
  NAND2_X1 U16572 ( .A1(n21313), .A2(n14690), .ZN(n21315) );
  NOR3_X1 U16573 ( .A1(n14688), .A2(n21308), .A3(n14690), .ZN(n15936) );
  INV_X1 U16574 ( .A(n15936), .ZN(n14689) );
  NAND3_X1 U16575 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21313), .ZN(n15934) );
  AOI21_X1 U16576 ( .B1(n21366), .B2(n15934), .A(n21401), .ZN(n21348) );
  INV_X1 U16577 ( .A(n21348), .ZN(n21321) );
  AOI21_X1 U16578 ( .B1(n16033), .B2(n14689), .A(n21321), .ZN(n21314) );
  OAI22_X1 U16579 ( .A1(n14691), .A2(n21315), .B1(n21314), .B2(n14690), .ZN(
        n14694) );
  INV_X1 U16580 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n14692) );
  OAI22_X1 U16581 ( .A1(n21414), .A2(n21471), .B1(n21419), .B2(n14692), .ZN(
        n14693) );
  AOI211_X1 U16582 ( .C1(n19954), .C2(n21422), .A(n14694), .B(n14693), .ZN(
        n14695) );
  INV_X1 U16583 ( .A(n14695), .ZN(P1_U3026) );
  INV_X1 U16584 ( .A(n15755), .ZN(n14700) );
  NAND2_X1 U16585 ( .A1(n14698), .A2(n14697), .ZN(n14699) );
  NAND2_X1 U16586 ( .A1(n14696), .A2(n14699), .ZN(n21500) );
  OAI222_X1 U16587 ( .A1(n15796), .A2(n14700), .B1(n15794), .B2(n11948), .C1(
        n15801), .C2(n21500), .ZN(P1_U2897) );
  INV_X1 U16588 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n14711) );
  OAI211_X1 U16589 ( .C1(n13169), .C2(n11406), .A(n16266), .B(n14701), .ZN(
        n14710) );
  NAND2_X1 U16590 ( .A1(n15285), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n14703) );
  NAND2_X1 U16591 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14702) );
  OAI211_X1 U16592 ( .C1(n15300), .C2(n14704), .A(n14703), .B(n14702), .ZN(
        n14705) );
  AOI21_X1 U16593 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n14705), .ZN(n14706) );
  AND2_X1 U16594 ( .A1(n14707), .A2(n14706), .ZN(n14708) );
  OR2_X1 U16595 ( .A1(n14708), .A2(n14854), .ZN(n16475) );
  INV_X1 U16596 ( .A(n16475), .ZN(n18282) );
  NAND2_X1 U16597 ( .A1(n18282), .A2(n11059), .ZN(n14709) );
  OAI211_X1 U16598 ( .C1(n11059), .C2(n14711), .A(n14710), .B(n14709), .ZN(
        P2_U2878) );
  AOI21_X1 U16599 ( .B1(n17106), .B2(n14712), .A(n14834), .ZN(n17097) );
  INV_X1 U16600 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15561) );
  INV_X1 U16601 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16452) );
  INV_X1 U16602 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18330) );
  INV_X1 U16603 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16094) );
  INV_X1 U16604 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16426) );
  INV_X1 U16605 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16413) );
  INV_X1 U16606 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16390) );
  INV_X1 U16607 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16091) );
  INV_X1 U16608 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16101) );
  INV_X1 U16609 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16355) );
  INV_X1 U16610 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16111) );
  XNOR2_X1 U16611 ( .A(n14713), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16343) );
  OAI22_X1 U16612 ( .A1(n14714), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n18247) );
  OAI22_X1 U16613 ( .A1(n14714), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13873), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16163) );
  AND2_X1 U16614 ( .A1(n18247), .A2(n16163), .ZN(n16149) );
  NAND2_X1 U16615 ( .A1(n16149), .A2(n16150), .ZN(n14835) );
  NAND2_X1 U16616 ( .A1(n18423), .A2(n14835), .ZN(n14715) );
  XNOR2_X1 U16617 ( .A(n17097), .B(n14715), .ZN(n14741) );
  NOR4_X1 U16618 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n15263), .ZN(n14716) );
  OR2_X1 U16619 ( .A1(n14718), .A2(n14717), .ZN(n14719) );
  NAND2_X1 U16620 ( .A1(n14719), .A2(n14846), .ZN(n17221) );
  INV_X1 U16621 ( .A(n17221), .ZN(n19470) );
  NAND2_X1 U16622 ( .A1(n18221), .A2(n11085), .ZN(n14737) );
  INV_X1 U16623 ( .A(n18222), .ZN(n21699) );
  NOR2_X1 U16624 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n21699), .ZN(n14725) );
  INV_X1 U16625 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n18489) );
  MUX2_X1 U16626 ( .A(n14722), .B(n14732), .S(n19381), .Z(n14723) );
  OAI21_X1 U16627 ( .B1(n14724), .B2(n14723), .A(n14842), .ZN(n15038) );
  OAI22_X1 U16628 ( .A1(n14142), .A2(n14726), .B1(P2_EBX_REG_31__SCAN_IN), 
        .B2(n14725), .ZN(n14728) );
  AND2_X1 U16629 ( .A1(n14728), .A2(n14727), .ZN(n14729) );
  NAND2_X1 U16630 ( .A1(n18221), .A2(n14729), .ZN(n18490) );
  NAND2_X1 U16631 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19214), .ZN(n18604) );
  NOR3_X1 U16632 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n17222), .A3(n18604), 
        .ZN(n18610) );
  INV_X1 U16633 ( .A(n18559), .ZN(n18521) );
  INV_X1 U16634 ( .A(n18482), .ZN(n18602) );
  NAND2_X1 U16635 ( .A1(n18521), .A2(n18602), .ZN(n14730) );
  OR2_X1 U16636 ( .A1(n18610), .A2(n14730), .ZN(n14731) );
  OAI22_X1 U16637 ( .A1(n18490), .A2(n14732), .B1(n17106), .B2(n18329), .ZN(
        n14733) );
  INV_X1 U16638 ( .A(n14733), .ZN(n14735) );
  NAND2_X1 U16639 ( .A1(n18473), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n14734) );
  OAI211_X1 U16640 ( .C1(n18494), .C2(n15038), .A(n14735), .B(n14734), .ZN(
        n14736) );
  AOI21_X1 U16641 ( .B1(n19470), .B2(n18500), .A(n14736), .ZN(n14739) );
  OR2_X1 U16642 ( .A1(n17101), .A2(n18478), .ZN(n14738) );
  OAI211_X1 U16643 ( .C1(n19239), .C2(n18241), .A(n14739), .B(n14738), .ZN(
        n14740) );
  AOI21_X1 U16644 ( .B1(n14741), .B2(n18482), .A(n14740), .ZN(n14742) );
  INV_X1 U16645 ( .A(n14742), .ZN(P2_U2852) );
  INV_X1 U16646 ( .A(n14696), .ZN(n14744) );
  OAI21_X1 U16647 ( .B1(n14744), .B2(n11396), .A(n14743), .ZN(n15094) );
  INV_X1 U16648 ( .A(n15090), .ZN(n14757) );
  INV_X1 U16649 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14750) );
  AND2_X1 U16650 ( .A1(n21483), .A2(n14745), .ZN(n21557) );
  INV_X1 U16651 ( .A(n21557), .ZN(n21485) );
  INV_X1 U16652 ( .A(n14746), .ZN(n14748) );
  INV_X1 U16653 ( .A(n14816), .ZN(n14747) );
  NAND3_X1 U16654 ( .A1(n21493), .A2(n14748), .A3(n14747), .ZN(n14749) );
  OAI211_X1 U16655 ( .C1(n21623), .C2(n14750), .A(n21485), .B(n14749), .ZN(
        n14756) );
  OAI21_X1 U16656 ( .B1(n14816), .B2(n21484), .A(n21483), .ZN(n14815) );
  INV_X1 U16657 ( .A(n19941), .ZN(n14797) );
  AOI21_X1 U16658 ( .B1(n14797), .B2(n19939), .A(n14751), .ZN(n14752) );
  NOR2_X1 U16659 ( .A1(n14752), .A2(n14942), .ZN(n21333) );
  AOI22_X1 U16660 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14815), .B1(n21590), 
        .B2(n21333), .ZN(n14753) );
  OAI21_X1 U16661 ( .B1(n14754), .B2(n21626), .A(n14753), .ZN(n14755) );
  AOI211_X1 U16662 ( .C1(n21634), .C2(n14757), .A(n14756), .B(n14755), .ZN(
        n14758) );
  OAI21_X1 U16663 ( .B1(n15094), .B2(n21630), .A(n14758), .ZN(P1_U2832) );
  AOI22_X1 U16664 ( .A1(n21333), .A2(n19925), .B1(n15724), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n14759) );
  OAI21_X1 U16665 ( .B1(n15094), .B2(n15726), .A(n14759), .ZN(P1_U2864) );
  OAI21_X1 U16666 ( .B1(n22202), .B2(n14793), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14761) );
  NAND2_X1 U16667 ( .A1(n21817), .A2(n14662), .ZN(n14760) );
  AOI21_X1 U16668 ( .B1(n14761), .B2(n14760), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n14764) );
  NOR2_X1 U16669 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14762), .ZN(
        n14765) );
  INV_X1 U16670 ( .A(n14766), .ZN(n14763) );
  NOR2_X1 U16671 ( .A1(n14763), .A2(n21922), .ZN(n21850) );
  NAND2_X1 U16672 ( .A1(n14789), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n14770) );
  INV_X1 U16673 ( .A(n14765), .ZN(n14791) );
  NOR2_X1 U16674 ( .A1(n21906), .A2(n21924), .ZN(n14767) );
  INV_X1 U16675 ( .A(n21830), .ZN(n21849) );
  NOR2_X1 U16676 ( .A1(n14766), .A2(n21922), .ZN(n21907) );
  AOI22_X1 U16677 ( .A1(n21817), .A2(n14767), .B1(n11386), .B2(n21907), .ZN(
        n14790) );
  OAI22_X1 U16678 ( .A1(n22034), .A2(n14791), .B1(n14790), .B2(n22043), .ZN(
        n14768) );
  AOI21_X1 U16679 ( .B1(n14793), .B2(n22040), .A(n14768), .ZN(n14769) );
  OAI211_X1 U16680 ( .C1(n14796), .C2(n22056), .A(n14770), .B(n14769), .ZN(
        P1_U3068) );
  NAND2_X1 U16681 ( .A1(n14789), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n14773) );
  OAI22_X1 U16682 ( .A1(n21852), .A2(n14791), .B1(n14790), .B2(n21889), .ZN(
        n14771) );
  AOI21_X1 U16683 ( .B1(n14793), .B2(n21881), .A(n14771), .ZN(n14772) );
  OAI211_X1 U16684 ( .C1(n14796), .C2(n21938), .A(n14773), .B(n14772), .ZN(
        P1_U3065) );
  NAND2_X1 U16685 ( .A1(n14789), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n14776) );
  OAI22_X1 U16686 ( .A1(n21956), .A2(n14791), .B1(n14790), .B2(n21965), .ZN(
        n14774) );
  AOI21_X1 U16687 ( .B1(n14793), .B2(n21962), .A(n14774), .ZN(n14775) );
  OAI211_X1 U16688 ( .C1(n14796), .C2(n21978), .A(n14776), .B(n14775), .ZN(
        P1_U3066) );
  NAND2_X1 U16689 ( .A1(n14789), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n14779) );
  OAI22_X1 U16690 ( .A1(n22115), .A2(n14791), .B1(n14790), .B2(n22124), .ZN(
        n14777) );
  AOI21_X1 U16691 ( .B1(n14793), .B2(n22121), .A(n14777), .ZN(n14778) );
  OAI211_X1 U16692 ( .C1(n14796), .C2(n22137), .A(n14779), .B(n14778), .ZN(
        P1_U3070) );
  NAND2_X1 U16693 ( .A1(n14789), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n14782) );
  OAI22_X1 U16694 ( .A1(n22228), .A2(n14791), .B1(n14790), .B2(n22247), .ZN(
        n14780) );
  AOI21_X1 U16695 ( .B1(n14793), .B2(n22242), .A(n14780), .ZN(n14781) );
  OAI211_X1 U16696 ( .C1(n14796), .C2(n22275), .A(n14782), .B(n14781), .ZN(
        P1_U3072) );
  NAND2_X1 U16697 ( .A1(n14789), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14785) );
  OAI22_X1 U16698 ( .A1(n22076), .A2(n14791), .B1(n14790), .B2(n22085), .ZN(
        n14783) );
  AOI21_X1 U16699 ( .B1(n14793), .B2(n22082), .A(n14783), .ZN(n14784) );
  OAI211_X1 U16700 ( .C1(n14796), .C2(n22098), .A(n14785), .B(n14784), .ZN(
        P1_U3069) );
  NAND2_X1 U16701 ( .A1(n14789), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n14788) );
  OAI22_X1 U16702 ( .A1(n21995), .A2(n14791), .B1(n14790), .B2(n22004), .ZN(
        n14786) );
  AOI21_X1 U16703 ( .B1(n14793), .B2(n22001), .A(n14786), .ZN(n14787) );
  OAI211_X1 U16704 ( .C1(n14796), .C2(n22017), .A(n14788), .B(n14787), .ZN(
        P1_U3067) );
  NAND2_X1 U16705 ( .A1(n14789), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n14795) );
  OAI22_X1 U16706 ( .A1(n22156), .A2(n14791), .B1(n14790), .B2(n22167), .ZN(
        n14792) );
  AOI21_X1 U16707 ( .B1(n14793), .B2(n22164), .A(n14792), .ZN(n14794) );
  OAI211_X1 U16708 ( .C1(n14796), .C2(n22180), .A(n14795), .B(n14794), .ZN(
        P1_U3071) );
  AOI21_X1 U16709 ( .B1(n14799), .B2(n14798), .A(n14797), .ZN(n21480) );
  INV_X1 U16710 ( .A(n21480), .ZN(n14802) );
  XOR2_X1 U16711 ( .A(n14800), .B(n14801), .Z(n21489) );
  INV_X1 U16712 ( .A(n21489), .ZN(n14806) );
  INV_X1 U16713 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21487) );
  OAI222_X1 U16714 ( .A1(n14802), .A2(n19942), .B1(n15726), .B2(n14806), .C1(
        n19946), .C2(n21487), .ZN(P1_U2866) );
  INV_X1 U16715 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14805) );
  OR2_X1 U16716 ( .A1(n15727), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14804) );
  INV_X1 U16717 ( .A(DATAI_8_), .ZN(n17041) );
  NAND2_X1 U16718 ( .A1(n15727), .A2(n17041), .ZN(n14803) );
  NAND2_X1 U16719 ( .A1(n14804), .A2(n14803), .ZN(n21734) );
  OAI222_X1 U16720 ( .A1(n15094), .A2(n15801), .B1(n15794), .B2(n14805), .C1(
        n21734), .C2(n15796), .ZN(P1_U2896) );
  INV_X1 U16721 ( .A(n15758), .ZN(n14807) );
  OAI222_X1 U16722 ( .A1(n15796), .A2(n14807), .B1(n15794), .B2(n11934), .C1(
        n15801), .C2(n14806), .ZN(P1_U2898) );
  AOI21_X1 U16723 ( .B1(n14810), .B2(n14743), .A(n14809), .ZN(n14811) );
  INV_X1 U16724 ( .A(n14811), .ZN(n15231) );
  XNOR2_X1 U16725 ( .A(n14942), .B(n14940), .ZN(n21345) );
  AOI22_X1 U16726 ( .A1(n21345), .A2(n19925), .B1(n15724), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n14812) );
  OAI21_X1 U16727 ( .B1(n15231), .B2(n15726), .A(n14812), .ZN(P1_U2863) );
  INV_X1 U16728 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15226) );
  OAI22_X1 U16729 ( .A1(n15226), .A2(n21626), .B1(n21613), .B2(n14813), .ZN(
        n14814) );
  AOI211_X1 U16730 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n14815), .A(n21557), .B(
        n14814), .ZN(n14821) );
  NAND2_X1 U16731 ( .A1(n14816), .A2(n21493), .ZN(n14818) );
  AOI22_X1 U16732 ( .A1(n21345), .A2(n21590), .B1(n21597), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n14817) );
  OAI21_X1 U16733 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(n14818), .A(n14817), .ZN(
        n14819) );
  INV_X1 U16734 ( .A(n14819), .ZN(n14820) );
  OAI211_X1 U16735 ( .C1(n15231), .C2(n21630), .A(n14821), .B(n14820), .ZN(
        P1_U2831) );
  INV_X1 U16736 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14824) );
  OR2_X1 U16737 ( .A1(n15727), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14823) );
  INV_X1 U16738 ( .A(DATAI_9_), .ZN(n16904) );
  NAND2_X1 U16739 ( .A1(n15727), .A2(n16904), .ZN(n14822) );
  NAND2_X1 U16740 ( .A1(n14823), .A2(n14822), .ZN(n15743) );
  OAI222_X1 U16741 ( .A1(n15231), .A2(n15801), .B1(n15794), .B2(n14824), .C1(
        n15743), .C2(n15796), .ZN(P1_U2895) );
  XNOR2_X1 U16742 ( .A(n14825), .B(n14948), .ZN(n14833) );
  INV_X1 U16743 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n16457) );
  NAND2_X1 U16744 ( .A1(n15556), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n14827) );
  NAND2_X1 U16745 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14826) );
  OAI211_X1 U16746 ( .C1(n15300), .C2(n16457), .A(n14827), .B(n14826), .ZN(
        n14828) );
  AOI21_X1 U16747 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n14828), .ZN(n14831) );
  INV_X1 U16748 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16705) );
  AOI22_X1 U16749 ( .A1(n15285), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n14830) );
  NAND2_X1 U16750 ( .A1(n15294), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n14829) );
  OAI211_X1 U16751 ( .C1(n15297), .C2(n16705), .A(n14830), .B(n14829), .ZN(
        n14853) );
  AOI21_X1 U16752 ( .B1(n14831), .B2(n14855), .A(n14901), .ZN(n18301) );
  INV_X1 U16753 ( .A(n18301), .ZN(n16697) );
  INV_X1 U16754 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n18299) );
  MUX2_X1 U16755 ( .A(n16697), .B(n18299), .S(n10963), .Z(n14832) );
  OAI21_X1 U16756 ( .B1(n14833), .B2(n16253), .A(n14832), .ZN(P2_U2876) );
  OAI21_X1 U16757 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n14834), .A(
        n14863), .ZN(n17112) );
  INV_X1 U16758 ( .A(n17112), .ZN(n14838) );
  NOR2_X1 U16759 ( .A1(n17097), .A2(n14835), .ZN(n14864) );
  NOR2_X1 U16760 ( .A1(n18436), .A2(n14864), .ZN(n14837) );
  AOI21_X1 U16761 ( .B1(n14838), .B2(n14837), .A(n18602), .ZN(n14836) );
  OAI21_X1 U16762 ( .B1(n14838), .B2(n14837), .A(n14836), .ZN(n14852) );
  MUX2_X1 U16763 ( .A(n14840), .B(n14839), .S(n19381), .Z(n14843) );
  OAI21_X1 U16764 ( .B1(n14843), .B2(n11149), .A(n11038), .ZN(n15129) );
  OAI21_X1 U16765 ( .B1(n14844), .B2(n18329), .A(n14141), .ZN(n14848) );
  XNOR2_X1 U16766 ( .A(n14846), .B(n14845), .ZN(n15061) );
  OAI22_X1 U16767 ( .A1(n18476), .A2(n15061), .B1(n13663), .B2(n18493), .ZN(
        n14847) );
  AOI211_X1 U16768 ( .C1(P2_EBX_REG_4__SCAN_IN), .C2(n18470), .A(n14848), .B(
        n14847), .ZN(n14849) );
  OAI21_X1 U16769 ( .B1(n15129), .B2(n18494), .A(n14849), .ZN(n14850) );
  AOI21_X1 U16770 ( .B1(n18501), .B2(n17108), .A(n14850), .ZN(n14851) );
  OAI211_X1 U16771 ( .C1(n19372), .C2(n18241), .A(n14852), .B(n14851), .ZN(
        P2_U2851) );
  OR2_X1 U16772 ( .A1(n14854), .A2(n14853), .ZN(n14856) );
  AND2_X1 U16773 ( .A1(n14856), .A2(n14855), .ZN(n18292) );
  INV_X1 U16774 ( .A(n18292), .ZN(n14862) );
  INV_X1 U16775 ( .A(n14701), .ZN(n14859) );
  INV_X1 U16776 ( .A(n14825), .ZN(n14857) );
  OAI211_X1 U16777 ( .C1(n14859), .C2(n14858), .A(n14857), .B(n16266), .ZN(
        n14861) );
  NAND2_X1 U16778 ( .A1(n10963), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14860) );
  OAI211_X1 U16779 ( .C1(n14862), .C2(n10963), .A(n14861), .B(n14860), .ZN(
        P2_U2877) );
  AOI21_X1 U16780 ( .B1(n16485), .B2(n14865), .A(n14866), .ZN(n18261) );
  AOI21_X1 U16781 ( .B1(n18249), .B2(n14863), .A(n10983), .ZN(n18255) );
  NAND2_X1 U16782 ( .A1(n14864), .A2(n17112), .ZN(n18253) );
  NOR2_X1 U16783 ( .A1(n18255), .A2(n18253), .ZN(n14883) );
  OAI21_X1 U16784 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10983), .A(
        n14865), .ZN(n17120) );
  NAND2_X1 U16785 ( .A1(n14883), .A2(n17120), .ZN(n18260) );
  NOR2_X1 U16786 ( .A1(n18261), .A2(n18260), .ZN(n15072) );
  NOR2_X1 U16787 ( .A1(n18436), .A2(n15072), .ZN(n14867) );
  OAI21_X1 U16788 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n14866), .A(
        n15071), .ZN(n17134) );
  XNOR2_X1 U16789 ( .A(n14867), .B(n17134), .ZN(n14868) );
  NAND2_X1 U16790 ( .A1(n14868), .A2(n18482), .ZN(n14878) );
  AOI21_X1 U16791 ( .B1(n14869), .B2(n16739), .A(n16723), .ZN(n19102) );
  AOI22_X1 U16792 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18498), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18473), .ZN(n14870) );
  OAI211_X1 U16793 ( .C1(n18490), .C2(n14872), .A(n14870), .B(n14141), .ZN(
        n14876) );
  MUX2_X1 U16794 ( .A(n18248), .B(n14871), .S(n15490), .Z(n15123) );
  MUX2_X1 U16795 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n15336), .S(n15490), .Z(
        n14886) );
  MUX2_X1 U16796 ( .A(n14644), .B(n11050), .S(n15490), .Z(n15345) );
  NOR2_X1 U16797 ( .A1(n15490), .A2(n14872), .ZN(n14873) );
  NAND2_X1 U16798 ( .A1(n15533), .A2(n14873), .ZN(n14874) );
  NAND2_X1 U16799 ( .A1(n15358), .A2(n14874), .ZN(n15343) );
  NOR2_X1 U16800 ( .A1(n15343), .A2(n18494), .ZN(n14875) );
  AOI211_X1 U16801 ( .C1(n18500), .C2(n19102), .A(n14876), .B(n14875), .ZN(
        n14877) );
  OAI211_X1 U16802 ( .C1(n18478), .C2(n14879), .A(n14878), .B(n14877), .ZN(
        P2_U2847) );
  INV_X1 U16803 ( .A(n14880), .ZN(n14881) );
  XNOR2_X1 U16804 ( .A(n14882), .B(n14881), .ZN(n16764) );
  INV_X1 U16805 ( .A(n16764), .ZN(n19328) );
  NOR2_X1 U16806 ( .A1(n18436), .A2(n14883), .ZN(n14884) );
  XNOR2_X1 U16807 ( .A(n14884), .B(n17120), .ZN(n14885) );
  NAND2_X1 U16808 ( .A1(n14885), .A2(n18482), .ZN(n14893) );
  INV_X1 U16809 ( .A(n17114), .ZN(n14891) );
  XNOR2_X1 U16810 ( .A(n15126), .B(n14886), .ZN(n15339) );
  NOR2_X1 U16811 ( .A1(n18494), .A2(n15339), .ZN(n14890) );
  NAND2_X1 U16812 ( .A1(n18470), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n14888) );
  AOI21_X1 U16813 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18498), .A(
        n18559), .ZN(n14887) );
  OAI211_X1 U16814 ( .C1(n18493), .C2(n17272), .A(n14888), .B(n14887), .ZN(
        n14889) );
  AOI211_X1 U16815 ( .C1(n14891), .C2(n18501), .A(n14890), .B(n14889), .ZN(
        n14892) );
  OAI211_X1 U16816 ( .C1(n19328), .C2(n18476), .A(n14893), .B(n14892), .ZN(
        P2_U2849) );
  INV_X1 U16817 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n16128) );
  AND2_X1 U16818 ( .A1(n14825), .A2(n14894), .ZN(n14950) );
  NAND2_X1 U16819 ( .A1(n14825), .A2(n14895), .ZN(n14919) );
  OAI211_X1 U16820 ( .C1(n14950), .C2(n14896), .A(n14919), .B(n16266), .ZN(
        n14910) );
  INV_X1 U16821 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n16143) );
  NAND2_X1 U16822 ( .A1(n15285), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14898) );
  NAND2_X1 U16823 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14897) );
  OAI211_X1 U16824 ( .C1(n15300), .C2(n16143), .A(n14898), .B(n14897), .ZN(
        n14899) );
  INV_X1 U16825 ( .A(n14899), .ZN(n14900) );
  OAI21_X1 U16826 ( .B1(n15297), .B2(n18530), .A(n14900), .ZN(n14946) );
  NAND2_X1 U16827 ( .A1(n15285), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n14903) );
  NAND2_X1 U16828 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14902) );
  OAI211_X1 U16829 ( .C1(n15300), .C2(n16453), .A(n14903), .B(n14902), .ZN(
        n14904) );
  AOI21_X1 U16830 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n14904), .ZN(n14906) );
  INV_X1 U16831 ( .A(n14915), .ZN(n14917) );
  NAND2_X1 U16832 ( .A1(n14905), .A2(n14906), .ZN(n14907) );
  NAND2_X1 U16833 ( .A1(n14917), .A2(n14907), .ZN(n16684) );
  INV_X1 U16834 ( .A(n16684), .ZN(n14908) );
  NAND2_X1 U16835 ( .A1(n11059), .A2(n14908), .ZN(n14909) );
  OAI211_X1 U16836 ( .C1(n11059), .C2(n16128), .A(n14910), .B(n14909), .ZN(
        P2_U2874) );
  NAND2_X1 U16837 ( .A1(n15556), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14912) );
  NAND2_X1 U16838 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14911) );
  OAI211_X1 U16839 ( .C1(n15300), .C2(n17274), .A(n14912), .B(n14911), .ZN(
        n14913) );
  AOI21_X1 U16840 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n14913), .ZN(n14918) );
  INV_X1 U16841 ( .A(n14918), .ZN(n14914) );
  NAND2_X1 U16842 ( .A1(n14915), .A2(n14914), .ZN(n14972) );
  INV_X1 U16843 ( .A(n14972), .ZN(n14916) );
  AOI21_X1 U16844 ( .B1(n14918), .B2(n14917), .A(n14916), .ZN(n16439) );
  INV_X1 U16845 ( .A(n16439), .ZN(n16672) );
  INV_X1 U16846 ( .A(n14919), .ZN(n14922) );
  OAI211_X1 U16847 ( .C1(n14922), .C2(n14921), .A(n16266), .B(n14920), .ZN(
        n14924) );
  NAND2_X1 U16848 ( .A1(n10963), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n14923) );
  OAI211_X1 U16849 ( .C1(n16672), .C2(n10963), .A(n14924), .B(n14923), .ZN(
        P2_U2873) );
  INV_X1 U16850 ( .A(n19575), .ZN(n14925) );
  XOR2_X1 U16851 ( .A(n19575), .B(n19142), .Z(n19578) );
  NOR2_X1 U16852 ( .A1(n19578), .A2(n19577), .ZN(n19576) );
  AOI21_X1 U16853 ( .B1(n14925), .B2(n19142), .A(n19576), .ZN(n14928) );
  XNOR2_X1 U16854 ( .A(n14927), .B(n14926), .ZN(n19523) );
  XNOR2_X1 U16855 ( .A(n14928), .B(n19523), .ZN(n19526) );
  NAND2_X1 U16856 ( .A1(n14928), .A2(n19523), .ZN(n14929) );
  OAI21_X1 U16857 ( .B1(n19526), .B2(n19238), .A(n14929), .ZN(n19472) );
  XNOR2_X1 U16858 ( .A(n19239), .B(n17221), .ZN(n19473) );
  NOR2_X1 U16859 ( .A1(n19472), .A2(n19473), .ZN(n19471) );
  NOR2_X1 U16860 ( .A1(n19110), .A2(n19470), .ZN(n14930) );
  OAI21_X1 U16861 ( .B1(n19471), .B2(n14930), .A(n15061), .ZN(n19374) );
  XOR2_X1 U16862 ( .A(n19372), .B(n19374), .Z(n14934) );
  INV_X1 U16863 ( .A(n15061), .ZN(n14931) );
  AOI22_X1 U16864 ( .A1(n19633), .A2(n14931), .B1(n19627), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n14933) );
  NAND2_X1 U16865 ( .A1(n19524), .A2(n19428), .ZN(n14932) );
  OAI211_X1 U16866 ( .C1(n14934), .C2(n19579), .A(n14933), .B(n14932), .ZN(
        P2_U2915) );
  OAI21_X1 U16867 ( .B1(n14809), .B2(n14936), .A(n14935), .ZN(n15930) );
  INV_X1 U16868 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14939) );
  OR2_X1 U16869 ( .A1(n15727), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14938) );
  INV_X1 U16870 ( .A(DATAI_10_), .ZN(n17035) );
  NAND2_X1 U16871 ( .A1(n15727), .A2(n17035), .ZN(n14937) );
  NAND2_X1 U16872 ( .A1(n14938), .A2(n14937), .ZN(n21747) );
  OAI222_X1 U16873 ( .A1(n15930), .A2(n15801), .B1(n15794), .B2(n14939), .C1(
        n21747), .C2(n15796), .ZN(P1_U2894) );
  INV_X1 U16874 ( .A(n14940), .ZN(n14941) );
  NAND2_X1 U16875 ( .A1(n14942), .A2(n14941), .ZN(n14944) );
  NAND2_X1 U16876 ( .A1(n14944), .A2(n14943), .ZN(n14945) );
  NAND2_X1 U16877 ( .A1(n14945), .A2(n19922), .ZN(n21354) );
  INV_X1 U16878 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14953) );
  OAI222_X1 U16879 ( .A1(n21354), .A2(n19942), .B1(n14953), .B2(n19946), .C1(
        n15726), .C2(n15930), .ZN(P1_U2862) );
  OAI21_X1 U16880 ( .B1(n14946), .B2(n14901), .A(n14905), .ZN(n16139) );
  AOI21_X1 U16881 ( .B1(n14825), .B2(n14948), .A(n14947), .ZN(n14949) );
  OR3_X1 U16882 ( .A1(n14950), .A2(n14949), .A3(n16253), .ZN(n14952) );
  NAND2_X1 U16883 ( .A1(n10963), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14951) );
  OAI211_X1 U16884 ( .C1(n16139), .C2(n10963), .A(n14952), .B(n14951), .ZN(
        P2_U2875) );
  INV_X1 U16885 ( .A(n15930), .ZN(n14963) );
  OAI22_X1 U16886 ( .A1(n21354), .A2(n21638), .B1(n21623), .B2(n14953), .ZN(
        n14954) );
  INV_X1 U16887 ( .A(n14954), .ZN(n14958) );
  INV_X1 U16888 ( .A(n14955), .ZN(n14956) );
  NAND3_X1 U16889 ( .A1(n14956), .A2(n19857), .A3(n21493), .ZN(n14957) );
  NAND2_X1 U16890 ( .A1(n14958), .A2(n14957), .ZN(n14962) );
  OAI21_X1 U16891 ( .B1(n15652), .B2(n21484), .A(n21483), .ZN(n21508) );
  NAND2_X1 U16892 ( .A1(n21508), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n14960) );
  AOI21_X1 U16893 ( .B1(n21615), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n21557), .ZN(n14959) );
  OAI211_X1 U16894 ( .C1(n15926), .C2(n21613), .A(n14960), .B(n14959), .ZN(
        n14961) );
  AOI211_X1 U16895 ( .C1(n14963), .C2(n21618), .A(n14962), .B(n14961), .ZN(
        n14964) );
  INV_X1 U16896 ( .A(n14964), .ZN(P1_U2830) );
  INV_X1 U16897 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14977) );
  INV_X1 U16898 ( .A(n14920), .ZN(n14966) );
  OAI211_X1 U16899 ( .C1(n14966), .C2(n14965), .A(n16266), .B(n11037), .ZN(
        n14976) );
  NAND2_X1 U16900 ( .A1(n15285), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14968) );
  NAND2_X1 U16901 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14967) );
  OAI211_X1 U16902 ( .C1(n15300), .C2(n14969), .A(n14968), .B(n14967), .ZN(
        n14970) );
  AOI21_X1 U16903 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n14970), .ZN(n14971) );
  NAND2_X1 U16904 ( .A1(n14972), .A2(n14971), .ZN(n14974) );
  INV_X1 U16905 ( .A(n15180), .ZN(n14973) );
  NAND2_X1 U16906 ( .A1(n11059), .A2(n18318), .ZN(n14975) );
  OAI211_X1 U16907 ( .C1(n11059), .C2(n14977), .A(n14976), .B(n14975), .ZN(
        P2_U2872) );
  AND2_X1 U16908 ( .A1(n14978), .A2(n18244), .ZN(n14984) );
  AND2_X2 U16909 ( .A1(n14982), .A2(n14988), .ZN(n19139) );
  INV_X1 U16910 ( .A(n14980), .ZN(n14981) );
  NOR2_X1 U16911 ( .A1(n14979), .A2(n14981), .ZN(n14985) );
  AND2_X2 U16912 ( .A1(n14983), .A2(n14988), .ZN(n19115) );
  AOI22_X1 U16913 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19139), .B1(
        n19115), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14993) );
  AND2_X2 U16914 ( .A1(n14983), .A2(n17101), .ZN(n19204) );
  AOI22_X1 U16915 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19232), .B1(
        n19204), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14992) );
  AOI22_X1 U16916 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n15095), .B1(
        n15096), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14991) );
  AOI22_X1 U16917 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19265), .B1(
        n19185), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14990) );
  AND4_X1 U16918 ( .A1(n14993), .A2(n14992), .A3(n14991), .A4(n14990), .ZN(
        n15013) );
  AND2_X1 U16919 ( .A1(n14995), .A2(n14994), .ZN(n15000) );
  OAI22_X1 U16920 ( .A1(n14997), .A2(n15104), .B1(n19154), .B2(n14996), .ZN(
        n15004) );
  INV_X1 U16921 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15001) );
  OAI22_X1 U16922 ( .A1(n15002), .A2(n15328), .B1(n15103), .B2(n15001), .ZN(
        n15003) );
  NOR2_X1 U16923 ( .A1(n15004), .A2(n15003), .ZN(n15012) );
  NOR2_X2 U16924 ( .A1(n15007), .A2(n10973), .ZN(n19274) );
  NAND2_X1 U16925 ( .A1(n14986), .A2(n15006), .ZN(n15009) );
  NOR2_X2 U16926 ( .A1(n15009), .A2(n16170), .ZN(n19196) );
  AOI22_X1 U16927 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19274), .B1(
        n19196), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15011) );
  INV_X1 U16928 ( .A(n15007), .ZN(n15008) );
  NOR2_X2 U16929 ( .A1(n15009), .A2(n10973), .ZN(n15110) );
  AOI22_X1 U16930 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n15109), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15010) );
  NAND4_X1 U16931 ( .A1(n15013), .A2(n15012), .A3(n15011), .A4(n15010), .ZN(
        n15017) );
  INV_X1 U16932 ( .A(n15014), .ZN(n15015) );
  NAND2_X1 U16933 ( .A1(n15015), .A2(n19585), .ZN(n15016) );
  AOI22_X1 U16934 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19232), .B1(
        n19139), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15021) );
  AOI22_X1 U16935 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19115), .B1(
        n19185), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15020) );
  AOI22_X1 U16936 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19265), .B1(
        n15096), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15019) );
  INV_X1 U16937 ( .A(n15103), .ZN(n19248) );
  AOI22_X1 U16938 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19248), .B1(
        n15095), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15018) );
  AND4_X1 U16939 ( .A1(n15021), .A2(n15020), .A3(n15019), .A4(n15018), .ZN(
        n15033) );
  INV_X1 U16940 ( .A(n15110), .ZN(n19170) );
  INV_X1 U16941 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15024) );
  AOI21_X1 U16942 ( .B1(n19204), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n19585), .ZN(n15023) );
  INV_X1 U16943 ( .A(n19154), .ZN(n19150) );
  NAND2_X1 U16944 ( .A1(n19150), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n15022) );
  OAI211_X1 U16945 ( .C1(n19170), .C2(n15024), .A(n15023), .B(n15022), .ZN(
        n15025) );
  INV_X1 U16946 ( .A(n15025), .ZN(n15032) );
  INV_X1 U16947 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19626) );
  NAND2_X1 U16948 ( .A1(n19212), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n15028) );
  INV_X1 U16949 ( .A(n15104), .ZN(n15026) );
  NAND2_X1 U16950 ( .A1(n15026), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n15027) );
  OAI211_X1 U16951 ( .C1(n19308), .C2(n19626), .A(n15028), .B(n15027), .ZN(
        n15029) );
  INV_X1 U16952 ( .A(n15029), .ZN(n15031) );
  AOI22_X1 U16953 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19274), .B1(
        n19196), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15030) );
  NAND4_X1 U16954 ( .A1(n15033), .A2(n15032), .A3(n15031), .A4(n15030), .ZN(
        n15037) );
  OR2_X1 U16955 ( .A1(n15035), .A2(n15034), .ZN(n15036) );
  INV_X1 U16956 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16776) );
  XNOR2_X1 U16957 ( .A(n15044), .B(n16776), .ZN(n16769) );
  NAND2_X1 U16958 ( .A1(n15040), .A2(n15039), .ZN(n15043) );
  INV_X1 U16959 ( .A(n16156), .ZN(n15041) );
  NAND2_X1 U16960 ( .A1(n15041), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15042) );
  NAND2_X1 U16961 ( .A1(n15043), .A2(n15042), .ZN(n16768) );
  NAND2_X1 U16962 ( .A1(n16769), .A2(n16768), .ZN(n15046) );
  NAND2_X1 U16963 ( .A1(n15044), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15045) );
  NAND2_X1 U16964 ( .A1(n15046), .A2(n15045), .ZN(n15128) );
  XNOR2_X1 U16965 ( .A(n15129), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15127) );
  XOR2_X1 U16966 ( .A(n15128), .B(n15127), .Z(n17109) );
  INV_X1 U16967 ( .A(n17109), .ZN(n15068) );
  NOR2_X1 U16968 ( .A1(n15047), .A2(n18593), .ZN(n15048) );
  OR2_X1 U16969 ( .A1(n15049), .A2(n15048), .ZN(n15050) );
  XNOR2_X1 U16970 ( .A(n15050), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16773) );
  NAND2_X1 U16971 ( .A1(n15050), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15051) );
  INV_X1 U16972 ( .A(n15052), .ZN(n15053) );
  NAND2_X1 U16973 ( .A1(n15054), .A2(n15053), .ZN(n15055) );
  NAND2_X1 U16974 ( .A1(n15119), .A2(n15055), .ZN(n15135) );
  XNOR2_X1 U16975 ( .A(n15133), .B(n15502), .ZN(n17107) );
  INV_X1 U16976 ( .A(n18567), .ZN(n18586) );
  NOR2_X1 U16977 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18586), .ZN(
        n15503) );
  INV_X1 U16978 ( .A(n15503), .ZN(n18571) );
  NAND2_X1 U16979 ( .A1(n18573), .A2(n18571), .ZN(n15058) );
  NAND2_X1 U16980 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18586), .ZN(
        n18570) );
  INV_X1 U16981 ( .A(n18570), .ZN(n15056) );
  NAND2_X1 U16982 ( .A1(n18568), .A2(n15056), .ZN(n15057) );
  NAND2_X1 U16983 ( .A1(n15058), .A2(n15057), .ZN(n16775) );
  NAND2_X1 U16984 ( .A1(n16775), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15142) );
  INV_X1 U16985 ( .A(n18566), .ZN(n15060) );
  NAND2_X1 U16986 ( .A1(n18568), .A2(n18570), .ZN(n18585) );
  NAND2_X1 U16987 ( .A1(n18573), .A2(n15503), .ZN(n15059) );
  AND3_X1 U16988 ( .A1(n15060), .A2(n18585), .A3(n15059), .ZN(n16778) );
  OAI21_X1 U16989 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18517), .A(
        n16778), .ZN(n15144) );
  NOR2_X1 U16990 ( .A1(n13663), .A2(n14141), .ZN(n15063) );
  NOR2_X1 U16991 ( .A1(n18579), .A2(n15061), .ZN(n15062) );
  AOI211_X1 U16992 ( .C1(n15144), .C2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n15063), .B(n15062), .ZN(n15065) );
  NAND2_X1 U16993 ( .A1(n17108), .A2(n18584), .ZN(n15064) );
  OAI211_X1 U16994 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n15142), .A(
        n15065), .B(n15064), .ZN(n15066) );
  AOI21_X1 U16995 ( .B1(n17107), .B2(n18556), .A(n15066), .ZN(n15067) );
  OAI21_X1 U16996 ( .B1(n15068), .B2(n16767), .A(n15067), .ZN(P2_U3042) );
  NOR2_X1 U16997 ( .A1(n15490), .A2(n14711), .ZN(n15357) );
  NAND2_X1 U16998 ( .A1(n19381), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15361) );
  NAND2_X1 U16999 ( .A1(n19381), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n15354) );
  INV_X1 U17000 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n16140) );
  NOR2_X1 U17001 ( .A1(n15490), .A2(n16140), .ZN(n15373) );
  NOR2_X1 U17002 ( .A1(n15490), .A2(n16128), .ZN(n15387) );
  NAND2_X1 U17003 ( .A1(n19381), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15069) );
  NOR2_X1 U17004 ( .A1(n15389), .A2(n15069), .ZN(n15070) );
  OR2_X1 U17005 ( .A1(n15392), .A2(n15070), .ZN(n15414) );
  AOI21_X1 U17006 ( .B1(n16452), .B2(n15075), .A(n15076), .ZN(n16122) );
  AOI21_X1 U17007 ( .B1(n18297), .B2(n15073), .A(n11040), .ZN(n16458) );
  AOI21_X1 U17008 ( .B1(n18275), .B2(n15071), .A(n15074), .ZN(n18281) );
  NAND2_X1 U17009 ( .A1(n15072), .A2(n17134), .ZN(n18279) );
  NOR2_X1 U17010 ( .A1(n18281), .A2(n18279), .ZN(n18289) );
  OAI21_X1 U17011 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n15074), .A(
        n15073), .ZN(n18290) );
  NAND2_X1 U17012 ( .A1(n18289), .A2(n18290), .ZN(n18307) );
  NOR2_X1 U17013 ( .A1(n16458), .A2(n18307), .ZN(n16137) );
  OAI21_X1 U17014 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n11040), .A(
        n15075), .ZN(n17145) );
  NAND2_X1 U17015 ( .A1(n16137), .A2(n17145), .ZN(n16121) );
  NOR2_X1 U17016 ( .A1(n16122), .A2(n16121), .ZN(n16123) );
  NAND2_X1 U17017 ( .A1(n18482), .A2(n18423), .ZN(n18505) );
  OAI21_X1 U17018 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n15076), .A(
        n15187), .ZN(n16442) );
  OAI22_X1 U17019 ( .A1(n16123), .A2(n18505), .B1(n16442), .B2(n18602), .ZN(
        n15078) );
  OR3_X1 U17020 ( .A1(n18436), .A2(n16123), .A3(n16442), .ZN(n15077) );
  NAND2_X1 U17021 ( .A1(n15078), .A2(n15077), .ZN(n15087) );
  NOR2_X1 U17022 ( .A1(n15080), .A2(n15079), .ZN(n15081) );
  NOR2_X1 U17023 ( .A1(n16651), .A2(n15081), .ZN(n19082) );
  INV_X1 U17024 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n15083) );
  AOI22_X1 U17025 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18498), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18473), .ZN(n15082) );
  OAI211_X1 U17026 ( .C1(n18490), .C2(n15083), .A(n15082), .B(n14141), .ZN(
        n15085) );
  NOR2_X1 U17027 ( .A1(n16672), .A2(n18478), .ZN(n15084) );
  AOI211_X1 U17028 ( .C1(n18500), .C2(n19082), .A(n15085), .B(n15084), .ZN(
        n15086) );
  OAI211_X1 U17029 ( .C1(n18494), .C2(n15414), .A(n15087), .B(n15086), .ZN(
        P2_U2841) );
  OAI21_X1 U17030 ( .B1(n11053), .B2(n15089), .A(n15088), .ZN(n21336) );
  NAND2_X1 U17031 ( .A1(n21336), .A2(n20020), .ZN(n15093) );
  NOR2_X1 U17032 ( .A1(n21419), .A2(n19855), .ZN(n21332) );
  NOR2_X1 U17033 ( .A1(n20024), .A2(n15090), .ZN(n15091) );
  AOI211_X1 U17034 ( .C1(n20014), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n21332), .B(n15091), .ZN(n15092) );
  OAI211_X1 U17035 ( .C1(n19975), .C2(n15094), .A(n15093), .B(n15092), .ZN(
        P1_U2991) );
  AOI22_X1 U17036 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19204), .B1(
        n19115), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15100) );
  AOI22_X1 U17037 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19232), .B1(
        n19139), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15099) );
  AOI22_X1 U17038 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19265), .B1(
        n19185), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15098) );
  AOI22_X1 U17039 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n15095), .B1(
        n15096), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15097) );
  OAI22_X1 U17040 ( .A1(n15102), .A2(n15328), .B1(n19154), .B2(n15101), .ZN(
        n15108) );
  OAI22_X1 U17041 ( .A1(n15106), .A2(n15103), .B1(n15104), .B2(n15105), .ZN(
        n15107) );
  NOR2_X1 U17042 ( .A1(n15108), .A2(n15107), .ZN(n15113) );
  AOI22_X1 U17043 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n15109), .B1(
        n19274), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15112) );
  AOI22_X1 U17044 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19196), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15111) );
  NAND4_X1 U17045 ( .A1(n15114), .A2(n15113), .A3(n15112), .A4(n15111), .ZN(
        n15117) );
  NAND2_X1 U17046 ( .A1(n19585), .A2(n15115), .ZN(n15116) );
  INV_X1 U17047 ( .A(n15120), .ZN(n15118) );
  NAND2_X1 U17048 ( .A1(n15119), .A2(n15118), .ZN(n15122) );
  INV_X1 U17049 ( .A(n15123), .ZN(n15124) );
  NAND2_X1 U17050 ( .A1(n11038), .A2(n15124), .ZN(n15125) );
  NAND2_X1 U17051 ( .A1(n15126), .A2(n15125), .ZN(n18250) );
  XNOR2_X1 U17052 ( .A(n15318), .B(n15501), .ZN(n15316) );
  NAND2_X1 U17053 ( .A1(n15128), .A2(n15127), .ZN(n15132) );
  INV_X1 U17054 ( .A(n15129), .ZN(n15130) );
  NAND2_X1 U17055 ( .A1(n15130), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15131) );
  NAND2_X1 U17056 ( .A1(n15132), .A2(n15131), .ZN(n15317) );
  XNOR2_X1 U17057 ( .A(n15316), .B(n15317), .ZN(n15159) );
  NAND2_X1 U17058 ( .A1(n15133), .A2(n15502), .ZN(n15138) );
  INV_X1 U17059 ( .A(n15134), .ZN(n15136) );
  NAND2_X1 U17060 ( .A1(n15136), .A2(n15135), .ZN(n15137) );
  OR2_X2 U17061 ( .A1(n15460), .A2(n15139), .ZN(n15469) );
  NAND2_X1 U17062 ( .A1(n15460), .A2(n15139), .ZN(n15140) );
  NAND2_X1 U17063 ( .A1(n15141), .A2(n15501), .ZN(n15153) );
  NAND3_X1 U17064 ( .A1(n15459), .A2(n18556), .A3(n15153), .ZN(n15152) );
  INV_X1 U17065 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n17271) );
  AOI221_X1 U17066 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n15502), .C2(n15501), .A(
        n15142), .ZN(n15143) );
  AOI21_X1 U17067 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n15144), .A(
        n15143), .ZN(n15145) );
  OAI21_X1 U17068 ( .B1(n18521), .B2(n17271), .A(n15145), .ZN(n15150) );
  OAI21_X1 U17069 ( .B1(n15148), .B2(n15147), .A(n15146), .ZN(n19377) );
  NOR2_X1 U17070 ( .A1(n19377), .A2(n18579), .ZN(n15149) );
  AOI211_X1 U17071 ( .C1(n18256), .C2(n18584), .A(n15150), .B(n15149), .ZN(
        n15151) );
  OAI211_X1 U17072 ( .C1(n15159), .C2(n16767), .A(n15152), .B(n15151), .ZN(
        P2_U3041) );
  NAND3_X1 U17073 ( .A1(n15459), .A2(n17203), .A3(n15153), .ZN(n15158) );
  OAI22_X1 U17074 ( .A1(n18249), .A2(n17151), .B1(n17271), .B2(n14141), .ZN(
        n15156) );
  NOR2_X1 U17075 ( .A1(n15154), .A2(n17207), .ZN(n15155) );
  AOI211_X1 U17076 ( .C1(n17163), .C2(n18255), .A(n15156), .B(n15155), .ZN(
        n15157) );
  OAI211_X1 U17077 ( .C1(n15159), .C2(n17156), .A(n15158), .B(n15157), .ZN(
        P2_U3009) );
  NAND2_X1 U17078 ( .A1(n14935), .A2(n15161), .ZN(n15162) );
  NAND2_X1 U17079 ( .A1(n15160), .A2(n15162), .ZN(n15170) );
  XNOR2_X1 U17080 ( .A(n15170), .B(n12013), .ZN(n21512) );
  INV_X1 U17081 ( .A(n15726), .ZN(n19932) );
  XNOR2_X1 U17082 ( .A(n19922), .B(n19921), .ZN(n21509) );
  OAI22_X1 U17083 ( .A1(n21509), .A2(n19942), .B1(n21506), .B2(n19946), .ZN(
        n15163) );
  AOI21_X1 U17084 ( .B1(n21512), .B2(n19932), .A(n15163), .ZN(n15164) );
  INV_X1 U17085 ( .A(n15164), .ZN(P1_U2861) );
  INV_X1 U17086 ( .A(n21512), .ZN(n19974) );
  OR2_X1 U17087 ( .A1(n15727), .A2(BUF1_REG_11__SCAN_IN), .ZN(n15167) );
  INV_X1 U17088 ( .A(DATAI_11_), .ZN(n15165) );
  NAND2_X1 U17089 ( .A1(n15727), .A2(n15165), .ZN(n15166) );
  NAND2_X1 U17090 ( .A1(n15167), .A2(n15166), .ZN(n21752) );
  OAI222_X1 U17091 ( .A1(n19974), .A2(n15801), .B1(n15794), .B2(n15168), .C1(
        n21752), .C2(n15796), .ZN(P1_U2893) );
  OAI21_X1 U17092 ( .B1(n15170), .B2(n15169), .A(n15160), .ZN(n15172) );
  NAND2_X1 U17093 ( .A1(n15172), .A2(n15171), .ZN(n15218) );
  OAI21_X1 U17094 ( .B1(n15172), .B2(n15171), .A(n15218), .ZN(n19919) );
  MUX2_X1 U17095 ( .A(BUF1_REG_12__SCAN_IN), .B(DATAI_12_), .S(n15727), .Z(
        n21757) );
  AOI22_X1 U17096 ( .A1(n15799), .A2(n21757), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15798), .ZN(n15173) );
  OAI21_X1 U17097 ( .B1(n19919), .B2(n15801), .A(n15173), .ZN(P1_U2892) );
  INV_X1 U17098 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16642) );
  NOR2_X1 U17099 ( .A1(n15300), .A2(n15174), .ZN(n15177) );
  INV_X1 U17100 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n15194) );
  INV_X1 U17101 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15175) );
  OAI22_X1 U17102 ( .A1(n15264), .A2(n15194), .B1(n15263), .B2(n15175), .ZN(
        n15176) );
  NOR2_X1 U17103 ( .A1(n15177), .A2(n15176), .ZN(n15178) );
  OAI21_X1 U17104 ( .B1(n15297), .B2(n16642), .A(n15178), .ZN(n15179) );
  OR2_X1 U17105 ( .A1(n15179), .A2(n15180), .ZN(n15181) );
  NAND2_X1 U17106 ( .A1(n15181), .A2(n11042), .ZN(n17155) );
  AOI21_X1 U17107 ( .B1(n15182), .B2(n11037), .A(n15209), .ZN(n19635) );
  NAND2_X1 U17108 ( .A1(n19635), .A2(n16266), .ZN(n15184) );
  NAND2_X1 U17109 ( .A1(n10963), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n15183) );
  OAI211_X1 U17110 ( .C1(n17155), .C2(n10963), .A(n15184), .B(n15183), .ZN(
        P2_U2871) );
  NAND2_X1 U17111 ( .A1(n19381), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n15391) );
  NOR2_X1 U17112 ( .A1(n15490), .A2(n15194), .ZN(n15185) );
  NAND2_X1 U17113 ( .A1(n15394), .A2(n15185), .ZN(n15186) );
  NAND2_X1 U17114 ( .A1(n11009), .A2(n15186), .ZN(n15382) );
  AOI21_X1 U17115 ( .B1(n18330), .B2(n15187), .A(n15188), .ZN(n18322) );
  NAND2_X1 U17116 ( .A1(n16123), .A2(n16442), .ZN(n18319) );
  NOR2_X1 U17117 ( .A1(n18322), .A2(n18319), .ZN(n18323) );
  NOR2_X1 U17118 ( .A1(n18436), .A2(n18323), .ZN(n15189) );
  OAI21_X1 U17119 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n15188), .A(
        n16093), .ZN(n17162) );
  XNOR2_X1 U17120 ( .A(n15189), .B(n17162), .ZN(n15190) );
  NAND2_X1 U17121 ( .A1(n15190), .A2(n18482), .ZN(n15198) );
  AOI21_X1 U17122 ( .B1(n15192), .B2(n16652), .A(n15191), .ZN(n19632) );
  AOI22_X1 U17123 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18498), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n18473), .ZN(n15193) );
  OAI211_X1 U17124 ( .C1(n18490), .C2(n15194), .A(n15193), .B(n14141), .ZN(
        n15196) );
  NOR2_X1 U17125 ( .A1(n18478), .A2(n17155), .ZN(n15195) );
  AOI211_X1 U17126 ( .C1(n18500), .C2(n19632), .A(n15196), .B(n15195), .ZN(
        n15197) );
  OAI211_X1 U17127 ( .C1(n18494), .C2(n15382), .A(n15198), .B(n15197), .ZN(
        P2_U2839) );
  OAI21_X1 U17128 ( .B1(n15199), .B2(n15201), .A(n15233), .ZN(n19988) );
  AOI22_X1 U17129 ( .A1(n15799), .A2(n21770), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15798), .ZN(n15202) );
  OAI21_X1 U17130 ( .B1(n19988), .B2(n15801), .A(n15202), .ZN(P1_U2890) );
  INV_X1 U17131 ( .A(n15203), .ZN(n15205) );
  INV_X1 U17132 ( .A(n15220), .ZN(n15204) );
  AOI21_X1 U17133 ( .B1(n15205), .B2(n15204), .A(n15238), .ZN(n21526) );
  AOI22_X1 U17134 ( .A1(n21526), .A2(n19925), .B1(n15724), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n15206) );
  OAI21_X1 U17135 ( .B1(n19988), .B2(n15726), .A(n15206), .ZN(P1_U2858) );
  OAI21_X1 U17136 ( .B1(n15209), .B2(n15208), .A(n16264), .ZN(n16340) );
  NAND2_X1 U17137 ( .A1(n10963), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15215) );
  INV_X1 U17138 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n18335) );
  OAI22_X1 U17139 ( .A1(n15264), .A2(n18335), .B1(n15263), .B2(n16094), .ZN(
        n15212) );
  INV_X1 U17140 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15210) );
  NOR2_X1 U17141 ( .A1(n15297), .A2(n15210), .ZN(n15211) );
  AOI211_X1 U17142 ( .C1(n15294), .C2(P2_REIP_REG_17__SCAN_IN), .A(n15212), 
        .B(n15211), .ZN(n15213) );
  AOI21_X1 U17143 ( .B1(n15213), .B2(n11042), .A(n16260), .ZN(n18339) );
  NAND2_X1 U17144 ( .A1(n18339), .A2(n11059), .ZN(n15214) );
  OAI211_X1 U17145 ( .C1(n16340), .C2(n16253), .A(n15215), .B(n15214), .ZN(
        P2_U2870) );
  INV_X1 U17146 ( .A(n15216), .ZN(n15217) );
  AOI21_X1 U17147 ( .B1(n15218), .B2(n15217), .A(n15199), .ZN(n15919) );
  AND2_X1 U17148 ( .A1(n19923), .A2(n15219), .ZN(n15221) );
  OR2_X1 U17149 ( .A1(n15221), .A2(n15220), .ZN(n16068) );
  OAI22_X1 U17150 ( .A1(n16068), .A2(n19942), .B1(n15656), .B2(n19946), .ZN(
        n15222) );
  AOI21_X1 U17151 ( .B1(n15919), .B2(n19932), .A(n15222), .ZN(n15223) );
  INV_X1 U17152 ( .A(n15223), .ZN(P1_U2859) );
  INV_X1 U17153 ( .A(n15921), .ZN(n15923) );
  AOI21_X1 U17154 ( .B1(n15225), .B2(n15224), .A(n15923), .ZN(n21350) );
  NAND2_X1 U17155 ( .A1(n21350), .A2(n20020), .ZN(n15230) );
  NAND2_X1 U17156 ( .A1(n14073), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n21343) );
  OAI21_X1 U17157 ( .B1(n15898), .B2(n15226), .A(n21343), .ZN(n15227) );
  AOI21_X1 U17158 ( .B1(n19989), .B2(n15228), .A(n15227), .ZN(n15229) );
  OAI211_X1 U17159 ( .C1(n19975), .C2(n15231), .A(n15230), .B(n15229), .ZN(
        P1_U2990) );
  AOI21_X1 U17160 ( .B1(n15234), .B2(n15233), .A(n11353), .ZN(n15907) );
  INV_X1 U17161 ( .A(n15907), .ZN(n15797) );
  OAI21_X1 U17162 ( .B1(n21601), .B2(n19866), .A(n15235), .ZN(n15245) );
  INV_X1 U17163 ( .A(n15236), .ZN(n15244) );
  OR2_X1 U17164 ( .A1(n15238), .A2(n15237), .ZN(n15239) );
  NAND2_X1 U17165 ( .A1(n15644), .A2(n15239), .ZN(n16056) );
  INV_X1 U17166 ( .A(n15905), .ZN(n15240) );
  AOI22_X1 U17167 ( .A1(n21615), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n21634), .B2(n15240), .ZN(n15242) );
  AOI21_X1 U17168 ( .B1(n21597), .B2(P1_EBX_REG_15__SCAN_IN), .A(n21557), .ZN(
        n15241) );
  OAI211_X1 U17169 ( .C1(n16056), .C2(n21638), .A(n15242), .B(n15241), .ZN(
        n15243) );
  AOI21_X1 U17170 ( .B1(n15245), .B2(n15244), .A(n15243), .ZN(n15246) );
  OAI21_X1 U17171 ( .B1(n15797), .B2(n21630), .A(n15246), .ZN(P1_U2825) );
  INV_X1 U17172 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15247) );
  OAI22_X1 U17173 ( .A1(n16056), .A2(n19942), .B1(n15247), .B2(n19946), .ZN(
        n15248) );
  AOI21_X1 U17174 ( .B1(n15907), .B2(n19932), .A(n15248), .ZN(n15249) );
  INV_X1 U17175 ( .A(n15249), .ZN(P1_U2857) );
  INV_X1 U17176 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15407) );
  INV_X1 U17177 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15252) );
  NAND2_X1 U17178 ( .A1(n15285), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15251) );
  NAND2_X1 U17179 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15250) );
  OAI211_X1 U17180 ( .C1(n15300), .C2(n15252), .A(n15251), .B(n15250), .ZN(
        n15253) );
  INV_X1 U17181 ( .A(n15253), .ZN(n15254) );
  OAI21_X1 U17182 ( .B1(n15297), .B2(n15407), .A(n15254), .ZN(n16261) );
  NAND2_X1 U17183 ( .A1(n15556), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15256) );
  NAND2_X1 U17184 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15255) );
  OAI211_X1 U17185 ( .C1(n15300), .C2(n17276), .A(n15256), .B(n15255), .ZN(
        n15257) );
  AOI21_X1 U17186 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15257), .ZN(n16254) );
  INV_X1 U17187 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18538) );
  NAND2_X1 U17188 ( .A1(n15556), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15259) );
  NAND2_X1 U17189 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15258) );
  OAI211_X1 U17190 ( .C1(n15300), .C2(n15260), .A(n15259), .B(n15258), .ZN(
        n15261) );
  INV_X1 U17191 ( .A(n15261), .ZN(n15262) );
  OAI21_X1 U17192 ( .B1(n15297), .B2(n18538), .A(n15262), .ZN(n16248) );
  NAND2_X1 U17193 ( .A1(n16247), .A2(n16248), .ZN(n16249) );
  INV_X1 U17194 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n18381) );
  OAI22_X1 U17195 ( .A1(n15264), .A2(n18381), .B1(n15263), .B2(n16413), .ZN(
        n15266) );
  INV_X1 U17196 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16588) );
  NOR2_X1 U17197 ( .A1(n15297), .A2(n16588), .ZN(n15265) );
  AOI211_X1 U17198 ( .C1(n15294), .C2(P2_REIP_REG_21__SCAN_IN), .A(n15266), 
        .B(n15265), .ZN(n16240) );
  INV_X1 U17199 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15425) );
  INV_X1 U17200 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n15269) );
  NAND2_X1 U17201 ( .A1(n15285), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15268) );
  NAND2_X1 U17202 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15267) );
  OAI211_X1 U17203 ( .C1(n15300), .C2(n15269), .A(n15268), .B(n15267), .ZN(
        n15270) );
  INV_X1 U17204 ( .A(n15270), .ZN(n15271) );
  OAI21_X1 U17205 ( .B1(n15297), .B2(n15425), .A(n15271), .ZN(n16231) );
  NAND2_X1 U17206 ( .A1(n15556), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15273) );
  NAND2_X1 U17207 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15272) );
  OAI211_X1 U17208 ( .C1(n15300), .C2(n17278), .A(n15273), .B(n15272), .ZN(
        n15274) );
  AOI21_X1 U17209 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15274), .ZN(n16225) );
  NAND2_X1 U17210 ( .A1(n15285), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15276) );
  NAND2_X1 U17211 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15275) );
  OAI211_X1 U17212 ( .C1(n15300), .C2(n15277), .A(n15276), .B(n15275), .ZN(
        n15278) );
  AOI21_X1 U17213 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15278), .ZN(n16217) );
  INV_X1 U17214 ( .A(n16217), .ZN(n15279) );
  NAND2_X1 U17215 ( .A1(n15285), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15281) );
  NAND2_X1 U17216 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15280) );
  OAI211_X1 U17217 ( .C1(n15300), .C2(n17279), .A(n15281), .B(n15280), .ZN(
        n15282) );
  AOI21_X1 U17218 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15282), .ZN(n16210) );
  INV_X1 U17219 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16525) );
  AOI22_X1 U17220 ( .A1(n15556), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n15284) );
  NAND2_X1 U17221 ( .A1(n15294), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15283) );
  OAI211_X1 U17222 ( .C1(n15297), .C2(n16525), .A(n15284), .B(n15283), .ZN(
        n16199) );
  NAND2_X1 U17223 ( .A1(n15285), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15287) );
  NAND2_X1 U17224 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15286) );
  OAI211_X1 U17225 ( .C1(n15300), .C2(n18448), .A(n15287), .B(n15286), .ZN(
        n15288) );
  AOI21_X1 U17226 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15288), .ZN(n16193) );
  NAND2_X1 U17227 ( .A1(n15556), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15290) );
  NAND2_X1 U17228 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15289) );
  OAI211_X1 U17229 ( .C1(n15300), .C2(n15291), .A(n15290), .B(n15289), .ZN(
        n15292) );
  AOI21_X1 U17230 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15292), .ZN(n16180) );
  INV_X1 U17231 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16491) );
  AOI22_X1 U17232 ( .A1(n15556), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n15296) );
  NAND2_X1 U17233 ( .A1(n15294), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15295) );
  OAI211_X1 U17234 ( .C1(n15297), .C2(n16491), .A(n15296), .B(n15295), .ZN(
        n15455) );
  NAND2_X1 U17235 ( .A1(n15293), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15299) );
  AOI22_X1 U17236 ( .A1(n15556), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n15298) );
  OAI211_X1 U17237 ( .C1(n15300), .C2(n17283), .A(n15299), .B(n15298), .ZN(
        n15554) );
  NOR2_X1 U17238 ( .A1(n16110), .A2(n10963), .ZN(n15301) );
  AOI21_X1 U17239 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n10963), .A(n15301), .ZN(
        n15302) );
  OAI21_X1 U17240 ( .B1(n15303), .B2(n16253), .A(n15302), .ZN(P2_U2857) );
  NOR2_X1 U17241 ( .A1(n15490), .A2(n18335), .ZN(n15383) );
  INV_X1 U17242 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n18347) );
  NAND2_X1 U17243 ( .A1(n19381), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15379) );
  NAND2_X1 U17244 ( .A1(n19381), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15396) );
  INV_X1 U17245 ( .A(n15396), .ZN(n15304) );
  NAND2_X1 U17246 ( .A1(n19381), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15399) );
  NAND2_X1 U17247 ( .A1(n19381), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15423) );
  INV_X1 U17248 ( .A(n15423), .ZN(n15305) );
  NAND2_X1 U17249 ( .A1(n19381), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15428) );
  NAND2_X1 U17250 ( .A1(n19381), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15432) );
  INV_X1 U17251 ( .A(n15432), .ZN(n15306) );
  NAND2_X1 U17252 ( .A1(n19381), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15436) );
  INV_X1 U17253 ( .A(n15440), .ZN(n15308) );
  NAND2_X1 U17254 ( .A1(n19381), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15439) );
  NAND2_X1 U17255 ( .A1(n19381), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15312) );
  NAND2_X1 U17256 ( .A1(n19381), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15445) );
  INV_X1 U17257 ( .A(n15445), .ZN(n15309) );
  NAND2_X1 U17258 ( .A1(n19381), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15489) );
  XNOR2_X1 U17259 ( .A(n15488), .B(n15489), .ZN(n15310) );
  INV_X1 U17260 ( .A(n15310), .ZN(n18472) );
  AOI21_X1 U17261 ( .B1(n18472), .B2(n11050), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15486) );
  NOR2_X1 U17262 ( .A1(n15486), .A2(n15534), .ZN(n15451) );
  INV_X1 U17263 ( .A(n15311), .ZN(n15314) );
  INV_X1 U17264 ( .A(n15312), .ZN(n15313) );
  NAND2_X1 U17265 ( .A1(n15314), .A2(n15313), .ZN(n15315) );
  NAND2_X1 U17266 ( .A1(n15444), .A2(n15315), .ZN(n18449) );
  NAND2_X1 U17267 ( .A1(n15317), .A2(n15316), .ZN(n15320) );
  NAND2_X1 U17268 ( .A1(n15318), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15319) );
  NAND2_X1 U17269 ( .A1(n15320), .A2(n15319), .ZN(n16752) );
  AOI22_X1 U17270 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19204), .B1(
        n19115), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15324) );
  AOI22_X1 U17271 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19232), .B1(
        n19139), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n15323) );
  AOI22_X1 U17272 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19185), .B1(
        n15096), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15322) );
  AOI22_X1 U17273 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n15095), .B1(
        n19265), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15321) );
  INV_X1 U17274 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n15326) );
  OAI22_X1 U17275 ( .A1(n15326), .A2(n15103), .B1(n19154), .B2(n15325), .ZN(
        n15331) );
  INV_X1 U17276 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15329) );
  OAI22_X1 U17277 ( .A1(n15329), .A2(n15328), .B1(n15104), .B2(n15327), .ZN(
        n15330) );
  NOR2_X1 U17278 ( .A1(n15331), .A2(n15330), .ZN(n15334) );
  AOI22_X1 U17279 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19274), .B1(
        n15110), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15333) );
  AOI22_X1 U17280 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n15109), .B1(
        n19196), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15332) );
  NAND4_X1 U17281 ( .A1(n15335), .A2(n15334), .A3(n15333), .A4(n15332), .ZN(
        n15338) );
  NAND2_X1 U17282 ( .A1(n19585), .A2(n15336), .ZN(n15337) );
  NAND2_X1 U17283 ( .A1(n15458), .A2(n10966), .ZN(n15340) );
  NAND2_X1 U17284 ( .A1(n15340), .A2(n15339), .ZN(n15341) );
  INV_X1 U17285 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16757) );
  XNOR2_X1 U17286 ( .A(n15341), .B(n16757), .ZN(n16753) );
  NAND2_X1 U17287 ( .A1(n15341), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15342) );
  NOR2_X1 U17288 ( .A1(n15343), .A2(n10966), .ZN(n15347) );
  NAND2_X1 U17289 ( .A1(n15347), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17122) );
  INV_X1 U17290 ( .A(n15344), .ZN(n15346) );
  XNOR2_X1 U17291 ( .A(n15346), .B(n15345), .ZN(n18267) );
  NAND2_X1 U17292 ( .A1(n18267), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17123) );
  NAND2_X1 U17293 ( .A1(n17122), .A2(n17123), .ZN(n15352) );
  INV_X1 U17294 ( .A(n15347), .ZN(n15349) );
  NAND2_X1 U17295 ( .A1(n15349), .A2(n15348), .ZN(n17121) );
  INV_X1 U17296 ( .A(n18267), .ZN(n15350) );
  NAND2_X1 U17297 ( .A1(n15350), .A2(n16745), .ZN(n17125) );
  AND2_X1 U17298 ( .A1(n17121), .A2(n17125), .ZN(n15351) );
  INV_X1 U17299 ( .A(n15353), .ZN(n15365) );
  XNOR2_X1 U17300 ( .A(n15365), .B(n15354), .ZN(n18296) );
  NAND2_X1 U17301 ( .A1(n18296), .A2(n11050), .ZN(n15355) );
  INV_X1 U17302 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15369) );
  NAND2_X1 U17303 ( .A1(n15355), .A2(n15369), .ZN(n16463) );
  INV_X1 U17304 ( .A(n15356), .ZN(n15363) );
  NAND2_X1 U17305 ( .A1(n15358), .A2(n15357), .ZN(n15359) );
  NAND2_X1 U17306 ( .A1(n15363), .A2(n15359), .ZN(n18276) );
  NOR2_X1 U17307 ( .A1(n18276), .A2(n10966), .ZN(n15366) );
  INV_X1 U17308 ( .A(n15366), .ZN(n15360) );
  INV_X1 U17309 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16730) );
  NAND2_X1 U17310 ( .A1(n15360), .A2(n16730), .ZN(n16470) );
  INV_X1 U17311 ( .A(n15361), .ZN(n15362) );
  NAND2_X1 U17312 ( .A1(n15363), .A2(n15362), .ZN(n15364) );
  AND2_X1 U17313 ( .A1(n15365), .A2(n15364), .ZN(n15368) );
  INV_X1 U17314 ( .A(n15368), .ZN(n18287) );
  OAI21_X1 U17315 ( .B1(n18287), .B2(n10966), .A(n16705), .ZN(n16714) );
  NAND3_X1 U17316 ( .A1(n16463), .A2(n16470), .A3(n16714), .ZN(n15372) );
  NAND2_X1 U17317 ( .A1(n15366), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16711) );
  NOR2_X1 U17318 ( .A1(n10966), .A2(n16705), .ZN(n15367) );
  NAND2_X1 U17319 ( .A1(n15368), .A2(n15367), .ZN(n16713) );
  NAND2_X1 U17320 ( .A1(n16711), .A2(n16713), .ZN(n16461) );
  NOR2_X1 U17321 ( .A1(n10966), .A2(n15369), .ZN(n15370) );
  AND2_X1 U17322 ( .A1(n18296), .A2(n15370), .ZN(n16464) );
  NOR2_X1 U17323 ( .A1(n16461), .A2(n16464), .ZN(n15371) );
  NAND2_X1 U17324 ( .A1(n15374), .A2(n15373), .ZN(n15375) );
  NAND2_X1 U17325 ( .A1(n15388), .A2(n15375), .ZN(n16144) );
  OR2_X1 U17326 ( .A1(n10966), .A2(n18530), .ZN(n15376) );
  OAI21_X1 U17327 ( .B1(n16144), .B2(n10966), .A(n18530), .ZN(n17139) );
  AND2_X1 U17328 ( .A1(n15385), .A2(n15377), .ZN(n15378) );
  NOR2_X1 U17329 ( .A1(n15380), .A2(n15378), .ZN(n18349) );
  NAND2_X1 U17330 ( .A1(n18349), .A2(n11050), .ZN(n15408) );
  NAND2_X1 U17331 ( .A1(n15408), .A2(n15407), .ZN(n17174) );
  INV_X1 U17332 ( .A(n17174), .ZN(n16421) );
  OR2_X1 U17333 ( .A1(n15380), .A2(n15379), .ZN(n15381) );
  AND2_X1 U17334 ( .A1(n15381), .A2(n15397), .ZN(n18361) );
  AOI21_X1 U17335 ( .B1(n18361), .B2(n11050), .A(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16420) );
  NOR2_X1 U17336 ( .A1(n16421), .A2(n16420), .ZN(n16404) );
  XNOR2_X1 U17337 ( .A(n15410), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16633) );
  NAND2_X1 U17338 ( .A1(n11009), .A2(n15383), .ZN(n15384) );
  AND2_X1 U17339 ( .A1(n15385), .A2(n15384), .ZN(n18337) );
  NAND2_X1 U17340 ( .A1(n18337), .A2(n11050), .ZN(n15386) );
  NAND2_X1 U17341 ( .A1(n15386), .A2(n15210), .ZN(n16613) );
  INV_X1 U17342 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16667) );
  OAI21_X1 U17343 ( .B1(n15414), .B2(n10966), .A(n16667), .ZN(n16645) );
  AND2_X1 U17344 ( .A1(n15388), .A2(n15387), .ZN(n15390) );
  OR2_X1 U17345 ( .A1(n15390), .A2(n15389), .ZN(n16135) );
  NOR2_X1 U17346 ( .A1(n16135), .A2(n10966), .ZN(n15417) );
  OR2_X1 U17347 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15417), .ZN(
        n16435) );
  OR2_X1 U17348 ( .A1(n15392), .A2(n15391), .ZN(n15393) );
  NAND2_X1 U17349 ( .A1(n15394), .A2(n15393), .ZN(n18314) );
  NOR2_X1 U17350 ( .A1(n18314), .A2(n10966), .ZN(n15413) );
  OR2_X1 U17351 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15413), .ZN(
        n16647) );
  AND2_X1 U17352 ( .A1(n16435), .A2(n16647), .ZN(n15395) );
  AND2_X1 U17353 ( .A1(n16645), .A2(n15395), .ZN(n16399) );
  AND3_X1 U17354 ( .A1(n16633), .A2(n16613), .A3(n16399), .ZN(n15405) );
  XNOR2_X1 U17355 ( .A(n15397), .B(n15396), .ZN(n18372) );
  NAND2_X1 U17356 ( .A1(n18372), .A2(n11050), .ZN(n16407) );
  NAND2_X1 U17357 ( .A1(n16407), .A2(n18538), .ZN(n15404) );
  INV_X1 U17358 ( .A(n15398), .ZN(n15401) );
  INV_X1 U17359 ( .A(n15399), .ZN(n15400) );
  NAND2_X1 U17360 ( .A1(n15401), .A2(n15400), .ZN(n15402) );
  NAND2_X1 U17361 ( .A1(n15424), .A2(n15402), .ZN(n18382) );
  OR2_X1 U17362 ( .A1(n18382), .A2(n10966), .ZN(n15403) );
  NAND2_X1 U17363 ( .A1(n15403), .A2(n16588), .ZN(n16409) );
  INV_X1 U17364 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18539) );
  NOR2_X1 U17365 ( .A1(n10966), .A2(n18539), .ZN(n15406) );
  AND2_X1 U17366 ( .A1(n18361), .A2(n15406), .ZN(n16419) );
  INV_X1 U17367 ( .A(n16419), .ZN(n15409) );
  OR2_X1 U17368 ( .A1(n15408), .A2(n15407), .ZN(n17175) );
  NAND2_X1 U17369 ( .A1(n15409), .A2(n17175), .ZN(n16405) );
  INV_X1 U17370 ( .A(n16405), .ZN(n15420) );
  INV_X1 U17371 ( .A(n15410), .ZN(n15411) );
  NAND2_X1 U17372 ( .A1(n15411), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16611) );
  NOR2_X1 U17373 ( .A1(n10966), .A2(n15210), .ZN(n15412) );
  NAND2_X1 U17374 ( .A1(n18337), .A2(n15412), .ZN(n16612) );
  NAND2_X1 U17375 ( .A1(n15413), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16646) );
  INV_X1 U17376 ( .A(n15414), .ZN(n15416) );
  NOR2_X1 U17377 ( .A1(n10966), .A2(n16667), .ZN(n15415) );
  NAND2_X1 U17378 ( .A1(n15416), .A2(n15415), .ZN(n16436) );
  NAND2_X1 U17379 ( .A1(n15417), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16434) );
  AND2_X1 U17380 ( .A1(n16436), .A2(n16434), .ZN(n15418) );
  AND2_X1 U17381 ( .A1(n16646), .A2(n15418), .ZN(n16400) );
  OR2_X1 U17382 ( .A1(n10966), .A2(n16588), .ZN(n15419) );
  OR2_X1 U17383 ( .A1(n18382), .A2(n15419), .ZN(n16410) );
  AND4_X1 U17384 ( .A1(n15420), .A2(n16403), .A3(n16400), .A4(n16410), .ZN(
        n15422) );
  OR2_X1 U17385 ( .A1(n16407), .A2(n18538), .ZN(n15421) );
  XNOR2_X1 U17386 ( .A(n15424), .B(n15423), .ZN(n18392) );
  NAND2_X1 U17387 ( .A1(n18392), .A2(n11050), .ZN(n15426) );
  NOR2_X1 U17388 ( .A1(n15426), .A2(n15425), .ZN(n16570) );
  NAND2_X1 U17389 ( .A1(n15426), .A2(n15425), .ZN(n16568) );
  INV_X1 U17390 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16557) );
  INV_X1 U17391 ( .A(n15427), .ZN(n15429) );
  XNOR2_X1 U17392 ( .A(n15429), .B(n15428), .ZN(n18401) );
  NAND2_X1 U17393 ( .A1(n18401), .A2(n11050), .ZN(n16394) );
  OAI21_X1 U17394 ( .B1(n16396), .B2(n16557), .A(n16394), .ZN(n15431) );
  NAND2_X1 U17395 ( .A1(n16396), .A2(n16557), .ZN(n15430) );
  NAND2_X1 U17396 ( .A1(n15431), .A2(n15430), .ZN(n16548) );
  XNOR2_X1 U17397 ( .A(n15433), .B(n15432), .ZN(n18412) );
  NAND2_X1 U17398 ( .A1(n18412), .A2(n11050), .ZN(n15434) );
  XNOR2_X1 U17399 ( .A(n15434), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16547) );
  INV_X1 U17400 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16550) );
  NAND2_X1 U17401 ( .A1(n15434), .A2(n16550), .ZN(n15435) );
  XNOR2_X1 U17402 ( .A(n15437), .B(n15436), .ZN(n18432) );
  AOI21_X1 U17403 ( .B1(n18432), .B2(n11050), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16383) );
  INV_X1 U17404 ( .A(n16383), .ZN(n15438) );
  XNOR2_X1 U17405 ( .A(n15440), .B(n15439), .ZN(n18444) );
  NAND2_X1 U17406 ( .A1(n18444), .A2(n11050), .ZN(n15441) );
  NAND2_X1 U17407 ( .A1(n15441), .A2(n16525), .ZN(n15443) );
  NOR2_X1 U17408 ( .A1(n10966), .A2(n16525), .ZN(n15442) );
  NAND2_X1 U17409 ( .A1(n18444), .A2(n15442), .ZN(n15450) );
  NAND2_X1 U17410 ( .A1(n15443), .A2(n15450), .ZN(n16370) );
  OAI21_X1 U17411 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16349), .A(
        n16368), .ZN(n15447) );
  XOR2_X1 U17412 ( .A(n15445), .B(n15444), .Z(n18459) );
  OAI21_X1 U17413 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n16351), .ZN(n15446) );
  INV_X1 U17414 ( .A(n16351), .ZN(n15448) );
  INV_X1 U17415 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16508) );
  INV_X1 U17416 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16538) );
  NOR2_X1 U17417 ( .A1(n10966), .A2(n16538), .ZN(n15449) );
  NAND2_X1 U17418 ( .A1(n18432), .A2(n15449), .ZN(n16381) );
  NAND2_X1 U17419 ( .A1(n15450), .A2(n16381), .ZN(n16348) );
  XOR2_X1 U17420 ( .A(n15451), .B(n15487), .Z(n16502) );
  INV_X1 U17421 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15454) );
  INV_X1 U17422 ( .A(n15452), .ZN(n16105) );
  INV_X1 U17423 ( .A(n15496), .ZN(n15453) );
  AOI21_X1 U17424 ( .B1(n15454), .B2(n16105), .A(n15453), .ZN(n16107) );
  NOR2_X1 U17425 ( .A1(n11007), .A2(n15455), .ZN(n15456) );
  NOR2_X1 U17426 ( .A1(n18521), .A2(n17282), .ZN(n16496) );
  AOI21_X1 U17427 ( .B1(n17200), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16496), .ZN(n15457) );
  OAI21_X1 U17428 ( .B1(n18479), .B2(n17207), .A(n15457), .ZN(n15484) );
  INV_X1 U17429 ( .A(n15460), .ZN(n15468) );
  INV_X1 U17430 ( .A(n15139), .ZN(n15461) );
  OAI21_X1 U17431 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n15461), .A(
        n11129), .ZN(n15465) );
  INV_X1 U17432 ( .A(n15473), .ZN(n15462) );
  MUX2_X1 U17433 ( .A(n15462), .B(n15501), .S(n15139), .Z(n15463) );
  OAI21_X1 U17434 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n15458), .A(
        n15463), .ZN(n15464) );
  NAND2_X1 U17435 ( .A1(n15459), .A2(n15469), .ZN(n15470) );
  NAND2_X1 U17436 ( .A1(n15470), .A2(n15458), .ZN(n15471) );
  XNOR2_X1 U17437 ( .A(n15475), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16482) );
  INV_X1 U17438 ( .A(n15475), .ZN(n15476) );
  NAND2_X1 U17439 ( .A1(n15476), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15477) );
  NAND2_X1 U17440 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16623) );
  NAND2_X1 U17441 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16432) );
  NAND3_X1 U17442 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18520) );
  NOR2_X1 U17443 ( .A1(n16432), .A2(n18520), .ZN(n16668) );
  NAND2_X1 U17444 ( .A1(n16668), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16654) );
  INV_X1 U17445 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16661) );
  OR2_X1 U17446 ( .A1(n16654), .A2(n16661), .ZN(n16624) );
  NOR2_X1 U17447 ( .A1(n16623), .A2(n16624), .ZN(n17165) );
  NAND2_X1 U17448 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17165), .ZN(
        n16602) );
  INV_X1 U17449 ( .A(n16602), .ZN(n16598) );
  AND3_X1 U17450 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n16598), .ZN(n16587) );
  NAND2_X1 U17451 ( .A1(n16587), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15511) );
  INV_X1 U17452 ( .A(n15511), .ZN(n15481) );
  AND2_X1 U17453 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15512) );
  AND2_X1 U17454 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15515) );
  INV_X1 U17455 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16493) );
  INV_X1 U17456 ( .A(n16354), .ZN(n16521) );
  NOR2_X1 U17457 ( .A1(n16521), .A2(n16508), .ZN(n15482) );
  NAND3_X1 U17458 ( .A1(n16354), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15495) );
  OAI21_X1 U17459 ( .B1(n15482), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15495), .ZN(n16490) );
  NOR2_X1 U17460 ( .A1(n16490), .A2(n17152), .ZN(n15483) );
  OAI21_X1 U17461 ( .B1(n16502), .B2(n17156), .A(n15485), .ZN(P2_U2985) );
  INV_X1 U17462 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n16112) );
  INV_X1 U17463 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15517) );
  AOI21_X1 U17464 ( .B1(n15491), .B2(n11050), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15542) );
  XNOR2_X1 U17465 ( .A(n15492), .B(n11391), .ZN(n15530) );
  AND2_X1 U17466 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15518) );
  AND2_X1 U17467 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15494) );
  NAND2_X1 U17468 ( .A1(n15518), .A2(n15494), .ZN(n15549) );
  NOR2_X2 U17469 ( .A1(n15493), .A2(n15549), .ZN(n15548) );
  AOI21_X1 U17470 ( .B1(n15495), .B2(n15517), .A(n15548), .ZN(n15528) );
  XOR2_X1 U17471 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n15496), .Z(
        n16108) );
  NOR2_X1 U17472 ( .A1(n18521), .A2(n17283), .ZN(n15520) );
  NOR2_X1 U17473 ( .A1(n16110), .A2(n17207), .ZN(n15497) );
  OAI21_X1 U17474 ( .B1(n16108), .B2(n17198), .A(n15498), .ZN(n15499) );
  AOI21_X1 U17475 ( .B1(n15528), .B2(n17203), .A(n15499), .ZN(n15500) );
  OAI21_X1 U17476 ( .B1(n15530), .B2(n17156), .A(n15500), .ZN(P2_U2984) );
  NAND2_X1 U17477 ( .A1(n16113), .A2(n18553), .ZN(n15526) );
  NOR2_X1 U17478 ( .A1(n16110), .A2(n18512), .ZN(n15524) );
  OR2_X1 U17479 ( .A1(n18517), .A2(n15515), .ZN(n15513) );
  NOR3_X1 U17480 ( .A1(n16776), .A2(n15502), .A3(n15501), .ZN(n16744) );
  NAND2_X1 U17481 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16744), .ZN(
        n15504) );
  NAND2_X1 U17482 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18560) );
  NOR3_X1 U17483 ( .A1(n15503), .A2(n15504), .A3(n18560), .ZN(n15507) );
  NAND2_X1 U17484 ( .A1(n18573), .A2(n15507), .ZN(n15506) );
  OR2_X1 U17485 ( .A1(n15504), .A2(n18570), .ZN(n16742) );
  NOR2_X1 U17486 ( .A1(n18560), .A2(n16742), .ZN(n16597) );
  NAND2_X1 U17487 ( .A1(n18568), .A2(n16597), .ZN(n15505) );
  NAND2_X1 U17488 ( .A1(n15506), .A2(n15505), .ZN(n16728) );
  NOR3_X1 U17489 ( .A1(n15425), .A2(n16557), .A3(n16575), .ZN(n15514) );
  AND2_X1 U17490 ( .A1(n16550), .A2(n15514), .ZN(n16552) );
  INV_X1 U17491 ( .A(n15507), .ZN(n15508) );
  AOI21_X1 U17492 ( .B1(n18573), .B2(n15508), .A(n18566), .ZN(n16600) );
  INV_X1 U17493 ( .A(n16600), .ZN(n15510) );
  INV_X1 U17494 ( .A(n16597), .ZN(n15509) );
  AND2_X1 U17495 ( .A1(n18568), .A2(n15509), .ZN(n16616) );
  NOR2_X1 U17496 ( .A1(n15510), .A2(n16616), .ZN(n16731) );
  INV_X1 U17497 ( .A(n16731), .ZN(n18518) );
  AOI21_X1 U17498 ( .B1(n15511), .B2(n18519), .A(n18518), .ZN(n16574) );
  OAI21_X1 U17499 ( .B1(n15512), .B2(n16575), .A(n16574), .ZN(n16562) );
  NOR2_X1 U17500 ( .A1(n16552), .A2(n16562), .ZN(n16537) );
  NAND2_X1 U17501 ( .A1(n15513), .A2(n16537), .ZN(n16519) );
  AOI21_X1 U17502 ( .B1(n15549), .B2(n18519), .A(n16519), .ZN(n15562) );
  OR2_X1 U17503 ( .A1(n15562), .A2(n15517), .ZN(n15522) );
  NAND2_X1 U17504 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15514), .ZN(
        n16536) );
  INV_X1 U17505 ( .A(n16536), .ZN(n15516) );
  NAND2_X1 U17506 ( .A1(n15516), .A2(n15515), .ZN(n16492) );
  INV_X1 U17507 ( .A(n16492), .ZN(n15519) );
  NOR2_X1 U17508 ( .A1(n11397), .A2(n15520), .ZN(n15521) );
  NAND2_X1 U17509 ( .A1(n15522), .A2(n15521), .ZN(n15523) );
  NAND2_X1 U17510 ( .A1(n15526), .A2(n15525), .ZN(n15527) );
  AOI21_X1 U17511 ( .B1(n15528), .B2(n18556), .A(n15527), .ZN(n15529) );
  OAI21_X1 U17512 ( .B1(n15530), .B2(n16767), .A(n15529), .ZN(P2_U3016) );
  NOR2_X1 U17513 ( .A1(n15531), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15532) );
  MUX2_X1 U17514 ( .A(n15533), .B(n15532), .S(n19381), .Z(n18491) );
  NAND2_X1 U17515 ( .A1(n18491), .A2(n11050), .ZN(n15539) );
  XNOR2_X1 U17516 ( .A(n15539), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15544) );
  INV_X1 U17517 ( .A(n15544), .ZN(n15537) );
  OR2_X1 U17518 ( .A1(n15535), .A2(n15534), .ZN(n15538) );
  INV_X1 U17519 ( .A(n15538), .ZN(n15536) );
  NAND2_X1 U17520 ( .A1(n15537), .A2(n15536), .ZN(n15547) );
  NAND2_X1 U17521 ( .A1(n15538), .A2(n15561), .ZN(n15541) );
  NAND2_X1 U17522 ( .A1(n15542), .A2(n15561), .ZN(n15540) );
  MUX2_X1 U17523 ( .A(n15541), .B(n15540), .S(n15539), .Z(n15546) );
  INV_X1 U17524 ( .A(n15542), .ZN(n15543) );
  NAND3_X1 U17525 ( .A1(n11017), .A2(n15544), .A3(n15543), .ZN(n15545) );
  OAI211_X1 U17526 ( .C1(n11017), .C2(n15547), .A(n15546), .B(n15545), .ZN(
        n16347) );
  XOR2_X1 U17527 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n15548), .Z(
        n16345) );
  AOI222_X1 U17528 ( .A1(n13682), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n15550), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n13655), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15551) );
  INV_X1 U17529 ( .A(n15551), .ZN(n15552) );
  NAND2_X1 U17530 ( .A1(n15555), .A2(n15554), .ZN(n15560) );
  INV_X1 U17531 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n18492) );
  AOI22_X1 U17532 ( .A1(n15556), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n15557) );
  OAI21_X1 U17533 ( .B1(n15300), .B2(n18492), .A(n15557), .ZN(n15558) );
  AOI21_X1 U17534 ( .B1(n15293), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n15558), .ZN(n15559) );
  OR2_X1 U17535 ( .A1(n15562), .A2(n15561), .ZN(n15564) );
  NOR2_X1 U17536 ( .A1(n18521), .A2(n18492), .ZN(n16342) );
  AND2_X1 U17537 ( .A1(n15564), .A2(n15563), .ZN(n15565) );
  INV_X1 U17538 ( .A(n16868), .ZN(n15569) );
  INV_X1 U17539 ( .A(n15566), .ZN(n15568) );
  NAND3_X1 U17540 ( .A1(n15569), .A2(n15568), .A3(n15567), .ZN(n15570) );
  NAND2_X1 U17541 ( .A1(n13821), .A2(n15570), .ZN(n15574) );
  INV_X1 U17542 ( .A(n15571), .ZN(n15572) );
  NAND2_X1 U17543 ( .A1(n11577), .A2(n15572), .ZN(n15573) );
  OAI211_X1 U17544 ( .C1(n13821), .C2(n15575), .A(n15574), .B(n15573), .ZN(
        n15577) );
  NAND2_X1 U17545 ( .A1(n15577), .A2(n15576), .ZN(n16869) );
  INV_X1 U17546 ( .A(n16869), .ZN(n15583) );
  NAND3_X1 U17547 ( .A1(n15579), .A2(n21692), .A3(n15578), .ZN(n15580) );
  NAND2_X1 U17548 ( .A1(n15580), .A2(n21683), .ZN(n21273) );
  NAND2_X1 U17549 ( .A1(n15581), .A2(n21273), .ZN(n16872) );
  AND2_X1 U17550 ( .A1(n16872), .A2(n15582), .ZN(n21641) );
  MUX2_X1 U17551 ( .A(P1_MORE_REG_SCAN_IN), .B(n15583), .S(n21641), .Z(
        P1_U3484) );
  INV_X1 U17552 ( .A(n15598), .ZN(n15586) );
  INV_X1 U17553 ( .A(n10978), .ZN(n15584) );
  OAI22_X1 U17554 ( .A1(n15586), .A2(n10954), .B1(n15585), .B2(n15584), .ZN(
        n15588) );
  XNOR2_X1 U17555 ( .A(n15588), .B(n15587), .ZN(n15963) );
  AOI22_X1 U17556 ( .A1(n21615), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        n21597), .B2(P1_EBX_REG_30__SCAN_IN), .ZN(n15589) );
  OAI21_X1 U17557 ( .B1(n21613), .B2(n15809), .A(n15589), .ZN(n15593) );
  AOI21_X1 U17558 ( .B1(n15807), .B2(n15591), .A(n15590), .ZN(n15592) );
  INV_X1 U17559 ( .A(n15597), .ZN(n15613) );
  OAI21_X1 U17560 ( .B1(n10978), .B2(n15599), .A(n15598), .ZN(n15972) );
  AOI22_X1 U17561 ( .A1(n21615), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n21597), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n15601) );
  NAND2_X1 U17562 ( .A1(n21634), .A2(n15815), .ZN(n15600) );
  OAI211_X1 U17563 ( .C1(n15972), .C2(n21638), .A(n15601), .B(n15600), .ZN(
        n15603) );
  NOR3_X1 U17564 ( .A1(n15613), .A2(n21601), .A3(n19888), .ZN(n15602) );
  AOI211_X1 U17565 ( .C1(n15613), .C2(n19888), .A(n15603), .B(n15602), .ZN(
        n15604) );
  OAI21_X1 U17566 ( .B1(n15825), .B2(n21630), .A(n15604), .ZN(P1_U2811) );
  AOI21_X1 U17567 ( .B1(n15606), .B2(n15605), .A(n15595), .ZN(n15835) );
  INV_X1 U17568 ( .A(n15835), .ZN(n15735) );
  NAND2_X1 U17569 ( .A1(n11173), .A2(n15607), .ZN(n15609) );
  AOI21_X1 U17570 ( .B1(n15610), .B2(n15609), .A(n10978), .ZN(n15979) );
  AOI22_X1 U17571 ( .A1(n21615), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n21597), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n15611) );
  OAI21_X1 U17572 ( .B1(n21613), .B2(n15833), .A(n15611), .ZN(n15616) );
  AOI21_X1 U17573 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n21627), .A(n15612), 
        .ZN(n15614) );
  NOR2_X1 U17574 ( .A1(n15614), .A2(n15613), .ZN(n15615) );
  AOI211_X1 U17575 ( .C1(n21590), .C2(n15979), .A(n15616), .B(n15615), .ZN(
        n15617) );
  OAI21_X1 U17576 ( .B1(n15735), .B2(n21630), .A(n15617), .ZN(P1_U2812) );
  INV_X1 U17577 ( .A(n15605), .ZN(n15620) );
  AOI21_X1 U17578 ( .B1(n15621), .B2(n15619), .A(n15620), .ZN(n15843) );
  INV_X1 U17579 ( .A(n15843), .ZN(n15739) );
  INV_X1 U17580 ( .A(n15612), .ZN(n15627) );
  OAI21_X1 U17581 ( .B1(n21601), .B2(n19884), .A(n15638), .ZN(n15626) );
  XNOR2_X1 U17582 ( .A(n15634), .B(n15622), .ZN(n15993) );
  INV_X1 U17583 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15666) );
  OAI22_X1 U17584 ( .A1(n21626), .A2(n15841), .B1(n21623), .B2(n15666), .ZN(
        n15623) );
  AOI21_X1 U17585 ( .B1(n15839), .B2(n21634), .A(n15623), .ZN(n15624) );
  OAI21_X1 U17586 ( .B1(n15993), .B2(n21638), .A(n15624), .ZN(n15625) );
  AOI21_X1 U17587 ( .B1(n15627), .B2(n15626), .A(n15625), .ZN(n15628) );
  OAI21_X1 U17588 ( .B1(n15739), .B2(n21630), .A(n15628), .ZN(P1_U2813) );
  OAI21_X1 U17589 ( .B1(n15629), .B2(n15630), .A(n15619), .ZN(n15853) );
  INV_X1 U17590 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15845) );
  INV_X1 U17591 ( .A(n21629), .ZN(n15631) );
  OAI21_X1 U17592 ( .B1(n21601), .B2(n15845), .A(n15631), .ZN(n15639) );
  NAND2_X1 U17593 ( .A1(n11043), .A2(n15632), .ZN(n15633) );
  NAND2_X1 U17594 ( .A1(n15634), .A2(n15633), .ZN(n16005) );
  NOR2_X1 U17595 ( .A1(n16005), .A2(n21638), .ZN(n15637) );
  AOI22_X1 U17596 ( .A1(n21615), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n21597), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n15635) );
  OAI21_X1 U17597 ( .B1(n21613), .B2(n15846), .A(n15635), .ZN(n15636) );
  AOI211_X1 U17598 ( .C1(n15639), .C2(n15638), .A(n15637), .B(n15636), .ZN(
        n15640) );
  OAI21_X1 U17599 ( .B1(n15853), .B2(n21630), .A(n15640), .ZN(P1_U2814) );
  AOI21_X1 U17600 ( .B1(n15642), .B2(n15232), .A(n15641), .ZN(n19997) );
  INV_X1 U17601 ( .A(n19997), .ZN(n15793) );
  INV_X1 U17602 ( .A(n15720), .ZN(n15643) );
  AOI21_X1 U17603 ( .B1(n15645), .B2(n15644), .A(n15643), .ZN(n21387) );
  AOI22_X1 U17604 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n21615), .B1(
        n21597), .B2(P1_EBX_REG_16__SCAN_IN), .ZN(n15646) );
  OAI21_X1 U17605 ( .B1(n20000), .B2(n21613), .A(n15646), .ZN(n15647) );
  AOI211_X1 U17606 ( .C1(n21387), .C2(n21590), .A(n15647), .B(n21557), .ZN(
        n15651) );
  INV_X1 U17607 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15648) );
  NOR2_X1 U17608 ( .A1(n21601), .A2(n15648), .ZN(n15649) );
  OAI21_X1 U17609 ( .B1(n15236), .B2(n15649), .A(n21540), .ZN(n15650) );
  OAI211_X1 U17610 ( .C1(n15793), .C2(n21630), .A(n15651), .B(n15650), .ZN(
        P1_U2824) );
  INV_X1 U17611 ( .A(n15919), .ZN(n15802) );
  NAND4_X1 U17612 ( .A1(n15652), .A2(P1_REIP_REG_11__SCAN_IN), .A3(
        P1_REIP_REG_12__SCAN_IN), .A4(n21483), .ZN(n15653) );
  AND2_X1 U17613 ( .A1(n15653), .A2(n21627), .ZN(n21518) );
  INV_X1 U17614 ( .A(n15917), .ZN(n15654) );
  AOI22_X1 U17615 ( .A1(n15654), .A2(n21634), .B1(n21615), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15655) );
  OAI211_X1 U17616 ( .C1(n15656), .C2(n21623), .A(n15655), .B(n21485), .ZN(
        n15659) );
  OAI22_X1 U17617 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15657), .B1(n21638), 
        .B2(n16068), .ZN(n15658) );
  AOI211_X1 U17618 ( .C1(n21518), .C2(P1_REIP_REG_13__SCAN_IN), .A(n15659), 
        .B(n15658), .ZN(n15660) );
  OAI21_X1 U17619 ( .B1(n15802), .B2(n21630), .A(n15660), .ZN(P1_U2827) );
  INV_X1 U17620 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15661) );
  OAI22_X1 U17621 ( .A1(n15931), .A2(n19942), .B1(n15661), .B2(n19946), .ZN(
        P1_U2841) );
  AOI22_X1 U17622 ( .A1(n15963), .A2(n19925), .B1(n15724), .B2(
        P1_EBX_REG_30__SCAN_IN), .ZN(n15662) );
  OAI21_X1 U17623 ( .B1(n15663), .B2(n15726), .A(n15662), .ZN(P1_U2842) );
  INV_X1 U17624 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15664) );
  OAI222_X1 U17625 ( .A1(n15664), .A2(n19946), .B1(n19942), .B2(n15972), .C1(
        n15825), .C2(n15726), .ZN(P1_U2843) );
  AOI22_X1 U17626 ( .A1(n15979), .A2(n19925), .B1(n15724), .B2(
        P1_EBX_REG_28__SCAN_IN), .ZN(n15665) );
  OAI21_X1 U17627 ( .B1(n15735), .B2(n15726), .A(n15665), .ZN(P1_U2844) );
  OAI222_X1 U17628 ( .A1(n15666), .A2(n19946), .B1(n19942), .B2(n15993), .C1(
        n15726), .C2(n15739), .ZN(P1_U2845) );
  INV_X1 U17629 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15667) );
  OAI222_X1 U17630 ( .A1(n15667), .A2(n19946), .B1(n19942), .B2(n16005), .C1(
        n15853), .C2(n15726), .ZN(P1_U2846) );
  INV_X1 U17631 ( .A(n15629), .ZN(n15669) );
  OAI21_X1 U17632 ( .B1(n15670), .B2(n15668), .A(n15669), .ZN(n21631) );
  INV_X1 U17633 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21624) );
  OR2_X1 U17634 ( .A1(n15671), .A2(n15672), .ZN(n15673) );
  NAND2_X1 U17635 ( .A1(n11043), .A2(n15673), .ZN(n21637) );
  OAI222_X1 U17636 ( .A1(n15726), .A2(n21631), .B1(n19946), .B2(n21624), .C1(
        n21637), .C2(n19942), .ZN(P1_U2847) );
  INV_X1 U17637 ( .A(n15674), .ZN(n15686) );
  INV_X1 U17638 ( .A(n15675), .ZN(n15677) );
  INV_X1 U17639 ( .A(n15676), .ZN(n15747) );
  OAI21_X1 U17640 ( .B1(n15686), .B2(n15677), .A(n15747), .ZN(n21603) );
  INV_X1 U17641 ( .A(n19929), .ZN(n15680) );
  NAND2_X1 U17642 ( .A1(n15689), .A2(n15678), .ZN(n15679) );
  NAND2_X1 U17643 ( .A1(n15680), .A2(n15679), .ZN(n21602) );
  INV_X1 U17644 ( .A(n21602), .ZN(n15681) );
  AOI22_X1 U17645 ( .A1(n15681), .A2(n19925), .B1(n15724), .B2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n15682) );
  OAI21_X1 U17646 ( .B1(n21603), .B2(n15726), .A(n15682), .ZN(P1_U2849) );
  INV_X1 U17647 ( .A(n15683), .ZN(n15688) );
  INV_X1 U17648 ( .A(n15685), .ZN(n15687) );
  INV_X1 U17649 ( .A(n21591), .ZN(n15761) );
  INV_X1 U17650 ( .A(n15689), .ZN(n15690) );
  AOI21_X1 U17651 ( .B1(n15691), .B2(n15698), .A(n15690), .ZN(n21589) );
  AOI22_X1 U17652 ( .A1(n21589), .A2(n19925), .B1(n15724), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n15692) );
  OAI21_X1 U17653 ( .B1(n15761), .B2(n15726), .A(n15692), .ZN(P1_U2850) );
  AOI21_X1 U17654 ( .B1(n15695), .B2(n15694), .A(n15685), .ZN(n21582) );
  OR2_X1 U17655 ( .A1(n19936), .A2(n15696), .ZN(n15697) );
  NAND2_X1 U17656 ( .A1(n15698), .A2(n15697), .ZN(n21585) );
  INV_X1 U17657 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n21576) );
  OAI22_X1 U17658 ( .A1(n21585), .A2(n19942), .B1(n21576), .B2(n19946), .ZN(
        n15699) );
  AOI21_X1 U17659 ( .B1(n21582), .B2(n19932), .A(n15699), .ZN(n15700) );
  INV_X1 U17660 ( .A(n15700), .ZN(P1_U2851) );
  INV_X1 U17661 ( .A(n15701), .ZN(n15704) );
  OAI21_X1 U17662 ( .B1(n15704), .B2(n11062), .A(n15766), .ZN(n21559) );
  NOR2_X1 U17663 ( .A1(n15713), .A2(n15706), .ZN(n15707) );
  OR2_X1 U17664 ( .A1(n15705), .A2(n15707), .ZN(n21555) );
  INV_X1 U17665 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n21554) );
  OAI22_X1 U17666 ( .A1(n21555), .A2(n19942), .B1(n21554), .B2(n19946), .ZN(
        n15708) );
  INV_X1 U17667 ( .A(n15708), .ZN(n15709) );
  OAI21_X1 U17668 ( .B1(n21559), .B2(n15726), .A(n15709), .ZN(P1_U2853) );
  OR2_X1 U17669 ( .A1(n15710), .A2(n15711), .ZN(n15712) );
  AND2_X1 U17670 ( .A1(n15701), .A2(n15712), .ZN(n21548) );
  INV_X1 U17671 ( .A(n21548), .ZN(n15780) );
  AOI21_X1 U17672 ( .B1(n15714), .B2(n11046), .A(n15713), .ZN(n21549) );
  AOI22_X1 U17673 ( .A1(n21549), .A2(n19925), .B1(n15724), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n15715) );
  OAI21_X1 U17674 ( .B1(n15780), .B2(n15726), .A(n15715), .ZN(P1_U2854) );
  INV_X1 U17675 ( .A(n15716), .ZN(n15718) );
  INV_X1 U17676 ( .A(n15641), .ZN(n15717) );
  AOI21_X1 U17677 ( .B1(n15718), .B2(n15717), .A(n15710), .ZN(n21542) );
  NAND2_X1 U17678 ( .A1(n15720), .A2(n15719), .ZN(n15721) );
  NAND2_X1 U17679 ( .A1(n11046), .A2(n15721), .ZN(n21545) );
  OAI22_X1 U17680 ( .A1(n21545), .A2(n19942), .B1(n21534), .B2(n19946), .ZN(
        n15722) );
  AOI21_X1 U17681 ( .B1(n21542), .B2(n19932), .A(n15722), .ZN(n15723) );
  INV_X1 U17682 ( .A(n15723), .ZN(P1_U2855) );
  AOI22_X1 U17683 ( .A1(n21387), .A2(n19925), .B1(n15724), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n15725) );
  OAI21_X1 U17684 ( .B1(n15793), .B2(n15726), .A(n15725), .ZN(P1_U2856) );
  AOI22_X1 U17685 ( .A1(n15776), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n15798), .ZN(n15729) );
  MUX2_X1 U17686 ( .A(BUF1_REG_13__SCAN_IN), .B(DATAI_13_), .S(n15727), .Z(
        n21763) );
  AOI22_X1 U17687 ( .A1(n15790), .A2(n21763), .B1(n15788), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15728) );
  OAI211_X1 U17688 ( .C1(n15825), .C2(n15801), .A(n15729), .B(n15728), .ZN(
        P1_U2875) );
  OAI22_X1 U17689 ( .A1(n15786), .A2(n15731), .B1(n15730), .B2(n15794), .ZN(
        n15732) );
  INV_X1 U17690 ( .A(n15732), .ZN(n15734) );
  AOI22_X1 U17691 ( .A1(n15790), .A2(n21757), .B1(n15788), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15733) );
  OAI211_X1 U17692 ( .C1(n15735), .C2(n15801), .A(n15734), .B(n15733), .ZN(
        P1_U2876) );
  AOI22_X1 U17693 ( .A1(n15776), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n15798), .ZN(n15738) );
  INV_X1 U17694 ( .A(n21752), .ZN(n15736) );
  AOI22_X1 U17695 ( .A1(n15790), .A2(n15736), .B1(n15788), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15737) );
  OAI211_X1 U17696 ( .C1(n15739), .C2(n15801), .A(n15738), .B(n15737), .ZN(
        P1_U2877) );
  AOI22_X1 U17697 ( .A1(n15776), .A2(DATAI_26_), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n15798), .ZN(n15742) );
  INV_X1 U17698 ( .A(n21747), .ZN(n15740) );
  AOI22_X1 U17699 ( .A1(n15790), .A2(n15740), .B1(n15788), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15741) );
  OAI211_X1 U17700 ( .C1(n15853), .C2(n15801), .A(n15742), .B(n15741), .ZN(
        P1_U2878) );
  AOI22_X1 U17701 ( .A1(n15776), .A2(DATAI_25_), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n15798), .ZN(n15745) );
  INV_X1 U17702 ( .A(n15743), .ZN(n21739) );
  AOI22_X1 U17703 ( .A1(n15790), .A2(n21739), .B1(n15788), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15744) );
  OAI211_X1 U17704 ( .C1(n21631), .C2(n15801), .A(n15745), .B(n15744), .ZN(
        P1_U2879) );
  AND2_X1 U17705 ( .A1(n15747), .A2(n15746), .ZN(n15748) );
  NOR2_X1 U17706 ( .A1(n15668), .A2(n15748), .ZN(n21619) );
  INV_X1 U17707 ( .A(n21619), .ZN(n15753) );
  OAI22_X1 U17708 ( .A1(n15786), .A2(n17010), .B1(n21736), .B2(n15794), .ZN(
        n15751) );
  INV_X1 U17709 ( .A(n15790), .ZN(n15749) );
  NOR2_X1 U17710 ( .A1(n15749), .A2(n21734), .ZN(n15750) );
  AOI211_X1 U17711 ( .C1(BUF1_REG_24__SCAN_IN), .C2(n15788), .A(n15751), .B(
        n15750), .ZN(n15752) );
  OAI21_X1 U17712 ( .B1(n15753), .B2(n15801), .A(n15752), .ZN(P1_U2880) );
  OAI22_X1 U17713 ( .A1(n15786), .A2(n14397), .B1(n14634), .B2(n15794), .ZN(
        n15754) );
  INV_X1 U17714 ( .A(n15754), .ZN(n15757) );
  AOI22_X1 U17715 ( .A1(n15790), .A2(n15755), .B1(n15788), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15756) );
  OAI211_X1 U17716 ( .C1(n21603), .C2(n15801), .A(n15757), .B(n15756), .ZN(
        P1_U2881) );
  AOI22_X1 U17717 ( .A1(n15776), .A2(DATAI_22_), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n15798), .ZN(n15760) );
  AOI22_X1 U17718 ( .A1(n15790), .A2(n15758), .B1(n15788), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15759) );
  OAI211_X1 U17719 ( .C1(n15761), .C2(n15801), .A(n15760), .B(n15759), .ZN(
        P1_U2882) );
  INV_X1 U17720 ( .A(n21582), .ZN(n15875) );
  AOI22_X1 U17721 ( .A1(n15776), .A2(DATAI_21_), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n15798), .ZN(n15764) );
  AOI22_X1 U17722 ( .A1(n15790), .A2(n15762), .B1(n15788), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n15763) );
  OAI211_X1 U17723 ( .C1(n15875), .C2(n15801), .A(n15764), .B(n15763), .ZN(
        P1_U2883) );
  NAND2_X1 U17724 ( .A1(n15766), .A2(n15765), .ZN(n15767) );
  NAND2_X1 U17725 ( .A1(n15694), .A2(n15767), .ZN(n21569) );
  OAI22_X1 U17726 ( .A1(n15786), .A2(n17021), .B1(n15768), .B2(n15794), .ZN(
        n15769) );
  INV_X1 U17727 ( .A(n15769), .ZN(n15772) );
  AOI22_X1 U17728 ( .A1(n15790), .A2(n15770), .B1(n15788), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n15771) );
  OAI211_X1 U17729 ( .C1(n21569), .C2(n15801), .A(n15772), .B(n15771), .ZN(
        P1_U2884) );
  AOI22_X1 U17730 ( .A1(n15776), .A2(DATAI_19_), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n15798), .ZN(n15775) );
  AOI22_X1 U17731 ( .A1(n15790), .A2(n15773), .B1(n15788), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n15774) );
  OAI211_X1 U17732 ( .C1(n21559), .C2(n15801), .A(n15775), .B(n15774), .ZN(
        P1_U2885) );
  AOI22_X1 U17733 ( .A1(n15776), .A2(DATAI_18_), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n15798), .ZN(n15779) );
  AOI22_X1 U17734 ( .A1(n15790), .A2(n15777), .B1(n15788), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15778) );
  OAI211_X1 U17735 ( .C1(n15780), .C2(n15801), .A(n15779), .B(n15778), .ZN(
        P1_U2886) );
  INV_X1 U17736 ( .A(n21542), .ZN(n15901) );
  OAI22_X1 U17737 ( .A1(n15786), .A2(n14409), .B1(n14239), .B2(n15794), .ZN(
        n15781) );
  INV_X1 U17738 ( .A(n15781), .ZN(n15784) );
  AOI22_X1 U17739 ( .A1(n15790), .A2(n15782), .B1(n15788), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n15783) );
  OAI211_X1 U17740 ( .C1(n15901), .C2(n15801), .A(n15784), .B(n15783), .ZN(
        P1_U2887) );
  OAI22_X1 U17741 ( .A1(n15786), .A2(n17026), .B1(n15785), .B2(n15794), .ZN(
        n15787) );
  INV_X1 U17742 ( .A(n15787), .ZN(n15792) );
  AOI22_X1 U17743 ( .A1(n15790), .A2(n15789), .B1(n15788), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n15791) );
  OAI211_X1 U17744 ( .C1(n15793), .C2(n15801), .A(n15792), .B(n15791), .ZN(
        P1_U2888) );
  OAI222_X1 U17745 ( .A1(n15797), .A2(n15801), .B1(n15796), .B2(n15795), .C1(
        n15794), .C2(n19844), .ZN(P1_U2889) );
  AOI22_X1 U17746 ( .A1(n15799), .A2(n21763), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15798), .ZN(n15800) );
  OAI21_X1 U17747 ( .B1(n15802), .B2(n15801), .A(n15800), .ZN(P1_U2891) );
  NAND2_X1 U17748 ( .A1(n19993), .A2(n15981), .ZN(n15803) );
  NAND2_X1 U17749 ( .A1(n15980), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15960) );
  MUX2_X1 U17750 ( .A(n15803), .B(n15960), .S(n15838), .Z(n15805) );
  INV_X1 U17751 ( .A(n15820), .ZN(n15804) );
  XNOR2_X1 U17752 ( .A(n15806), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15966) );
  NOR2_X1 U17753 ( .A1(n21419), .A2(n15807), .ZN(n15962) );
  AOI21_X1 U17754 ( .B1(n20014), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15962), .ZN(n15808) );
  OAI21_X1 U17755 ( .B1(n20024), .B2(n15809), .A(n15808), .ZN(n15810) );
  AOI21_X1 U17756 ( .B1(n15811), .B2(n20021), .A(n15810), .ZN(n15812) );
  OAI21_X1 U17757 ( .B1(n15966), .B2(n21639), .A(n15812), .ZN(P1_U2969) );
  NAND2_X1 U17758 ( .A1(n14073), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15971) );
  OAI21_X1 U17759 ( .B1(n15898), .B2(n15813), .A(n15971), .ZN(n15814) );
  AOI21_X1 U17760 ( .B1(n15815), .B2(n19989), .A(n15814), .ZN(n15824) );
  AOI21_X1 U17761 ( .B1(n15820), .B2(n15816), .A(n15818), .ZN(n15822) );
  INV_X1 U17762 ( .A(n15817), .ZN(n15821) );
  INV_X1 U17763 ( .A(n15818), .ZN(n15819) );
  NAND2_X1 U17764 ( .A1(n15967), .A2(n20020), .ZN(n15823) );
  OAI211_X1 U17765 ( .C1(n15825), .C2(n19975), .A(n15824), .B(n15823), .ZN(
        P1_U2970) );
  NAND2_X1 U17766 ( .A1(n20018), .A2(n15848), .ZN(n15830) );
  OAI21_X1 U17767 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15827), .A(
        n15830), .ZN(n15829) );
  MUX2_X1 U17768 ( .A(n15990), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n20015), .Z(n15828) );
  OAI211_X1 U17769 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15830), .A(
        n15829), .B(n15828), .ZN(n15831) );
  XOR2_X1 U17770 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n15831), .Z(
        n15988) );
  NAND2_X1 U17771 ( .A1(n14073), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15984) );
  NAND2_X1 U17772 ( .A1(n20014), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15832) );
  OAI211_X1 U17773 ( .C1(n20024), .C2(n15833), .A(n15984), .B(n15832), .ZN(
        n15834) );
  AOI21_X1 U17774 ( .B1(n15835), .B2(n20021), .A(n15834), .ZN(n15836) );
  OAI21_X1 U17775 ( .B1(n21639), .B2(n15988), .A(n15836), .ZN(P1_U2971) );
  XNOR2_X1 U17776 ( .A(n12852), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15837) );
  XNOR2_X1 U17777 ( .A(n15838), .B(n15837), .ZN(n15997) );
  NAND2_X1 U17778 ( .A1(n19989), .A2(n15839), .ZN(n15840) );
  NAND2_X1 U17779 ( .A1(n14073), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15992) );
  OAI211_X1 U17780 ( .C1(n15898), .C2(n15841), .A(n15840), .B(n15992), .ZN(
        n15842) );
  AOI21_X1 U17781 ( .B1(n15843), .B2(n20021), .A(n15842), .ZN(n15844) );
  OAI21_X1 U17782 ( .B1(n15997), .B2(n21639), .A(n15844), .ZN(P1_U2972) );
  NOR2_X1 U17783 ( .A1(n21419), .A2(n15845), .ZN(n16002) );
  NOR2_X1 U17784 ( .A1(n20024), .A2(n15846), .ZN(n15847) );
  AOI211_X1 U17785 ( .C1(n20014), .C2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16002), .B(n15847), .ZN(n15852) );
  NAND3_X1 U17786 ( .A1(n15849), .A2(n15854), .A3(n15848), .ZN(n15850) );
  XNOR2_X1 U17787 ( .A(n15850), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16007) );
  NAND2_X1 U17788 ( .A1(n16007), .A2(n20020), .ZN(n15851) );
  OAI211_X1 U17789 ( .C1(n15853), .C2(n19975), .A(n15852), .B(n15851), .ZN(
        P1_U2973) );
  NOR2_X1 U17790 ( .A1(n20018), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15855) );
  NAND2_X1 U17791 ( .A1(n19993), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15864) );
  OAI211_X1 U17792 ( .C1(n15855), .C2(n15951), .A(n15854), .B(n15864), .ZN(
        n15856) );
  XNOR2_X1 U17793 ( .A(n15856), .B(n16011), .ZN(n16016) );
  INV_X1 U17794 ( .A(n21631), .ZN(n15860) );
  INV_X1 U17795 ( .A(n21635), .ZN(n15858) );
  AOI22_X1 U17796 ( .A1(n20014), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n14073), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n15857) );
  OAI21_X1 U17797 ( .B1(n20024), .B2(n15858), .A(n15857), .ZN(n15859) );
  AOI21_X1 U17798 ( .B1(n15860), .B2(n20021), .A(n15859), .ZN(n15861) );
  OAI21_X1 U17799 ( .B1(n21639), .B2(n16016), .A(n15861), .ZN(P1_U2974) );
  NOR2_X1 U17800 ( .A1(n21419), .A2(n21600), .ZN(n16020) );
  INV_X1 U17801 ( .A(n21598), .ZN(n15862) );
  NOR2_X1 U17802 ( .A1(n20024), .A2(n15862), .ZN(n15863) );
  AOI211_X1 U17803 ( .C1(n20014), .C2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16020), .B(n15863), .ZN(n15867) );
  OAI21_X1 U17804 ( .B1(n19993), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15864), .ZN(n15865) );
  XNOR2_X1 U17805 ( .A(n20018), .B(n15865), .ZN(n16017) );
  NAND2_X1 U17806 ( .A1(n16017), .A2(n20020), .ZN(n15866) );
  OAI211_X1 U17807 ( .C1(n21603), .C2(n19975), .A(n15867), .B(n15866), .ZN(
        P1_U2976) );
  INV_X1 U17808 ( .A(n15868), .ZN(n15882) );
  XNOR2_X1 U17809 ( .A(n19971), .B(n16041), .ZN(n15881) );
  AOI21_X1 U17810 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n20001), .A(
        n21398), .ZN(n15869) );
  MUX2_X1 U17811 ( .A(n15876), .B(n20001), .S(n19993), .Z(n20002) );
  XNOR2_X1 U17812 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n15870), .ZN(
        n21416) );
  INV_X1 U17813 ( .A(n21416), .ZN(n15871) );
  OAI22_X1 U17814 ( .A1(n21639), .A2(n15871), .B1(n21419), .B2(n21592), .ZN(
        n15872) );
  AOI21_X1 U17815 ( .B1(n20014), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15872), .ZN(n15874) );
  NAND2_X1 U17816 ( .A1(n19989), .A2(n21580), .ZN(n15873) );
  OAI211_X1 U17817 ( .C1(n15875), .C2(n19975), .A(n15874), .B(n15873), .ZN(
        P1_U2978) );
  XNOR2_X1 U17818 ( .A(n12852), .B(n15876), .ZN(n15877) );
  XNOR2_X1 U17819 ( .A(n20001), .B(n15877), .ZN(n16025) );
  NAND2_X1 U17820 ( .A1(n16025), .A2(n20020), .ZN(n15880) );
  NOR2_X1 U17821 ( .A1(n21419), .A2(n19870), .ZN(n16029) );
  NOR2_X1 U17822 ( .A1(n20024), .A2(n21564), .ZN(n15878) );
  AOI211_X1 U17823 ( .C1(n20014), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16029), .B(n15878), .ZN(n15879) );
  OAI211_X1 U17824 ( .C1(n19975), .C2(n21559), .A(n15880), .B(n15879), .ZN(
        P1_U2980) );
  XNOR2_X1 U17825 ( .A(n15882), .B(n15881), .ZN(n16045) );
  NAND2_X1 U17826 ( .A1(n14073), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16037) );
  NAND2_X1 U17827 ( .A1(n20014), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15883) );
  OAI211_X1 U17828 ( .C1(n20024), .C2(n15884), .A(n16037), .B(n15883), .ZN(
        n15885) );
  AOI21_X1 U17829 ( .B1(n21548), .B2(n20021), .A(n15885), .ZN(n15886) );
  OAI21_X1 U17830 ( .B1(n16045), .B2(n21639), .A(n15886), .ZN(P1_U2981) );
  NAND2_X1 U17831 ( .A1(n14073), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16047) );
  OR2_X1 U17832 ( .A1(n15887), .A2(n15888), .ZN(n19982) );
  OR2_X1 U17833 ( .A1(n20015), .A2(n16058), .ZN(n19994) );
  OAI211_X1 U17834 ( .C1(n20015), .C2(n21287), .A(n19994), .B(n19983), .ZN(
        n15889) );
  AOI21_X1 U17835 ( .B1(n15890), .B2(n19982), .A(n15889), .ZN(n15891) );
  INV_X1 U17836 ( .A(n16046), .ZN(n21384) );
  NOR2_X1 U17837 ( .A1(n15891), .A2(n21384), .ZN(n15894) );
  INV_X1 U17838 ( .A(n15891), .ZN(n15892) );
  NOR2_X1 U17839 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15892), .ZN(
        n15893) );
  MUX2_X1 U17840 ( .A(n15894), .B(n15893), .S(n19993), .Z(n15895) );
  XNOR2_X1 U17841 ( .A(n15896), .B(n15895), .ZN(n16050) );
  NAND2_X1 U17842 ( .A1(n20020), .A2(n16050), .ZN(n15897) );
  OAI211_X1 U17843 ( .C1(n15898), .C2(n21535), .A(n16047), .B(n15897), .ZN(
        n15899) );
  AOI21_X1 U17844 ( .B1(n19989), .B2(n21537), .A(n15899), .ZN(n15900) );
  OAI21_X1 U17845 ( .B1(n15901), .B2(n19975), .A(n15900), .ZN(P1_U2982) );
  NOR2_X1 U17846 ( .A1(n11032), .A2(n15902), .ZN(n19992) );
  OAI21_X1 U17847 ( .B1(n19993), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n19994), .ZN(n15903) );
  XNOR2_X1 U17848 ( .A(n19992), .B(n15903), .ZN(n16060) );
  NAND2_X1 U17849 ( .A1(n20014), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15904) );
  NAND2_X1 U17850 ( .A1(n14073), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n16054) );
  OAI211_X1 U17851 ( .C1(n20024), .C2(n15905), .A(n15904), .B(n16054), .ZN(
        n15906) );
  AOI21_X1 U17852 ( .B1(n15907), .B2(n20021), .A(n15906), .ZN(n15908) );
  OAI21_X1 U17853 ( .B1(n16060), .B2(n21639), .A(n15908), .ZN(P1_U2984) );
  INV_X1 U17854 ( .A(n15909), .ZN(n15910) );
  AOI21_X1 U17855 ( .B1(n15887), .B2(n15911), .A(n15910), .ZN(n19978) );
  AND2_X1 U17856 ( .A1(n15912), .A2(n15913), .ZN(n19977) );
  NAND2_X1 U17857 ( .A1(n19978), .A2(n19977), .ZN(n19976) );
  NAND2_X1 U17858 ( .A1(n19976), .A2(n15913), .ZN(n15915) );
  XNOR2_X1 U17859 ( .A(n15915), .B(n15914), .ZN(n16072) );
  AOI22_X1 U17860 ( .A1(n20014), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n14073), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n15916) );
  OAI21_X1 U17861 ( .B1(n20024), .B2(n15917), .A(n15916), .ZN(n15918) );
  AOI21_X1 U17862 ( .B1(n15919), .B2(n20021), .A(n15918), .ZN(n15920) );
  OAI21_X1 U17863 ( .B1(n16072), .B2(n21639), .A(n15920), .ZN(P1_U2986) );
  MUX2_X1 U17864 ( .A(n15921), .B(n15887), .S(n19993), .Z(n15922) );
  AOI21_X1 U17865 ( .B1(n15923), .B2(n20015), .A(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15925) );
  NOR3_X1 U17866 ( .A1(n19972), .A2(n15887), .A3(n19971), .ZN(n19970) );
  INV_X1 U17867 ( .A(n19970), .ZN(n15924) );
  OAI21_X1 U17868 ( .B1(n19972), .B2(n15925), .A(n15924), .ZN(n21357) );
  NAND2_X1 U17869 ( .A1(n21357), .A2(n20020), .ZN(n15929) );
  NOR2_X1 U17870 ( .A1(n21419), .A2(n19857), .ZN(n21355) );
  NOR2_X1 U17871 ( .A1(n20024), .A2(n15926), .ZN(n15927) );
  AOI211_X1 U17872 ( .C1(n20014), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n21355), .B(n15927), .ZN(n15928) );
  OAI211_X1 U17873 ( .C1(n19975), .C2(n15930), .A(n15929), .B(n15928), .ZN(
        P1_U2989) );
  NOR2_X1 U17874 ( .A1(n15931), .A2(n21414), .ZN(n15956) );
  NOR2_X1 U17875 ( .A1(n21406), .A2(n21408), .ZN(n15948) );
  NAND2_X1 U17876 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15937) );
  INV_X1 U17877 ( .A(n15937), .ZN(n21342) );
  NAND3_X1 U17878 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n21342), .ZN(n21346) );
  NOR2_X1 U17879 ( .A1(n15933), .A2(n15932), .ZN(n15938) );
  INV_X1 U17880 ( .A(n15938), .ZN(n21353) );
  NOR3_X1 U17881 ( .A1(n21346), .A2(n21353), .A3(n15934), .ZN(n21364) );
  NAND3_X1 U17882 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n21364), .ZN(n16061) );
  NAND2_X1 U17883 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16039) );
  OR3_X1 U17884 ( .A1(n16041), .A2(n16040), .A3(n16039), .ZN(n16024) );
  NOR2_X1 U17885 ( .A1(n16061), .A2(n16024), .ZN(n15949) );
  INV_X1 U17886 ( .A(n15949), .ZN(n15935) );
  AOI21_X1 U17887 ( .B1(n21366), .B2(n15935), .A(n21401), .ZN(n16026) );
  NAND2_X1 U17888 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15936), .ZN(
        n21322) );
  NOR2_X1 U17889 ( .A1(n15937), .A2(n21322), .ZN(n21349) );
  NAND2_X1 U17890 ( .A1(n15938), .A2(n21349), .ZN(n16023) );
  NOR2_X1 U17891 ( .A1(n11614), .A2(n16023), .ZN(n21369) );
  NAND2_X1 U17892 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21369), .ZN(
        n16064) );
  NOR2_X1 U17893 ( .A1(n16024), .A2(n16064), .ZN(n16027) );
  NAND2_X1 U17894 ( .A1(n15948), .A2(n16027), .ZN(n15950) );
  OAI21_X1 U17895 ( .B1(n15939), .B2(n15950), .A(n16033), .ZN(n15940) );
  OAI211_X1 U17896 ( .C1(n15941), .C2(n15948), .A(n16026), .B(n15940), .ZN(
        n21426) );
  OAI22_X1 U17897 ( .A1(n15943), .A2(n16062), .B1(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15942), .ZN(n15944) );
  AOI211_X1 U17898 ( .C1(n21429), .C2(n15945), .A(n21426), .B(n15944), .ZN(
        n16010) );
  NAND3_X1 U17899 ( .A1(n16010), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15978) );
  NAND2_X1 U17900 ( .A1(n16010), .A2(n16032), .ZN(n15977) );
  OAI21_X1 U17901 ( .B1(n15978), .B2(n15960), .A(n15977), .ZN(n15959) );
  INV_X1 U17902 ( .A(n15977), .ZN(n15947) );
  AOI211_X1 U17903 ( .C1(n15959), .C2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15947), .B(n15946), .ZN(n15955) );
  NAND2_X1 U17904 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16000) );
  NAND3_X1 U17905 ( .A1(n15949), .A2(n15948), .A3(n21301), .ZN(n21425) );
  OAI21_X1 U17906 ( .B1(n15950), .B2(n21368), .A(n21425), .ZN(n21428) );
  NAND2_X1 U17907 ( .A1(n15951), .A2(n21428), .ZN(n16012) );
  OR2_X1 U17908 ( .A1(n16000), .A2(n16012), .ZN(n15968) );
  NOR4_X1 U17909 ( .A1(n15960), .A2(n15952), .A3(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A4(n15968), .ZN(n15953) );
  NOR4_X1 U17910 ( .A1(n15956), .A2(n15955), .A3(n15954), .A4(n15953), .ZN(
        n15957) );
  OAI21_X1 U17911 ( .B1(n15958), .B2(n21382), .A(n15957), .ZN(P1_U3000) );
  INV_X1 U17912 ( .A(n15959), .ZN(n15974) );
  NOR3_X1 U17913 ( .A1(n15960), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15968), .ZN(n15961) );
  AOI211_X1 U17914 ( .C1(n15974), .C2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15962), .B(n15961), .ZN(n15965) );
  NAND2_X1 U17915 ( .A1(n15963), .A2(n21421), .ZN(n15964) );
  OAI211_X1 U17916 ( .C1(n15966), .C2(n21382), .A(n15965), .B(n15964), .ZN(
        P1_U3001) );
  INV_X1 U17917 ( .A(n15967), .ZN(n15976) );
  INV_X1 U17918 ( .A(n15968), .ZN(n15989) );
  NAND3_X1 U17919 ( .A1(n15980), .A2(n15989), .A3(n15969), .ZN(n15970) );
  OAI211_X1 U17920 ( .C1(n15972), .C2(n21414), .A(n15971), .B(n15970), .ZN(
        n15973) );
  AOI21_X1 U17921 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15974), .A(
        n15973), .ZN(n15975) );
  OAI21_X1 U17922 ( .B1(n15976), .B2(n21382), .A(n15975), .ZN(P1_U3002) );
  AND2_X1 U17923 ( .A1(n15978), .A2(n15977), .ZN(n15995) );
  INV_X1 U17924 ( .A(n15979), .ZN(n15985) );
  NOR2_X1 U17925 ( .A1(n15981), .A2(n15980), .ZN(n15982) );
  NAND2_X1 U17926 ( .A1(n15989), .A2(n15982), .ZN(n15983) );
  OAI211_X1 U17927 ( .C1(n15985), .C2(n21414), .A(n15984), .B(n15983), .ZN(
        n15986) );
  AOI21_X1 U17928 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n15995), .A(
        n15986), .ZN(n15987) );
  OAI21_X1 U17929 ( .B1(n15988), .B2(n21382), .A(n15987), .ZN(P1_U3003) );
  NAND2_X1 U17930 ( .A1(n15990), .A2(n15989), .ZN(n15991) );
  OAI211_X1 U17931 ( .C1(n15993), .C2(n21414), .A(n15992), .B(n15991), .ZN(
        n15994) );
  AOI21_X1 U17932 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15995), .A(
        n15994), .ZN(n15996) );
  OAI21_X1 U17933 ( .B1(n15997), .B2(n21382), .A(n15996), .ZN(P1_U3004) );
  INV_X1 U17934 ( .A(n16010), .ZN(n16001) );
  AOI21_X1 U17935 ( .B1(n16011), .B2(n15998), .A(n16012), .ZN(n15999) );
  AOI22_X1 U17936 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n16001), .B1(
        n16000), .B2(n15999), .ZN(n16004) );
  INV_X1 U17937 ( .A(n16002), .ZN(n16003) );
  OAI211_X1 U17938 ( .C1(n16005), .C2(n21414), .A(n16004), .B(n16003), .ZN(
        n16006) );
  AOI21_X1 U17939 ( .B1(n16007), .B2(n21422), .A(n16006), .ZN(n16008) );
  INV_X1 U17940 ( .A(n16008), .ZN(P1_U3005) );
  INV_X1 U17941 ( .A(n21637), .ZN(n16014) );
  NAND2_X1 U17942 ( .A1(n14073), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n16009) );
  OAI221_X1 U17943 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16012), 
        .C1(n16011), .C2(n16010), .A(n16009), .ZN(n16013) );
  AOI21_X1 U17944 ( .B1(n16014), .B2(n21421), .A(n16013), .ZN(n16015) );
  OAI21_X1 U17945 ( .B1(n16016), .B2(n21382), .A(n16015), .ZN(P1_U3006) );
  NAND2_X1 U17946 ( .A1(n16017), .A2(n21422), .ZN(n16022) );
  INV_X1 U17947 ( .A(n21428), .ZN(n16018) );
  NOR2_X1 U17948 ( .A1(n16018), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16019) );
  AOI211_X1 U17949 ( .C1(n21426), .C2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16020), .B(n16019), .ZN(n16021) );
  OAI211_X1 U17950 ( .C1(n21414), .C2(n21602), .A(n16022), .B(n16021), .ZN(
        P1_U3008) );
  NAND2_X1 U17951 ( .A1(n21364), .A2(n21301), .ZN(n21371) );
  OAI21_X1 U17952 ( .B1(n16023), .B2(n21368), .A(n21371), .ZN(n21378) );
  NAND3_X1 U17953 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n21378), .ZN(n21281) );
  NOR2_X1 U17954 ( .A1(n16024), .A2(n21281), .ZN(n21404) );
  INV_X1 U17955 ( .A(n21404), .ZN(n21407) );
  NAND2_X1 U17956 ( .A1(n16025), .A2(n21422), .ZN(n16031) );
  OAI21_X1 U17957 ( .B1(n16027), .B2(n21368), .A(n16026), .ZN(n21403) );
  NOR2_X1 U17958 ( .A1(n21555), .A2(n21414), .ZN(n16028) );
  AOI211_X1 U17959 ( .C1(n21403), .C2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16029), .B(n16028), .ZN(n16030) );
  OAI211_X1 U17960 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n21407), .A(
        n16031), .B(n16030), .ZN(P1_U3012) );
  INV_X1 U17961 ( .A(n16032), .ZN(n21400) );
  INV_X1 U17962 ( .A(n21401), .ZN(n16035) );
  AOI22_X1 U17963 ( .A1(n16033), .A2(n16064), .B1(n21366), .B2(n16061), .ZN(
        n16034) );
  NAND2_X1 U17964 ( .A1(n16035), .A2(n16034), .ZN(n21283) );
  AOI21_X1 U17965 ( .B1(n21400), .B2(n16039), .A(n21283), .ZN(n16036) );
  INV_X1 U17966 ( .A(n16036), .ZN(n21386) );
  AOI21_X1 U17967 ( .B1(n16040), .B2(n21400), .A(n21386), .ZN(n16052) );
  OAI21_X1 U17968 ( .B1(n16052), .B2(n16041), .A(n16037), .ZN(n16038) );
  AOI21_X1 U17969 ( .B1(n21549), .B2(n21421), .A(n16038), .ZN(n16044) );
  NOR2_X1 U17970 ( .A1(n16039), .A2(n21281), .ZN(n21385) );
  INV_X1 U17971 ( .A(n16040), .ZN(n16042) );
  NAND3_X1 U17972 ( .A1(n21385), .A2(n16042), .A3(n16041), .ZN(n16043) );
  OAI211_X1 U17973 ( .C1(n16045), .C2(n21382), .A(n16044), .B(n16043), .ZN(
        P1_U3013) );
  AOI21_X1 U17974 ( .B1(n21385), .B2(n16046), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16053) );
  INV_X1 U17975 ( .A(n16047), .ZN(n16049) );
  NOR2_X1 U17976 ( .A1(n21545), .A2(n21414), .ZN(n16048) );
  AOI211_X1 U17977 ( .C1(n21422), .C2(n16050), .A(n16049), .B(n16048), .ZN(
        n16051) );
  OAI21_X1 U17978 ( .B1(n16053), .B2(n16052), .A(n16051), .ZN(P1_U3014) );
  NAND2_X1 U17979 ( .A1(n21386), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16055) );
  OAI211_X1 U17980 ( .C1(n21414), .C2(n16056), .A(n16055), .B(n16054), .ZN(
        n16057) );
  AOI21_X1 U17981 ( .B1(n21385), .B2(n16058), .A(n16057), .ZN(n16059) );
  OAI21_X1 U17982 ( .B1(n16060), .B2(n21382), .A(n16059), .ZN(P1_U3016) );
  INV_X1 U17983 ( .A(n16061), .ZN(n16067) );
  NOR2_X1 U17984 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16062), .ZN(
        n21284) );
  NAND3_X1 U17985 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16063), .A3(
        n16067), .ZN(n16065) );
  AOI211_X1 U17986 ( .C1(n16065), .C2(n21368), .A(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n16064), .ZN(n21285) );
  NOR2_X1 U17987 ( .A1(n21419), .A2(n19861), .ZN(n16066) );
  AOI211_X1 U17988 ( .C1(n16067), .C2(n21284), .A(n21285), .B(n16066), .ZN(
        n16071) );
  INV_X1 U17989 ( .A(n16068), .ZN(n16069) );
  AOI22_X1 U17990 ( .A1(n21283), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n21421), .B2(n16069), .ZN(n16070) );
  OAI211_X1 U17991 ( .C1(n16072), .C2(n21382), .A(n16071), .B(n16070), .ZN(
        P1_U3018) );
  OAI21_X1 U17992 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n16073), .A(n21862), 
        .ZN(n16074) );
  OAI21_X1 U17993 ( .B1(n16075), .B2(n14662), .A(n16074), .ZN(n16076) );
  MUX2_X1 U17994 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n16076), .S(
        n16887), .Z(P1_U3477) );
  INV_X1 U17995 ( .A(n16085), .ZN(n16078) );
  INV_X1 U17996 ( .A(n11421), .ZN(n16077) );
  NAND3_X1 U17997 ( .A1(n16079), .A2(n16078), .A3(n16077), .ZN(n16080) );
  OAI21_X1 U17998 ( .B1(n16081), .B2(n11531), .A(n16080), .ZN(n16082) );
  AOI21_X1 U17999 ( .B1(n21906), .B2(n16083), .A(n16082), .ZN(n16855) );
  INV_X1 U18000 ( .A(n16084), .ZN(n16088) );
  INV_X1 U18001 ( .A(n21658), .ZN(n21643) );
  NOR3_X1 U18002 ( .A1(n11421), .A2(n16085), .A3(n21643), .ZN(n16086) );
  AOI21_X1 U18003 ( .B1(n16088), .B2(n16087), .A(n16086), .ZN(n16089) );
  OAI21_X1 U18004 ( .B1(n16855), .B2(n21645), .A(n16089), .ZN(n16090) );
  MUX2_X1 U18005 ( .A(n11531), .B(n16090), .S(n21647), .Z(P1_U3473) );
  AOI21_X1 U18006 ( .B1(n16092), .B2(n16091), .A(n11058), .ZN(n18424) );
  OAI21_X1 U18007 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n16099), .A(
        n16092), .ZN(n18416) );
  AOI21_X1 U18008 ( .B1(n16426), .B2(n16095), .A(n11039), .ZN(n18357) );
  AOI21_X1 U18009 ( .B1(n16094), .B2(n16093), .A(n16096), .ZN(n18333) );
  NAND2_X1 U18010 ( .A1(n18323), .A2(n17162), .ZN(n18331) );
  NOR2_X1 U18011 ( .A1(n18333), .A2(n18331), .ZN(n18343) );
  OAI21_X1 U18012 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16096), .A(
        n16095), .ZN(n18344) );
  NAND2_X1 U18013 ( .A1(n18343), .A2(n18344), .ZN(n18355) );
  NOR2_X1 U18014 ( .A1(n18357), .A2(n18355), .ZN(n18367) );
  OAI21_X1 U18015 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11039), .A(
        n16097), .ZN(n18369) );
  AOI21_X1 U18016 ( .B1(n16413), .B2(n16097), .A(n16098), .ZN(n18385) );
  NAND2_X1 U18017 ( .A1(n18423), .A2(n18387), .ZN(n18396) );
  OAI21_X1 U18018 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16098), .A(
        n16100), .ZN(n18395) );
  NAND2_X1 U18019 ( .A1(n18423), .A2(n18394), .ZN(n18407) );
  AOI21_X1 U18020 ( .B1(n16390), .B2(n16100), .A(n16099), .ZN(n16393) );
  INV_X1 U18021 ( .A(n16393), .ZN(n18406) );
  NAND2_X1 U18022 ( .A1(n18423), .A2(n18405), .ZN(n18417) );
  NAND2_X1 U18023 ( .A1(n18416), .A2(n18417), .ZN(n18422) );
  NOR2_X1 U18024 ( .A1(n18424), .A2(n18422), .ZN(n18435) );
  OAI21_X1 U18025 ( .B1(n11058), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16102), .ZN(n18438) );
  AOI21_X1 U18026 ( .B1(n18435), .B2(n18438), .A(n18436), .ZN(n18452) );
  NAND2_X1 U18027 ( .A1(n16102), .A2(n16101), .ZN(n16103) );
  AND2_X1 U18028 ( .A1(n16104), .A2(n16103), .ZN(n18451) );
  NAND2_X1 U18029 ( .A1(n18423), .A2(n18454), .ZN(n18465) );
  INV_X1 U18030 ( .A(n16104), .ZN(n16106) );
  OAI21_X1 U18031 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16106), .A(
        n16105), .ZN(n18464) );
  NAND2_X1 U18032 ( .A1(n18423), .A2(n18463), .ZN(n18484) );
  INV_X1 U18033 ( .A(n16107), .ZN(n18483) );
  NAND2_X1 U18034 ( .A1(n18423), .A2(n18481), .ZN(n16109) );
  OAI211_X1 U18035 ( .C1(n16109), .C2(n16108), .A(n18482), .B(n18506), .ZN(
        n16119) );
  INV_X1 U18036 ( .A(n16110), .ZN(n16117) );
  OAI22_X1 U18037 ( .A1(n18490), .A2(n16112), .B1(n16111), .B2(n18329), .ZN(
        n16116) );
  INV_X1 U18038 ( .A(n16113), .ZN(n16114) );
  OAI22_X1 U18039 ( .A1(n16114), .A2(n18476), .B1(n17283), .B2(n18493), .ZN(
        n16115) );
  AOI211_X1 U18040 ( .C1(n16117), .C2(n18501), .A(n16116), .B(n16115), .ZN(
        n16118) );
  OAI211_X1 U18041 ( .C1(n16120), .C2(n18494), .A(n16119), .B(n16118), .ZN(
        P2_U2825) );
  INV_X1 U18042 ( .A(n16121), .ZN(n16125) );
  INV_X1 U18043 ( .A(n16122), .ZN(n16451) );
  NOR2_X1 U18044 ( .A1(n16123), .A2(n18505), .ZN(n16124) );
  OAI21_X1 U18045 ( .B1(n16125), .B2(n16451), .A(n16124), .ZN(n16134) );
  XOR2_X1 U18046 ( .A(n11036), .B(n16126), .Z(n19086) );
  NOR2_X1 U18047 ( .A1(n18423), .A2(n18602), .ZN(n18321) );
  INV_X1 U18048 ( .A(n18321), .ZN(n18313) );
  AOI22_X1 U18049 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18498), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n18473), .ZN(n16127) );
  OAI211_X1 U18050 ( .C1(n16451), .C2(n18313), .A(n16127), .B(n14141), .ZN(
        n16130) );
  NOR2_X1 U18051 ( .A1(n18490), .A2(n16128), .ZN(n16129) );
  AOI211_X1 U18052 ( .C1(n18500), .C2(n19086), .A(n16130), .B(n16129), .ZN(
        n16131) );
  OAI21_X1 U18053 ( .B1(n16684), .B2(n18478), .A(n16131), .ZN(n16132) );
  INV_X1 U18054 ( .A(n16132), .ZN(n16133) );
  OAI211_X1 U18055 ( .C1(n16135), .C2(n18494), .A(n16134), .B(n16133), .ZN(
        P2_U2842) );
  AOI21_X1 U18056 ( .B1(n16689), .B2(n16136), .A(n11036), .ZN(n18524) );
  INV_X1 U18057 ( .A(n18524), .ZN(n19092) );
  NOR2_X1 U18058 ( .A1(n18436), .A2(n16137), .ZN(n18308) );
  XNOR2_X1 U18059 ( .A(n18308), .B(n17145), .ZN(n16138) );
  NAND2_X1 U18060 ( .A1(n16138), .A2(n18482), .ZN(n16148) );
  INV_X1 U18061 ( .A(n16139), .ZN(n18526) );
  NOR2_X1 U18062 ( .A1(n18490), .A2(n16140), .ZN(n16141) );
  AOI211_X1 U18063 ( .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n18474), .A(
        n18559), .B(n16141), .ZN(n16142) );
  OAI21_X1 U18064 ( .B1(n16143), .B2(n18493), .A(n16142), .ZN(n16146) );
  NOR2_X1 U18065 ( .A1(n16144), .A2(n18494), .ZN(n16145) );
  AOI211_X1 U18066 ( .C1(n18501), .C2(n18526), .A(n16146), .B(n16145), .ZN(
        n16147) );
  OAI211_X1 U18067 ( .C1(n18476), .C2(n19092), .A(n16148), .B(n16147), .ZN(
        P2_U2843) );
  NOR2_X1 U18068 ( .A1(n18436), .A2(n16149), .ZN(n16162) );
  XNOR2_X1 U18069 ( .A(n16162), .B(n16150), .ZN(n16151) );
  NAND2_X1 U18070 ( .A1(n16151), .A2(n18482), .ZN(n16161) );
  OAI22_X1 U18071 ( .A1(n18490), .A2(n13879), .B1(n16152), .B2(n18329), .ZN(
        n16153) );
  INV_X1 U18072 ( .A(n16153), .ZN(n16155) );
  NAND2_X1 U18073 ( .A1(n18473), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n16154) );
  OAI211_X1 U18074 ( .C1(n18494), .C2(n16156), .A(n16155), .B(n16154), .ZN(
        n16159) );
  NOR2_X1 U18075 ( .A1(n16157), .A2(n18478), .ZN(n16158) );
  AOI211_X1 U18076 ( .C1(n18500), .C2(n19523), .A(n16159), .B(n16158), .ZN(
        n16160) );
  OAI211_X1 U18077 ( .C1(n18241), .C2(n19238), .A(n16161), .B(n16160), .ZN(
        P2_U2853) );
  OAI21_X1 U18078 ( .B1(n18247), .B2(n16163), .A(n16162), .ZN(n16788) );
  OAI22_X1 U18079 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18313), .B1(
        n16788), .B2(n18602), .ZN(n16164) );
  INV_X1 U18080 ( .A(n16164), .ZN(n16172) );
  INV_X1 U18081 ( .A(n16165), .ZN(n16168) );
  AOI22_X1 U18082 ( .A1(n18473), .A2(P2_REIP_REG_1__SCAN_IN), .B1(n18500), 
        .B2(n19575), .ZN(n16167) );
  AOI22_X1 U18083 ( .A1(n18470), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18474), .ZN(n16166) );
  OAI211_X1 U18084 ( .C1(n18494), .C2(n16168), .A(n16167), .B(n16166), .ZN(
        n16169) );
  AOI21_X1 U18085 ( .B1(n16170), .B2(n18501), .A(n16169), .ZN(n16171) );
  OAI211_X1 U18086 ( .C1(n19142), .C2(n18241), .A(n16172), .B(n16171), .ZN(
        P2_U2854) );
  NAND2_X1 U18087 ( .A1(n18502), .A2(n11059), .ZN(n16173) );
  OAI21_X1 U18088 ( .B1(n11059), .B2(n18489), .A(n16173), .ZN(P2_U2856) );
  XNOR2_X1 U18089 ( .A(n16176), .B(n16175), .ZN(n16177) );
  XNOR2_X1 U18090 ( .A(n16174), .B(n16177), .ZN(n16274) );
  NOR2_X1 U18091 ( .A1(n18479), .A2(n10963), .ZN(n16178) );
  AOI21_X1 U18092 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n10963), .A(n16178), .ZN(
        n16179) );
  OAI21_X1 U18093 ( .B1(n16274), .B2(n16253), .A(n16179), .ZN(P2_U2858) );
  AOI21_X1 U18094 ( .B1(n16180), .B2(n16195), .A(n11007), .ZN(n18462) );
  INV_X1 U18095 ( .A(n18462), .ZN(n16186) );
  NOR2_X1 U18096 ( .A1(n16187), .A2(n16181), .ZN(n16183) );
  XNOR2_X1 U18097 ( .A(n16183), .B(n16182), .ZN(n16275) );
  NAND2_X1 U18098 ( .A1(n16275), .A2(n16266), .ZN(n16185) );
  NAND2_X1 U18099 ( .A1(n10963), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16184) );
  OAI211_X1 U18100 ( .C1(n10963), .C2(n16186), .A(n16185), .B(n16184), .ZN(
        P2_U2859) );
  INV_X1 U18101 ( .A(n16187), .ZN(n16189) );
  NAND2_X1 U18102 ( .A1(n16189), .A2(n16188), .ZN(n16190) );
  XOR2_X1 U18103 ( .A(n16191), .B(n16190), .Z(n16292) );
  NAND2_X1 U18104 ( .A1(n16192), .A2(n16193), .ZN(n16194) );
  NAND2_X1 U18105 ( .A1(n16195), .A2(n16194), .ZN(n16514) );
  NOR2_X1 U18106 ( .A1(n16514), .A2(n10963), .ZN(n16196) );
  AOI21_X1 U18107 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n10963), .A(n16196), .ZN(
        n16197) );
  OAI21_X1 U18108 ( .B1(n16292), .B2(n16253), .A(n16197), .ZN(P2_U2860) );
  OR2_X1 U18109 ( .A1(n16198), .A2(n16199), .ZN(n16200) );
  NAND2_X1 U18110 ( .A1(n16192), .A2(n16200), .ZN(n18442) );
  AOI21_X1 U18111 ( .B1(n16203), .B2(n16202), .A(n16201), .ZN(n16299) );
  NAND2_X1 U18112 ( .A1(n16299), .A2(n16266), .ZN(n16205) );
  NAND2_X1 U18113 ( .A1(n10963), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16204) );
  OAI211_X1 U18114 ( .C1(n18442), .C2(n10963), .A(n16205), .B(n16204), .ZN(
        P2_U2861) );
  INV_X1 U18115 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16215) );
  OAI21_X1 U18116 ( .B1(n16208), .B2(n16207), .A(n16206), .ZN(n16307) );
  OR2_X1 U18117 ( .A1(n16307), .A2(n16253), .ZN(n16214) );
  AND2_X1 U18118 ( .A1(n16209), .A2(n16210), .ZN(n16211) );
  OR2_X1 U18119 ( .A1(n16211), .A2(n16198), .ZN(n18430) );
  INV_X1 U18120 ( .A(n18430), .ZN(n16212) );
  NAND2_X1 U18121 ( .A1(n16212), .A2(n11059), .ZN(n16213) );
  OAI211_X1 U18122 ( .C1(n11059), .C2(n16215), .A(n16214), .B(n16213), .ZN(
        P2_U2862) );
  NAND2_X1 U18123 ( .A1(n16227), .A2(n16217), .ZN(n16218) );
  NAND2_X1 U18124 ( .A1(n16209), .A2(n16218), .ZN(n18413) );
  AOI21_X1 U18125 ( .B1(n16220), .B2(n16219), .A(n11018), .ZN(n16312) );
  NAND2_X1 U18126 ( .A1(n16312), .A2(n16266), .ZN(n16222) );
  NAND2_X1 U18127 ( .A1(n10963), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16221) );
  OAI211_X1 U18128 ( .C1(n18413), .C2(n10963), .A(n16222), .B(n16221), .ZN(
        P2_U2863) );
  XNOR2_X1 U18129 ( .A(n16234), .B(n16224), .ZN(n16320) );
  NAND2_X1 U18130 ( .A1(n16233), .A2(n16225), .ZN(n16226) );
  NAND2_X1 U18131 ( .A1(n16227), .A2(n16226), .ZN(n18402) );
  NOR2_X1 U18132 ( .A1(n10963), .A2(n18402), .ZN(n16228) );
  AOI21_X1 U18133 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n10963), .A(n16228), .ZN(
        n16229) );
  OAI21_X1 U18134 ( .B1(n16320), .B2(n16253), .A(n16229), .ZN(P2_U2864) );
  OR2_X1 U18135 ( .A1(n16231), .A2(n16230), .ZN(n16232) );
  AND2_X1 U18136 ( .A1(n16233), .A2(n16232), .ZN(n18393) );
  INV_X1 U18137 ( .A(n18393), .ZN(n16579) );
  AOI21_X1 U18138 ( .B1(n16235), .B2(n16238), .A(n16234), .ZN(n19323) );
  NAND2_X1 U18139 ( .A1(n19323), .A2(n16266), .ZN(n16237) );
  NAND2_X1 U18140 ( .A1(n10963), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16236) );
  OAI211_X1 U18141 ( .C1(n16579), .C2(n10963), .A(n16237), .B(n16236), .ZN(
        P2_U2865) );
  OAI21_X1 U18142 ( .B1(n16246), .B2(n16239), .A(n16238), .ZN(n16327) );
  AOI21_X1 U18143 ( .B1(n16240), .B2(n16249), .A(n16230), .ZN(n18386) );
  INV_X1 U18144 ( .A(n18386), .ZN(n16591) );
  NOR2_X1 U18145 ( .A1(n16591), .A2(n10963), .ZN(n16241) );
  AOI21_X1 U18146 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n10963), .A(n16241), .ZN(
        n16242) );
  OAI21_X1 U18147 ( .B1(n16327), .B2(n16253), .A(n16242), .ZN(P2_U2866) );
  NOR2_X1 U18148 ( .A1(n16243), .A2(n16244), .ZN(n16245) );
  OR2_X1 U18149 ( .A1(n16246), .A2(n16245), .ZN(n19423) );
  OR2_X1 U18150 ( .A1(n16248), .A2(n16247), .ZN(n16250) );
  AND2_X1 U18151 ( .A1(n16250), .A2(n16249), .ZN(n18533) );
  NAND2_X1 U18152 ( .A1(n11059), .A2(n18533), .ZN(n16252) );
  NAND2_X1 U18153 ( .A1(n10963), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n16251) );
  OAI211_X1 U18154 ( .C1(n19423), .C2(n16253), .A(n16252), .B(n16251), .ZN(
        P2_U2867) );
  AOI21_X1 U18155 ( .B1(n16254), .B2(n10984), .A(n16247), .ZN(n18363) );
  INV_X1 U18156 ( .A(n18363), .ZN(n16259) );
  INV_X1 U18157 ( .A(n16255), .ZN(n16263) );
  AOI21_X1 U18158 ( .B1(n16256), .B2(n16263), .A(n16243), .ZN(n16332) );
  NAND2_X1 U18159 ( .A1(n16332), .A2(n16266), .ZN(n16258) );
  NAND2_X1 U18160 ( .A1(n10963), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n16257) );
  OAI211_X1 U18161 ( .C1(n16259), .C2(n10963), .A(n16258), .B(n16257), .ZN(
        P2_U2868) );
  OR2_X1 U18162 ( .A1(n16261), .A2(n16260), .ZN(n16262) );
  AND2_X1 U18163 ( .A1(n16262), .A2(n10984), .ZN(n18548) );
  INV_X1 U18164 ( .A(n18548), .ZN(n16269) );
  AOI21_X1 U18165 ( .B1(n16265), .B2(n16264), .A(n16255), .ZN(n19519) );
  NAND2_X1 U18166 ( .A1(n19519), .A2(n16266), .ZN(n16268) );
  NAND2_X1 U18167 ( .A1(n10963), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n16267) );
  OAI211_X1 U18168 ( .C1(n16269), .C2(n10963), .A(n16268), .B(n16267), .ZN(
        P2_U2869) );
  AOI22_X1 U18169 ( .A1(n19630), .A2(BUF2_REG_29__SCAN_IN), .B1(n19631), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n16271) );
  XNOR2_X1 U18170 ( .A(n16278), .B(n11069), .ZN(n18475) );
  AOI22_X1 U18171 ( .A1(n19633), .A2(n18475), .B1(n19627), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n16270) );
  OAI211_X1 U18172 ( .C1(n19087), .C2(n16337), .A(n16271), .B(n16270), .ZN(
        n16272) );
  INV_X1 U18173 ( .A(n16272), .ZN(n16273) );
  OAI21_X1 U18174 ( .B1(n16274), .B2(n19579), .A(n16273), .ZN(P2_U2890) );
  NAND2_X1 U18175 ( .A1(n16275), .A2(n19634), .ZN(n16282) );
  AND2_X1 U18176 ( .A1(n16286), .A2(n16276), .ZN(n16277) );
  NOR2_X1 U18177 ( .A1(n16278), .A2(n16277), .ZN(n18461) );
  AOI22_X1 U18178 ( .A1(n19633), .A2(n18461), .B1(n19627), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16281) );
  AOI22_X1 U18179 ( .A1(n19630), .A2(BUF2_REG_28__SCAN_IN), .B1(n19631), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n16280) );
  INV_X1 U18180 ( .A(n16337), .ZN(n19629) );
  NAND2_X1 U18181 ( .A1(n19629), .A2(n19090), .ZN(n16279) );
  NAND4_X1 U18182 ( .A1(n16282), .A2(n16281), .A3(n16280), .A4(n16279), .ZN(
        P2_U2891) );
  AOI22_X1 U18183 ( .A1(n19630), .A2(BUF2_REG_27__SCAN_IN), .B1(n19631), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n16289) );
  NAND2_X1 U18184 ( .A1(n16284), .A2(n16283), .ZN(n16285) );
  NAND2_X1 U18185 ( .A1(n16286), .A2(n16285), .ZN(n18458) );
  INV_X1 U18186 ( .A(n18458), .ZN(n16287) );
  AOI22_X1 U18187 ( .A1(n19633), .A2(n16287), .B1(n19627), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16288) );
  OAI211_X1 U18188 ( .C1(n19093), .C2(n16337), .A(n16289), .B(n16288), .ZN(
        n16290) );
  INV_X1 U18189 ( .A(n16290), .ZN(n16291) );
  OAI21_X1 U18190 ( .B1(n16292), .B2(n19579), .A(n16291), .ZN(P2_U2892) );
  AOI22_X1 U18191 ( .A1(n19630), .A2(BUF2_REG_26__SCAN_IN), .B1(n19631), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n16297) );
  INV_X1 U18192 ( .A(n16294), .ZN(n16295) );
  XNOR2_X1 U18193 ( .A(n16293), .B(n16295), .ZN(n18439) );
  AOI22_X1 U18194 ( .A1(n19633), .A2(n18439), .B1(n19627), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16296) );
  OAI211_X1 U18195 ( .C1(n19096), .C2(n16337), .A(n16297), .B(n16296), .ZN(
        n16298) );
  AOI21_X1 U18196 ( .B1(n16299), .B2(n19634), .A(n16298), .ZN(n16300) );
  INV_X1 U18197 ( .A(n16300), .ZN(P2_U2893) );
  AOI22_X1 U18198 ( .A1(n19630), .A2(BUF2_REG_25__SCAN_IN), .B1(n19631), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n16304) );
  AND2_X1 U18199 ( .A1(n11005), .A2(n16301), .ZN(n16302) );
  NOR2_X1 U18200 ( .A1(n16293), .A2(n16302), .ZN(n18428) );
  AOI22_X1 U18201 ( .A1(n19633), .A2(n18428), .B1(n19627), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16303) );
  OAI211_X1 U18202 ( .C1(n19099), .C2(n16337), .A(n16304), .B(n16303), .ZN(
        n16305) );
  INV_X1 U18203 ( .A(n16305), .ZN(n16306) );
  OAI21_X1 U18204 ( .B1(n16307), .B2(n19579), .A(n16306), .ZN(P2_U2894) );
  AOI22_X1 U18205 ( .A1(n19630), .A2(BUF2_REG_24__SCAN_IN), .B1(n19631), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n16310) );
  XNOR2_X1 U18206 ( .A(n16308), .B(n10987), .ZN(n18414) );
  AOI22_X1 U18207 ( .A1(n19633), .A2(n18414), .B1(n19627), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16309) );
  OAI211_X1 U18208 ( .C1(n19103), .C2(n16337), .A(n16310), .B(n16309), .ZN(
        n16311) );
  AOI21_X1 U18209 ( .B1(n16312), .B2(n19634), .A(n16311), .ZN(n16313) );
  INV_X1 U18210 ( .A(n16313), .ZN(P2_U2895) );
  AOI22_X1 U18211 ( .A1(n19630), .A2(BUF2_REG_23__SCAN_IN), .B1(n19631), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16317) );
  OAI21_X1 U18212 ( .B1(n16315), .B2(n16314), .A(n10987), .ZN(n16558) );
  INV_X1 U18213 ( .A(n16558), .ZN(n18403) );
  AOI22_X1 U18214 ( .A1(n19633), .A2(n18403), .B1(n19627), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16316) );
  OAI211_X1 U18215 ( .C1(n19113), .C2(n16337), .A(n16317), .B(n16316), .ZN(
        n16318) );
  INV_X1 U18216 ( .A(n16318), .ZN(n16319) );
  OAI21_X1 U18217 ( .B1(n16320), .B2(n19579), .A(n16319), .ZN(P2_U2896) );
  AOI22_X1 U18218 ( .A1(n19630), .A2(BUF2_REG_21__SCAN_IN), .B1(n19631), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n16324) );
  OAI21_X1 U18219 ( .B1(n16321), .B2(n18370), .A(n16576), .ZN(n18391) );
  INV_X1 U18220 ( .A(n18391), .ZN(n16322) );
  AOI22_X1 U18221 ( .A1(n19633), .A2(n16322), .B1(n19627), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16323) );
  OAI211_X1 U18222 ( .C1(n19379), .C2(n16337), .A(n16324), .B(n16323), .ZN(
        n16325) );
  INV_X1 U18223 ( .A(n16325), .ZN(n16326) );
  OAI21_X1 U18224 ( .B1(n16327), .B2(n19579), .A(n16326), .ZN(P2_U2898) );
  AOI22_X1 U18225 ( .A1(n19630), .A2(BUF2_REG_19__SCAN_IN), .B1(n19631), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n16330) );
  OAI21_X1 U18226 ( .B1(n16328), .B2(n18350), .A(n11006), .ZN(n16605) );
  INV_X1 U18227 ( .A(n16605), .ZN(n18362) );
  AOI22_X1 U18228 ( .A1(n19633), .A2(n18362), .B1(n19627), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16329) );
  OAI211_X1 U18229 ( .C1(n19477), .C2(n16337), .A(n16330), .B(n16329), .ZN(
        n16331) );
  AOI21_X1 U18230 ( .B1(n16332), .B2(n19634), .A(n16331), .ZN(n16333) );
  INV_X1 U18231 ( .A(n16333), .ZN(P2_U2900) );
  AOI22_X1 U18232 ( .A1(n19630), .A2(BUF2_REG_17__SCAN_IN), .B1(n19631), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n16336) );
  OAI21_X1 U18233 ( .B1(n16334), .B2(n15191), .A(n11044), .ZN(n16628) );
  INV_X1 U18234 ( .A(n16628), .ZN(n18338) );
  AOI22_X1 U18235 ( .A1(n19633), .A2(n18338), .B1(n19627), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16335) );
  OAI211_X1 U18236 ( .C1(n19584), .C2(n16337), .A(n16336), .B(n16335), .ZN(
        n16338) );
  INV_X1 U18237 ( .A(n16338), .ZN(n16339) );
  OAI21_X1 U18238 ( .B1(n16340), .B2(n19579), .A(n16339), .ZN(P2_U2902) );
  OAI21_X1 U18239 ( .B1(n16347), .B2(n17156), .A(n16346), .ZN(P2_U2983) );
  NAND2_X1 U18240 ( .A1(n16350), .A2(n16349), .ZN(n16360) );
  OAI21_X1 U18241 ( .B1(n16362), .B2(n16493), .A(n16360), .ZN(n16353) );
  XNOR2_X1 U18242 ( .A(n16351), .B(n16508), .ZN(n16352) );
  XNOR2_X1 U18243 ( .A(n16353), .B(n16352), .ZN(n16513) );
  XNOR2_X1 U18244 ( .A(n16354), .B(n16508), .ZN(n16511) );
  NAND2_X1 U18245 ( .A1(n18559), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n16503) );
  OAI21_X1 U18246 ( .B1(n17151), .B2(n16355), .A(n16503), .ZN(n16356) );
  AOI21_X1 U18247 ( .B1(n18462), .B2(n17190), .A(n16356), .ZN(n16357) );
  OAI21_X1 U18248 ( .B1(n18464), .B2(n17198), .A(n16357), .ZN(n16358) );
  AOI21_X1 U18249 ( .B1(n16511), .B2(n17203), .A(n16358), .ZN(n16359) );
  OAI21_X1 U18250 ( .B1(n16513), .B2(n17156), .A(n16359), .ZN(P2_U2986) );
  INV_X1 U18251 ( .A(n16360), .ZN(n16361) );
  NOR2_X1 U18252 ( .A1(n16362), .A2(n16361), .ZN(n16363) );
  XNOR2_X1 U18253 ( .A(n16363), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16524) );
  NOR2_X1 U18254 ( .A1(n18521), .A2(n18448), .ZN(n16515) );
  AOI21_X1 U18255 ( .B1(n17200), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16515), .ZN(n16364) );
  OAI21_X1 U18256 ( .B1(n16514), .B2(n17207), .A(n16364), .ZN(n16365) );
  AOI21_X1 U18257 ( .B1(n18451), .B2(n17163), .A(n16365), .ZN(n16367) );
  NAND2_X1 U18258 ( .A1(n15493), .A2(n16493), .ZN(n16520) );
  NAND3_X1 U18259 ( .A1(n16521), .A2(n17203), .A3(n16520), .ZN(n16366) );
  OAI211_X1 U18260 ( .C1(n16524), .C2(n17156), .A(n16367), .B(n16366), .ZN(
        P2_U2987) );
  INV_X1 U18261 ( .A(n16368), .ZN(n16373) );
  NAND2_X1 U18262 ( .A1(n16369), .A2(n16381), .ZN(n16371) );
  MUX2_X1 U18263 ( .A(n16381), .B(n16371), .S(n16370), .Z(n16372) );
  NAND2_X1 U18264 ( .A1(n16373), .A2(n16372), .ZN(n16535) );
  INV_X1 U18265 ( .A(n15493), .ZN(n16376) );
  AOI21_X1 U18266 ( .B1(n16374), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16375) );
  NOR2_X1 U18267 ( .A1(n16376), .A2(n16375), .ZN(n16533) );
  NOR2_X1 U18268 ( .A1(n18521), .A2(n17280), .ZN(n16527) );
  NOR2_X1 U18269 ( .A1(n18442), .A2(n17207), .ZN(n16377) );
  AOI211_X1 U18270 ( .C1(n17200), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16527), .B(n16377), .ZN(n16378) );
  OAI21_X1 U18271 ( .B1(n18438), .B2(n17198), .A(n16378), .ZN(n16379) );
  AOI21_X1 U18272 ( .B1(n16533), .B2(n17203), .A(n16379), .ZN(n16380) );
  OAI21_X1 U18273 ( .B1(n16535), .B2(n17156), .A(n16380), .ZN(P2_U2988) );
  INV_X1 U18274 ( .A(n16381), .ZN(n16382) );
  NOR2_X1 U18275 ( .A1(n16383), .A2(n16382), .ZN(n16385) );
  XOR2_X1 U18276 ( .A(n16385), .B(n16384), .Z(n16546) );
  XOR2_X1 U18277 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n16374), .Z(
        n16544) );
  NAND2_X1 U18278 ( .A1(n18424), .A2(n17163), .ZN(n16387) );
  NOR2_X1 U18279 ( .A1(n18521), .A2(n17279), .ZN(n16540) );
  AOI21_X1 U18280 ( .B1(n17200), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16540), .ZN(n16386) );
  OAI211_X1 U18281 ( .C1(n17207), .C2(n18430), .A(n16387), .B(n16386), .ZN(
        n16388) );
  AOI21_X1 U18282 ( .B1(n16544), .B2(n17203), .A(n16388), .ZN(n16389) );
  OAI21_X1 U18283 ( .B1(n16546), .B2(n17156), .A(n16389), .ZN(P2_U2989) );
  AND2_X1 U18284 ( .A1(n16567), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17193) );
  OAI21_X1 U18285 ( .B1(n17193), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16549), .ZN(n16566) );
  OAI22_X1 U18286 ( .A1(n16390), .A2(n17151), .B1(n17278), .B2(n18521), .ZN(
        n16392) );
  NOR2_X1 U18287 ( .A1(n17207), .A2(n18402), .ZN(n16391) );
  AOI211_X1 U18288 ( .C1(n16393), .C2(n17163), .A(n16392), .B(n16391), .ZN(
        n16398) );
  XNOR2_X1 U18289 ( .A(n16394), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16395) );
  XNOR2_X1 U18290 ( .A(n16396), .B(n16395), .ZN(n16563) );
  NAND2_X1 U18291 ( .A1(n16563), .A2(n17202), .ZN(n16397) );
  OAI211_X1 U18292 ( .C1(n16566), .C2(n17152), .A(n16398), .B(n16397), .ZN(
        P2_U2991) );
  INV_X1 U18293 ( .A(n16399), .ZN(n16401) );
  NAND2_X1 U18294 ( .A1(n16633), .A2(n16634), .ZN(n16635) );
  INV_X1 U18295 ( .A(n16613), .ZN(n16402) );
  NOR2_X1 U18296 ( .A1(n16407), .A2(n16406), .ZN(n16408) );
  NOR2_X1 U18297 ( .A1(n16408), .A2(n17183), .ZN(n16412) );
  NAND2_X1 U18298 ( .A1(n16410), .A2(n16409), .ZN(n16411) );
  XNOR2_X1 U18299 ( .A(n16412), .B(n16411), .ZN(n16595) );
  OAI22_X1 U18300 ( .A1(n16413), .A2(n17151), .B1(n17277), .B2(n18521), .ZN(
        n16415) );
  NOR2_X1 U18301 ( .A1(n16591), .A2(n17207), .ZN(n16414) );
  AOI211_X1 U18302 ( .C1(n18385), .C2(n17163), .A(n16415), .B(n16414), .ZN(
        n16418) );
  NAND2_X1 U18303 ( .A1(n16416), .A2(n16587), .ZN(n17184) );
  AOI21_X1 U18304 ( .B1(n16588), .B2(n17184), .A(n16567), .ZN(n16593) );
  NAND2_X1 U18305 ( .A1(n16593), .A2(n17203), .ZN(n16417) );
  OAI211_X1 U18306 ( .C1(n16595), .C2(n17156), .A(n16418), .B(n16417), .ZN(
        P2_U2993) );
  NOR2_X1 U18307 ( .A1(n16420), .A2(n16419), .ZN(n16424) );
  INV_X1 U18308 ( .A(n17176), .ZN(n16422) );
  AOI21_X1 U18309 ( .B1(n17175), .B2(n16422), .A(n16421), .ZN(n16423) );
  XNOR2_X1 U18310 ( .A(n16424), .B(n16423), .ZN(n16610) );
  NAND2_X1 U18311 ( .A1(n16416), .A2(n16598), .ZN(n17178) );
  NAND3_X1 U18312 ( .A1(n16416), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16598), .ZN(n17186) );
  INV_X1 U18313 ( .A(n17186), .ZN(n16425) );
  AOI21_X1 U18314 ( .B1(n18539), .B2(n17178), .A(n16425), .ZN(n16607) );
  INV_X1 U18315 ( .A(n18357), .ZN(n16429) );
  OAI22_X1 U18316 ( .A1(n16426), .A2(n17151), .B1(n17276), .B2(n14141), .ZN(
        n16427) );
  AOI21_X1 U18317 ( .B1(n17190), .B2(n18363), .A(n16427), .ZN(n16428) );
  OAI21_X1 U18318 ( .B1(n17198), .B2(n16429), .A(n16428), .ZN(n16430) );
  AOI21_X1 U18319 ( .B1(n16607), .B2(n17203), .A(n16430), .ZN(n16431) );
  OAI21_X1 U18320 ( .B1(n16610), .B2(n17156), .A(n16431), .ZN(P2_U2995) );
  NAND2_X1 U18321 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16692) );
  NOR2_X1 U18322 ( .A1(n17142), .A2(n16432), .ZN(n16445) );
  INV_X1 U18323 ( .A(n16654), .ZN(n16433) );
  NAND2_X1 U18324 ( .A1(n16416), .A2(n16433), .ZN(n16662) );
  OAI21_X1 U18325 ( .B1(n16445), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16662), .ZN(n16677) );
  AND2_X1 U18326 ( .A1(n16434), .A2(n16435), .ZN(n16449) );
  NAND2_X1 U18327 ( .A1(n16450), .A2(n16449), .ZN(n16448) );
  NAND2_X1 U18328 ( .A1(n16448), .A2(n16435), .ZN(n16438) );
  AND2_X1 U18329 ( .A1(n16645), .A2(n16436), .ZN(n16437) );
  NAND2_X1 U18330 ( .A1(n16438), .A2(n16437), .ZN(n16644) );
  OAI21_X1 U18331 ( .B1(n16438), .B2(n16437), .A(n16644), .ZN(n16675) );
  NAND2_X1 U18332 ( .A1(n16439), .A2(n17190), .ZN(n16441) );
  NOR2_X1 U18333 ( .A1(n14141), .A2(n17274), .ZN(n16669) );
  AOI21_X1 U18334 ( .B1(n17200), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16669), .ZN(n16440) );
  OAI211_X1 U18335 ( .C1(n16442), .C2(n17198), .A(n16441), .B(n16440), .ZN(
        n16443) );
  AOI21_X1 U18336 ( .B1(n16675), .B2(n17202), .A(n16443), .ZN(n16444) );
  OAI21_X1 U18337 ( .B1(n16677), .B2(n17152), .A(n16444), .ZN(P2_U3000) );
  INV_X1 U18338 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18530) );
  NOR2_X1 U18339 ( .A1(n17142), .A2(n18530), .ZN(n16447) );
  INV_X1 U18340 ( .A(n16445), .ZN(n16446) );
  OAI21_X1 U18341 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16447), .A(
        n16446), .ZN(n16688) );
  OAI21_X1 U18342 ( .B1(n16450), .B2(n16449), .A(n16448), .ZN(n16686) );
  OAI22_X1 U18343 ( .A1(n16452), .A2(n17151), .B1(n17198), .B2(n16451), .ZN(
        n16455) );
  OAI22_X1 U18344 ( .A1(n17207), .A2(n16684), .B1(n18521), .B2(n16453), .ZN(
        n16454) );
  AOI211_X1 U18345 ( .C1(n16686), .C2(n17202), .A(n16455), .B(n16454), .ZN(
        n16456) );
  OAI21_X1 U18346 ( .B1(n16688), .B2(n17152), .A(n16456), .ZN(P2_U3001) );
  OAI21_X1 U18347 ( .B1(n16704), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17142), .ZN(n16703) );
  NOR2_X1 U18348 ( .A1(n14141), .A2(n16457), .ZN(n16693) );
  INV_X1 U18349 ( .A(n16458), .ZN(n18312) );
  OAI22_X1 U18350 ( .A1(n18297), .A2(n17151), .B1(n17198), .B2(n18312), .ZN(
        n16459) );
  AOI211_X1 U18351 ( .C1(n17190), .C2(n18301), .A(n16693), .B(n16459), .ZN(
        n16469) );
  INV_X1 U18352 ( .A(n16460), .ZN(n16472) );
  NAND2_X1 U18353 ( .A1(n16472), .A2(n16470), .ZN(n16712) );
  INV_X1 U18354 ( .A(n16712), .ZN(n16462) );
  AOI21_X1 U18355 ( .B1(n16462), .B2(n16714), .A(n16461), .ZN(n16467) );
  INV_X1 U18356 ( .A(n16463), .ZN(n16465) );
  NOR2_X1 U18357 ( .A1(n16465), .A2(n16464), .ZN(n16466) );
  XNOR2_X1 U18358 ( .A(n16467), .B(n16466), .ZN(n16700) );
  NAND2_X1 U18359 ( .A1(n16700), .A2(n17202), .ZN(n16468) );
  OAI211_X1 U18360 ( .C1(n16703), .C2(n17152), .A(n16469), .B(n16468), .ZN(
        P2_U3003) );
  INV_X1 U18361 ( .A(n16711), .ZN(n16473) );
  AND2_X1 U18362 ( .A1(n16711), .A2(n16470), .ZN(n16471) );
  OAI22_X1 U18363 ( .A1(n16712), .A2(n16473), .B1(n16472), .B2(n16471), .ZN(
        n16735) );
  NAND2_X1 U18364 ( .A1(n17167), .A2(n16730), .ZN(n16722) );
  NAND2_X1 U18365 ( .A1(n16416), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16721) );
  NAND3_X1 U18366 ( .A1(n16722), .A2(n17203), .A3(n16721), .ZN(n16479) );
  INV_X1 U18367 ( .A(n18281), .ZN(n16474) );
  OAI22_X1 U18368 ( .A1(n18275), .A2(n17151), .B1(n17198), .B2(n16474), .ZN(
        n16477) );
  NOR2_X1 U18369 ( .A1(n16475), .A2(n17207), .ZN(n16476) );
  AOI211_X1 U18370 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n18559), .A(n16477), .B(
        n16476), .ZN(n16478) );
  OAI211_X1 U18371 ( .C1(n17156), .C2(n16735), .A(n16479), .B(n16478), .ZN(
        P2_U3005) );
  NAND2_X1 U18372 ( .A1(n17123), .A2(n17125), .ZN(n16481) );
  XOR2_X1 U18373 ( .A(n16481), .B(n16480), .Z(n16751) );
  OR2_X1 U18374 ( .A1(n16483), .A2(n16482), .ZN(n16736) );
  NAND3_X1 U18375 ( .A1(n16736), .A2(n17203), .A3(n16484), .ZN(n16489) );
  OAI22_X1 U18376 ( .A1(n16485), .A2(n17151), .B1(n18265), .B2(n18521), .ZN(
        n16487) );
  NOR2_X1 U18377 ( .A1(n18269), .A2(n17207), .ZN(n16486) );
  AOI211_X1 U18378 ( .C1(n17163), .C2(n18261), .A(n16487), .B(n16486), .ZN(
        n16488) );
  OAI211_X1 U18379 ( .C1(n16751), .C2(n17156), .A(n16489), .B(n16488), .ZN(
        P2_U3007) );
  INV_X1 U18380 ( .A(n16490), .ZN(n16500) );
  NOR2_X1 U18381 ( .A1(n16492), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16517) );
  NOR2_X1 U18382 ( .A1(n16517), .A2(n16519), .ZN(n16509) );
  NOR2_X1 U18383 ( .A1(n16509), .A2(n16491), .ZN(n16499) );
  XNOR2_X1 U18384 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16494) );
  OR2_X1 U18385 ( .A1(n16493), .A2(n16492), .ZN(n16505) );
  NOR2_X1 U18386 ( .A1(n16494), .A2(n16505), .ZN(n16495) );
  AOI211_X1 U18387 ( .C1(n18553), .C2(n18475), .A(n16496), .B(n16495), .ZN(
        n16497) );
  OAI21_X1 U18388 ( .B1(n18479), .B2(n18512), .A(n16497), .ZN(n16498) );
  AOI211_X1 U18389 ( .C1(n16500), .C2(n18556), .A(n16499), .B(n16498), .ZN(
        n16501) );
  OAI21_X1 U18390 ( .B1(n16502), .B2(n16767), .A(n16501), .ZN(P2_U3017) );
  NAND2_X1 U18391 ( .A1(n18553), .A2(n18461), .ZN(n16504) );
  OAI211_X1 U18392 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n16505), .A(
        n16504), .B(n16503), .ZN(n16506) );
  AOI21_X1 U18393 ( .B1(n18462), .B2(n18584), .A(n16506), .ZN(n16507) );
  OAI21_X1 U18394 ( .B1(n16509), .B2(n16508), .A(n16507), .ZN(n16510) );
  AOI21_X1 U18395 ( .B1(n16511), .B2(n18556), .A(n16510), .ZN(n16512) );
  OAI21_X1 U18396 ( .B1(n16513), .B2(n16767), .A(n16512), .ZN(P2_U3018) );
  INV_X1 U18397 ( .A(n16514), .ZN(n18453) );
  AOI21_X1 U18398 ( .B1(n18453), .B2(n18584), .A(n16515), .ZN(n16516) );
  OAI21_X1 U18399 ( .B1(n18579), .B2(n18458), .A(n16516), .ZN(n16518) );
  AOI211_X1 U18400 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n16519), .A(
        n16518), .B(n16517), .ZN(n16523) );
  NAND3_X1 U18401 ( .A1(n16521), .A2(n18556), .A3(n16520), .ZN(n16522) );
  OAI211_X1 U18402 ( .C1(n16524), .C2(n16767), .A(n16523), .B(n16522), .ZN(
        P2_U3019) );
  XNOR2_X1 U18403 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16531) );
  INV_X1 U18404 ( .A(n18442), .ZN(n16528) );
  NOR2_X1 U18405 ( .A1(n16525), .A2(n16537), .ZN(n16526) );
  AOI211_X1 U18406 ( .C1(n16528), .C2(n18584), .A(n16527), .B(n16526), .ZN(
        n16530) );
  NAND2_X1 U18407 ( .A1(n18553), .A2(n18439), .ZN(n16529) );
  OAI211_X1 U18408 ( .C1(n16536), .C2(n16531), .A(n16530), .B(n16529), .ZN(
        n16532) );
  AOI21_X1 U18409 ( .B1(n16533), .B2(n18556), .A(n16532), .ZN(n16534) );
  OAI21_X1 U18410 ( .B1(n16535), .B2(n16767), .A(n16534), .ZN(P2_U3020) );
  NOR2_X1 U18411 ( .A1(n16536), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16543) );
  NOR2_X1 U18412 ( .A1(n16538), .A2(n16537), .ZN(n16539) );
  AOI211_X1 U18413 ( .C1(n18553), .C2(n18428), .A(n16540), .B(n16539), .ZN(
        n16541) );
  OAI21_X1 U18414 ( .B1(n18512), .B2(n18430), .A(n16541), .ZN(n16542) );
  AOI211_X1 U18415 ( .C1(n16544), .C2(n18556), .A(n16543), .B(n16542), .ZN(
        n16545) );
  OAI21_X1 U18416 ( .B1(n16767), .B2(n16546), .A(n16545), .ZN(P2_U3021) );
  XNOR2_X1 U18417 ( .A(n16548), .B(n16547), .ZN(n17201) );
  INV_X1 U18418 ( .A(n17201), .ZN(n16556) );
  AOI21_X1 U18419 ( .B1(n16550), .B2(n16549), .A(n16374), .ZN(n17204) );
  NAND2_X1 U18420 ( .A1(n17204), .A2(n18556), .ZN(n16555) );
  AOI22_X1 U18421 ( .A1(n18553), .A2(n18414), .B1(n18559), .B2(
        P2_REIP_REG_24__SCAN_IN), .ZN(n16551) );
  OAI21_X1 U18422 ( .B1(n18512), .B2(n18413), .A(n16551), .ZN(n16553) );
  AOI211_X1 U18423 ( .C1(n16562), .C2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16553), .B(n16552), .ZN(n16554) );
  OAI211_X1 U18424 ( .C1(n16556), .C2(n16767), .A(n16555), .B(n16554), .ZN(
        P2_U3022) );
  OAI21_X1 U18425 ( .B1(n15425), .B2(n16575), .A(n16557), .ZN(n16561) );
  NOR2_X1 U18426 ( .A1(n18579), .A2(n16558), .ZN(n16560) );
  OAI22_X1 U18427 ( .A1(n18512), .A2(n18402), .B1(n17278), .B2(n18521), .ZN(
        n16559) );
  AOI211_X1 U18428 ( .C1(n16562), .C2(n16561), .A(n16560), .B(n16559), .ZN(
        n16565) );
  NAND2_X1 U18429 ( .A1(n16563), .A2(n18582), .ZN(n16564) );
  OAI211_X1 U18430 ( .C1(n16566), .C2(n18576), .A(n16565), .B(n16564), .ZN(
        P2_U3023) );
  OR2_X1 U18431 ( .A1(n16567), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17189) );
  NAND2_X1 U18432 ( .A1(n17189), .A2(n18556), .ZN(n16583) );
  INV_X1 U18433 ( .A(n16568), .ZN(n16569) );
  OR2_X1 U18434 ( .A1(n16570), .A2(n16569), .ZN(n16571) );
  XNOR2_X1 U18435 ( .A(n16572), .B(n16571), .ZN(n17191) );
  NAND2_X1 U18436 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n18559), .ZN(n16573) );
  OAI221_X1 U18437 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16575), 
        .C1(n15425), .C2(n16574), .A(n16573), .ZN(n16581) );
  AOI21_X1 U18438 ( .B1(n16577), .B2(n16576), .A(n16314), .ZN(n19322) );
  INV_X1 U18439 ( .A(n19322), .ZN(n16578) );
  OAI22_X1 U18440 ( .A1(n18512), .A2(n16579), .B1(n18579), .B2(n16578), .ZN(
        n16580) );
  AOI211_X1 U18441 ( .C1(n17191), .C2(n18582), .A(n16581), .B(n16580), .ZN(
        n16582) );
  OAI21_X1 U18442 ( .B1(n17193), .B2(n16583), .A(n16582), .ZN(P2_U3024) );
  OAI21_X1 U18443 ( .B1(n16587), .B2(n18517), .A(n16731), .ZN(n16586) );
  NOR2_X1 U18444 ( .A1(n17277), .A2(n14141), .ZN(n16585) );
  NOR2_X1 U18445 ( .A1(n18579), .A2(n18391), .ZN(n16584) );
  AOI211_X1 U18446 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n16586), .A(
        n16585), .B(n16584), .ZN(n16590) );
  NAND3_X1 U18447 ( .A1(n16728), .A2(n16588), .A3(n16587), .ZN(n16589) );
  OAI211_X1 U18448 ( .C1(n16591), .C2(n18512), .A(n16590), .B(n16589), .ZN(
        n16592) );
  AOI21_X1 U18449 ( .B1(n16593), .B2(n18556), .A(n16592), .ZN(n16594) );
  OAI21_X1 U18450 ( .B1(n16595), .B2(n16767), .A(n16594), .ZN(P2_U3025) );
  NOR3_X1 U18451 ( .A1(n18568), .A2(n16661), .A3(n16623), .ZN(n16596) );
  AOI211_X1 U18452 ( .C1(n16598), .C2(n16597), .A(n18517), .B(n16596), .ZN(
        n16601) );
  NAND2_X1 U18453 ( .A1(n18573), .A2(n16654), .ZN(n16599) );
  NAND2_X1 U18454 ( .A1(n16600), .A2(n16599), .ZN(n16621) );
  NOR2_X1 U18455 ( .A1(n16601), .A2(n16621), .ZN(n18546) );
  NAND3_X1 U18456 ( .A1(n17165), .A2(n15407), .A3(n16728), .ZN(n18545) );
  NAND2_X1 U18457 ( .A1(n18546), .A2(n18545), .ZN(n18532) );
  NAND2_X1 U18458 ( .A1(n18584), .A2(n18363), .ZN(n16604) );
  NOR2_X1 U18459 ( .A1(n16694), .A2(n16602), .ZN(n18537) );
  AOI22_X1 U18460 ( .A1(n18559), .A2(P2_REIP_REG_19__SCAN_IN), .B1(n18537), 
        .B2(n18539), .ZN(n16603) );
  OAI211_X1 U18461 ( .C1(n16605), .C2(n18579), .A(n16604), .B(n16603), .ZN(
        n16606) );
  AOI21_X1 U18462 ( .B1(n18532), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16606), .ZN(n16609) );
  NAND2_X1 U18463 ( .A1(n16607), .A2(n18556), .ZN(n16608) );
  OAI211_X1 U18464 ( .C1(n16610), .C2(n16767), .A(n16609), .B(n16608), .ZN(
        P2_U3027) );
  NAND2_X1 U18465 ( .A1(n16611), .A2(n16635), .ZN(n16615) );
  NAND2_X1 U18466 ( .A1(n16613), .A2(n16612), .ZN(n16614) );
  XNOR2_X1 U18467 ( .A(n16615), .B(n16614), .ZN(n17164) );
  INV_X1 U18468 ( .A(n16624), .ZN(n16619) );
  NAND2_X1 U18469 ( .A1(n16416), .A2(n16619), .ZN(n17153) );
  INV_X1 U18470 ( .A(n18573), .ZN(n16743) );
  NAND2_X1 U18471 ( .A1(n16743), .A2(n18576), .ZN(n16622) );
  INV_X1 U18472 ( .A(n18568), .ZN(n16618) );
  INV_X1 U18473 ( .A(n16616), .ZN(n16617) );
  OAI21_X1 U18474 ( .B1(n16619), .B2(n16618), .A(n16617), .ZN(n16620) );
  OR2_X1 U18475 ( .A1(n16621), .A2(n16620), .ZN(n16660) );
  AOI21_X1 U18476 ( .B1(n17153), .B2(n16622), .A(n16660), .ZN(n16643) );
  OAI21_X1 U18477 ( .B1(n18519), .B2(n18556), .A(n16623), .ZN(n16626) );
  OAI22_X1 U18478 ( .A1(n17153), .A2(n18576), .B1(n16694), .B2(n16624), .ZN(
        n16632) );
  AOI21_X1 U18479 ( .B1(n16632), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16625) );
  AOI21_X1 U18480 ( .B1(n16643), .B2(n16626), .A(n16625), .ZN(n16630) );
  NAND2_X1 U18481 ( .A1(n18584), .A2(n18339), .ZN(n16627) );
  NAND2_X1 U18482 ( .A1(n18559), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n17170) );
  OAI211_X1 U18483 ( .C1(n16628), .C2(n18579), .A(n16627), .B(n17170), .ZN(
        n16629) );
  AOI211_X1 U18484 ( .C1(n17164), .C2(n18582), .A(n16630), .B(n16629), .ZN(
        n16631) );
  INV_X1 U18485 ( .A(n16631), .ZN(P2_U3029) );
  NAND2_X1 U18486 ( .A1(n16632), .A2(n16642), .ZN(n16641) );
  OR2_X1 U18487 ( .A1(n16634), .A2(n16633), .ZN(n16636) );
  AND2_X1 U18488 ( .A1(n16636), .A2(n16635), .ZN(n17154) );
  NAND2_X1 U18489 ( .A1(n18553), .A2(n19632), .ZN(n16638) );
  NAND2_X1 U18490 ( .A1(n18559), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16637) );
  OAI211_X1 U18491 ( .C1(n18512), .C2(n17155), .A(n16638), .B(n16637), .ZN(
        n16639) );
  AOI21_X1 U18492 ( .B1(n17154), .B2(n18582), .A(n16639), .ZN(n16640) );
  OAI211_X1 U18493 ( .C1(n16643), .C2(n16642), .A(n16641), .B(n16640), .ZN(
        P2_U3030) );
  NAND2_X1 U18494 ( .A1(n16645), .A2(n16644), .ZN(n16649) );
  NAND2_X1 U18495 ( .A1(n16647), .A2(n16646), .ZN(n16648) );
  XNOR2_X1 U18496 ( .A(n16649), .B(n16648), .ZN(n17147) );
  OR2_X1 U18497 ( .A1(n16651), .A2(n16650), .ZN(n16653) );
  NAND2_X1 U18498 ( .A1(n16653), .A2(n16652), .ZN(n19081) );
  NAND2_X1 U18499 ( .A1(n18584), .A2(n18318), .ZN(n16658) );
  NOR2_X1 U18500 ( .A1(n16694), .A2(n16654), .ZN(n16656) );
  NOR2_X1 U18501 ( .A1(n14969), .A2(n14141), .ZN(n16655) );
  AOI21_X1 U18502 ( .B1(n16661), .B2(n16656), .A(n16655), .ZN(n16657) );
  OAI211_X1 U18503 ( .C1(n19081), .C2(n18579), .A(n16658), .B(n16657), .ZN(
        n16659) );
  AOI21_X1 U18504 ( .B1(n16660), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16659), .ZN(n16665) );
  NAND2_X1 U18505 ( .A1(n16662), .A2(n16661), .ZN(n16663) );
  NAND2_X1 U18506 ( .A1(n16663), .A2(n17153), .ZN(n17146) );
  OR2_X1 U18507 ( .A1(n17146), .A2(n18576), .ZN(n16664) );
  OAI211_X1 U18508 ( .C1(n17147), .C2(n16767), .A(n16665), .B(n16664), .ZN(
        P2_U3031) );
  NOR3_X1 U18509 ( .A1(n16694), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n18520), .ZN(n18523) );
  AOI211_X1 U18510 ( .C1(n18520), .C2(n18519), .A(n18523), .B(n18518), .ZN(
        n16680) );
  NOR2_X1 U18511 ( .A1(n16694), .A2(n18520), .ZN(n16666) );
  INV_X1 U18512 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16679) );
  NAND2_X1 U18513 ( .A1(n16666), .A2(n16679), .ZN(n16678) );
  AOI21_X1 U18514 ( .B1(n16680), .B2(n16678), .A(n16667), .ZN(n16674) );
  NAND3_X1 U18515 ( .A1(n16728), .A2(n16668), .A3(n16667), .ZN(n16671) );
  AOI21_X1 U18516 ( .B1(n18553), .B2(n19082), .A(n16669), .ZN(n16670) );
  OAI211_X1 U18517 ( .C1(n16672), .C2(n18512), .A(n16671), .B(n16670), .ZN(
        n16673) );
  AOI211_X1 U18518 ( .C1(n16675), .C2(n18582), .A(n16674), .B(n16673), .ZN(
        n16676) );
  OAI21_X1 U18519 ( .B1(n16677), .B2(n18576), .A(n16676), .ZN(P2_U3032) );
  OAI22_X1 U18520 ( .A1(n16680), .A2(n16679), .B1(n18530), .B2(n16678), .ZN(
        n16682) );
  NOR2_X1 U18521 ( .A1(n14141), .A2(n16453), .ZN(n16681) );
  AOI211_X1 U18522 ( .C1(n18553), .C2(n19086), .A(n16682), .B(n16681), .ZN(
        n16683) );
  OAI21_X1 U18523 ( .B1(n18512), .B2(n16684), .A(n16683), .ZN(n16685) );
  AOI21_X1 U18524 ( .B1(n16686), .B2(n18582), .A(n16685), .ZN(n16687) );
  OAI21_X1 U18525 ( .B1(n16688), .B2(n18576), .A(n16687), .ZN(P2_U3033) );
  OAI21_X1 U18526 ( .B1(n16691), .B2(n16690), .A(n16689), .ZN(n19095) );
  INV_X1 U18527 ( .A(n19095), .ZN(n18306) );
  NOR3_X1 U18528 ( .A1(n16694), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n16692), .ZN(n16699) );
  INV_X1 U18529 ( .A(n16693), .ZN(n16696) );
  NOR3_X1 U18530 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16694), .A3(
        n16730), .ZN(n16706) );
  OAI21_X1 U18531 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18517), .A(
        n16731), .ZN(n16708) );
  OAI21_X1 U18532 ( .B1(n16706), .B2(n16708), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16695) );
  OAI211_X1 U18533 ( .C1(n18512), .C2(n16697), .A(n16696), .B(n16695), .ZN(
        n16698) );
  AOI211_X1 U18534 ( .C1(n18306), .C2(n18553), .A(n16699), .B(n16698), .ZN(
        n16702) );
  NAND2_X1 U18535 ( .A1(n16700), .A2(n18582), .ZN(n16701) );
  OAI211_X1 U18536 ( .C1(n16703), .C2(n18576), .A(n16702), .B(n16701), .ZN(
        P2_U3035) );
  AOI21_X1 U18537 ( .B1(n16705), .B2(n16721), .A(n16704), .ZN(n17135) );
  NAND2_X1 U18538 ( .A1(n17135), .A2(n18556), .ZN(n16720) );
  NOR2_X1 U18539 ( .A1(n13733), .A2(n14141), .ZN(n16707) );
  AOI211_X1 U18540 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16708), .A(
        n16707), .B(n16706), .ZN(n16719) );
  XNOR2_X1 U18541 ( .A(n16709), .B(n16725), .ZN(n19098) );
  NOR2_X1 U18542 ( .A1(n18579), .A2(n19098), .ZN(n16710) );
  AOI21_X1 U18543 ( .B1(n18292), .B2(n18584), .A(n16710), .ZN(n16718) );
  NAND2_X1 U18544 ( .A1(n16712), .A2(n16711), .ZN(n16716) );
  NAND2_X1 U18545 ( .A1(n16714), .A2(n16713), .ZN(n16715) );
  XNOR2_X1 U18546 ( .A(n16716), .B(n16715), .ZN(n17136) );
  NAND2_X1 U18547 ( .A1(n17136), .A2(n18582), .ZN(n16717) );
  NAND4_X1 U18548 ( .A1(n16720), .A2(n16719), .A3(n16718), .A4(n16717), .ZN(
        P2_U3036) );
  NAND3_X1 U18549 ( .A1(n16722), .A2(n18556), .A3(n16721), .ZN(n16734) );
  OR2_X1 U18550 ( .A1(n16724), .A2(n16723), .ZN(n16726) );
  NAND2_X1 U18551 ( .A1(n16726), .A2(n16725), .ZN(n19101) );
  OAI22_X1 U18552 ( .A1(n18579), .A2(n19101), .B1(n14704), .B2(n14141), .ZN(
        n16727) );
  AOI21_X1 U18553 ( .B1(n16728), .B2(n16730), .A(n16727), .ZN(n16729) );
  OAI21_X1 U18554 ( .B1(n16731), .B2(n16730), .A(n16729), .ZN(n16732) );
  AOI21_X1 U18555 ( .B1(n18584), .B2(n18282), .A(n16732), .ZN(n16733) );
  OAI211_X1 U18556 ( .C1(n16735), .C2(n16767), .A(n16734), .B(n16733), .ZN(
        P2_U3037) );
  NAND3_X1 U18557 ( .A1(n16736), .A2(n18556), .A3(n16484), .ZN(n16750) );
  OR2_X1 U18558 ( .A1(n16738), .A2(n16737), .ZN(n16740) );
  NAND2_X1 U18559 ( .A1(n16740), .A2(n16739), .ZN(n19107) );
  INV_X1 U18560 ( .A(n19107), .ZN(n18271) );
  AOI21_X1 U18561 ( .B1(n18571), .B2(n16744), .A(n16743), .ZN(n16741) );
  AOI211_X1 U18562 ( .C1(n18568), .C2(n16742), .A(n18566), .B(n16741), .ZN(
        n16758) );
  OAI21_X1 U18563 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16743), .A(
        n16758), .ZN(n18554) );
  NAND2_X1 U18564 ( .A1(n18554), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16747) );
  NAND2_X1 U18565 ( .A1(n16744), .A2(n16775), .ZN(n16761) );
  NOR2_X1 U18566 ( .A1(n16757), .A2(n16761), .ZN(n18561) );
  AOI22_X1 U18567 ( .A1(n18559), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n16745), 
        .B2(n18561), .ZN(n16746) );
  OAI211_X1 U18568 ( .C1(n18269), .C2(n18512), .A(n16747), .B(n16746), .ZN(
        n16748) );
  AOI21_X1 U18569 ( .B1(n18271), .B2(n18553), .A(n16748), .ZN(n16749) );
  OAI211_X1 U18570 ( .C1(n16751), .C2(n16767), .A(n16750), .B(n16749), .ZN(
        P2_U3039) );
  XNOR2_X1 U18571 ( .A(n16753), .B(n16752), .ZN(n17115) );
  NOR2_X1 U18572 ( .A1(n16754), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17113) );
  INV_X1 U18573 ( .A(n17113), .ZN(n16756) );
  NAND3_X1 U18574 ( .A1(n16756), .A2(n18556), .A3(n16755), .ZN(n16766) );
  NOR2_X1 U18575 ( .A1(n17114), .A2(n18512), .ZN(n16763) );
  OR2_X1 U18576 ( .A1(n16758), .A2(n16757), .ZN(n16760) );
  NAND2_X1 U18577 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n18559), .ZN(n16759) );
  OAI211_X1 U18578 ( .C1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16761), .A(
        n16760), .B(n16759), .ZN(n16762) );
  AOI211_X1 U18579 ( .C1(n16764), .C2(n18553), .A(n16763), .B(n16762), .ZN(
        n16765) );
  OAI211_X1 U18580 ( .C1(n17115), .C2(n16767), .A(n16766), .B(n16765), .ZN(
        P2_U3040) );
  XOR2_X1 U18581 ( .A(n16769), .B(n16768), .Z(n17103) );
  NAND2_X1 U18582 ( .A1(n17103), .A2(n18582), .ZN(n16782) );
  OR2_X1 U18583 ( .A1(n18512), .A2(n17101), .ZN(n16771) );
  NAND2_X1 U18584 ( .A1(n18559), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16770) );
  OAI211_X1 U18585 ( .C1(n17221), .C2(n18579), .A(n16771), .B(n16770), .ZN(
        n16772) );
  INV_X1 U18586 ( .A(n16772), .ZN(n16781) );
  NAND2_X1 U18587 ( .A1(n16774), .A2(n16773), .ZN(n17098) );
  NAND3_X1 U18588 ( .A1(n17099), .A2(n18556), .A3(n17098), .ZN(n16780) );
  INV_X1 U18589 ( .A(n16775), .ZN(n16777) );
  MUX2_X1 U18590 ( .A(n16778), .B(n16777), .S(n16776), .Z(n16779) );
  NAND4_X1 U18591 ( .A1(n16782), .A2(n16781), .A3(n16780), .A4(n16779), .ZN(
        P2_U3043) );
  AOI221_X1 U18592 ( .B1(n18423), .B2(n18247), .C1(n18436), .C2(n16783), .A(
        n15263), .ZN(n16796) );
  INV_X1 U18593 ( .A(n16796), .ZN(n16790) );
  OAI21_X1 U18594 ( .B1(n16784), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n15263), 
        .ZN(n16785) );
  AOI22_X1 U18595 ( .A1(n16790), .A2(n16785), .B1(n19123), .B2(n16794), .ZN(
        n16787) );
  NAND2_X1 U18596 ( .A1(n16799), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16786) );
  OAI21_X1 U18597 ( .B1(n16787), .B2(n16799), .A(n16786), .ZN(P2_U3601) );
  OAI21_X1 U18598 ( .B1(n18423), .B2(n16789), .A(n16788), .ZN(n16795) );
  OAI222_X1 U18599 ( .A1(n18606), .A2(n19142), .B1(n16791), .B2(n18596), .C1(
        n16790), .C2(n16795), .ZN(n16793) );
  MUX2_X1 U18600 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16793), .S(
        n16792), .Z(P2_U3600) );
  AOI222_X1 U18601 ( .A1(n16797), .A2(n17213), .B1(n16796), .B2(n16795), .C1(
        n19525), .C2(n16794), .ZN(n16800) );
  NAND2_X1 U18602 ( .A1(n16799), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16798) );
  OAI21_X1 U18603 ( .B1(n16800), .B2(n16799), .A(n16798), .ZN(P2_U3599) );
  NAND2_X1 U18604 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18672) );
  NAND2_X1 U18605 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18047) );
  INV_X1 U18606 ( .A(n18047), .ZN(n17722) );
  NAND2_X1 U18607 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n17692) );
  NAND2_X1 U18608 ( .A1(n21252), .A2(n17692), .ZN(n20096) );
  NOR2_X1 U18609 ( .A1(n17722), .A2(n20096), .ZN(n16804) );
  NAND2_X1 U18610 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n21216), .ZN(n17694) );
  INV_X1 U18611 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21234) );
  OAI21_X1 U18612 ( .B1(n20821), .B2(n20794), .A(n21234), .ZN(n16801) );
  INV_X1 U18613 ( .A(n16801), .ZN(n16811) );
  NAND2_X1 U18614 ( .A1(n16811), .A2(n17598), .ZN(n17693) );
  NOR2_X1 U18615 ( .A1(n17690), .A2(n17692), .ZN(n21249) );
  OAI21_X1 U18616 ( .B1(n17693), .B2(P3_FLUSH_REG_SCAN_IN), .A(n21249), .ZN(
        n16803) );
  INV_X1 U18617 ( .A(n21255), .ZN(n16802) );
  NOR2_X1 U18618 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21252), .ZN(
        n21254) );
  AOI21_X1 U18619 ( .B1(n16802), .B2(n17692), .A(n21254), .ZN(n18654) );
  NOR2_X1 U18620 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18654), .ZN(n18932) );
  INV_X1 U18621 ( .A(n18932), .ZN(n18979) );
  NAND2_X1 U18622 ( .A1(n16803), .A2(n18979), .ZN(n18096) );
  NAND2_X1 U18623 ( .A1(n17694), .A2(n18096), .ZN(n18097) );
  AOI221_X1 U18624 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18672), .C1(n16804), 
        .C2(n18672), .A(n18097), .ZN(n18094) );
  INV_X1 U18625 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21672) );
  NOR3_X1 U18626 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n21672), .ZN(n18693) );
  AOI21_X1 U18627 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n16804), .ZN(n16805) );
  INV_X1 U18628 ( .A(n16805), .ZN(n18095) );
  OAI221_X1 U18629 ( .B1(n18693), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18693), .C2(n18095), .A(n18096), .ZN(n18092) );
  AOI22_X1 U18630 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18094), .B1(
        n18092), .B2(n18652), .ZN(P3_U2865) );
  NOR2_X1 U18631 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21252), .ZN(n21248) );
  INV_X1 U18632 ( .A(n16806), .ZN(n16809) );
  NAND2_X1 U18633 ( .A1(n17696), .A2(n16807), .ZN(n17293) );
  INV_X1 U18634 ( .A(n20155), .ZN(n20100) );
  NOR2_X1 U18635 ( .A1(n21206), .A2(n20100), .ZN(n16824) );
  INV_X1 U18636 ( .A(n21207), .ZN(n21200) );
  OAI211_X1 U18637 ( .C1(n16824), .C2(n20593), .A(n21723), .B(n21200), .ZN(
        n16808) );
  NAND3_X1 U18638 ( .A1(n16809), .A2(n17293), .A3(n16808), .ZN(n21233) );
  NOR2_X1 U18639 ( .A1(n21224), .A2(n21263), .ZN(n16810) );
  NOR2_X1 U18640 ( .A1(n16811), .A2(n21204), .ZN(n21238) );
  INV_X1 U18641 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20785) );
  NAND2_X1 U18642 ( .A1(n20785), .A2(n21252), .ZN(n20790) );
  INV_X1 U18643 ( .A(n20790), .ZN(n20824) );
  NAND3_X1 U18644 ( .A1(n20826), .A2(n21238), .A3(n20824), .ZN(n16812) );
  OAI21_X1 U18645 ( .B1(n20826), .B2(n21234), .A(n16812), .ZN(P3_U3284) );
  NAND2_X1 U18646 ( .A1(n16814), .A2(n16813), .ZN(n16816) );
  OAI22_X1 U18647 ( .A1(n16817), .A2(n16816), .B1(n16815), .B2(n21647), .ZN(
        P1_U3468) );
  INV_X1 U18648 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21715) );
  OAI21_X1 U18649 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n21715), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18171) );
  NAND2_X1 U18650 ( .A1(n21724), .A2(n18171), .ZN(n16819) );
  INV_X1 U18651 ( .A(n16819), .ZN(n21675) );
  NOR2_X1 U18652 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n21676) );
  OAI21_X1 U18653 ( .B1(BS16), .B2(n21676), .A(n21675), .ZN(n21673) );
  OAI21_X1 U18654 ( .B1(P3_DATAWIDTH_REG_0__SCAN_IN), .B2(n21675), .A(n21673), 
        .ZN(n16818) );
  INV_X1 U18655 ( .A(n16818), .ZN(P3_U3280) );
  AND2_X1 U18656 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n16819), .ZN(P3_U3028) );
  AND2_X1 U18657 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n16819), .ZN(P3_U3027) );
  AND2_X1 U18658 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n16819), .ZN(P3_U3026) );
  AND2_X1 U18659 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n16819), .ZN(P3_U3025) );
  AND2_X1 U18660 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n16819), .ZN(P3_U3024) );
  AND2_X1 U18661 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n16819), .ZN(P3_U3023) );
  AND2_X1 U18662 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n16819), .ZN(P3_U3022) );
  AND2_X1 U18663 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n16819), .ZN(P3_U3021) );
  AND2_X1 U18664 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n16819), .ZN(
        P3_U3020) );
  AND2_X1 U18665 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n16819), .ZN(
        P3_U3019) );
  AND2_X1 U18666 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n16819), .ZN(
        P3_U3018) );
  AND2_X1 U18667 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n16819), .ZN(
        P3_U3017) );
  AND2_X1 U18668 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n16819), .ZN(
        P3_U3016) );
  AND2_X1 U18669 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n16819), .ZN(
        P3_U3015) );
  AND2_X1 U18670 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n16819), .ZN(
        P3_U3014) );
  AND2_X1 U18671 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n16819), .ZN(
        P3_U3013) );
  AND2_X1 U18672 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n16819), .ZN(
        P3_U3012) );
  AND2_X1 U18673 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n16819), .ZN(
        P3_U3011) );
  AND2_X1 U18674 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n16819), .ZN(
        P3_U3010) );
  AND2_X1 U18675 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n16819), .ZN(
        P3_U3009) );
  AND2_X1 U18676 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n16819), .ZN(
        P3_U3008) );
  AND2_X1 U18677 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n16819), .ZN(
        P3_U3007) );
  AND2_X1 U18678 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n16819), .ZN(
        P3_U3006) );
  AND2_X1 U18679 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n16819), .ZN(
        P3_U3005) );
  AND2_X1 U18680 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n16819), .ZN(
        P3_U3004) );
  AND2_X1 U18681 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n16819), .ZN(
        P3_U3003) );
  AND2_X1 U18682 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n16819), .ZN(
        P3_U3002) );
  AND2_X1 U18683 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n16819), .ZN(
        P3_U3001) );
  AND2_X1 U18684 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n16819), .ZN(
        P3_U3000) );
  AND2_X1 U18685 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n16819), .ZN(
        P3_U2999) );
  AOI21_X1 U18686 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n16821)
         );
  INV_X1 U18687 ( .A(n21723), .ZN(n21679) );
  INV_X1 U18688 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n16823) );
  NAND4_X1 U18689 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(n21679), .A4(n16823), .ZN(n21245) );
  INV_X1 U18690 ( .A(n21245), .ZN(n16820) );
  AOI211_X1 U18691 ( .C1(n18047), .C2(n16821), .A(n21249), .B(n16820), .ZN(
        P3_U2998) );
  NOR2_X1 U18692 ( .A1(n16822), .A2(n18096), .ZN(P3_U2867) );
  NOR2_X1 U18693 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n16823), .ZN(n17839) );
  INV_X1 U18694 ( .A(n17839), .ZN(n18086) );
  OR2_X1 U18695 ( .A1(n20785), .A2(n18086), .ZN(n20097) );
  AND2_X1 U18697 ( .A1(n18159), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U18698 ( .A1(n17691), .A2(n20157), .ZN(n16827) );
  OAI22_X1 U18699 ( .A1(P3_READREQUEST_REG_SCAN_IN), .A2(n16827), .B1(n20102), 
        .B2(n20157), .ZN(n16826) );
  INV_X1 U18700 ( .A(n16826), .ZN(P3_U3298) );
  NOR2_X1 U18701 ( .A1(n20592), .A2(n20157), .ZN(n20584) );
  NOR2_X1 U18702 ( .A1(P3_MEMORYFETCH_REG_SCAN_IN), .A2(n16827), .ZN(n16828)
         );
  NOR2_X1 U18703 ( .A1(n20584), .A2(n16828), .ZN(P3_U3299) );
  AND2_X1 U18704 ( .A1(n21713), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21705) );
  AOI21_X1 U18705 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21705), .A(n16829), 
        .ZN(n16831) );
  INV_X1 U18706 ( .A(n16831), .ZN(n21671) );
  NOR2_X1 U18707 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n21700) );
  OAI21_X1 U18708 ( .B1(BS16), .B2(n21700), .A(n21671), .ZN(n21669) );
  OAI21_X1 U18709 ( .B1(n21671), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n21669), 
        .ZN(n16830) );
  INV_X1 U18710 ( .A(n16830), .ZN(P2_U3591) );
  INV_X1 U18711 ( .A(n21671), .ZN(n17239) );
  AND2_X1 U18712 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17239), .ZN(P2_U3208) );
  AND2_X1 U18713 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17239), .ZN(P2_U3207) );
  AND2_X1 U18714 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17239), .ZN(P2_U3206) );
  AND2_X1 U18715 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17239), .ZN(P2_U3205) );
  AND2_X1 U18716 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17239), .ZN(P2_U3204) );
  AND2_X1 U18717 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17239), .ZN(P2_U3203) );
  AND2_X1 U18718 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17239), .ZN(P2_U3202) );
  AND2_X1 U18719 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17239), .ZN(P2_U3201) );
  AND2_X1 U18720 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n16831), .ZN(
        P2_U3200) );
  AND2_X1 U18721 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n16831), .ZN(
        P2_U3199) );
  AND2_X1 U18722 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n16831), .ZN(
        P2_U3198) );
  AND2_X1 U18723 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n16831), .ZN(
        P2_U3197) );
  AND2_X1 U18724 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n16831), .ZN(
        P2_U3196) );
  AND2_X1 U18725 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n16831), .ZN(
        P2_U3195) );
  AND2_X1 U18726 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n16831), .ZN(
        P2_U3194) );
  AND2_X1 U18727 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17239), .ZN(
        P2_U3193) );
  AND2_X1 U18728 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17239), .ZN(
        P2_U3192) );
  AND2_X1 U18729 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17239), .ZN(
        P2_U3191) );
  AND2_X1 U18730 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17239), .ZN(
        P2_U3190) );
  AND2_X1 U18731 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17239), .ZN(
        P2_U3189) );
  AND2_X1 U18732 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17239), .ZN(
        P2_U3188) );
  AND2_X1 U18733 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17239), .ZN(
        P2_U3187) );
  AND2_X1 U18734 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17239), .ZN(
        P2_U3186) );
  AND2_X1 U18735 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17239), .ZN(
        P2_U3185) );
  AND2_X1 U18736 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17239), .ZN(
        P2_U3184) );
  AND2_X1 U18737 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17239), .ZN(
        P2_U3183) );
  AND2_X1 U18738 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17239), .ZN(
        P2_U3182) );
  AND2_X1 U18739 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17239), .ZN(
        P2_U3181) );
  AND2_X1 U18740 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17239), .ZN(
        P2_U3180) );
  AND2_X1 U18741 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17239), .ZN(
        P2_U3179) );
  NAND2_X1 U18742 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18222), .ZN(n18597) );
  AOI21_X1 U18743 ( .B1(n16832), .B2(n14714), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16834) );
  AOI221_X1 U18744 ( .B1(n18597), .B2(n16834), .C1(n15263), .C2(n16834), .A(
        n16833), .ZN(P2_U3178) );
  AOI21_X1 U18745 ( .B1(n15263), .B2(n19214), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18605) );
  NAND2_X1 U18746 ( .A1(n16835), .A2(n18605), .ZN(n19116) );
  OAI221_X1 U18747 ( .B1(n16837), .B2(n18624), .C1(n16837), .C2(n16836), .A(
        n19639), .ZN(n17228) );
  NOR2_X1 U18748 ( .A1(n16838), .A2(n17228), .ZN(P2_U3047) );
  AND2_X1 U18749 ( .A1(n17254), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U18750 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16842) );
  NOR4_X1 U18751 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16841) );
  NOR4_X1 U18752 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16840) );
  NOR4_X1 U18753 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16839) );
  NAND4_X1 U18754 ( .A1(n16842), .A2(n16841), .A3(n16840), .A4(n16839), .ZN(
        n16848) );
  NOR4_X1 U18755 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16846) );
  AOI211_X1 U18756 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16845) );
  NOR4_X1 U18757 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16844) );
  NOR4_X1 U18758 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16843) );
  NAND4_X1 U18759 ( .A1(n16846), .A2(n16845), .A3(n16844), .A4(n16843), .ZN(
        n16847) );
  NOR2_X1 U18760 ( .A1(n16848), .A2(n16847), .ZN(n17235) );
  INV_X1 U18761 ( .A(n17235), .ZN(n17234) );
  NOR2_X1 U18762 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17234), .ZN(n17229) );
  OR3_X1 U18763 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17233) );
  INV_X1 U18764 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17288) );
  AOI22_X1 U18765 ( .A1(n17229), .A2(n17233), .B1(n17234), .B2(n17288), .ZN(
        P2_U2821) );
  INV_X1 U18766 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U18767 ( .A1(n17229), .A2(n18240), .B1(n17234), .B2(n17286), .ZN(
        P2_U2820) );
  INV_X1 U18768 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21696) );
  NAND2_X1 U18769 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21696), .ZN(n22276) );
  NAND2_X1 U18770 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21684), .ZN(n16889) );
  NAND2_X1 U18771 ( .A1(n22276), .A2(n16889), .ZN(n16850) );
  INV_X1 U18772 ( .A(n16850), .ZN(n21668) );
  OAI221_X1 U18773 ( .B1(n11585), .B2(BS16), .C1(n21690), .C2(BS16), .A(n21668), .ZN(n21666) );
  OAI21_X1 U18774 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21668), .A(n21666), 
        .ZN(n16849) );
  INV_X1 U18775 ( .A(n16849), .ZN(P1_U3464) );
  AND2_X1 U18776 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n16850), .ZN(P1_U3193) );
  AND2_X1 U18777 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n16850), .ZN(P1_U3192) );
  AND2_X1 U18778 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n16850), .ZN(P1_U3191) );
  AND2_X1 U18779 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n16850), .ZN(P1_U3190) );
  AND2_X1 U18780 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n16850), .ZN(P1_U3189) );
  AND2_X1 U18781 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n16850), .ZN(P1_U3188) );
  AND2_X1 U18782 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n16850), .ZN(P1_U3187) );
  AND2_X1 U18783 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n16850), .ZN(P1_U3186) );
  AND2_X1 U18784 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n16850), .ZN(
        P1_U3185) );
  AND2_X1 U18785 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n16850), .ZN(
        P1_U3184) );
  AND2_X1 U18786 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n16850), .ZN(
        P1_U3183) );
  AND2_X1 U18787 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n16850), .ZN(
        P1_U3182) );
  AND2_X1 U18788 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n16850), .ZN(
        P1_U3181) );
  AND2_X1 U18789 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n16850), .ZN(
        P1_U3180) );
  AND2_X1 U18790 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n16850), .ZN(
        P1_U3179) );
  AND2_X1 U18791 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n16850), .ZN(
        P1_U3178) );
  AND2_X1 U18792 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n16850), .ZN(
        P1_U3177) );
  AND2_X1 U18793 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n16850), .ZN(
        P1_U3176) );
  AND2_X1 U18794 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n16850), .ZN(
        P1_U3175) );
  AND2_X1 U18795 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n16850), .ZN(
        P1_U3174) );
  AND2_X1 U18796 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n16850), .ZN(
        P1_U3173) );
  AND2_X1 U18797 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n16850), .ZN(
        P1_U3172) );
  AND2_X1 U18798 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n16850), .ZN(
        P1_U3171) );
  AND2_X1 U18799 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n16850), .ZN(
        P1_U3170) );
  AND2_X1 U18800 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n16850), .ZN(
        P1_U3169) );
  AND2_X1 U18801 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n16850), .ZN(
        P1_U3168) );
  AND2_X1 U18802 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n16850), .ZN(
        P1_U3167) );
  AND2_X1 U18803 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n16850), .ZN(
        P1_U3166) );
  AND2_X1 U18804 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n16850), .ZN(
        P1_U3165) );
  AND2_X1 U18805 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n16850), .ZN(
        P1_U3164) );
  INV_X1 U18806 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17073) );
  INV_X1 U18807 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21640) );
  AND2_X1 U18808 ( .A1(n17073), .A2(n21640), .ZN(n16871) );
  NOR2_X1 U18809 ( .A1(n16860), .A2(n16851), .ZN(n16863) );
  NOR2_X1 U18810 ( .A1(n16852), .A2(n21892), .ZN(n16853) );
  AND2_X1 U18811 ( .A1(n16854), .A2(n16853), .ZN(n16857) );
  INV_X1 U18812 ( .A(n16857), .ZN(n16859) );
  OAI22_X1 U18813 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16857), .B1(
        n16856), .B2(n16855), .ZN(n16858) );
  OAI21_X1 U18814 ( .B1(n16859), .B2(n21880), .A(n16858), .ZN(n16862) );
  INV_X1 U18815 ( .A(n16860), .ZN(n16861) );
  OAI22_X1 U18816 ( .A1(n16863), .A2(n16862), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16861), .ZN(n16864) );
  AOI222_X1 U18817 ( .A1(n16865), .A2(n11834), .B1(n16865), .B2(n16864), .C1(
        n11834), .C2(n16864), .ZN(n16866) );
  NOR2_X1 U18818 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16866), .ZN(
        n16867) );
  NOR2_X1 U18819 ( .A1(n16868), .A2(n16867), .ZN(n16870) );
  OAI211_X1 U18820 ( .C1(n16872), .C2(n16871), .A(n16870), .B(n16869), .ZN(
        n16873) );
  NOR2_X1 U18821 ( .A1(n16874), .A2(n16873), .ZN(n21665) );
  INV_X1 U18822 ( .A(n21665), .ZN(n16881) );
  OR2_X1 U18823 ( .A1(n16875), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n16879) );
  OAI21_X1 U18824 ( .B1(n21683), .B2(n16877), .A(n16876), .ZN(n16878) );
  OAI21_X1 U18825 ( .B1(n16880), .B2(n16879), .A(n16878), .ZN(n16883) );
  AOI221_X1 U18826 ( .B1(n21655), .B2(n16886), .C1(n16881), .C2(n16886), .A(
        n16883), .ZN(n21657) );
  NOR2_X1 U18827 ( .A1(n21657), .A2(n21655), .ZN(n21656) );
  OAI211_X1 U18828 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21683), .A(n21656), 
        .B(n16882), .ZN(n21661) );
  NOR2_X1 U18829 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21655), .ZN(n21651) );
  AOI21_X1 U18830 ( .B1(n21691), .B2(n21651), .A(n16886), .ZN(n21650) );
  AND3_X1 U18831 ( .A1(n21650), .A2(n16884), .A3(n16883), .ZN(n16885) );
  AOI21_X1 U18832 ( .B1(n16886), .B2(n21661), .A(n16885), .ZN(P1_U3162) );
  NOR2_X1 U18833 ( .A1(n16888), .A2(n16887), .ZN(P1_U3032) );
  AND2_X1 U18834 ( .A1(n19841), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OAI21_X1 U18835 ( .B1(n16889), .B2(P1_ADS_N_REG_SCAN_IN), .A(n22276), .ZN(
        n16890) );
  INV_X1 U18836 ( .A(n16890), .ZN(P1_U2802) );
  AOI222_X1 U18837 ( .A1(P1_EAX_REG_9__SCAN_IN), .A2(n19820), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n19841), .C1(n21278), .C2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n17095) );
  INV_X1 U18838 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n19872) );
  OAI22_X1 U18839 ( .A1(n19872), .A2(keyinput_63), .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_62), .ZN(n16891) );
  AOI221_X1 U18840 ( .B1(n19872), .B2(keyinput_63), .C1(keyinput_62), .C2(
        P1_REIP_REG_21__SCAN_IN), .A(n16891), .ZN(n16986) );
  INV_X1 U18841 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U18842 ( .A1(n19881), .A2(keyinput_58), .B1(n19877), .B2(
        keyinput_59), .ZN(n16892) );
  OAI221_X1 U18843 ( .B1(n19881), .B2(keyinput_58), .C1(n19877), .C2(
        keyinput_59), .A(n16892), .ZN(n16984) );
  AOI22_X1 U18844 ( .A1(n19884), .A2(keyinput_56), .B1(n15807), .B2(
        keyinput_53), .ZN(n16893) );
  OAI221_X1 U18845 ( .B1(n19884), .B2(keyinput_56), .C1(n15807), .C2(
        keyinput_53), .A(n16893), .ZN(n16896) );
  AOI22_X1 U18846 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_54), .B1(n19891), .B2(keyinput_52), .ZN(n16894) );
  OAI221_X1 U18847 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_54), .C1(
        n19891), .C2(keyinput_52), .A(n16894), .ZN(n16895) );
  AOI211_X1 U18848 ( .C1(keyinput_55), .C2(P1_REIP_REG_28__SCAN_IN), .A(n16896), .B(n16895), .ZN(n16897) );
  OAI21_X1 U18849 ( .B1(keyinput_55), .B2(P1_REIP_REG_28__SCAN_IN), .A(n16897), 
        .ZN(n16980) );
  INV_X1 U18850 ( .A(keyinput_51), .ZN(n16978) );
  INV_X1 U18851 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19895) );
  INV_X1 U18852 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19910) );
  INV_X1 U18853 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19914) );
  AOI22_X1 U18854 ( .A1(P1_BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_48), .B1(
        n19914), .B2(keyinput_49), .ZN(n16898) );
  OAI221_X1 U18855 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_48), .C1(
        n19914), .C2(keyinput_49), .A(n16898), .ZN(n16975) );
  INV_X1 U18856 ( .A(keyinput_47), .ZN(n16973) );
  INV_X1 U18857 ( .A(keyinput_46), .ZN(n16971) );
  INV_X1 U18858 ( .A(keyinput_45), .ZN(n16969) );
  INV_X1 U18859 ( .A(keyinput_44), .ZN(n16967) );
  INV_X1 U18860 ( .A(keyinput_43), .ZN(n16965) );
  INV_X1 U18861 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n17067) );
  INV_X1 U18862 ( .A(keyinput_42), .ZN(n16963) );
  INV_X1 U18863 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20026) );
  AOI22_X1 U18864 ( .A1(keyinput_39), .A2(P1_ADS_N_REG_SCAN_IN), .B1(n16996), 
        .B2(keyinput_40), .ZN(n16899) );
  OAI221_X1 U18865 ( .B1(keyinput_39), .B2(P1_ADS_N_REG_SCAN_IN), .C1(n16996), 
        .C2(keyinput_40), .A(n16899), .ZN(n16960) );
  INV_X1 U18866 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n17059) );
  INV_X1 U18867 ( .A(keyinput_38), .ZN(n16958) );
  OAI22_X1 U18868 ( .A1(READY1), .A2(keyinput_36), .B1(READY2), .B2(
        keyinput_37), .ZN(n16900) );
  AOI221_X1 U18869 ( .B1(READY1), .B2(keyinput_36), .C1(keyinput_37), .C2(
        READY2), .A(n16900), .ZN(n16955) );
  INV_X1 U18870 ( .A(DATAI_7_), .ZN(n16902) );
  OAI22_X1 U18871 ( .A1(n16902), .A2(keyinput_25), .B1(DATAI_6_), .B2(
        keyinput_26), .ZN(n16901) );
  AOI221_X1 U18872 ( .B1(n16902), .B2(keyinput_25), .C1(keyinput_26), .C2(
        DATAI_6_), .A(n16901), .ZN(n16943) );
  AOI22_X1 U18873 ( .A1(n16904), .A2(keyinput_23), .B1(n17035), .B2(
        keyinput_22), .ZN(n16903) );
  OAI221_X1 U18874 ( .B1(n16904), .B2(keyinput_23), .C1(n17035), .C2(
        keyinput_22), .A(n16903), .ZN(n16939) );
  AOI22_X1 U18875 ( .A1(DATAI_19_), .A2(keyinput_13), .B1(n17002), .B2(
        keyinput_14), .ZN(n16905) );
  OAI221_X1 U18876 ( .B1(DATAI_19_), .B2(keyinput_13), .C1(n17002), .C2(
        keyinput_14), .A(n16905), .ZN(n16927) );
  INV_X1 U18877 ( .A(keyinput_12), .ZN(n16925) );
  INV_X1 U18878 ( .A(keyinput_11), .ZN(n16923) );
  XNOR2_X1 U18879 ( .A(keyinput_6), .B(n16906), .ZN(n16921) );
  OAI22_X1 U18880 ( .A1(DATAI_31_), .A2(keyinput_1), .B1(
        P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_0), .ZN(n16907) );
  AOI221_X1 U18881 ( .B1(DATAI_31_), .B2(keyinput_1), .C1(keyinput_0), .C2(
        P1_MEMORYFETCH_REG_SCAN_IN), .A(n16907), .ZN(n16914) );
  AOI22_X1 U18882 ( .A1(n16910), .A2(keyinput_3), .B1(n16909), .B2(keyinput_2), 
        .ZN(n16908) );
  OAI221_X1 U18883 ( .B1(n16910), .B2(keyinput_3), .C1(n16909), .C2(keyinput_2), .A(n16908), .ZN(n16913) );
  OAI22_X1 U18884 ( .A1(DATAI_28_), .A2(keyinput_4), .B1(DATAI_27_), .B2(
        keyinput_5), .ZN(n16911) );
  AOI221_X1 U18885 ( .B1(DATAI_28_), .B2(keyinput_4), .C1(keyinput_5), .C2(
        DATAI_27_), .A(n16911), .ZN(n16912) );
  OAI21_X1 U18886 ( .B1(n16914), .B2(n16913), .A(n16912), .ZN(n16920) );
  AOI22_X1 U18887 ( .A1(n17010), .A2(keyinput_8), .B1(keyinput_10), .B2(n16916), .ZN(n16915) );
  OAI221_X1 U18888 ( .B1(n17010), .B2(keyinput_8), .C1(n16916), .C2(
        keyinput_10), .A(n16915), .ZN(n16919) );
  AOI22_X1 U18889 ( .A1(DATAI_23_), .A2(keyinput_9), .B1(DATAI_25_), .B2(
        keyinput_7), .ZN(n16917) );
  OAI221_X1 U18890 ( .B1(DATAI_23_), .B2(keyinput_9), .C1(DATAI_25_), .C2(
        keyinput_7), .A(n16917), .ZN(n16918) );
  AOI211_X1 U18891 ( .C1(n16921), .C2(n16920), .A(n16919), .B(n16918), .ZN(
        n16922) );
  AOI221_X1 U18892 ( .B1(DATAI_21_), .B2(keyinput_11), .C1(n17017), .C2(n16923), .A(n16922), .ZN(n16924) );
  AOI221_X1 U18893 ( .B1(DATAI_20_), .B2(keyinput_12), .C1(n17021), .C2(n16925), .A(n16924), .ZN(n16926) );
  OAI22_X1 U18894 ( .A1(n16927), .A2(n16926), .B1(DATAI_17_), .B2(keyinput_15), 
        .ZN(n16928) );
  AOI21_X1 U18895 ( .B1(DATAI_17_), .B2(keyinput_15), .A(n16928), .ZN(n16936)
         );
  OAI22_X1 U18896 ( .A1(DATAI_16_), .A2(keyinput_16), .B1(keyinput_17), .B2(
        DATAI_15_), .ZN(n16929) );
  AOI221_X1 U18897 ( .B1(DATAI_16_), .B2(keyinput_16), .C1(DATAI_15_), .C2(
        keyinput_17), .A(n16929), .ZN(n16935) );
  INV_X1 U18898 ( .A(DATAI_13_), .ZN(n16931) );
  AOI22_X1 U18899 ( .A1(DATAI_14_), .A2(keyinput_18), .B1(n16931), .B2(
        keyinput_19), .ZN(n16930) );
  OAI221_X1 U18900 ( .B1(DATAI_14_), .B2(keyinput_18), .C1(n16931), .C2(
        keyinput_19), .A(n16930), .ZN(n16934) );
  AOI22_X1 U18901 ( .A1(DATAI_11_), .A2(keyinput_21), .B1(DATAI_12_), .B2(
        keyinput_20), .ZN(n16932) );
  OAI221_X1 U18902 ( .B1(DATAI_11_), .B2(keyinput_21), .C1(DATAI_12_), .C2(
        keyinput_20), .A(n16932), .ZN(n16933) );
  AOI211_X1 U18903 ( .C1(n16936), .C2(n16935), .A(n16934), .B(n16933), .ZN(
        n16938) );
  NAND2_X1 U18904 ( .A1(DATAI_8_), .A2(keyinput_24), .ZN(n16937) );
  OAI221_X1 U18905 ( .B1(n16939), .B2(n16938), .C1(DATAI_8_), .C2(keyinput_24), 
        .A(n16937), .ZN(n16942) );
  INV_X1 U18906 ( .A(DATAI_4_), .ZN(n16998) );
  INV_X1 U18907 ( .A(DATAI_5_), .ZN(n16999) );
  AOI22_X1 U18908 ( .A1(n16998), .A2(keyinput_28), .B1(n16999), .B2(
        keyinput_27), .ZN(n16940) );
  OAI221_X1 U18909 ( .B1(n16998), .B2(keyinput_28), .C1(n16999), .C2(
        keyinput_27), .A(n16940), .ZN(n16941) );
  AOI21_X1 U18910 ( .B1(n16943), .B2(n16942), .A(n16941), .ZN(n16948) );
  INV_X1 U18911 ( .A(DATAI_1_), .ZN(n16945) );
  OAI22_X1 U18912 ( .A1(n16945), .A2(keyinput_31), .B1(DATAI_2_), .B2(
        keyinput_30), .ZN(n16944) );
  AOI221_X1 U18913 ( .B1(n16945), .B2(keyinput_31), .C1(keyinput_30), .C2(
        DATAI_2_), .A(n16944), .ZN(n16946) );
  OAI21_X1 U18914 ( .B1(keyinput_29), .B2(DATAI_3_), .A(n16946), .ZN(n16947)
         );
  AOI211_X1 U18915 ( .C1(keyinput_29), .C2(DATAI_3_), .A(n16948), .B(n16947), 
        .ZN(n16952) );
  AOI22_X1 U18916 ( .A1(HOLD), .A2(keyinput_33), .B1(n16950), .B2(keyinput_32), 
        .ZN(n16949) );
  OAI221_X1 U18917 ( .B1(HOLD), .B2(keyinput_33), .C1(n16950), .C2(keyinput_32), .A(n16949), .ZN(n16951) );
  AOI211_X1 U18918 ( .C1(NA), .C2(keyinput_34), .A(n16952), .B(n16951), .ZN(
        n16953) );
  OAI21_X1 U18919 ( .B1(NA), .B2(keyinput_34), .A(n16953), .ZN(n16954) );
  OAI211_X1 U18920 ( .C1(BS16), .C2(keyinput_35), .A(n16955), .B(n16954), .ZN(
        n16956) );
  AOI21_X1 U18921 ( .B1(BS16), .B2(keyinput_35), .A(n16956), .ZN(n16957) );
  AOI221_X1 U18922 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_38), .C1(
        n17059), .C2(n16958), .A(n16957), .ZN(n16959) );
  OAI22_X1 U18923 ( .A1(n16960), .A2(n16959), .B1(keyinput_41), .B2(
        P1_M_IO_N_REG_SCAN_IN), .ZN(n16961) );
  AOI21_X1 U18924 ( .B1(keyinput_41), .B2(P1_M_IO_N_REG_SCAN_IN), .A(n16961), 
        .ZN(n16962) );
  AOI221_X1 U18925 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(n16963), .C1(n20026), .C2(
        keyinput_42), .A(n16962), .ZN(n16964) );
  AOI221_X1 U18926 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n16965), .C1(
        n17067), .C2(keyinput_43), .A(n16964), .ZN(n16966) );
  AOI221_X1 U18927 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n16967), .C1(n14439), 
        .C2(keyinput_44), .A(n16966), .ZN(n16968) );
  AOI221_X1 U18928 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_45), .C1(n17073), 
        .C2(n16969), .A(n16968), .ZN(n16970) );
  AOI221_X1 U18929 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_46), .C1(n21640), 
        .C2(n16971), .A(n16970), .ZN(n16972) );
  AOI221_X1 U18930 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_47), .C1(n20095), 
        .C2(n16973), .A(n16972), .ZN(n16974) );
  OAI22_X1 U18931 ( .A1(keyinput_50), .A2(n19910), .B1(n16975), .B2(n16974), 
        .ZN(n16976) );
  AOI21_X1 U18932 ( .B1(keyinput_50), .B2(n19910), .A(n16976), .ZN(n16977) );
  AOI221_X1 U18933 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(n16978), .C1(
        n19895), .C2(keyinput_51), .A(n16977), .ZN(n16979) );
  OAI22_X1 U18934 ( .A1(n16980), .A2(n16979), .B1(keyinput_57), .B2(
        P1_REIP_REG_26__SCAN_IN), .ZN(n16981) );
  AOI21_X1 U18935 ( .B1(keyinput_57), .B2(P1_REIP_REG_26__SCAN_IN), .A(n16981), 
        .ZN(n16983) );
  NAND2_X1 U18936 ( .A1(n21600), .A2(keyinput_60), .ZN(n16982) );
  OAI221_X1 U18937 ( .B1(n16984), .B2(n16983), .C1(n21600), .C2(keyinput_60), 
        .A(n16982), .ZN(n16985) );
  OAI211_X1 U18938 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(keyinput_61), .A(n16986), .B(n16985), .ZN(n16987) );
  AOI21_X1 U18939 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_61), .A(n16987), 
        .ZN(n17093) );
  AOI22_X1 U18940 ( .A1(n19877), .A2(keyinput_123), .B1(keyinput_122), .B2(
        n19881), .ZN(n16988) );
  OAI221_X1 U18941 ( .B1(n19877), .B2(keyinput_123), .C1(n19881), .C2(
        keyinput_122), .A(n16988), .ZN(n17087) );
  INV_X1 U18942 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U18943 ( .A1(n15807), .A2(keyinput_117), .B1(keyinput_119), .B2(
        n19887), .ZN(n16989) );
  OAI221_X1 U18944 ( .B1(n15807), .B2(keyinput_117), .C1(n19887), .C2(
        keyinput_119), .A(n16989), .ZN(n16992) );
  AOI22_X1 U18945 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_118), .B1(
        n19884), .B2(keyinput_120), .ZN(n16990) );
  OAI221_X1 U18946 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_118), .C1(
        n19884), .C2(keyinput_120), .A(n16990), .ZN(n16991) );
  AOI211_X1 U18947 ( .C1(keyinput_116), .C2(P1_REIP_REG_31__SCAN_IN), .A(
        n16992), .B(n16991), .ZN(n16993) );
  OAI21_X1 U18948 ( .B1(keyinput_116), .B2(P1_REIP_REG_31__SCAN_IN), .A(n16993), .ZN(n17084) );
  INV_X1 U18949 ( .A(keyinput_115), .ZN(n17082) );
  INV_X1 U18950 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19917) );
  AOI22_X1 U18951 ( .A1(n19914), .A2(keyinput_113), .B1(keyinput_112), .B2(
        n19917), .ZN(n16994) );
  OAI221_X1 U18952 ( .B1(n19914), .B2(keyinput_113), .C1(n19917), .C2(
        keyinput_112), .A(n16994), .ZN(n17079) );
  INV_X1 U18953 ( .A(keyinput_111), .ZN(n17077) );
  INV_X1 U18954 ( .A(keyinput_110), .ZN(n17075) );
  INV_X1 U18955 ( .A(keyinput_109), .ZN(n17072) );
  INV_X1 U18956 ( .A(keyinput_108), .ZN(n17070) );
  INV_X1 U18957 ( .A(keyinput_107), .ZN(n17068) );
  INV_X1 U18958 ( .A(keyinput_106), .ZN(n17065) );
  AOI22_X1 U18959 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(keyinput_103), .B1(n16996), 
        .B2(keyinput_104), .ZN(n16995) );
  OAI221_X1 U18960 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_103), .C1(n16996), 
        .C2(keyinput_104), .A(n16995), .ZN(n17062) );
  INV_X1 U18961 ( .A(keyinput_102), .ZN(n17060) );
  INV_X1 U18962 ( .A(DATAI_3_), .ZN(n17046) );
  OAI22_X1 U18963 ( .A1(n16999), .A2(keyinput_91), .B1(n16998), .B2(
        keyinput_92), .ZN(n16997) );
  AOI221_X1 U18964 ( .B1(n16999), .B2(keyinput_91), .C1(keyinput_92), .C2(
        n16998), .A(n16997), .ZN(n17044) );
  AOI22_X1 U18965 ( .A1(n17002), .A2(keyinput_78), .B1(n17001), .B2(
        keyinput_77), .ZN(n17000) );
  OAI221_X1 U18966 ( .B1(n17002), .B2(keyinput_78), .C1(n17001), .C2(
        keyinput_77), .A(n17000), .ZN(n17023) );
  INV_X1 U18967 ( .A(keyinput_76), .ZN(n17020) );
  INV_X1 U18968 ( .A(keyinput_75), .ZN(n17018) );
  OAI22_X1 U18969 ( .A1(DATAI_31_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n17003) );
  AOI221_X1 U18970 ( .B1(DATAI_31_), .B2(keyinput_65), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_64), .A(n17003), .ZN(n17008)
         );
  AOI22_X1 U18971 ( .A1(DATAI_29_), .A2(keyinput_67), .B1(DATAI_30_), .B2(
        keyinput_66), .ZN(n17004) );
  OAI221_X1 U18972 ( .B1(DATAI_29_), .B2(keyinput_67), .C1(DATAI_30_), .C2(
        keyinput_66), .A(n17004), .ZN(n17007) );
  OAI22_X1 U18973 ( .A1(DATAI_28_), .A2(keyinput_68), .B1(DATAI_27_), .B2(
        keyinput_69), .ZN(n17005) );
  AOI221_X1 U18974 ( .B1(DATAI_28_), .B2(keyinput_68), .C1(keyinput_69), .C2(
        DATAI_27_), .A(n17005), .ZN(n17006) );
  OAI21_X1 U18975 ( .B1(n17008), .B2(n17007), .A(n17006), .ZN(n17015) );
  XNOR2_X1 U18976 ( .A(DATAI_26_), .B(keyinput_70), .ZN(n17014) );
  AOI22_X1 U18977 ( .A1(DATAI_23_), .A2(keyinput_73), .B1(n17010), .B2(
        keyinput_72), .ZN(n17009) );
  OAI221_X1 U18978 ( .B1(DATAI_23_), .B2(keyinput_73), .C1(n17010), .C2(
        keyinput_72), .A(n17009), .ZN(n17013) );
  AOI22_X1 U18979 ( .A1(DATAI_22_), .A2(keyinput_74), .B1(DATAI_25_), .B2(
        keyinput_71), .ZN(n17011) );
  OAI221_X1 U18980 ( .B1(DATAI_22_), .B2(keyinput_74), .C1(DATAI_25_), .C2(
        keyinput_71), .A(n17011), .ZN(n17012) );
  AOI211_X1 U18981 ( .C1(n17015), .C2(n17014), .A(n17013), .B(n17012), .ZN(
        n17016) );
  AOI221_X1 U18982 ( .B1(DATAI_21_), .B2(n17018), .C1(n17017), .C2(keyinput_75), .A(n17016), .ZN(n17019) );
  AOI221_X1 U18983 ( .B1(DATAI_20_), .B2(keyinput_76), .C1(n17021), .C2(n17020), .A(n17019), .ZN(n17022) );
  OAI22_X1 U18984 ( .A1(n17023), .A2(n17022), .B1(DATAI_15_), .B2(keyinput_81), 
        .ZN(n17024) );
  AOI21_X1 U18985 ( .B1(DATAI_15_), .B2(keyinput_81), .A(n17024), .ZN(n17033)
         );
  OAI22_X1 U18986 ( .A1(n17026), .A2(keyinput_80), .B1(keyinput_79), .B2(
        DATAI_17_), .ZN(n17025) );
  AOI221_X1 U18987 ( .B1(n17026), .B2(keyinput_80), .C1(DATAI_17_), .C2(
        keyinput_79), .A(n17025), .ZN(n17032) );
  INV_X1 U18988 ( .A(DATAI_12_), .ZN(n17028) );
  AOI22_X1 U18989 ( .A1(DATAI_11_), .A2(keyinput_85), .B1(n17028), .B2(
        keyinput_84), .ZN(n17027) );
  OAI221_X1 U18990 ( .B1(DATAI_11_), .B2(keyinput_85), .C1(n17028), .C2(
        keyinput_84), .A(n17027), .ZN(n17031) );
  AOI22_X1 U18991 ( .A1(DATAI_13_), .A2(keyinput_83), .B1(DATAI_14_), .B2(
        keyinput_82), .ZN(n17029) );
  OAI221_X1 U18992 ( .B1(DATAI_13_), .B2(keyinput_83), .C1(DATAI_14_), .C2(
        keyinput_82), .A(n17029), .ZN(n17030) );
  AOI211_X1 U18993 ( .C1(n17033), .C2(n17032), .A(n17031), .B(n17030), .ZN(
        n17037) );
  AOI22_X1 U18994 ( .A1(DATAI_9_), .A2(keyinput_87), .B1(n17035), .B2(
        keyinput_86), .ZN(n17034) );
  OAI221_X1 U18995 ( .B1(DATAI_9_), .B2(keyinput_87), .C1(n17035), .C2(
        keyinput_86), .A(n17034), .ZN(n17036) );
  OAI22_X1 U18996 ( .A1(n17037), .A2(n17036), .B1(keyinput_88), .B2(n17041), 
        .ZN(n17042) );
  INV_X1 U18997 ( .A(DATAI_6_), .ZN(n17039) );
  OAI22_X1 U18998 ( .A1(n17039), .A2(keyinput_90), .B1(DATAI_7_), .B2(
        keyinput_89), .ZN(n17038) );
  AOI221_X1 U18999 ( .B1(n17039), .B2(keyinput_90), .C1(keyinput_89), .C2(
        DATAI_7_), .A(n17038), .ZN(n17040) );
  OAI221_X1 U19000 ( .B1(n17042), .B2(keyinput_88), .C1(n17042), .C2(n17041), 
        .A(n17040), .ZN(n17043) );
  AOI22_X1 U19001 ( .A1(n17044), .A2(n17043), .B1(keyinput_93), .B2(n17046), 
        .ZN(n17045) );
  OAI21_X1 U19002 ( .B1(keyinput_93), .B2(n17046), .A(n17045), .ZN(n17049) );
  AOI22_X1 U19003 ( .A1(DATAI_1_), .A2(keyinput_95), .B1(DATAI_2_), .B2(
        keyinput_94), .ZN(n17047) );
  OAI221_X1 U19004 ( .B1(DATAI_1_), .B2(keyinput_95), .C1(DATAI_2_), .C2(
        keyinput_94), .A(n17047), .ZN(n17048) );
  OAI22_X1 U19005 ( .A1(n17049), .A2(n17048), .B1(NA), .B2(keyinput_98), .ZN(
        n17050) );
  AOI21_X1 U19006 ( .B1(NA), .B2(keyinput_98), .A(n17050), .ZN(n17057) );
  OAI22_X1 U19007 ( .A1(DATAI_0_), .A2(keyinput_96), .B1(HOLD), .B2(
        keyinput_97), .ZN(n17051) );
  AOI221_X1 U19008 ( .B1(DATAI_0_), .B2(keyinput_96), .C1(keyinput_97), .C2(
        HOLD), .A(n17051), .ZN(n17056) );
  XOR2_X1 U19009 ( .A(READY2), .B(keyinput_101), .Z(n17055) );
  INV_X1 U19010 ( .A(READY1), .ZN(n17053) );
  AOI22_X1 U19011 ( .A1(BS16), .A2(keyinput_99), .B1(n17053), .B2(keyinput_100), .ZN(n17052) );
  OAI221_X1 U19012 ( .B1(BS16), .B2(keyinput_99), .C1(n17053), .C2(
        keyinput_100), .A(n17052), .ZN(n17054) );
  AOI211_X1 U19013 ( .C1(n17057), .C2(n17056), .A(n17055), .B(n17054), .ZN(
        n17058) );
  AOI221_X1 U19014 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(n17060), .C1(n17059), 
        .C2(keyinput_102), .A(n17058), .ZN(n17061) );
  OAI22_X1 U19015 ( .A1(keyinput_105), .A2(n22277), .B1(n17062), .B2(n17061), 
        .ZN(n17063) );
  AOI21_X1 U19016 ( .B1(keyinput_105), .B2(n22277), .A(n17063), .ZN(n17064) );
  AOI221_X1 U19017 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(n17065), .C1(n20026), .C2(
        keyinput_106), .A(n17064), .ZN(n17066) );
  AOI221_X1 U19018 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n17068), .C1(
        n17067), .C2(keyinput_107), .A(n17066), .ZN(n17069) );
  AOI221_X1 U19019 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_108), .C1(
        n14439), .C2(n17070), .A(n17069), .ZN(n17071) );
  AOI221_X1 U19020 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_109), .C1(n17073), 
        .C2(n17072), .A(n17071), .ZN(n17074) );
  AOI221_X1 U19021 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_110), .C1(n21640), 
        .C2(n17075), .A(n17074), .ZN(n17076) );
  AOI221_X1 U19022 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_111), .C1(n20095), 
        .C2(n17077), .A(n17076), .ZN(n17078) );
  OAI22_X1 U19023 ( .A1(keyinput_114), .A2(n19910), .B1(n17079), .B2(n17078), 
        .ZN(n17080) );
  AOI21_X1 U19024 ( .B1(keyinput_114), .B2(n19910), .A(n17080), .ZN(n17081) );
  AOI221_X1 U19025 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_115), 
        .C1(n19895), .C2(n17082), .A(n17081), .ZN(n17083) );
  OAI22_X1 U19026 ( .A1(n17084), .A2(n17083), .B1(keyinput_121), .B2(
        P1_REIP_REG_26__SCAN_IN), .ZN(n17085) );
  AOI21_X1 U19027 ( .B1(keyinput_121), .B2(P1_REIP_REG_26__SCAN_IN), .A(n17085), .ZN(n17086) );
  OAI22_X1 U19028 ( .A1(n17087), .A2(n17086), .B1(keyinput_124), .B2(
        P1_REIP_REG_23__SCAN_IN), .ZN(n17088) );
  AOI21_X1 U19029 ( .B1(keyinput_124), .B2(P1_REIP_REG_23__SCAN_IN), .A(n17088), .ZN(n17092) );
  XNOR2_X1 U19030 ( .A(P1_REIP_REG_22__SCAN_IN), .B(keyinput_125), .ZN(n17091)
         );
  AOI22_X1 U19031 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_127), .B1(
        n21592), .B2(keyinput_126), .ZN(n17089) );
  OAI221_X1 U19032 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_127), .C1(
        n21592), .C2(keyinput_126), .A(n17089), .ZN(n17090) );
  NOR4_X1 U19033 ( .A1(n17093), .A2(n17092), .A3(n17091), .A4(n17090), .ZN(
        n17094) );
  XNOR2_X1 U19034 ( .A(n17095), .B(n17094), .ZN(P1_U2927) );
  INV_X1 U19035 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17096) );
  OAI22_X1 U19036 ( .A1(n18221), .A2(n17096), .B1(n18596), .B2(n18604), .ZN(
        P2_U2816) );
  AOI22_X1 U19037 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n18559), .B1(n17163), 
        .B2(n17097), .ZN(n17105) );
  NAND3_X1 U19038 ( .A1(n17099), .A2(n17098), .A3(n17203), .ZN(n17100) );
  OAI21_X1 U19039 ( .B1(n17207), .B2(n17101), .A(n17100), .ZN(n17102) );
  AOI21_X1 U19040 ( .B1(n17103), .B2(n17202), .A(n17102), .ZN(n17104) );
  OAI211_X1 U19041 ( .C1(n17106), .C2(n17151), .A(n17105), .B(n17104), .ZN(
        P2_U3011) );
  AOI22_X1 U19042 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17200), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n18559), .ZN(n17111) );
  AOI222_X1 U19043 ( .A1(n17109), .A2(n17202), .B1(n17190), .B2(n17108), .C1(
        n17107), .C2(n17203), .ZN(n17110) );
  OAI211_X1 U19044 ( .C1(n17198), .C2(n17112), .A(n17111), .B(n17110), .ZN(
        P2_U3010) );
  AOI22_X1 U19045 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17200), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n18559), .ZN(n17119) );
  NOR2_X1 U19046 ( .A1(n17113), .A2(n17152), .ZN(n17117) );
  OAI22_X1 U19047 ( .A1(n17115), .A2(n17156), .B1(n17207), .B2(n17114), .ZN(
        n17116) );
  AOI21_X1 U19048 ( .B1(n17117), .B2(n16755), .A(n17116), .ZN(n17118) );
  OAI211_X1 U19049 ( .C1(n17198), .C2(n17120), .A(n17119), .B(n17118), .ZN(
        P2_U3008) );
  AOI22_X1 U19050 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17200), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18559), .ZN(n17133) );
  NAND2_X1 U19051 ( .A1(n17122), .A2(n17121), .ZN(n17127) );
  INV_X1 U19052 ( .A(n17123), .ZN(n17124) );
  AOI21_X1 U19053 ( .B1(n16480), .B2(n17125), .A(n17124), .ZN(n17126) );
  XOR2_X1 U19054 ( .A(n17127), .B(n17126), .Z(n18558) );
  OAI21_X1 U19055 ( .B1(n17130), .B2(n17129), .A(n17128), .ZN(n17131) );
  INV_X1 U19056 ( .A(n17131), .ZN(n18555) );
  AOI222_X1 U19057 ( .A1(n18558), .A2(n17202), .B1(n17190), .B2(n18557), .C1(
        n17203), .C2(n18555), .ZN(n17132) );
  OAI211_X1 U19058 ( .C1(n17198), .C2(n17134), .A(n17133), .B(n17132), .ZN(
        P2_U3006) );
  AOI22_X1 U19059 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17200), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n18559), .ZN(n17138) );
  AOI222_X1 U19060 ( .A1(n17136), .A2(n17202), .B1(n17190), .B2(n18292), .C1(
        n17203), .C2(n17135), .ZN(n17137) );
  OAI211_X1 U19061 ( .C1(n17198), .C2(n18290), .A(n17138), .B(n17137), .ZN(
        P2_U3004) );
  AOI22_X1 U19062 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17200), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18559), .ZN(n17144) );
  NAND2_X1 U19063 ( .A1(n11060), .A2(n17139), .ZN(n17140) );
  XNOR2_X1 U19064 ( .A(n17141), .B(n17140), .ZN(n18527) );
  AOI222_X1 U19065 ( .A1(n18527), .A2(n17202), .B1(n17190), .B2(n18526), .C1(
        n18525), .C2(n17203), .ZN(n17143) );
  OAI211_X1 U19066 ( .C1(n17198), .C2(n17145), .A(n17144), .B(n17143), .ZN(
        P2_U3002) );
  AOI22_X1 U19067 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n18559), .B1(n17163), 
        .B2(n18322), .ZN(n17150) );
  OAI22_X1 U19068 ( .A1(n17147), .A2(n17156), .B1(n17152), .B2(n17146), .ZN(
        n17148) );
  AOI21_X1 U19069 ( .B1(n17190), .B2(n18318), .A(n17148), .ZN(n17149) );
  OAI211_X1 U19070 ( .C1(n18330), .C2(n17151), .A(n17150), .B(n17149), .ZN(
        P2_U2999) );
  AOI22_X1 U19071 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17200), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n18559), .ZN(n17161) );
  NOR2_X1 U19072 ( .A1(n17153), .A2(n16642), .ZN(n17169) );
  AOI211_X1 U19073 ( .C1(n16642), .C2(n17153), .A(n17152), .B(n17169), .ZN(
        n17159) );
  INV_X1 U19074 ( .A(n17154), .ZN(n17157) );
  OAI22_X1 U19075 ( .A1(n17157), .A2(n17156), .B1(n17207), .B2(n17155), .ZN(
        n17158) );
  NOR2_X1 U19076 ( .A1(n17159), .A2(n17158), .ZN(n17160) );
  OAI211_X1 U19077 ( .C1(n17198), .C2(n17162), .A(n17161), .B(n17160), .ZN(
        P2_U2998) );
  AOI22_X1 U19078 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17200), .B1(
        n17163), .B2(n18333), .ZN(n17173) );
  AOI22_X1 U19079 ( .A1(n17164), .A2(n17202), .B1(n17190), .B2(n18339), .ZN(
        n17172) );
  INV_X1 U19080 ( .A(n17165), .ZN(n17166) );
  NOR2_X1 U19081 ( .A1(n17167), .A2(n17166), .ZN(n17179) );
  INV_X1 U19082 ( .A(n17179), .ZN(n17168) );
  OAI211_X1 U19083 ( .C1(n17169), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n17168), .B(n17203), .ZN(n17171) );
  NAND4_X1 U19084 ( .A1(n17173), .A2(n17172), .A3(n17171), .A4(n17170), .ZN(
        P2_U2997) );
  AOI22_X1 U19085 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17200), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n18559), .ZN(n17182) );
  NAND2_X1 U19086 ( .A1(n17175), .A2(n17174), .ZN(n17177) );
  XNOR2_X1 U19087 ( .A(n17177), .B(n17176), .ZN(n18549) );
  OAI21_X1 U19088 ( .B1(n17179), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17178), .ZN(n18552) );
  INV_X1 U19089 ( .A(n18552), .ZN(n17180) );
  AOI222_X1 U19090 ( .A1(n18549), .A2(n17202), .B1(n17203), .B2(n17180), .C1(
        n17190), .C2(n18548), .ZN(n17181) );
  OAI211_X1 U19091 ( .C1(n17198), .C2(n18344), .A(n17182), .B(n17181), .ZN(
        P2_U2996) );
  AOI22_X1 U19092 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17200), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18559), .ZN(n17188) );
  INV_X1 U19093 ( .A(n17184), .ZN(n17185) );
  AOI21_X1 U19094 ( .B1(n18538), .B2(n17186), .A(n17185), .ZN(n18534) );
  OAI211_X1 U19095 ( .C1(n17198), .C2(n18369), .A(n17188), .B(n17187), .ZN(
        P2_U2994) );
  AOI22_X1 U19096 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17200), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18559), .ZN(n17197) );
  NAND2_X1 U19097 ( .A1(n17189), .A2(n17203), .ZN(n17194) );
  AOI22_X1 U19098 ( .A1(n17191), .A2(n17202), .B1(n17190), .B2(n18393), .ZN(
        n17192) );
  OAI21_X1 U19099 ( .B1(n17194), .B2(n17193), .A(n17192), .ZN(n17195) );
  INV_X1 U19100 ( .A(n17195), .ZN(n17196) );
  OAI211_X1 U19101 ( .C1(n17198), .C2(n18395), .A(n17197), .B(n17196), .ZN(
        P2_U2992) );
  OAI22_X1 U19102 ( .A1(n15277), .A2(n14141), .B1(n17198), .B2(n18416), .ZN(
        n17199) );
  AOI21_X1 U19103 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17200), .A(
        n17199), .ZN(n17206) );
  AOI22_X1 U19104 ( .A1(n17204), .A2(n17203), .B1(n17202), .B2(n17201), .ZN(
        n17205) );
  OAI211_X1 U19105 ( .C1(n17207), .C2(n18413), .A(n17206), .B(n17205), .ZN(
        P2_U2990) );
  INV_X1 U19106 ( .A(n17228), .ZN(n17220) );
  NOR2_X1 U19107 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n17208), .ZN(n18220) );
  NOR2_X1 U19108 ( .A1(n17209), .A2(n19214), .ZN(n18612) );
  NOR2_X1 U19109 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n17222), .ZN(
        n17210) );
  OR2_X1 U19110 ( .A1(n18612), .A2(n17210), .ZN(n17211) );
  AOI21_X1 U19111 ( .B1(n19123), .B2(n18220), .A(n17211), .ZN(n17212) );
  AOI22_X1 U19112 ( .A1(n17220), .A2(n19288), .B1(n17212), .B2(n17228), .ZN(
        P2_U3605) );
  OR2_X1 U19113 ( .A1(n19142), .A2(n13854), .ZN(n19259) );
  AOI21_X1 U19114 ( .B1(n19259), .B2(n19304), .A(n17213), .ZN(n17223) );
  INV_X1 U19115 ( .A(n19259), .ZN(n17224) );
  NAND3_X1 U19116 ( .A1(n19238), .A2(n19304), .A3(n17224), .ZN(n17214) );
  OAI21_X1 U19117 ( .B1(n17223), .B2(n19238), .A(n17214), .ZN(n17215) );
  AOI21_X1 U19118 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19523), .A(n17215), 
        .ZN(n17216) );
  AOI22_X1 U19119 ( .A1(n17220), .A2(n19256), .B1(n17216), .B2(n17228), .ZN(
        P2_U3603) );
  NAND2_X1 U19120 ( .A1(n19304), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17217) );
  AOI21_X1 U19121 ( .B1(n19142), .B2(n17217), .A(n17223), .ZN(n17218) );
  AOI21_X1 U19122 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19575), .A(n17218), 
        .ZN(n17219) );
  AOI22_X1 U19123 ( .A1(n17220), .A2(n19260), .B1(n17219), .B2(n17228), .ZN(
        P2_U3604) );
  OAI22_X1 U19124 ( .A1(n19239), .A2(n17223), .B1(n17222), .B2(n17221), .ZN(
        n17226) );
  NAND2_X1 U19125 ( .A1(n19225), .A2(n17224), .ZN(n19203) );
  INV_X1 U19126 ( .A(n19178), .ZN(n19179) );
  AOI21_X1 U19127 ( .B1(n19203), .B2(n19179), .A(n19290), .ZN(n17225) );
  OAI21_X1 U19128 ( .B1(n17226), .B2(n17225), .A(n17228), .ZN(n17227) );
  OAI21_X1 U19129 ( .B1(n17228), .B2(n19255), .A(n17227), .ZN(P2_U3602) );
  INV_X1 U19130 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21670) );
  NAND2_X1 U19131 ( .A1(n17229), .A2(n21670), .ZN(n17232) );
  OAI21_X1 U19132 ( .B1(n13869), .B2(n18240), .A(n17235), .ZN(n17230) );
  OAI21_X1 U19133 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17235), .A(n17230), 
        .ZN(n17231) );
  OAI221_X1 U19134 ( .B1(n17232), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17232), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17231), .ZN(P2_U2822) );
  INV_X1 U19135 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17290) );
  OAI221_X1 U19136 ( .B1(n17235), .B2(n17290), .C1(n17234), .C2(n17233), .A(
        n17232), .ZN(P2_U2823) );
  INV_X1 U19137 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n17236) );
  AOI22_X1 U19138 ( .A1(n17281), .A2(n17237), .B1(n17236), .B2(n21702), .ZN(
        P2_U3611) );
  INV_X1 U19139 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17238) );
  AOI22_X1 U19140 ( .A1(n17281), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17238), 
        .B2(n21702), .ZN(P2_U3608) );
  INV_X1 U19141 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n17240) );
  OAI21_X1 U19142 ( .B1(n17269), .B2(n17240), .A(n17239), .ZN(P2_U2815) );
  AOI22_X1 U19143 ( .A1(n17265), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17254), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17242) );
  OAI21_X1 U19144 ( .B1(n13593), .B2(n17267), .A(n17242), .ZN(P2_U2951) );
  INV_X1 U19145 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17244) );
  AOI22_X1 U19146 ( .A1(n17265), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17254), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17243) );
  OAI21_X1 U19147 ( .B1(n17244), .B2(n17267), .A(n17243), .ZN(P2_U2950) );
  INV_X1 U19148 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19530) );
  AOI22_X1 U19149 ( .A1(n17265), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17254), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17245) );
  OAI21_X1 U19150 ( .B1(n19530), .B2(n17267), .A(n17245), .ZN(P2_U2949) );
  INV_X1 U19151 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U19152 ( .A1(n17256), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17246) );
  OAI21_X1 U19153 ( .B1(n17247), .B2(n17267), .A(n17246), .ZN(P2_U2948) );
  INV_X1 U19154 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17249) );
  AOI22_X1 U19155 ( .A1(n17265), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17254), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17248) );
  OAI21_X1 U19156 ( .B1(n17249), .B2(n17267), .A(n17248), .ZN(P2_U2947) );
  INV_X1 U19157 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19370) );
  AOI22_X1 U19158 ( .A1(n17256), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17254), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17250) );
  OAI21_X1 U19159 ( .B1(n19370), .B2(n17267), .A(n17250), .ZN(P2_U2946) );
  INV_X1 U19160 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19327) );
  AOI22_X1 U19161 ( .A1(n17256), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17251) );
  OAI21_X1 U19162 ( .B1(n19327), .B2(n17267), .A(n17251), .ZN(P2_U2945) );
  INV_X1 U19163 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19106) );
  AOI22_X1 U19164 ( .A1(n17256), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17254), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17252) );
  OAI21_X1 U19165 ( .B1(n19106), .B2(n17267), .A(n17252), .ZN(P2_U2944) );
  INV_X1 U19166 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19104) );
  AOI22_X1 U19167 ( .A1(n17256), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17254), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17253) );
  OAI21_X1 U19168 ( .B1(n19104), .B2(n17267), .A(n17253), .ZN(P2_U2943) );
  INV_X1 U19169 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19100) );
  AOI22_X1 U19170 ( .A1(n17265), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17254), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17255) );
  OAI21_X1 U19171 ( .B1(n19100), .B2(n17267), .A(n17255), .ZN(P2_U2942) );
  INV_X1 U19172 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19097) );
  AOI22_X1 U19173 ( .A1(n17256), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17257) );
  OAI21_X1 U19174 ( .B1(n19097), .B2(n17267), .A(n17257), .ZN(P2_U2941) );
  INV_X1 U19175 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19094) );
  AOI22_X1 U19176 ( .A1(n17265), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17258) );
  OAI21_X1 U19177 ( .B1(n19094), .B2(n17267), .A(n17258), .ZN(P2_U2940) );
  AOI22_X1 U19178 ( .A1(n17265), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17259) );
  OAI21_X1 U19179 ( .B1(n17260), .B2(n17267), .A(n17259), .ZN(P2_U2939) );
  INV_X1 U19180 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19088) );
  AOI22_X1 U19181 ( .A1(n17265), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17261) );
  OAI21_X1 U19182 ( .B1(n19088), .B2(n17267), .A(n17261), .ZN(P2_U2938) );
  AOI22_X1 U19183 ( .A1(n17265), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17262) );
  OAI21_X1 U19184 ( .B1(n17263), .B2(n17267), .A(n17262), .ZN(P2_U2937) );
  AOI22_X1 U19185 ( .A1(n17265), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17264), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17266) );
  OAI21_X1 U19186 ( .B1(n19080), .B2(n17267), .A(n17266), .ZN(P2_U2936) );
  AOI21_X1 U19187 ( .B1(n17269), .B2(n17268), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n17270) );
  AOI21_X1 U19188 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n17281), .A(n17270), 
        .ZN(P2_U2817) );
  AND2_X1 U19189 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17281), .ZN(n21704) );
  OAI222_X1 U19190 ( .A1(n17284), .A2(n18577), .B1(n19757), .B2(n17281), .C1(
        n13869), .C2(n10969), .ZN(P2_U3212) );
  INV_X1 U19191 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19759) );
  OAI222_X1 U19192 ( .A1(n17284), .A2(n13662), .B1(n19759), .B2(n17281), .C1(
        n18577), .C2(n10969), .ZN(P2_U3213) );
  INV_X1 U19193 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19761) );
  OAI222_X1 U19194 ( .A1(n17284), .A2(n13663), .B1(n19761), .B2(n17281), .C1(
        n13662), .C2(n10969), .ZN(P2_U3214) );
  INV_X1 U19195 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19763) );
  OAI222_X1 U19196 ( .A1(n17284), .A2(n17271), .B1(n19763), .B2(n17281), .C1(
        n13663), .C2(n10969), .ZN(P2_U3215) );
  INV_X1 U19197 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19765) );
  OAI222_X1 U19198 ( .A1(n17284), .A2(n17272), .B1(n19765), .B2(n17281), .C1(
        n17271), .C2(n10969), .ZN(P2_U3216) );
  INV_X1 U19199 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19767) );
  OAI222_X1 U19200 ( .A1(n17284), .A2(n18265), .B1(n19767), .B2(n17281), .C1(
        n17272), .C2(n10969), .ZN(P2_U3217) );
  INV_X1 U19201 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n17273) );
  INV_X1 U19202 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19769) );
  OAI222_X1 U19203 ( .A1(n17284), .A2(n17273), .B1(n19769), .B2(n17281), .C1(
        n18265), .C2(n10969), .ZN(P2_U3218) );
  INV_X1 U19204 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19771) );
  OAI222_X1 U19205 ( .A1(n17284), .A2(n14704), .B1(n19771), .B2(n17281), .C1(
        n17273), .C2(n10969), .ZN(P2_U3219) );
  INV_X1 U19206 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19773) );
  OAI222_X1 U19207 ( .A1(n10969), .A2(n14704), .B1(n19773), .B2(n17281), .C1(
        n13733), .C2(n17284), .ZN(P2_U3220) );
  INV_X1 U19208 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19775) );
  OAI222_X1 U19209 ( .A1(n10969), .A2(n13733), .B1(n19775), .B2(n17281), .C1(
        n16457), .C2(n17284), .ZN(P2_U3221) );
  INV_X1 U19210 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19777) );
  OAI222_X1 U19211 ( .A1(n10969), .A2(n16457), .B1(n19777), .B2(n17281), .C1(
        n16143), .C2(n17284), .ZN(P2_U3222) );
  INV_X1 U19212 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19779) );
  OAI222_X1 U19213 ( .A1(n10969), .A2(n16143), .B1(n19779), .B2(n17281), .C1(
        n16453), .C2(n17284), .ZN(P2_U3223) );
  INV_X1 U19214 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19781) );
  OAI222_X1 U19215 ( .A1(n10969), .A2(n16453), .B1(n19781), .B2(n17281), .C1(
        n17274), .C2(n17284), .ZN(P2_U3224) );
  INV_X1 U19216 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19783) );
  OAI222_X1 U19217 ( .A1(n10969), .A2(n17274), .B1(n19783), .B2(n17281), .C1(
        n14969), .C2(n17284), .ZN(P2_U3225) );
  INV_X1 U19218 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19785) );
  OAI222_X1 U19219 ( .A1(n10969), .A2(n14969), .B1(n19785), .B2(n17281), .C1(
        n15174), .C2(n17284), .ZN(P2_U3226) );
  INV_X1 U19220 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19787) );
  OAI222_X1 U19221 ( .A1(n10969), .A2(n15174), .B1(n19787), .B2(n17281), .C1(
        n17275), .C2(n17284), .ZN(P2_U3227) );
  INV_X1 U19222 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19789) );
  OAI222_X1 U19223 ( .A1(n10969), .A2(n17275), .B1(n19789), .B2(n17281), .C1(
        n15252), .C2(n17284), .ZN(P2_U3228) );
  INV_X1 U19224 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19791) );
  OAI222_X1 U19225 ( .A1(n17284), .A2(n17276), .B1(n19791), .B2(n17281), .C1(
        n15252), .C2(n10969), .ZN(P2_U3229) );
  INV_X1 U19226 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19793) );
  OAI222_X1 U19227 ( .A1(n10969), .A2(n17276), .B1(n19793), .B2(n17281), .C1(
        n15260), .C2(n17284), .ZN(P2_U3230) );
  INV_X1 U19228 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19795) );
  OAI222_X1 U19229 ( .A1(n17284), .A2(n17277), .B1(n19795), .B2(n17281), .C1(
        n15260), .C2(n10969), .ZN(P2_U3231) );
  INV_X1 U19230 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19797) );
  OAI222_X1 U19231 ( .A1(n17284), .A2(n15269), .B1(n19797), .B2(n17281), .C1(
        n17277), .C2(n10969), .ZN(P2_U3232) );
  INV_X1 U19232 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19799) );
  OAI222_X1 U19233 ( .A1(n17284), .A2(n17278), .B1(n19799), .B2(n17281), .C1(
        n15269), .C2(n10969), .ZN(P2_U3233) );
  INV_X1 U19234 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19801) );
  OAI222_X1 U19235 ( .A1(n17284), .A2(n15277), .B1(n19801), .B2(n17281), .C1(
        n17278), .C2(n10969), .ZN(P2_U3234) );
  INV_X1 U19236 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19803) );
  OAI222_X1 U19237 ( .A1(n17284), .A2(n17279), .B1(n19803), .B2(n17281), .C1(
        n15277), .C2(n10969), .ZN(P2_U3235) );
  INV_X1 U19238 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19806) );
  OAI222_X1 U19239 ( .A1(n10969), .A2(n17279), .B1(n19806), .B2(n17281), .C1(
        n17280), .C2(n17284), .ZN(P2_U3236) );
  INV_X1 U19240 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19808) );
  OAI222_X1 U19241 ( .A1(n17284), .A2(n18448), .B1(n19808), .B2(n17281), .C1(
        n17280), .C2(n10969), .ZN(P2_U3237) );
  INV_X1 U19242 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19810) );
  OAI222_X1 U19243 ( .A1(n10969), .A2(n18448), .B1(n19810), .B2(n17281), .C1(
        n15291), .C2(n17284), .ZN(P2_U3238) );
  INV_X1 U19244 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19812) );
  OAI222_X1 U19245 ( .A1(n10969), .A2(n15291), .B1(n19812), .B2(n17281), .C1(
        n17282), .C2(n17284), .ZN(P2_U3239) );
  INV_X1 U19246 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19814) );
  OAI222_X1 U19247 ( .A1(n10969), .A2(n17282), .B1(n19814), .B2(n17281), .C1(
        n17283), .C2(n17284), .ZN(P2_U3240) );
  INV_X1 U19248 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19817) );
  OAI222_X1 U19249 ( .A1(n17284), .A2(n18492), .B1(n19817), .B2(n17281), .C1(
        n17283), .C2(n10969), .ZN(P2_U3241) );
  INV_X1 U19250 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n17285) );
  AOI22_X1 U19251 ( .A1(n17281), .A2(n17286), .B1(n17285), .B2(n21702), .ZN(
        P2_U3588) );
  INV_X1 U19252 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U19253 ( .A1(n17281), .A2(n17288), .B1(n17287), .B2(n21702), .ZN(
        P2_U3587) );
  MUX2_X1 U19254 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n17281), .Z(P2_U3586) );
  INV_X1 U19255 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U19256 ( .A1(n17281), .A2(n17290), .B1(n17289), .B2(n21702), .ZN(
        P2_U3585) );
  NAND3_X1 U19257 ( .A1(n20667), .A2(n18811), .A3(n17291), .ZN(n17292) );
  NAND3_X1 U19258 ( .A1(n20595), .A2(n12661), .A3(n20592), .ZN(n17684) );
  INV_X1 U19259 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20173) );
  NAND2_X1 U19260 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17300) );
  NOR2_X1 U19261 ( .A1(n20173), .A2(n17300), .ZN(n17294) );
  NAND3_X1 U19262 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17294), .ZN(n17434) );
  NOR2_X1 U19263 ( .A1(n17684), .A2(n17434), .ZN(n17322) );
  INV_X1 U19264 ( .A(n17322), .ZN(n17313) );
  NOR2_X1 U19265 ( .A1(n20693), .A2(n17313), .ZN(n17320) );
  INV_X2 U19266 ( .A(n17685), .ZN(n17682) );
  NAND2_X1 U19267 ( .A1(n20667), .A2(n17438), .ZN(n17687) );
  INV_X1 U19268 ( .A(n17687), .ZN(n17680) );
  NAND2_X1 U19269 ( .A1(n17294), .A2(n17680), .ZN(n17301) );
  NOR2_X1 U19270 ( .A1(n20190), .A2(n17301), .ZN(n17299) );
  AOI21_X1 U19271 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17682), .A(n17299), .ZN(
        n17296) );
  OAI22_X1 U19272 ( .A1(n17320), .A2(n17296), .B1(n17295), .B2(n17682), .ZN(
        P3_U2699) );
  INV_X1 U19273 ( .A(n17301), .ZN(n17297) );
  AOI21_X1 U19274 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17682), .A(n17297), .ZN(
        n17298) );
  OAI22_X1 U19275 ( .A1(n17299), .A2(n17298), .B1(n17509), .B2(n17682), .ZN(
        P3_U2700) );
  INV_X1 U19276 ( .A(n17300), .ZN(n17679) );
  OAI221_X1 U19277 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n17438), .C1(
        P3_EBX_REG_2__SCAN_IN), .C2(n17679), .A(n17301), .ZN(n17302) );
  AOI22_X1 U19278 ( .A1(n17685), .A2(n17405), .B1(n17302), .B2(n17682), .ZN(
        P3_U2701) );
  AOI22_X1 U19279 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17306) );
  AOI22_X1 U19280 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17656), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17305) );
  AOI22_X1 U19281 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17304) );
  AOI22_X1 U19282 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17303) );
  NAND4_X1 U19283 ( .A1(n17306), .A2(n17305), .A3(n17304), .A4(n17303), .ZN(
        n17312) );
  AOI22_X1 U19284 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U19285 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U19286 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U19287 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17307) );
  NAND4_X1 U19288 ( .A1(n17310), .A2(n17309), .A3(n17308), .A4(n17307), .ZN(
        n17311) );
  NOR2_X1 U19289 ( .A1(n17312), .A2(n17311), .ZN(n20766) );
  NAND3_X1 U19290 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n17435) );
  NOR2_X1 U19291 ( .A1(n17435), .A2(n17313), .ZN(n17317) );
  OAI21_X1 U19292 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17317), .A(n17682), .ZN(
        n17314) );
  OAI22_X1 U19293 ( .A1(n20766), .A2(n17682), .B1(n17431), .B2(n17314), .ZN(
        P3_U2695) );
  AND3_X1 U19294 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17320), .ZN(n17319) );
  AOI21_X1 U19295 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17682), .A(n17319), .ZN(
        n17316) );
  OAI22_X1 U19296 ( .A1(n17317), .A2(n17316), .B1(n17315), .B2(n17682), .ZN(
        P3_U2696) );
  AOI22_X1 U19297 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17682), .B1(
        P3_EBX_REG_5__SCAN_IN), .B2(n17320), .ZN(n17318) );
  OAI22_X1 U19298 ( .A1(n17319), .A2(n17318), .B1(n17597), .B2(n17682), .ZN(
        P3_U2697) );
  NAND2_X1 U19299 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17320), .ZN(n17321) );
  OAI21_X1 U19300 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17322), .A(n17321), .ZN(
        n17323) );
  AOI22_X1 U19301 ( .A1(n17685), .A2(n17522), .B1(n17323), .B2(n17682), .ZN(
        P3_U2698) );
  INV_X1 U19302 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20358) );
  INV_X1 U19303 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20336) );
  INV_X1 U19304 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17363) );
  INV_X1 U19305 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20304) );
  NOR3_X1 U19306 ( .A1(n20336), .A2(n17363), .A3(n20304), .ZN(n17437) );
  NAND2_X1 U19307 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17431), .ZN(n17430) );
  INV_X1 U19308 ( .A(n17430), .ZN(n17417) );
  NAND2_X1 U19309 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17417), .ZN(n17416) );
  INV_X1 U19310 ( .A(n17416), .ZN(n17401) );
  NAND3_X1 U19311 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17437), .A3(n17401), 
        .ZN(n17348) );
  NOR2_X1 U19312 ( .A1(n20358), .A2(n17348), .ZN(n17324) );
  NAND2_X1 U19313 ( .A1(n20667), .A2(n17324), .ZN(n17337) );
  NOR2_X1 U19314 ( .A1(n17685), .A2(n17324), .ZN(n17349) );
  AOI22_X1 U19315 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17656), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17335) );
  AOI22_X1 U19316 ( .A1(n12529), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U19317 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17325) );
  OAI21_X1 U19318 ( .B1(n17598), .B2(n17326), .A(n17325), .ZN(n17332) );
  AOI22_X1 U19319 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U19320 ( .A1(n10980), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U19321 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U19322 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17327) );
  NAND4_X1 U19323 ( .A1(n17330), .A2(n17329), .A3(n17328), .A4(n17327), .ZN(
        n17331) );
  AOI211_X1 U19324 ( .C1(n17668), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n17332), .B(n17331), .ZN(n17333) );
  NAND3_X1 U19325 ( .A1(n17335), .A2(n17334), .A3(n17333), .ZN(n20742) );
  AOI22_X1 U19326 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17349), .B1(n17685), 
        .B2(n20742), .ZN(n17336) );
  OAI21_X1 U19327 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17337), .A(n17336), .ZN(
        P3_U2687) );
  AOI22_X1 U19328 ( .A1(n12529), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17341) );
  AOI22_X1 U19329 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17640), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17340) );
  AOI22_X1 U19330 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17339) );
  AOI22_X1 U19331 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17338) );
  NAND4_X1 U19332 ( .A1(n17341), .A2(n17340), .A3(n17339), .A4(n17338), .ZN(
        n17347) );
  AOI22_X1 U19333 ( .A1(n10980), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17345) );
  AOI22_X1 U19334 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17344) );
  AOI22_X1 U19335 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17343) );
  AOI22_X1 U19336 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17342) );
  NAND4_X1 U19337 ( .A1(n17345), .A2(n17344), .A3(n17343), .A4(n17342), .ZN(
        n17346) );
  NOR2_X1 U19338 ( .A1(n17347), .A2(n17346), .ZN(n20760) );
  INV_X1 U19339 ( .A(n17348), .ZN(n17350) );
  OAI21_X1 U19340 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17350), .A(n17349), .ZN(
        n17351) );
  OAI21_X1 U19341 ( .B1(n20760), .B2(n17682), .A(n17351), .ZN(P3_U2688) );
  AOI22_X1 U19342 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17362) );
  AOI22_X1 U19343 ( .A1(n12529), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12465), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17361) );
  AOI22_X1 U19344 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17352) );
  OAI21_X1 U19345 ( .B1(n17406), .B2(n17522), .A(n17352), .ZN(n17359) );
  AOI22_X1 U19346 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17536), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U19347 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17356) );
  AOI22_X1 U19348 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17640), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17355) );
  AOI22_X1 U19349 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17354) );
  NAND4_X1 U19350 ( .A1(n17357), .A2(n17356), .A3(n17355), .A4(n17354), .ZN(
        n17358) );
  AOI211_X1 U19351 ( .C1(n17657), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n17359), .B(n17358), .ZN(n17360) );
  NAND3_X1 U19352 ( .A1(n17362), .A2(n17361), .A3(n17360), .ZN(n20603) );
  INV_X1 U19353 ( .A(n20603), .ZN(n17365) );
  NOR3_X1 U19354 ( .A1(n17416), .A2(n17363), .A3(n20304), .ZN(n17390) );
  AOI21_X1 U19355 ( .B1(n17437), .B2(n17401), .A(n17685), .ZN(n17376) );
  OAI21_X1 U19356 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17390), .A(n17376), .ZN(
        n17364) );
  OAI21_X1 U19357 ( .B1(n17365), .B2(n17682), .A(n17364), .ZN(P3_U2690) );
  NAND3_X1 U19358 ( .A1(n20667), .A2(n17437), .A3(n17401), .ZN(n17378) );
  AOI22_X1 U19359 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17375) );
  AOI22_X1 U19360 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10980), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17374) );
  AOI22_X1 U19361 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17366) );
  OAI21_X1 U19362 ( .B1(n17406), .B2(n17597), .A(n17366), .ZN(n17372) );
  AOI22_X1 U19363 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17536), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17370) );
  AOI22_X1 U19364 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U19365 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17368) );
  AOI22_X1 U19366 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17640), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17367) );
  NAND4_X1 U19367 ( .A1(n17370), .A2(n17369), .A3(n17368), .A4(n17367), .ZN(
        n17371) );
  AOI211_X1 U19368 ( .C1(n17489), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17372), .B(n17371), .ZN(n17373) );
  NAND3_X1 U19369 ( .A1(n17375), .A2(n17374), .A3(n17373), .ZN(n20750) );
  AOI22_X1 U19370 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17376), .B1(n17685), 
        .B2(n20750), .ZN(n17377) );
  OAI21_X1 U19371 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17378), .A(n17377), .ZN(
        P3_U2689) );
  NOR2_X1 U19372 ( .A1(n20304), .A2(n17416), .ZN(n17403) );
  OAI21_X1 U19373 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17403), .A(n17682), .ZN(
        n17389) );
  AOI22_X1 U19374 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17667), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U19375 ( .A1(n17664), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U19376 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17627), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U19377 ( .A1(n17659), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17379) );
  NAND4_X1 U19378 ( .A1(n17382), .A2(n17381), .A3(n17380), .A4(n17379), .ZN(
        n17388) );
  AOI22_X1 U19379 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U19380 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U19381 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U19382 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10980), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17383) );
  NAND4_X1 U19383 ( .A1(n17386), .A2(n17385), .A3(n17384), .A4(n17383), .ZN(
        n17387) );
  NOR2_X1 U19384 ( .A1(n17388), .A2(n17387), .ZN(n20607) );
  OAI22_X1 U19385 ( .A1(n17390), .A2(n17389), .B1(n20607), .B2(n17682), .ZN(
        P3_U2691) );
  AOI22_X1 U19386 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17394) );
  AOI22_X1 U19387 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17393) );
  AOI22_X1 U19388 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U19389 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17391) );
  NAND4_X1 U19390 ( .A1(n17394), .A2(n17393), .A3(n17392), .A4(n17391), .ZN(
        n17400) );
  AOI22_X1 U19391 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17398) );
  AOI22_X1 U19392 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17668), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U19393 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U19394 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17395) );
  NAND4_X1 U19395 ( .A1(n17398), .A2(n17397), .A3(n17396), .A4(n17395), .ZN(
        n17399) );
  NOR2_X1 U19396 ( .A1(n17400), .A2(n17399), .ZN(n20611) );
  OAI21_X1 U19397 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17401), .A(n17682), .ZN(
        n17402) );
  OAI22_X1 U19398 ( .A1(n20611), .A2(n17682), .B1(n17403), .B2(n17402), .ZN(
        P3_U2692) );
  AOI22_X1 U19399 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17415) );
  AOI22_X1 U19400 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17536), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17414) );
  AOI22_X1 U19401 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17404) );
  OAI21_X1 U19402 ( .B1(n17406), .B2(n17405), .A(n17404), .ZN(n17412) );
  AOI22_X1 U19403 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U19404 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17409) );
  AOI22_X1 U19405 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U19406 ( .A1(n17353), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17407) );
  NAND4_X1 U19407 ( .A1(n17410), .A2(n17409), .A3(n17408), .A4(n17407), .ZN(
        n17411) );
  AOI211_X1 U19408 ( .C1(n17656), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n17412), .B(n17411), .ZN(n17413) );
  NAND3_X1 U19409 ( .A1(n17415), .A2(n17414), .A3(n17413), .ZN(n20615) );
  INV_X1 U19410 ( .A(n20615), .ZN(n17419) );
  OAI21_X1 U19411 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17417), .A(n17416), .ZN(
        n17418) );
  AOI22_X1 U19412 ( .A1(n17685), .A2(n17419), .B1(n17418), .B2(n17682), .ZN(
        P3_U2693) );
  AOI22_X1 U19413 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17423) );
  AOI22_X1 U19414 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17664), .B1(
        n17668), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U19415 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17667), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17421) );
  AOI22_X1 U19416 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17627), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17628), .ZN(n17420) );
  NAND4_X1 U19417 ( .A1(n17423), .A2(n17422), .A3(n17421), .A4(n17420), .ZN(
        n17429) );
  AOI22_X1 U19418 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17642), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n10970), .ZN(n17427) );
  AOI22_X1 U19419 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17426) );
  AOI22_X1 U19420 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17425) );
  AOI22_X1 U19421 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17424) );
  NAND4_X1 U19422 ( .A1(n17427), .A2(n17426), .A3(n17425), .A4(n17424), .ZN(
        n17428) );
  NOR2_X1 U19423 ( .A1(n17429), .A2(n17428), .ZN(n20620) );
  OAI21_X1 U19424 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17431), .A(n17430), .ZN(
        n17432) );
  AOI22_X1 U19425 ( .A1(n17685), .A2(n20620), .B1(n17432), .B2(n17682), .ZN(
        P3_U2694) );
  INV_X1 U19426 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n20576) );
  INV_X1 U19427 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n20423) );
  INV_X1 U19428 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20390) );
  NAND4_X1 U19429 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_14__SCAN_IN), .A4(P3_EBX_REG_10__SCAN_IN), .ZN(n17433)
         );
  NOR3_X1 U19430 ( .A1(n17435), .A2(n17434), .A3(n17433), .ZN(n17436) );
  NAND4_X1 U19431 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n17437), .A4(n17436), .ZN(n17676) );
  NOR2_X1 U19432 ( .A1(n20390), .A2(n17676), .ZN(n17675) );
  NAND2_X1 U19433 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17654), .ZN(n17653) );
  INV_X1 U19434 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n20495) );
  INV_X1 U19435 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17560) );
  INV_X1 U19436 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20437) );
  NAND4_X1 U19437 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_28__SCAN_IN), 
        .A3(P3_EBX_REG_27__SCAN_IN), .A4(P3_EBX_REG_26__SCAN_IN), .ZN(n17439)
         );
  NOR4_X1 U19438 ( .A1(n20495), .A2(n17560), .A3(n20437), .A4(n17439), .ZN(
        n17440) );
  NAND4_X1 U19439 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n17546), .A4(n17440), .ZN(n17443) );
  NOR2_X1 U19440 ( .A1(n20576), .A2(n17443), .ZN(n17545) );
  NAND2_X1 U19441 ( .A1(n17682), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17442) );
  NAND2_X1 U19442 ( .A1(n17545), .A2(n20667), .ZN(n17441) );
  OAI22_X1 U19443 ( .A1(n17545), .A2(n17442), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17441), .ZN(P3_U2672) );
  NAND2_X1 U19444 ( .A1(n20576), .A2(n17443), .ZN(n17444) );
  NAND2_X1 U19445 ( .A1(n17444), .A2(n17682), .ZN(n17544) );
  AOI22_X1 U19446 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U19447 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17447) );
  AOI22_X1 U19448 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17446) );
  AOI22_X1 U19449 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17445) );
  NAND4_X1 U19450 ( .A1(n17448), .A2(n17447), .A3(n17446), .A4(n17445), .ZN(
        n17454) );
  AOI22_X1 U19451 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U19452 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U19453 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17667), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17450) );
  AOI22_X1 U19454 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17449) );
  NAND4_X1 U19455 ( .A1(n17452), .A2(n17451), .A3(n17450), .A4(n17449), .ZN(
        n17453) );
  NOR2_X1 U19456 ( .A1(n17454), .A2(n17453), .ZN(n17566) );
  AOI22_X1 U19457 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U19458 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17457) );
  AOI22_X1 U19459 ( .A1(n17664), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U19460 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17455) );
  NAND4_X1 U19461 ( .A1(n17458), .A2(n17457), .A3(n17456), .A4(n17455), .ZN(
        n17464) );
  AOI22_X1 U19462 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U19463 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17667), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17461) );
  AOI22_X1 U19464 ( .A1(n10980), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U19465 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17459) );
  NAND4_X1 U19466 ( .A1(n17462), .A2(n17461), .A3(n17460), .A4(n17459), .ZN(
        n17463) );
  NOR2_X1 U19467 ( .A1(n17464), .A2(n17463), .ZN(n17561) );
  AOI22_X1 U19468 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U19469 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17467) );
  AOI22_X1 U19470 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17466) );
  AOI22_X1 U19471 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17465) );
  NAND4_X1 U19472 ( .A1(n17468), .A2(n17467), .A3(n17466), .A4(n17465), .ZN(
        n17474) );
  AOI22_X1 U19473 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17472) );
  AOI22_X1 U19474 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17667), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17471) );
  AOI22_X1 U19475 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17470) );
  AOI22_X1 U19476 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17469) );
  NAND4_X1 U19477 ( .A1(n17472), .A2(n17471), .A3(n17470), .A4(n17469), .ZN(
        n17473) );
  NOR2_X1 U19478 ( .A1(n17474), .A2(n17473), .ZN(n17581) );
  AOI22_X1 U19479 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U19480 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17477) );
  AOI22_X1 U19481 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U19482 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17475) );
  NAND4_X1 U19483 ( .A1(n17478), .A2(n17477), .A3(n17476), .A4(n17475), .ZN(
        n17484) );
  AOI22_X1 U19484 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17657), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U19485 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17481) );
  AOI22_X1 U19486 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17480) );
  AOI22_X1 U19487 ( .A1(n17659), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17479) );
  NAND4_X1 U19488 ( .A1(n17482), .A2(n17481), .A3(n17480), .A4(n17479), .ZN(
        n17483) );
  NOR2_X1 U19489 ( .A1(n17484), .A2(n17483), .ZN(n17590) );
  AOI22_X1 U19490 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17488) );
  AOI22_X1 U19491 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17487) );
  AOI22_X1 U19492 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17627), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17486) );
  AOI22_X1 U19493 ( .A1(n17659), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17485) );
  NAND4_X1 U19494 ( .A1(n17488), .A2(n17487), .A3(n17486), .A4(n17485), .ZN(
        n17495) );
  AOI22_X1 U19495 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17493) );
  AOI22_X1 U19496 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17536), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U19497 ( .A1(n17641), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17491) );
  AOI22_X1 U19498 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17667), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17490) );
  NAND4_X1 U19499 ( .A1(n17493), .A2(n17492), .A3(n17491), .A4(n17490), .ZN(
        n17494) );
  NOR2_X1 U19500 ( .A1(n17495), .A2(n17494), .ZN(n17591) );
  NOR2_X1 U19501 ( .A1(n17590), .A2(n17591), .ZN(n17589) );
  AOI22_X1 U19502 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17656), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17507) );
  AOI22_X1 U19503 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17657), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17666), .ZN(n17506) );
  INV_X1 U19504 ( .A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17497) );
  AOI22_X1 U19505 ( .A1(n10980), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17628), .ZN(n17496) );
  OAI21_X1 U19506 ( .B1(n17497), .B2(n20196), .A(n17496), .ZN(n17504) );
  AOI22_X1 U19507 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17664), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17659), .ZN(n17502) );
  AOI22_X1 U19508 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17498), .ZN(n17501) );
  AOI22_X1 U19509 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17536), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17500) );
  AOI22_X1 U19510 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10970), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17499) );
  NAND4_X1 U19511 ( .A1(n17502), .A2(n17501), .A3(n17500), .A4(n17499), .ZN(
        n17503) );
  AOI211_X1 U19512 ( .C1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .C2(n17640), .A(
        n17504), .B(n17503), .ZN(n17505) );
  NAND3_X1 U19513 ( .A1(n17507), .A2(n17506), .A3(n17505), .ZN(n17586) );
  NAND2_X1 U19514 ( .A1(n17589), .A2(n17586), .ZN(n17585) );
  NOR2_X1 U19515 ( .A1(n17581), .A2(n17585), .ZN(n17580) );
  AOI22_X1 U19516 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17519) );
  AOI22_X1 U19517 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17518) );
  AOI22_X1 U19518 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17508) );
  OAI21_X1 U19519 ( .B1(n12572), .B2(n17509), .A(n17508), .ZN(n17516) );
  AOI22_X1 U19520 ( .A1(n17641), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17656), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17514) );
  AOI22_X1 U19521 ( .A1(n17510), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U19522 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17512) );
  AOI22_X1 U19523 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17511) );
  NAND4_X1 U19524 ( .A1(n17514), .A2(n17513), .A3(n17512), .A4(n17511), .ZN(
        n17515) );
  AOI211_X1 U19525 ( .C1(n17520), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n17516), .B(n17515), .ZN(n17517) );
  NAND3_X1 U19526 ( .A1(n17519), .A2(n17518), .A3(n17517), .ZN(n17577) );
  NAND2_X1 U19527 ( .A1(n17580), .A2(n17577), .ZN(n17576) );
  NOR2_X1 U19528 ( .A1(n17561), .A2(n17576), .ZN(n17573) );
  AOI22_X1 U19529 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17531) );
  AOI22_X1 U19530 ( .A1(n17641), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10980), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17530) );
  AOI22_X1 U19531 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17521) );
  OAI21_X1 U19532 ( .B1(n12572), .B2(n17522), .A(n17521), .ZN(n17528) );
  AOI22_X1 U19533 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17526) );
  AOI22_X1 U19534 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17525) );
  AOI22_X1 U19535 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17524) );
  AOI22_X1 U19536 ( .A1(n17628), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17523) );
  NAND4_X1 U19537 ( .A1(n17526), .A2(n17525), .A3(n17524), .A4(n17523), .ZN(
        n17527) );
  AOI211_X1 U19538 ( .C1(n17599), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n17528), .B(n17527), .ZN(n17529) );
  NAND3_X1 U19539 ( .A1(n17531), .A2(n17530), .A3(n17529), .ZN(n17572) );
  NAND2_X1 U19540 ( .A1(n17573), .A2(n17572), .ZN(n17571) );
  NOR2_X1 U19541 ( .A1(n17566), .A2(n17571), .ZN(n17565) );
  AOI22_X1 U19542 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17535) );
  AOI22_X1 U19543 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17666), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17534) );
  AOI22_X1 U19544 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17533) );
  AOI22_X1 U19545 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17532) );
  NAND4_X1 U19546 ( .A1(n17535), .A2(n17534), .A3(n17533), .A4(n17532), .ZN(
        n17542) );
  AOI22_X1 U19547 ( .A1(n17536), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17540) );
  AOI22_X1 U19548 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U19549 ( .A1(n17641), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17667), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17538) );
  AOI22_X1 U19550 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17537) );
  NAND4_X1 U19551 ( .A1(n17540), .A2(n17539), .A3(n17538), .A4(n17537), .ZN(
        n17541) );
  NOR2_X1 U19552 ( .A1(n17542), .A2(n17541), .ZN(n17543) );
  XOR2_X1 U19553 ( .A(n17565), .B(n17543), .Z(n20709) );
  OAI22_X1 U19554 ( .A1(n17545), .A2(n17544), .B1(n20709), .B2(n17682), .ZN(
        P3_U2673) );
  NAND2_X1 U19555 ( .A1(n20667), .A2(n17546), .ZN(n17559) );
  NOR2_X1 U19556 ( .A1(n17685), .A2(n17546), .ZN(n17623) );
  AOI22_X1 U19557 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17550) );
  AOI22_X1 U19558 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17549) );
  AOI22_X1 U19559 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17627), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17548) );
  AOI22_X1 U19560 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17547) );
  NAND4_X1 U19561 ( .A1(n17550), .A2(n17549), .A3(n17548), .A4(n17547), .ZN(
        n17556) );
  AOI22_X1 U19562 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U19563 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17553) );
  AOI22_X1 U19564 ( .A1(n17641), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17552) );
  AOI22_X1 U19565 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17551) );
  NAND4_X1 U19566 ( .A1(n17554), .A2(n17553), .A3(n17552), .A4(n17551), .ZN(
        n17555) );
  NOR2_X1 U19567 ( .A1(n17556), .A2(n17555), .ZN(n20658) );
  INV_X1 U19568 ( .A(n20658), .ZN(n17557) );
  AOI22_X1 U19569 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17623), .B1(n17685), 
        .B2(n17557), .ZN(n17558) );
  OAI21_X1 U19570 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17559), .A(n17558), .ZN(
        P3_U2682) );
  NOR2_X1 U19571 ( .A1(n20437), .A2(n17559), .ZN(n17595) );
  NAND2_X1 U19572 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17611), .ZN(n17588) );
  NOR3_X1 U19573 ( .A1(n20495), .A2(n17560), .A3(n17588), .ZN(n17584) );
  AND2_X1 U19574 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17584), .ZN(n17579) );
  NAND2_X1 U19575 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17579), .ZN(n17575) );
  INV_X1 U19576 ( .A(n17575), .ZN(n17568) );
  AOI21_X1 U19577 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17682), .A(n17579), .ZN(
        n17563) );
  AOI21_X1 U19578 ( .B1(n17561), .B2(n17576), .A(n17573), .ZN(n20726) );
  INV_X1 U19579 ( .A(n20726), .ZN(n17562) );
  OAI22_X1 U19580 ( .A1(n17568), .A2(n17563), .B1(n17562), .B2(n17682), .ZN(
        P3_U2676) );
  NAND2_X1 U19581 ( .A1(n17682), .A2(n17575), .ZN(n17564) );
  OAI21_X1 U19582 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17687), .A(n17564), .ZN(
        n17567) );
  AOI21_X1 U19583 ( .B1(n17566), .B2(n17571), .A(n17565), .ZN(n20714) );
  AOI22_X1 U19584 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17567), .B1(n20714), 
        .B2(n17685), .ZN(n17570) );
  INV_X1 U19585 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n20544) );
  NAND3_X1 U19586 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17568), .A3(n20544), 
        .ZN(n17569) );
  NAND2_X1 U19587 ( .A1(n17570), .A2(n17569), .ZN(P3_U2674) );
  OAI21_X1 U19588 ( .B1(n17573), .B2(n17572), .A(n17571), .ZN(n20720) );
  NAND3_X1 U19589 ( .A1(n17575), .A2(P3_EBX_REG_28__SCAN_IN), .A3(n17682), 
        .ZN(n17574) );
  OAI221_X1 U19590 ( .B1(n17575), .B2(P3_EBX_REG_28__SCAN_IN), .C1(n17682), 
        .C2(n20720), .A(n17574), .ZN(P3_U2675) );
  AOI21_X1 U19591 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17682), .A(n17584), .ZN(
        n17578) );
  OAI21_X1 U19592 ( .B1(n17580), .B2(n17577), .A(n17576), .ZN(n20703) );
  OAI22_X1 U19593 ( .A1(n17579), .A2(n17578), .B1(n20703), .B2(n17682), .ZN(
        P3_U2677) );
  INV_X1 U19594 ( .A(n17588), .ZN(n17594) );
  AOI22_X1 U19595 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17682), .B1(
        P3_EBX_REG_24__SCAN_IN), .B2(n17594), .ZN(n17583) );
  AOI21_X1 U19596 ( .B1(n17581), .B2(n17585), .A(n17580), .ZN(n20697) );
  INV_X1 U19597 ( .A(n20697), .ZN(n17582) );
  OAI22_X1 U19598 ( .A1(n17584), .A2(n17583), .B1(n17582), .B2(n17682), .ZN(
        P3_U2678) );
  OAI21_X1 U19599 ( .B1(n17589), .B2(n17586), .A(n17585), .ZN(n20733) );
  NAND3_X1 U19600 ( .A1(n17588), .A2(P3_EBX_REG_24__SCAN_IN), .A3(n17682), 
        .ZN(n17587) );
  OAI221_X1 U19601 ( .B1(n17588), .B2(P3_EBX_REG_24__SCAN_IN), .C1(n17682), 
        .C2(n20733), .A(n17587), .ZN(P3_U2679) );
  AOI21_X1 U19602 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17682), .A(n17611), .ZN(
        n17593) );
  AOI21_X1 U19603 ( .B1(n17591), .B2(n17590), .A(n17589), .ZN(n20734) );
  INV_X1 U19604 ( .A(n20734), .ZN(n17592) );
  OAI22_X1 U19605 ( .A1(n17594), .A2(n17593), .B1(n17592), .B2(n17682), .ZN(
        P3_U2680) );
  AOI21_X1 U19606 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17682), .A(n17595), .ZN(
        n17610) );
  AOI22_X1 U19607 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17667), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17608) );
  AOI22_X1 U19608 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17607) );
  AOI22_X1 U19609 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17666), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17596) );
  OAI21_X1 U19610 ( .B1(n17598), .B2(n17597), .A(n17596), .ZN(n17605) );
  AOI22_X1 U19611 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17603) );
  AOI22_X1 U19612 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17602) );
  AOI22_X1 U19613 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17601) );
  AOI22_X1 U19614 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17600) );
  NAND4_X1 U19615 ( .A1(n17603), .A2(n17602), .A3(n17601), .A4(n17600), .ZN(
        n17604) );
  AOI211_X1 U19616 ( .C1(n17668), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17605), .B(n17604), .ZN(n17606) );
  NAND3_X1 U19617 ( .A1(n17608), .A2(n17607), .A3(n17606), .ZN(n20666) );
  INV_X1 U19618 ( .A(n20666), .ZN(n17609) );
  OAI22_X1 U19619 ( .A1(n17611), .A2(n17610), .B1(n17609), .B2(n17682), .ZN(
        P3_U2681) );
  AOI22_X1 U19620 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17616) );
  AOI22_X1 U19621 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17615) );
  AOI22_X1 U19622 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17614) );
  AOI22_X1 U19623 ( .A1(n17627), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17612), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17613) );
  NAND4_X1 U19624 ( .A1(n17616), .A2(n17615), .A3(n17614), .A4(n17613), .ZN(
        n17622) );
  AOI22_X1 U19625 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17620) );
  AOI22_X1 U19626 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17657), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17619) );
  AOI22_X1 U19627 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17666), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17618) );
  AOI22_X1 U19628 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17617) );
  NAND4_X1 U19629 ( .A1(n17620), .A2(n17619), .A3(n17618), .A4(n17617), .ZN(
        n17621) );
  NOR2_X1 U19630 ( .A1(n17622), .A2(n17621), .ZN(n20665) );
  INV_X1 U19631 ( .A(n17653), .ZN(n17624) );
  OAI21_X1 U19632 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17624), .A(n17623), .ZN(
        n17625) );
  OAI21_X1 U19633 ( .B1(n20665), .B2(n17682), .A(n17625), .ZN(P3_U2683) );
  OAI21_X1 U19634 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17626), .A(n17682), .ZN(
        n17639) );
  AOI22_X1 U19635 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17632) );
  AOI22_X1 U19636 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17631) );
  AOI22_X1 U19637 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17353), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17630) );
  AOI22_X1 U19638 ( .A1(n17641), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17629) );
  NAND4_X1 U19639 ( .A1(n17632), .A2(n17631), .A3(n17630), .A4(n17629), .ZN(
        n17638) );
  AOI22_X1 U19640 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10960), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17636) );
  AOI22_X1 U19641 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17635) );
  AOI22_X1 U19642 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17634) );
  AOI22_X1 U19643 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17633) );
  NAND4_X1 U19644 ( .A1(n17636), .A2(n17635), .A3(n17634), .A4(n17633), .ZN(
        n17637) );
  NOR2_X1 U19645 ( .A1(n17638), .A2(n17637), .ZN(n20684) );
  OAI22_X1 U19646 ( .A1(n17654), .A2(n17639), .B1(n20684), .B2(n17682), .ZN(
        P3_U2685) );
  AOI22_X1 U19647 ( .A1(n17641), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17640), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17646) );
  AOI22_X1 U19648 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17645) );
  AOI22_X1 U19649 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10980), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17644) );
  AOI22_X1 U19650 ( .A1(n17353), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17628), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17643) );
  NAND4_X1 U19651 ( .A1(n17646), .A2(n17645), .A3(n17644), .A4(n17643), .ZN(
        n17652) );
  AOI22_X1 U19652 ( .A1(n17498), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17659), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17650) );
  AOI22_X1 U19653 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10970), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17649) );
  AOI22_X1 U19654 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17664), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17648) );
  AOI22_X1 U19655 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17666), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17647) );
  NAND4_X1 U19656 ( .A1(n17650), .A2(n17649), .A3(n17648), .A4(n17647), .ZN(
        n17651) );
  NOR2_X1 U19657 ( .A1(n17652), .A2(n17651), .ZN(n20680) );
  OAI21_X1 U19658 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17654), .A(n17653), .ZN(
        n17655) );
  AOI22_X1 U19659 ( .A1(n17685), .A2(n20680), .B1(n17655), .B2(n17682), .ZN(
        P3_U2684) );
  AOI22_X1 U19660 ( .A1(n17657), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17656), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17663) );
  AOI22_X1 U19661 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10970), .B1(
        n17642), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17662) );
  AOI22_X1 U19662 ( .A1(n17599), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17659), .ZN(n17661) );
  AOI22_X1 U19663 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17627), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17628), .ZN(n17660) );
  NAND4_X1 U19664 ( .A1(n17663), .A2(n17662), .A3(n17661), .A4(n17660), .ZN(
        n17674) );
  AOI22_X1 U19665 ( .A1(n17665), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17664), .ZN(n17672) );
  AOI22_X1 U19666 ( .A1(n17667), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17666), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17671) );
  AOI22_X1 U19667 ( .A1(n17668), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17520), .ZN(n17670) );
  AOI22_X1 U19668 ( .A1(n10960), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17498), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17669) );
  NAND4_X1 U19669 ( .A1(n17672), .A2(n17671), .A3(n17670), .A4(n17669), .ZN(
        n17673) );
  NOR2_X1 U19670 ( .A1(n17674), .A2(n17673), .ZN(n20690) );
  AOI211_X1 U19671 ( .C1(n20390), .C2(n17676), .A(n17675), .B(n17687), .ZN(
        n17677) );
  AOI21_X1 U19672 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17684), .A(n17677), .ZN(
        n17678) );
  OAI21_X1 U19673 ( .B1(n20690), .B2(n17682), .A(n17678), .ZN(P3_U2686) );
  INV_X1 U19674 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17683) );
  NOR2_X1 U19675 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n20174) );
  NOR2_X1 U19676 ( .A1(n20174), .A2(n17679), .ZN(n20162) );
  AOI22_X1 U19677 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n17684), .B1(n17680), .B2(
        n20162), .ZN(n17681) );
  OAI21_X1 U19678 ( .B1(n17683), .B2(n17682), .A(n17681), .ZN(P3_U2702) );
  AOI22_X1 U19679 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17685), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17684), .ZN(n17686) );
  OAI21_X1 U19680 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17687), .A(n17686), .ZN(
        P3_U2703) );
  OAI21_X1 U19681 ( .B1(n21198), .B2(n20108), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17689) );
  OAI21_X1 U19682 ( .B1(n17691), .B2(n17690), .A(n17689), .ZN(P3_U2634) );
  INV_X1 U19683 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21271) );
  AOI21_X1 U19684 ( .B1(n21271), .B2(n17693), .A(n17692), .ZN(n21258) );
  INV_X1 U19685 ( .A(n17694), .ZN(n18653) );
  OAI21_X1 U19686 ( .B1(n21258), .B2(n18653), .A(n18096), .ZN(n17695) );
  OAI221_X1 U19687 ( .B1(n21216), .B2(n20096), .C1(n21216), .C2(n18096), .A(
        n17695), .ZN(P3_U2863) );
  INV_X1 U19688 ( .A(n17957), .ZN(n20938) );
  INV_X1 U19689 ( .A(n21263), .ZN(n21266) );
  INV_X1 U19690 ( .A(n17696), .ZN(n21211) );
  NOR2_X4 U19691 ( .A1(n20158), .A2(n21270), .ZN(n18081) );
  OAI22_X2 U19692 ( .A1(n20938), .A2(n18091), .B1(n18002), .B2(n21130), .ZN(
        n17975) );
  NAND2_X1 U19693 ( .A1(n20832), .A2(n17975), .ZN(n17764) );
  AOI22_X1 U19694 ( .A1(n21129), .A2(n10982), .B1(n20989), .B2(n17952), .ZN(
        n17741) );
  INV_X1 U19695 ( .A(n17741), .ZN(n17727) );
  AOI21_X1 U19696 ( .B1(n17928), .B2(n21132), .A(n17727), .ZN(n17933) );
  NAND2_X1 U19697 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18005) );
  NAND2_X1 U19698 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17959) );
  NOR2_X2 U19699 ( .A1(n18005), .A2(n17959), .ZN(n20288) );
  NAND2_X1 U19700 ( .A1(n20288), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17944) );
  NOR2_X1 U19701 ( .A1(n20316), .A2(n20323), .ZN(n20322) );
  NAND2_X1 U19702 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17735) );
  INV_X1 U19703 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20163) );
  NOR2_X1 U19704 ( .A1(n17925), .A2(n20163), .ZN(n17698) );
  AOI21_X1 U19705 ( .B1(n17722), .B2(n17925), .A(n18059), .ZN(n17930) );
  OAI21_X1 U19706 ( .B1(n17698), .B2(n18086), .A(n17930), .ZN(n17710) );
  NAND2_X1 U19707 ( .A1(n18932), .A2(n18693), .ZN(n18773) );
  INV_X1 U19708 ( .A(n17879), .ZN(n17724) );
  NOR3_X1 U19709 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17724), .A3(
        n17925), .ZN(n17711) );
  INV_X1 U19710 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21143) );
  INV_X1 U19711 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20402) );
  NAND2_X1 U19712 ( .A1(n17713), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17708) );
  OAI21_X1 U19713 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17698), .A(
        n17708), .ZN(n20405) );
  OAI22_X1 U19714 ( .A1(n10961), .A2(n21143), .B1(n17897), .B2(n20405), .ZN(
        n17699) );
  AOI211_X1 U19715 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17710), .A(
        n17711), .B(n17699), .ZN(n17702) );
  AOI21_X1 U19716 ( .B1(n17971), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17788), .ZN(n17700) );
  XOR2_X1 U19717 ( .A(n17705), .B(n17700), .Z(n21141) );
  NOR2_X1 U19718 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21132), .ZN(
        n21140) );
  AOI22_X1 U19719 ( .A1(n18004), .A2(n21141), .B1(n17928), .B2(n21140), .ZN(
        n17701) );
  OAI211_X1 U19720 ( .C1(n17933), .C2(n17703), .A(n17702), .B(n17701), .ZN(
        P3_U2812) );
  NAND2_X1 U19721 ( .A1(n17704), .A2(n17928), .ZN(n17838) );
  NAND2_X1 U19722 ( .A1(n17704), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n20834) );
  OR2_X1 U19723 ( .A1(n20989), .A2(n20834), .ZN(n21109) );
  OR2_X1 U19724 ( .A1(n21129), .A2(n20834), .ZN(n21110) );
  AOI22_X1 U19725 ( .A1(n17952), .A2(n21109), .B1(n10982), .B2(n21110), .ZN(
        n17791) );
  AND2_X1 U19726 ( .A1(n17788), .A2(n17705), .ZN(n17779) );
  AND3_X1 U19727 ( .A1(n17971), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17706), .ZN(n17787) );
  NOR2_X1 U19728 ( .A1(n17779), .A2(n17787), .ZN(n17707) );
  XNOR2_X1 U19729 ( .A(n17707), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21117) );
  INV_X1 U19730 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20416) );
  NOR2_X1 U19731 ( .A1(n10961), .A2(n20416), .ZN(n21116) );
  INV_X1 U19732 ( .A(n17708), .ZN(n17709) );
  NAND2_X1 U19733 ( .A1(n17713), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17766) );
  INV_X1 U19734 ( .A(n17766), .ZN(n17794) );
  NAND2_X1 U19735 ( .A1(n17794), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17795) );
  OAI21_X1 U19736 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17709), .A(
        n17795), .ZN(n20403) );
  OAI21_X1 U19737 ( .B1(n17711), .B2(n17710), .A(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17715) );
  INV_X1 U19738 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17712) );
  NAND3_X1 U19739 ( .A1(n17713), .A2(n17712), .A3(n17879), .ZN(n17714) );
  OAI211_X1 U19740 ( .C1(n20403), .C2(n17897), .A(n17715), .B(n17714), .ZN(
        n17716) );
  AOI211_X1 U19741 ( .C1(n18004), .C2(n21117), .A(n21116), .B(n17716), .ZN(
        n17717) );
  OAI221_X1 U19742 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17838), 
        .C1(n21120), .C2(n17791), .A(n17717), .ZN(P3_U2811) );
  NAND2_X1 U19743 ( .A1(n20998), .A2(n12545), .ZN(n17730) );
  INV_X1 U19744 ( .A(n17984), .ZN(n17970) );
  NOR2_X1 U19745 ( .A1(n17719), .A2(n17970), .ZN(n17937) );
  NOR2_X1 U19746 ( .A1(n17955), .A2(n17720), .ZN(n17938) );
  AOI22_X1 U19747 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17937), .B1(
        n17938), .B2(n17950), .ZN(n17721) );
  XNOR2_X1 U19748 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17721), .ZN(
        n20992) );
  NOR2_X1 U19749 ( .A1(n17723), .A2(n20163), .ZN(n20349) );
  NAND2_X1 U19750 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20349), .ZN(
        n17733) );
  OAI21_X1 U19751 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20349), .A(
        n17733), .ZN(n20348) );
  AOI21_X1 U19752 ( .B1(n17722), .B2(n17723), .A(n18059), .ZN(n17945) );
  OAI21_X1 U19753 ( .B1(n20349), .B2(n18086), .A(n17945), .ZN(n17734) );
  NOR2_X1 U19754 ( .A1(n17724), .A2(n17723), .ZN(n17736) );
  INV_X1 U19755 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20362) );
  AOI22_X1 U19756 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17734), .B1(
        n17736), .B2(n20362), .ZN(n17725) );
  NAND2_X1 U19757 ( .A1(n21189), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n21000) );
  OAI211_X1 U19758 ( .C1(n17897), .C2(n20348), .A(n17725), .B(n21000), .ZN(
        n17726) );
  AOI21_X1 U19759 ( .B1(n18004), .B2(n20992), .A(n17726), .ZN(n17729) );
  OAI21_X1 U19760 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n20988), .A(
        n17727), .ZN(n17728) );
  OAI211_X1 U19761 ( .C1(n17730), .C2(n18091), .A(n17729), .B(n17728), .ZN(
        P3_U2815) );
  AOI22_X1 U19762 ( .A1(n17971), .A2(n21155), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17869), .ZN(n17731) );
  XNOR2_X1 U19763 ( .A(n17732), .B(n17731), .ZN(n21157) );
  INV_X1 U19764 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n21159) );
  INV_X1 U19765 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20369) );
  NAND2_X1 U19766 ( .A1(n17929), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20380) );
  INV_X1 U19767 ( .A(n20380), .ZN(n17926) );
  AOI21_X1 U19768 ( .B1(n20369), .B2(n17733), .A(n17926), .ZN(n20367) );
  AOI22_X1 U19769 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17734), .B1(
        n17917), .B2(n20367), .ZN(n17738) );
  OAI211_X1 U19770 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17736), .B(n17735), .ZN(n17737) );
  OAI211_X1 U19771 ( .C1(n21159), .C2(n10961), .A(n17738), .B(n17737), .ZN(
        n17739) );
  AOI21_X1 U19772 ( .B1(n18004), .B2(n21157), .A(n17739), .ZN(n17740) );
  OAI221_X1 U19773 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17764), 
        .C1(n21155), .C2(n17741), .A(n17740), .ZN(P3_U2814) );
  NAND2_X1 U19774 ( .A1(n20958), .A2(n20957), .ZN(n17742) );
  NAND2_X1 U19775 ( .A1(n20957), .A2(n17957), .ZN(n20961) );
  AOI22_X1 U19776 ( .A1(n17952), .A2(n17742), .B1(n10982), .B2(n20961), .ZN(
        n17761) );
  NAND2_X1 U19777 ( .A1(n17743), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17960) );
  NOR2_X1 U19778 ( .A1(n20316), .A2(n17960), .ZN(n17940) );
  AOI21_X1 U19779 ( .B1(n20316), .B2(n17960), .A(n17940), .ZN(n20314) );
  NAND2_X1 U19780 ( .A1(n17743), .A2(n17879), .ZN(n17752) );
  OAI21_X1 U19781 ( .B1(n17743), .B2(n18047), .A(n18087), .ZN(n17744) );
  AOI21_X1 U19782 ( .B1(n17839), .B2(n17960), .A(n17744), .ZN(n17753) );
  NAND2_X1 U19783 ( .A1(n21189), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n20966) );
  OAI221_X1 U19784 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17752), .C1(
        n20316), .C2(n17753), .A(n20966), .ZN(n17745) );
  AOI21_X1 U19785 ( .B1(n17917), .B2(n20314), .A(n17745), .ZN(n17750) );
  INV_X1 U19786 ( .A(n20946), .ZN(n20940) );
  NAND2_X1 U19787 ( .A1(n20940), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n20951) );
  NOR2_X1 U19788 ( .A1(n11268), .A2(n20951), .ZN(n17746) );
  MUX2_X1 U19789 ( .A(n17746), .B(n11054), .S(n17869), .Z(n17747) );
  XNOR2_X1 U19790 ( .A(n20968), .B(n17747), .ZN(n20965) );
  NOR2_X1 U19791 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n20951), .ZN(
        n17748) );
  AOI22_X1 U19792 ( .A1(n18004), .A2(n20965), .B1(n17748), .B2(n17975), .ZN(
        n17749) );
  OAI211_X1 U19793 ( .C1(n17761), .C2(n20968), .A(n17750), .B(n17749), .ZN(
        P3_U2818) );
  INV_X1 U19794 ( .A(n17940), .ZN(n17751) );
  AOI22_X1 U19795 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17940), .B1(
        n17751), .B2(n20323), .ZN(n20328) );
  AOI211_X1 U19796 ( .C1(n20316), .C2(n20323), .A(n20322), .B(n17752), .ZN(
        n17755) );
  NAND2_X1 U19797 ( .A1(n21189), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n21171) );
  OAI21_X1 U19798 ( .B1(n17753), .B2(n20323), .A(n21171), .ZN(n17754) );
  AOI211_X1 U19799 ( .C1(n17917), .C2(n20328), .A(n17755), .B(n17754), .ZN(
        n17760) );
  AOI22_X1 U19800 ( .A1(n17984), .A2(n20957), .B1(n17756), .B2(n17869), .ZN(
        n17757) );
  XNOR2_X1 U19801 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17757), .ZN(
        n21170) );
  NAND2_X1 U19802 ( .A1(n20957), .A2(n21166), .ZN(n21173) );
  INV_X1 U19803 ( .A(n21173), .ZN(n17758) );
  AOI22_X1 U19804 ( .A1(n18004), .A2(n21170), .B1(n17758), .B2(n17975), .ZN(
        n17759) );
  OAI211_X1 U19805 ( .C1(n17761), .C2(n21166), .A(n17760), .B(n17759), .ZN(
        P3_U2817) );
  AOI21_X1 U19806 ( .B1(n17763), .B2(n17762), .A(n17785), .ZN(n17807) );
  XNOR2_X1 U19807 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17807), .ZN(
        n21012) );
  NOR2_X1 U19808 ( .A1(n17765), .A2(n17764), .ZN(n17902) );
  INV_X1 U19809 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21094) );
  NOR2_X1 U19810 ( .A1(n17765), .A2(n21129), .ZN(n20838) );
  NOR2_X1 U19811 ( .A1(n17765), .A2(n20989), .ZN(n20837) );
  OAI22_X1 U19812 ( .A1(n20838), .A2(n18091), .B1(n20837), .B2(n18002), .ZN(
        n17782) );
  INV_X1 U19813 ( .A(n17881), .ZN(n17862) );
  INV_X1 U19814 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n20424) );
  AOI21_X1 U19815 ( .B1(n17839), .B2(n17795), .A(n18059), .ZN(n17767) );
  OAI21_X1 U19816 ( .B1(n17768), .B2(n18047), .A(n17767), .ZN(n17793) );
  AOI21_X1 U19817 ( .B1(n17862), .B2(n20424), .A(n17793), .ZN(n17775) );
  INV_X1 U19818 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n20458) );
  NAND3_X1 U19819 ( .A1(n17768), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17769) );
  NOR2_X1 U19820 ( .A1(n17802), .A2(n20163), .ZN(n17803) );
  AOI21_X1 U19821 ( .B1(n20458), .B2(n17769), .A(n17803), .ZN(n20452) );
  AOI22_X1 U19822 ( .A1(n21161), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n17917), 
        .B2(n20452), .ZN(n17771) );
  INV_X1 U19823 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17777) );
  AND2_X1 U19824 ( .A1(n17879), .A2(n17768), .ZN(n17778) );
  OAI221_X1 U19825 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n20458), .C2(n17777), .A(
        n17778), .ZN(n17770) );
  OAI211_X1 U19826 ( .C1(n17775), .C2(n20458), .A(n17771), .B(n17770), .ZN(
        n17772) );
  AOI221_X1 U19827 ( .B1(n17902), .B2(n21094), .C1(n17782), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17772), .ZN(n17773) );
  OAI21_X1 U19828 ( .B1(n17967), .B2(n21012), .A(n17773), .ZN(P3_U2808) );
  NAND2_X1 U19829 ( .A1(n20841), .A2(n21007), .ZN(n20845) );
  INV_X1 U19830 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20442) );
  NOR2_X1 U19831 ( .A1(n10961), .A2(n20442), .ZN(n20830) );
  NAND2_X1 U19832 ( .A1(n17768), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17774) );
  XOR2_X1 U19833 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n17774), .Z(
        n20431) );
  OAI22_X1 U19834 ( .A1(n17775), .A2(n17777), .B1(n17897), .B2(n20431), .ZN(
        n17776) );
  AOI211_X1 U19835 ( .C1(n17778), .C2(n17777), .A(n20830), .B(n17776), .ZN(
        n17784) );
  AOI22_X1 U19836 ( .A1(n20841), .A2(n17787), .B1(n17780), .B2(n17779), .ZN(
        n17781) );
  XNOR2_X1 U19837 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17781), .ZN(
        n20831) );
  AOI22_X1 U19838 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17782), .B1(
        n18004), .B2(n20831), .ZN(n17783) );
  OAI211_X1 U19839 ( .C1(n20845), .C2(n17838), .A(n17784), .B(n17783), .ZN(
        P3_U2809) );
  INV_X1 U19840 ( .A(n17785), .ZN(n17786) );
  OAI221_X1 U19841 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17788), 
        .C1(n21120), .C2(n17787), .A(n17786), .ZN(n17789) );
  XNOR2_X1 U19842 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17789), .ZN(
        n21123) );
  NAND2_X1 U19843 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17790), .ZN(
        n21128) );
  OAI22_X1 U19844 ( .A1(n17791), .A2(n17790), .B1(n17838), .B2(n21128), .ZN(
        n17792) );
  AOI21_X1 U19845 ( .B1(n18004), .B2(n21123), .A(n17792), .ZN(n17798) );
  NAND2_X1 U19846 ( .A1(n21189), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n21125) );
  INV_X2 U19847 ( .A(n18773), .ZN(n18978) );
  OAI221_X1 U19848 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17794), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18978), .A(n17793), .ZN(
        n17797) );
  AOI22_X1 U19849 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17768), .B1(
        n20424), .B2(n17795), .ZN(n20421) );
  OAI21_X1 U19850 ( .B1(n17917), .B2(n17862), .A(n20421), .ZN(n17796) );
  NAND4_X1 U19851 ( .A1(n17798), .A2(n21125), .A3(n17797), .A4(n17796), .ZN(
        P3_U2810) );
  NOR2_X1 U19852 ( .A1(n21084), .A2(n18002), .ZN(n17800) );
  NOR2_X1 U19853 ( .A1(n21087), .A2(n18091), .ZN(n17799) );
  AOI22_X1 U19854 ( .A1(n17800), .A2(n20837), .B1(n17799), .B2(n20838), .ZN(
        n17812) );
  INV_X1 U19855 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17818) );
  INV_X1 U19856 ( .A(n17815), .ZN(n17804) );
  NAND2_X1 U19857 ( .A1(n18978), .A2(n17804), .ZN(n17801) );
  OAI211_X1 U19858 ( .C1(n17803), .C2(n18086), .A(n18087), .B(n17801), .ZN(
        n17817) );
  OAI21_X1 U19859 ( .B1(n17802), .B2(n18773), .A(n17818), .ZN(n17806) );
  OAI22_X1 U19860 ( .A1(n20163), .A2(n17804), .B1(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17803), .ZN(n20463) );
  AOI21_X1 U19861 ( .B1(n17897), .B2(n17881), .A(n20463), .ZN(n17805) );
  INV_X1 U19862 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20468) );
  NOR2_X1 U19863 ( .A1(n10961), .A2(n20468), .ZN(n21095) );
  AOI211_X1 U19864 ( .C1(n17817), .C2(n17806), .A(n17805), .B(n21095), .ZN(
        n17811) );
  OAI22_X1 U19865 ( .A1(n21087), .A2(n18091), .B1(n21084), .B2(n18002), .ZN(
        n17835) );
  OAI221_X1 U19866 ( .B1(n17808), .B2(n17971), .C1(n17808), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17807), .ZN(n17809) );
  XNOR2_X1 U19867 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n17809), .ZN(
        n21096) );
  AOI22_X1 U19868 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17835), .B1(
        n18004), .B2(n21096), .ZN(n17810) );
  OAI211_X1 U19869 ( .C1(n17812), .C2(n21094), .A(n17811), .B(n17810), .ZN(
        P3_U2807) );
  NAND2_X1 U19870 ( .A1(n17869), .A2(n17833), .ZN(n17868) );
  OAI21_X1 U19871 ( .B1(n17869), .B2(n17813), .A(n17868), .ZN(n17814) );
  XNOR2_X1 U19872 ( .A(n17814), .B(n21016), .ZN(n21030) );
  INV_X1 U19873 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n20491) );
  NAND3_X1 U19874 ( .A1(n17815), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17816) );
  NOR2_X1 U19875 ( .A1(n17865), .A2(n20163), .ZN(n17864) );
  AOI21_X1 U19876 ( .B1(n20491), .B2(n17816), .A(n17864), .ZN(n20489) );
  INV_X1 U19877 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17830) );
  NAND2_X1 U19878 ( .A1(n17815), .A2(n17879), .ZN(n17831) );
  AOI221_X1 U19879 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n20491), .C2(n17830), .A(
        n17831), .ZN(n17820) );
  AOI21_X1 U19880 ( .B1(n17862), .B2(n17818), .A(n17817), .ZN(n17829) );
  INV_X1 U19881 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20501) );
  OAI22_X1 U19882 ( .A1(n17829), .A2(n20491), .B1(n10961), .B2(n20501), .ZN(
        n17819) );
  AOI211_X1 U19883 ( .C1(n20489), .C2(n17917), .A(n17820), .B(n17819), .ZN(
        n17826) );
  AOI21_X1 U19884 ( .B1(n21016), .B2(n17822), .A(n17821), .ZN(n21023) );
  AOI21_X1 U19885 ( .B1(n21016), .B2(n17824), .A(n17823), .ZN(n21026) );
  AOI22_X1 U19886 ( .A1(n17952), .A2(n21023), .B1(n10982), .B2(n21026), .ZN(
        n17825) );
  OAI211_X1 U19887 ( .C1(n17967), .C2(n21030), .A(n17826), .B(n17825), .ZN(
        P3_U2805) );
  OR3_X1 U19888 ( .A1(n21019), .A2(n17827), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21108) );
  NAND2_X1 U19889 ( .A1(n17815), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17828) );
  XNOR2_X1 U19890 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n17828), .ZN(
        n20477) );
  NAND2_X1 U19891 ( .A1(n21189), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n21106) );
  OAI221_X1 U19892 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17831), .C1(
        n17830), .C2(n17829), .A(n21106), .ZN(n17832) );
  AOI21_X1 U19893 ( .B1(n17917), .B2(n20477), .A(n17832), .ZN(n17837) );
  OAI21_X1 U19894 ( .B1(n17834), .B2(n21101), .A(n17833), .ZN(n21105) );
  AOI22_X1 U19895 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17835), .B1(
        n18004), .B2(n21105), .ZN(n17836) );
  OAI211_X1 U19896 ( .C1(n17838), .C2(n21108), .A(n17837), .B(n17836), .ZN(
        P3_U2806) );
  INV_X1 U19897 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20515) );
  AND2_X1 U19898 ( .A1(n11067), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17854) );
  NOR2_X1 U19899 ( .A1(n17907), .A2(n20163), .ZN(n17884) );
  INV_X1 U19900 ( .A(n17884), .ZN(n17916) );
  OAI21_X1 U19901 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17854), .A(
        n17916), .ZN(n20547) );
  INV_X1 U19902 ( .A(n20547), .ZN(n20534) );
  AND3_X1 U19903 ( .A1(n11200), .A2(n17879), .A3(n11067), .ZN(n17843) );
  OAI21_X1 U19904 ( .B1(n17865), .B2(n20163), .A(n17839), .ZN(n17840) );
  OAI211_X1 U19905 ( .C1(n11057), .C2(n18047), .A(n18087), .B(n17840), .ZN(
        n17867) );
  AOI21_X1 U19906 ( .B1(n17862), .B2(n20515), .A(n17867), .ZN(n17855) );
  NAND3_X1 U19907 ( .A1(n11057), .A2(n11201), .A3(n17879), .ZN(n17860) );
  OAI221_X1 U19908 ( .B1(n11200), .B2(n17855), .C1(n11200), .C2(n17860), .A(
        n17841), .ZN(n17842) );
  AOI211_X1 U19909 ( .C1(n17917), .C2(n20534), .A(n17843), .B(n17842), .ZN(
        n17851) );
  AOI22_X1 U19910 ( .A1(n10982), .A2(n21032), .B1(n17952), .B2(n21034), .ZN(
        n17873) );
  NAND2_X1 U19911 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17873), .ZN(
        n17857) );
  OAI211_X1 U19912 ( .C1(n17952), .C2(n10982), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17857), .ZN(n17850) );
  NAND3_X1 U19913 ( .A1(n17844), .A2(n17902), .A3(n12747), .ZN(n17849) );
  OAI211_X1 U19914 ( .C1(n17847), .C2(n17846), .A(n18004), .B(n17845), .ZN(
        n17848) );
  NAND4_X1 U19915 ( .A1(n17851), .A2(n17850), .A3(n17849), .A4(n17848), .ZN(
        P3_U2802) );
  OAI21_X1 U19916 ( .B1(n17971), .B2(n17853), .A(n17852), .ZN(n21053) );
  INV_X1 U19917 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20539) );
  NOR2_X1 U19918 ( .A1(n10961), .A2(n20539), .ZN(n21054) );
  NAND2_X1 U19919 ( .A1(n11057), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17863) );
  AOI21_X1 U19920 ( .B1(n11201), .B2(n17863), .A(n17854), .ZN(n20520) );
  OAI22_X1 U19921 ( .A1(n17855), .A2(n11201), .B1(n17897), .B2(n11195), .ZN(
        n17856) );
  AOI211_X1 U19922 ( .C1(n18004), .C2(n21053), .A(n21054), .B(n17856), .ZN(
        n17861) );
  INV_X1 U19923 ( .A(n17902), .ZN(n17872) );
  NOR2_X1 U19924 ( .A1(n21044), .A2(n17872), .ZN(n17858) );
  OAI21_X1 U19925 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17858), .A(
        n17857), .ZN(n17859) );
  NAND3_X1 U19926 ( .A1(n17861), .A2(n17860), .A3(n17859), .ZN(P3_U2803) );
  NOR2_X1 U19927 ( .A1(n17862), .A2(n17917), .ZN(n17927) );
  OAI21_X1 U19928 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17864), .A(
        n17863), .ZN(n20507) );
  OAI21_X1 U19929 ( .B1(n17865), .B2(n18773), .A(n20515), .ZN(n17866) );
  AOI22_X1 U19930 ( .A1(n21161), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17867), 
        .B2(n17866), .ZN(n17878) );
  OAI221_X1 U19931 ( .B1(n17870), .B2(n17869), .C1(n17870), .C2(n21016), .A(
        n17868), .ZN(n17871) );
  XNOR2_X1 U19932 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n17871), .ZN(
        n21041) );
  NOR2_X1 U19933 ( .A1(n21031), .A2(n17872), .ZN(n17875) );
  INV_X1 U19934 ( .A(n17873), .ZN(n17874) );
  MUX2_X1 U19935 ( .A(n17875), .B(n17874), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17876) );
  AOI21_X1 U19936 ( .B1(n18004), .B2(n21041), .A(n17876), .ZN(n17877) );
  OAI211_X1 U19937 ( .C1(n17927), .C2(n20507), .A(n17878), .B(n17877), .ZN(
        P3_U2804) );
  INV_X1 U19938 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20554) );
  NOR2_X2 U19939 ( .A1(n17907), .A2(n20554), .ZN(n17880) );
  NAND2_X1 U19940 ( .A1(n17880), .A2(n17879), .ZN(n17899) );
  INV_X1 U19941 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n20573) );
  XOR2_X1 U19942 ( .A(n20573), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n17885) );
  NOR2_X1 U19943 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17881), .ZN(
        n17918) );
  AOI21_X1 U19944 ( .B1(n18978), .B2(n17882), .A(n18059), .ZN(n17883) );
  OAI21_X1 U19945 ( .B1(n17884), .B2(n18086), .A(n17883), .ZN(n17909) );
  NOR2_X1 U19946 ( .A1(n17918), .A2(n17909), .ZN(n17898) );
  OAI22_X1 U19947 ( .A1(n17899), .A2(n17885), .B1(n17898), .B2(n20573), .ZN(
        n17886) );
  AOI211_X1 U19948 ( .C1(n10956), .C2(n17917), .A(n17887), .B(n17886), .ZN(
        n17893) );
  INV_X1 U19949 ( .A(n17888), .ZN(n17889) );
  AOI21_X1 U19950 ( .B1(n17891), .B2(n18004), .A(n17890), .ZN(n17892) );
  OAI211_X1 U19951 ( .C1(n17894), .C2(n18002), .A(n17893), .B(n17892), .ZN(
        P3_U2799) );
  AOI22_X1 U19952 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n17910), .B1(
        n17911), .B2(n21075), .ZN(n17895) );
  XNOR2_X1 U19953 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n17895), .ZN(
        n21083) );
  OAI22_X1 U19954 ( .A1(n21062), .A2(n18091), .B1(n21064), .B2(n18002), .ZN(
        n17914) );
  INV_X1 U19955 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n20557) );
  OAI21_X1 U19956 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17915), .A(
        n17896), .ZN(n20567) );
  OAI22_X1 U19957 ( .A1(n17898), .A2(n20557), .B1(n20567), .B2(n17897), .ZN(
        n17901) );
  INV_X1 U19958 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20569) );
  OAI22_X1 U19959 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n17899), .B1(
        n10961), .B2(n20569), .ZN(n17900) );
  AOI211_X1 U19960 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n17914), .A(
        n17901), .B(n17900), .ZN(n17906) );
  NAND4_X1 U19961 ( .A1(n17904), .A2(n17903), .A3(n17902), .A4(n21074), .ZN(
        n17905) );
  OAI211_X1 U19962 ( .C1(n21083), .C2(n17967), .A(n17906), .B(n17905), .ZN(
        P3_U2800) );
  OAI21_X1 U19963 ( .B1(n17907), .B2(n18773), .A(n20554), .ZN(n17908) );
  AOI22_X1 U19964 ( .A1(n21189), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n17909), 
        .B2(n17908), .ZN(n17922) );
  NOR2_X1 U19965 ( .A1(n21062), .A2(n18091), .ZN(n17913) );
  NAND2_X1 U19966 ( .A1(n17911), .A2(n17910), .ZN(n17912) );
  XNOR2_X1 U19967 ( .A(n17912), .B(n21075), .ZN(n21070) );
  AOI22_X1 U19968 ( .A1(n21061), .A2(n17913), .B1(n18004), .B2(n21070), .ZN(
        n17921) );
  OAI21_X1 U19969 ( .B1(n21058), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n17914), .ZN(n17920) );
  AOI21_X1 U19970 ( .B1(n17916), .B2(n20554), .A(n17915), .ZN(n20549) );
  OAI21_X1 U19971 ( .B1(n17918), .B2(n17917), .A(n20549), .ZN(n17919) );
  NAND4_X1 U19972 ( .A1(n17922), .A2(n17921), .A3(n17920), .A4(n17919), .ZN(
        P3_U2801) );
  AOI21_X1 U19973 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17924), .A(
        n17923), .ZN(n21151) );
  OAI22_X1 U19974 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17926), .B1(
        n20163), .B2(n17925), .ZN(n20382) );
  INV_X1 U19975 ( .A(n20382), .ZN(n17935) );
  INV_X1 U19976 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20394) );
  NOR2_X1 U19977 ( .A1(n10961), .A2(n20394), .ZN(n21145) );
  AOI21_X1 U19978 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17928), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17932) );
  AOI21_X1 U19979 ( .B1(n17929), .B2(n18978), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17931) );
  OAI22_X1 U19980 ( .A1(n17933), .A2(n17932), .B1(n17931), .B2(n17930), .ZN(
        n17934) );
  AOI211_X1 U19981 ( .C1(n17935), .C2(n18061), .A(n21145), .B(n17934), .ZN(
        n17936) );
  OAI21_X1 U19982 ( .B1(n21151), .B2(n17967), .A(n17936), .ZN(P3_U2813) );
  NOR2_X1 U19983 ( .A1(n17938), .A2(n17937), .ZN(n17939) );
  XNOR2_X1 U19984 ( .A(n17939), .B(n17950), .ZN(n20982) );
  INV_X1 U19985 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17942) );
  NAND2_X1 U19986 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17940), .ZN(
        n17941) );
  AOI21_X1 U19987 ( .B1(n17942), .B2(n17941), .A(n20349), .ZN(n20338) );
  NAND3_X1 U19988 ( .A1(n17943), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n18978), .ZN(n18015) );
  NOR2_X1 U19989 ( .A1(n17944), .A2(n18015), .ZN(n17962) );
  AOI21_X1 U19990 ( .B1(n20322), .B2(n17962), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17946) );
  INV_X1 U19991 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20340) );
  OAI22_X1 U19992 ( .A1(n17946), .A2(n17945), .B1(n10961), .B2(n20340), .ZN(
        n17947) );
  AOI21_X1 U19993 ( .B1(n20338), .B2(n18061), .A(n17947), .ZN(n17954) );
  AOI21_X1 U19994 ( .B1(n17950), .B2(n17948), .A(n20988), .ZN(n20975) );
  AOI21_X1 U19995 ( .B1(n17950), .B2(n17949), .A(n20998), .ZN(n20978) );
  AOI22_X1 U19996 ( .A1(n17952), .A2(n20975), .B1(n10982), .B2(n20978), .ZN(
        n17953) );
  OAI211_X1 U19997 ( .C1(n20982), .C2(n17967), .A(n17954), .B(n17953), .ZN(
        P3_U2816) );
  NOR2_X1 U19998 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17955), .ZN(
        n17985) );
  AOI22_X1 U19999 ( .A1(n20940), .A2(n17984), .B1(n17976), .B2(n17985), .ZN(
        n17956) );
  XNOR2_X1 U20000 ( .A(n17956), .B(n20956), .ZN(n20950) );
  OAI22_X1 U20001 ( .A1(n20958), .A2(n18002), .B1(n17957), .B2(n18091), .ZN(
        n17983) );
  INV_X1 U20002 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18183) );
  NOR2_X1 U20003 ( .A1(n10961), .A2(n18183), .ZN(n17964) );
  INV_X1 U20004 ( .A(n18015), .ZN(n17977) );
  NAND2_X1 U20005 ( .A1(n18087), .A2(n18047), .ZN(n18028) );
  AOI22_X1 U20006 ( .A1(n20288), .A2(n17977), .B1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18028), .ZN(n17961) );
  INV_X1 U20007 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17996) );
  INV_X1 U20008 ( .A(n18014), .ZN(n17995) );
  NAND3_X1 U20009 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17995), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20253) );
  NOR2_X1 U20010 ( .A1(n17996), .A2(n20253), .ZN(n20266) );
  INV_X1 U20011 ( .A(n20266), .ZN(n17958) );
  NOR2_X1 U20012 ( .A1(n17959), .A2(n17958), .ZN(n17968) );
  OAI21_X1 U20013 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17968), .A(
        n17960), .ZN(n20299) );
  OAI22_X1 U20014 ( .A1(n17962), .A2(n17961), .B1(n17927), .B2(n20299), .ZN(
        n17963) );
  AOI211_X1 U20015 ( .C1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n17983), .A(
        n17964), .B(n17963), .ZN(n17966) );
  OAI211_X1 U20016 ( .C1(n20940), .C2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n20951), .B(n17975), .ZN(n17965) );
  OAI211_X1 U20017 ( .C1(n20950), .C2(n17967), .A(n17966), .B(n17965), .ZN(
        P3_U2819) );
  INV_X1 U20018 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17969) );
  NAND2_X1 U20019 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n20266), .ZN(
        n20289) );
  AOI21_X1 U20020 ( .B1(n17969), .B2(n20289), .A(n17968), .ZN(n20292) );
  AOI22_X1 U20021 ( .A1(n21189), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n20292), 
        .B2(n18061), .ZN(n17982) );
  INV_X1 U20022 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21174) );
  AOI221_X1 U20023 ( .B1(n17971), .B2(n17970), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17970), .A(n21174), .ZN(
        n17974) );
  INV_X1 U20024 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21188) );
  AOI221_X1 U20025 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17984), .C1(
        n21188), .C2(n17985), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17972) );
  AOI22_X1 U20026 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17983), .B1(
        n18004), .B2(n21175), .ZN(n17981) );
  INV_X1 U20027 ( .A(n17975), .ZN(n17994) );
  OR3_X1 U20028 ( .A1(n20940), .A2(n17976), .A3(n17994), .ZN(n17980) );
  INV_X1 U20029 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20278) );
  NOR3_X1 U20030 ( .A1(n18005), .A2(n20278), .A3(n18015), .ZN(n17989) );
  NAND2_X1 U20031 ( .A1(n20288), .A2(n17977), .ZN(n17978) );
  OAI211_X1 U20032 ( .C1(n17989), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18028), .B(n17978), .ZN(n17979) );
  NAND4_X1 U20033 ( .A1(n17982), .A2(n17981), .A3(n17980), .A4(n17979), .ZN(
        P3_U2820) );
  INV_X1 U20034 ( .A(n17983), .ZN(n17993) );
  NOR2_X1 U20035 ( .A1(n17985), .A2(n17984), .ZN(n17986) );
  XNOR2_X1 U20036 ( .A(n17986), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n21193) );
  NAND2_X1 U20037 ( .A1(n21189), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n21195) );
  INV_X1 U20038 ( .A(n21195), .ZN(n17991) );
  NOR2_X1 U20039 ( .A1(n18005), .A2(n18015), .ZN(n17987) );
  AOI21_X1 U20040 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18028), .A(
        n17987), .ZN(n17988) );
  OAI21_X1 U20041 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n20266), .A(
        n20289), .ZN(n20268) );
  OAI22_X1 U20042 ( .A1(n17989), .A2(n17988), .B1(n17927), .B2(n20268), .ZN(
        n17990) );
  AOI211_X1 U20043 ( .C1(n18004), .C2(n21193), .A(n17991), .B(n17990), .ZN(
        n17992) );
  OAI221_X1 U20044 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17994), .C1(
        n21188), .C2(n17993), .A(n17992), .ZN(P3_U2821) );
  OAI21_X1 U20045 ( .B1(n17995), .B2(n18047), .A(n18087), .ZN(n18019) );
  AOI21_X1 U20046 ( .B1(n17996), .B2(n20253), .A(n20266), .ZN(n20255) );
  AOI22_X1 U20047 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18019), .B1(
        n20255), .B2(n18061), .ZN(n18009) );
  AOI21_X1 U20048 ( .B1(n17999), .B2(n17998), .A(n17997), .ZN(n20931) );
  OAI21_X1 U20049 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18001), .A(
        n18000), .ZN(n20930) );
  OAI22_X1 U20050 ( .A1(n20931), .A2(n18002), .B1(n18091), .B2(n20930), .ZN(
        n18003) );
  AOI21_X1 U20051 ( .B1(n18004), .B2(n20931), .A(n18003), .ZN(n18008) );
  NAND2_X1 U20052 ( .A1(n21189), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n20933) );
  INV_X1 U20053 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20247) );
  NOR2_X1 U20054 ( .A1(n20247), .A2(n18014), .ZN(n18006) );
  OAI211_X1 U20055 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18006), .A(
        n18978), .B(n18005), .ZN(n18007) );
  NAND4_X1 U20056 ( .A1(n18009), .A2(n18008), .A3(n20933), .A4(n18007), .ZN(
        P3_U2822) );
  OAI21_X1 U20057 ( .B1(n18012), .B2(n18011), .A(n18010), .ZN(n18013) );
  XNOR2_X1 U20058 ( .A(n18013), .B(n20927), .ZN(n20920) );
  NOR2_X1 U20059 ( .A1(n18014), .A2(n20163), .ZN(n20286) );
  OAI21_X1 U20060 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20286), .A(
        n20253), .ZN(n20238) );
  OAI22_X1 U20061 ( .A1(n17927), .A2(n20238), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18015), .ZN(n18016) );
  AOI21_X1 U20062 ( .B1(n21189), .B2(P3_REIP_REG_7__SCAN_IN), .A(n18016), .ZN(
        n18021) );
  AOI21_X1 U20063 ( .B1(n20927), .B2(n18018), .A(n18017), .ZN(n20919) );
  AOI22_X1 U20064 ( .A1(n18081), .A2(n20919), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18019), .ZN(n18020) );
  OAI211_X1 U20065 ( .C1(n18091), .C2(n20920), .A(n18021), .B(n18020), .ZN(
        P3_U2823) );
  OAI21_X1 U20066 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18023), .A(
        n18022), .ZN(n20914) );
  AOI21_X1 U20067 ( .B1(n11066), .B2(n18025), .A(n18024), .ZN(n20912) );
  NAND2_X1 U20068 ( .A1(n17943), .A2(n18978), .ZN(n18026) );
  INV_X1 U20069 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20908) );
  OAI22_X1 U20070 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18026), .B1(
        n10961), .B2(n20908), .ZN(n18027) );
  AOI21_X1 U20071 ( .B1(n18081), .B2(n20912), .A(n18027), .ZN(n18030) );
  INV_X1 U20072 ( .A(n18028), .ZN(n18083) );
  AOI21_X1 U20073 ( .B1(n18978), .B2(n17943), .A(n18083), .ZN(n18038) );
  INV_X1 U20074 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20237) );
  NAND2_X1 U20075 ( .A1(n17943), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20228) );
  AOI21_X1 U20076 ( .B1(n20237), .B2(n20228), .A(n20286), .ZN(n20229) );
  AOI22_X1 U20077 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18038), .B1(
        n20229), .B2(n18061), .ZN(n18029) );
  OAI211_X1 U20078 ( .C1(n18091), .C2(n20914), .A(n18030), .B(n18029), .ZN(
        P3_U2824) );
  OAI21_X1 U20079 ( .B1(n18033), .B2(n18032), .A(n18031), .ZN(n20898) );
  AOI21_X1 U20080 ( .B1(n20903), .B2(n18035), .A(n18034), .ZN(n20901) );
  AOI22_X1 U20081 ( .A1(n21189), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18081), 
        .B2(n20901), .ZN(n18040) );
  OAI21_X1 U20082 ( .B1(n18059), .B2(n20198), .A(n20221), .ZN(n18037) );
  NOR2_X1 U20083 ( .A1(n20198), .A2(n20163), .ZN(n18049) );
  OAI21_X1 U20084 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18049), .A(
        n20228), .ZN(n18036) );
  INV_X1 U20085 ( .A(n18036), .ZN(n20214) );
  AOI22_X1 U20086 ( .A1(n18038), .A2(n18037), .B1(n20214), .B2(n18061), .ZN(
        n18039) );
  OAI211_X1 U20087 ( .C1(n18091), .C2(n20898), .A(n18040), .B(n18039), .ZN(
        P3_U2825) );
  OAI21_X1 U20088 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18042), .A(
        n18041), .ZN(n20894) );
  AOI21_X1 U20089 ( .B1(n18045), .B2(n18044), .A(n18043), .ZN(n20890) );
  INV_X1 U20090 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20211) );
  NOR2_X1 U20091 ( .A1(n10961), .A2(n20211), .ZN(n20885) );
  AND3_X1 U20092 ( .A1(n11185), .A2(n18048), .A3(n18978), .ZN(n18046) );
  AOI211_X1 U20093 ( .C1(n18081), .C2(n20890), .A(n20885), .B(n18046), .ZN(
        n18051) );
  OAI21_X1 U20094 ( .B1(n18048), .B2(n18047), .A(n18087), .ZN(n18064) );
  NAND2_X1 U20095 ( .A1(n18048), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18060) );
  AOI21_X1 U20096 ( .B1(n11185), .B2(n18060), .A(n18049), .ZN(n20205) );
  AOI22_X1 U20097 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18064), .B1(
        n20205), .B2(n18061), .ZN(n18050) );
  OAI211_X1 U20098 ( .C1(n18091), .C2(n20894), .A(n18051), .B(n18050), .ZN(
        P3_U2826) );
  OAI21_X1 U20099 ( .B1(n18054), .B2(n18053), .A(n18052), .ZN(n20884) );
  AOI21_X1 U20100 ( .B1(n18057), .B2(n18056), .A(n18055), .ZN(n20882) );
  AOI22_X1 U20101 ( .A1(n21161), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18081), 
        .B2(n20882), .ZN(n18066) );
  OAI21_X1 U20102 ( .B1(n18059), .B2(n20183), .A(n18058), .ZN(n18063) );
  NOR2_X1 U20103 ( .A1(n20183), .A2(n20163), .ZN(n20171) );
  OAI21_X1 U20104 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20171), .A(
        n18060), .ZN(n20187) );
  INV_X1 U20105 ( .A(n20187), .ZN(n18062) );
  AOI22_X1 U20106 ( .A1(n18064), .A2(n18063), .B1(n18062), .B2(n18061), .ZN(
        n18065) );
  OAI211_X1 U20107 ( .C1(n18091), .C2(n20884), .A(n18066), .B(n18065), .ZN(
        P3_U2827) );
  AOI21_X1 U20108 ( .B1(n18069), .B2(n18068), .A(n18067), .ZN(n20864) );
  INV_X1 U20109 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20169) );
  NOR2_X1 U20110 ( .A1(n10961), .A2(n20169), .ZN(n20868) );
  AOI21_X1 U20111 ( .B1(n20183), .B2(n20163), .A(n20171), .ZN(n18070) );
  INV_X1 U20112 ( .A(n18070), .ZN(n20177) );
  OAI21_X1 U20113 ( .B1(n18073), .B2(n18072), .A(n18071), .ZN(n20870) );
  OAI22_X1 U20114 ( .A1(n17927), .A2(n20177), .B1(n18091), .B2(n20870), .ZN(
        n18074) );
  AOI211_X1 U20115 ( .C1(n18081), .C2(n20864), .A(n20868), .B(n18074), .ZN(
        n18075) );
  OAI221_X1 U20116 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18773), .C1(
        n20183), .C2(n18087), .A(n18075), .ZN(P3_U2828) );
  AOI21_X1 U20117 ( .B1(n18077), .B2(n18084), .A(n18076), .ZN(n20851) );
  AOI21_X1 U20118 ( .B1(n18085), .B2(n18079), .A(n18078), .ZN(n20854) );
  INV_X1 U20119 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20859) );
  OAI22_X1 U20120 ( .A1(n20854), .A2(n18091), .B1(n10961), .B2(n20859), .ZN(
        n18080) );
  AOI21_X1 U20121 ( .B1(n18081), .B2(n20851), .A(n18080), .ZN(n18082) );
  OAI221_X1 U20122 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17927), .C1(
        n20163), .C2(n18083), .A(n18082), .ZN(P3_U2829) );
  NAND2_X1 U20123 ( .A1(n18085), .A2(n18084), .ZN(n20848) );
  INV_X1 U20124 ( .A(n20848), .ZN(n20847) );
  NAND3_X1 U20125 ( .A1(n20785), .A2(n18087), .A3(n18086), .ZN(n18088) );
  AOI22_X1 U20126 ( .A1(n21161), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18088), .ZN(n18089) );
  OAI221_X1 U20127 ( .B1(n20847), .B2(n18091), .C1(n20848), .C2(n18090), .A(
        n18089), .ZN(P3_U2830) );
  INV_X1 U20128 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21228) );
  NOR2_X1 U20129 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18652), .ZN(
        n18698) );
  NOR2_X1 U20130 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n21228), .ZN(
        n18681) );
  NOR2_X1 U20131 ( .A1(n18698), .A2(n18681), .ZN(n18093) );
  OAI22_X1 U20132 ( .A1(n18094), .A2(n21228), .B1(n18093), .B2(n18092), .ZN(
        P3_U2866) );
  NAND2_X1 U20133 ( .A1(n18096), .A2(n18095), .ZN(n18099) );
  OAI21_X1 U20134 ( .B1(n18097), .B2(n18693), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18098) );
  OAI21_X1 U20135 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18099), .A(
        n18098), .ZN(P3_U2864) );
  NOR4_X1 U20136 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18103) );
  NOR4_X1 U20137 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18102) );
  NOR4_X1 U20138 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18101) );
  NOR4_X1 U20139 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18100) );
  NAND4_X1 U20140 ( .A1(n18103), .A2(n18102), .A3(n18101), .A4(n18100), .ZN(
        n18109) );
  NOR4_X1 U20141 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18107) );
  AOI211_X1 U20142 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18106) );
  NOR4_X1 U20143 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18105) );
  NOR4_X1 U20144 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18104) );
  NAND4_X1 U20145 ( .A1(n18107), .A2(n18106), .A3(n18105), .A4(n18104), .ZN(
        n18108) );
  NOR2_X1 U20146 ( .A1(n18109), .A2(n18108), .ZN(n18115) );
  INV_X1 U20147 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18211) );
  OAI21_X1 U20148 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18115), .ZN(n18110) );
  OAI21_X1 U20149 ( .B1(n18115), .B2(n18211), .A(n18110), .ZN(P3_U3293) );
  INV_X1 U20150 ( .A(n18115), .ZN(n18116) );
  INV_X1 U20151 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18216) );
  AOI21_X1 U20152 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18111) );
  AOI221_X1 U20153 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .C1(n20859), .C2(n18111), .A(n18116), .ZN(n18112) );
  AOI21_X1 U20154 ( .B1(n18116), .B2(n18216), .A(n18112), .ZN(P3_U3292) );
  INV_X1 U20155 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18213) );
  NOR2_X1 U20156 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18114) );
  INV_X1 U20157 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18113) );
  NAND3_X1 U20158 ( .A1(n18115), .A2(n18114), .A3(n18113), .ZN(n18117) );
  OAI221_X1 U20159 ( .B1(n18115), .B2(n18213), .C1(n18116), .C2(n20859), .A(
        n18117), .ZN(P3_U2638) );
  NAND2_X1 U20160 ( .A1(n18115), .A2(n20859), .ZN(n18119) );
  NAND2_X1 U20161 ( .A1(P3_BYTEENABLE_REG_3__SCAN_IN), .A2(n18116), .ZN(n18118) );
  OAI211_X1 U20162 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(n18119), .A(n18118), 
        .B(n18117), .ZN(P3_U2639) );
  INV_X1 U20163 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18120) );
  INV_X1 U20164 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18217) );
  AOI22_X1 U20165 ( .A1(n21682), .A2(n18120), .B1(n18217), .B2(n18214), .ZN(
        P3_U3297) );
  INV_X1 U20166 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18121) );
  AOI22_X1 U20167 ( .A1(n21682), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18121), 
        .B2(n18214), .ZN(P3_U3294) );
  AOI22_X1 U20168 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(n18214), .B1(n21676), .B2(
        n21678), .ZN(n18122) );
  OAI21_X1 U20169 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n21724), .A(n18122), 
        .ZN(P3_U2635) );
  INV_X1 U20170 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20780) );
  AOI22_X1 U20171 ( .A1(n21253), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18123) );
  OAI21_X1 U20172 ( .B1(n20780), .B2(n18144), .A(n18123), .ZN(P3_U2767) );
  INV_X1 U20173 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20769) );
  AOI22_X1 U20174 ( .A1(n21253), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18124) );
  OAI21_X1 U20175 ( .B1(n20769), .B2(n18144), .A(n18124), .ZN(P3_U2766) );
  INV_X1 U20176 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18126) );
  AOI22_X1 U20177 ( .A1(n21253), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18159), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18125) );
  OAI21_X1 U20178 ( .B1(n18126), .B2(n18144), .A(n18125), .ZN(P3_U2765) );
  INV_X1 U20179 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20132) );
  AOI22_X1 U20180 ( .A1(n21253), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18159), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18127) );
  OAI21_X1 U20181 ( .B1(n20132), .B2(n18144), .A(n18127), .ZN(P3_U2764) );
  INV_X1 U20182 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18129) );
  AOI22_X1 U20183 ( .A1(n21253), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18159), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18128) );
  OAI21_X1 U20184 ( .B1(n18129), .B2(n18144), .A(n18128), .ZN(P3_U2763) );
  INV_X1 U20185 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18131) );
  AOI22_X1 U20186 ( .A1(n21253), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18159), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18130) );
  OAI21_X1 U20187 ( .B1(n18131), .B2(n18144), .A(n18130), .ZN(P3_U2762) );
  INV_X1 U20188 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20625) );
  AOI22_X1 U20189 ( .A1(n21253), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18159), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18132) );
  OAI21_X1 U20190 ( .B1(n20625), .B2(n18144), .A(n18132), .ZN(P3_U2761) );
  INV_X1 U20191 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18134) );
  AOI22_X1 U20193 ( .A1(n21253), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18133) );
  OAI21_X1 U20194 ( .B1(n18134), .B2(n18144), .A(n18133), .ZN(P3_U2760) );
  INV_X1 U20195 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20762) );
  AOI22_X1 U20196 ( .A1(n21253), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18135) );
  OAI21_X1 U20197 ( .B1(n20762), .B2(n18144), .A(n18135), .ZN(P3_U2759) );
  INV_X1 U20198 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20598) );
  AOI22_X1 U20199 ( .A1(n21253), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18136) );
  OAI21_X1 U20200 ( .B1(n20598), .B2(n18144), .A(n18136), .ZN(P3_U2758) );
  INV_X1 U20201 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20140) );
  AOI22_X1 U20202 ( .A1(n21253), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18137) );
  OAI21_X1 U20203 ( .B1(n20140), .B2(n18144), .A(n18137), .ZN(P3_U2757) );
  INV_X1 U20204 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20599) );
  AOI22_X1 U20205 ( .A1(n21253), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18138) );
  OAI21_X1 U20206 ( .B1(n20599), .B2(n18144), .A(n18138), .ZN(P3_U2756) );
  INV_X1 U20207 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18140) );
  AOI22_X1 U20208 ( .A1(n21253), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18139) );
  OAI21_X1 U20209 ( .B1(n18140), .B2(n18144), .A(n18139), .ZN(P3_U2755) );
  INV_X1 U20210 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20147) );
  AOI22_X1 U20211 ( .A1(n21253), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18141) );
  OAI21_X1 U20212 ( .B1(n20147), .B2(n18144), .A(n18141), .ZN(P3_U2754) );
  INV_X1 U20213 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20149) );
  AOI22_X1 U20214 ( .A1(n21253), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18142) );
  OAI21_X1 U20215 ( .B1(n20149), .B2(n18144), .A(n18142), .ZN(P3_U2753) );
  INV_X1 U20216 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20756) );
  AOI22_X1 U20217 ( .A1(n21253), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18143) );
  OAI21_X1 U20218 ( .B1(n20756), .B2(n18144), .A(n18143), .ZN(P3_U2752) );
  INV_X1 U20219 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18147) );
  NAND2_X1 U20220 ( .A1(n18145), .A2(n20592), .ZN(n18170) );
  AOI22_X1 U20221 ( .A1(n21253), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18146) );
  OAI21_X1 U20222 ( .B1(n18147), .B2(n18170), .A(n18146), .ZN(P3_U2751) );
  INV_X1 U20223 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20654) );
  AOI22_X1 U20224 ( .A1(n21253), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18148) );
  OAI21_X1 U20225 ( .B1(n20654), .B2(n18170), .A(n18148), .ZN(P3_U2750) );
  INV_X1 U20226 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18150) );
  AOI22_X1 U20227 ( .A1(n21253), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18149) );
  OAI21_X1 U20228 ( .B1(n18150), .B2(n18170), .A(n18149), .ZN(P3_U2749) );
  INV_X1 U20229 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20676) );
  AOI22_X1 U20230 ( .A1(n21253), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18151) );
  OAI21_X1 U20231 ( .B1(n20676), .B2(n18170), .A(n18151), .ZN(P3_U2748) );
  INV_X1 U20232 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18153) );
  AOI22_X1 U20233 ( .A1(n21253), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18159), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18152) );
  OAI21_X1 U20234 ( .B1(n18153), .B2(n18170), .A(n18152), .ZN(P3_U2747) );
  INV_X1 U20235 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20661) );
  AOI22_X1 U20236 ( .A1(n21253), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18159), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18154) );
  OAI21_X1 U20237 ( .B1(n20661), .B2(n18170), .A(n18154), .ZN(P3_U2746) );
  INV_X1 U20238 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18156) );
  AOI22_X1 U20239 ( .A1(n21253), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18159), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18155) );
  OAI21_X1 U20240 ( .B1(n18156), .B2(n18170), .A(n18155), .ZN(P3_U2745) );
  INV_X1 U20241 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18158) );
  AOI22_X1 U20242 ( .A1(n21253), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18159), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18157) );
  OAI21_X1 U20243 ( .B1(n18158), .B2(n18170), .A(n18157), .ZN(P3_U2744) );
  INV_X1 U20244 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20118) );
  AOI22_X1 U20245 ( .A1(n21253), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18159), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18160) );
  OAI21_X1 U20246 ( .B1(n20118), .B2(n18170), .A(n18160), .ZN(P3_U2743) );
  INV_X1 U20247 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20694) );
  AOI22_X1 U20248 ( .A1(n21253), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18161) );
  OAI21_X1 U20249 ( .B1(n20694), .B2(n18170), .A(n18161), .ZN(P3_U2742) );
  INV_X1 U20250 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20121) );
  AOI22_X1 U20251 ( .A1(n21253), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18162) );
  OAI21_X1 U20252 ( .B1(n20121), .B2(n18170), .A(n18162), .ZN(P3_U2741) );
  INV_X1 U20253 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20723) );
  AOI22_X1 U20254 ( .A1(n21253), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18163) );
  OAI21_X1 U20255 ( .B1(n20723), .B2(n18170), .A(n18163), .ZN(P3_U2740) );
  INV_X1 U20256 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18165) );
  AOI22_X1 U20257 ( .A1(n21253), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18164) );
  OAI21_X1 U20258 ( .B1(n18165), .B2(n18170), .A(n18164), .ZN(P3_U2739) );
  INV_X1 U20259 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20711) );
  AOI22_X1 U20260 ( .A1(n21253), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18166) );
  OAI21_X1 U20261 ( .B1(n20711), .B2(n18170), .A(n18166), .ZN(P3_U2738) );
  INV_X1 U20262 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20126) );
  AOI22_X1 U20263 ( .A1(n21253), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18167), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18169) );
  OAI21_X1 U20264 ( .B1(n20126), .B2(n18170), .A(n18169), .ZN(P3_U2737) );
  NOR2_X1 U20265 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18171), .ZN(n18172) );
  NOR2_X1 U20266 ( .A1(n21682), .A2(n18172), .ZN(P3_U2633) );
  NAND2_X1 U20267 ( .A1(n21682), .A2(n21726), .ZN(n18209) );
  AOI22_X1 U20268 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n21724), .ZN(n18173) );
  OAI21_X1 U20269 ( .B1(n20169), .B2(n18209), .A(n18173), .ZN(P3_U3032) );
  INV_X1 U20270 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20879) );
  AOI22_X1 U20271 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n21724), .ZN(n18174) );
  OAI21_X1 U20272 ( .B1(n20879), .B2(n18209), .A(n18174), .ZN(P3_U3033) );
  AOI22_X1 U20273 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n21724), .ZN(n18175) );
  OAI21_X1 U20274 ( .B1(n20211), .B2(n18209), .A(n18175), .ZN(P3_U3034) );
  INV_X1 U20275 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20899) );
  AOI22_X1 U20276 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n21724), .ZN(n18176) );
  OAI21_X1 U20277 ( .B1(n20899), .B2(n18209), .A(n18176), .ZN(P3_U3035) );
  AOI22_X1 U20278 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n21724), .ZN(n18177) );
  OAI21_X1 U20279 ( .B1(n20908), .B2(n18209), .A(n18177), .ZN(P3_U3036) );
  INV_X1 U20280 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20252) );
  AOI22_X1 U20281 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n21724), .ZN(n18178) );
  OAI21_X1 U20282 ( .B1(n20252), .B2(n18209), .A(n18178), .ZN(P3_U3037) );
  INV_X1 U20283 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20258) );
  AOI22_X1 U20284 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n21724), .ZN(n18179) );
  OAI21_X1 U20285 ( .B1(n20258), .B2(n18209), .A(n18179), .ZN(P3_U3038) );
  INV_X1 U20286 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20269) );
  AOI22_X1 U20287 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n18214), .ZN(n18180) );
  OAI21_X1 U20288 ( .B1(n20269), .B2(n18209), .A(n18180), .ZN(P3_U3039) );
  INV_X1 U20289 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20297) );
  AOI22_X1 U20290 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_8__SCAN_IN), .B2(n18214), .ZN(n18181) );
  OAI21_X1 U20291 ( .B1(n20297), .B2(n18209), .A(n18181), .ZN(P3_U3040) );
  AOI22_X1 U20292 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_9__SCAN_IN), .B2(n18214), .ZN(n18182) );
  OAI21_X1 U20293 ( .B1(n18183), .B2(n18209), .A(n18182), .ZN(P3_U3041) );
  INV_X1 U20294 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20320) );
  AOI22_X1 U20295 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_10__SCAN_IN), .B2(n21724), .ZN(n18184) );
  OAI21_X1 U20296 ( .B1(n20320), .B2(n18209), .A(n18184), .ZN(P3_U3042) );
  INV_X1 U20297 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20330) );
  AOI22_X1 U20298 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18194), .B1(
        P3_ADDRESS_REG_11__SCAN_IN), .B2(n21724), .ZN(n18185) );
  OAI21_X1 U20299 ( .B1(n20330), .B2(n18209), .A(n18185), .ZN(P3_U3043) );
  INV_X1 U20300 ( .A(n18209), .ZN(n18203) );
  INV_X1 U20301 ( .A(n18203), .ZN(n18199) );
  AOI22_X1 U20302 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n18194), .B1(
        P3_ADDRESS_REG_12__SCAN_IN), .B2(n21724), .ZN(n18186) );
  OAI21_X1 U20303 ( .B1(n20340), .B2(n18199), .A(n18186), .ZN(P3_U3044) );
  INV_X1 U20304 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20376) );
  AOI22_X1 U20305 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n18194), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n21724), .ZN(n18187) );
  OAI21_X1 U20306 ( .B1(n20376), .B2(n18199), .A(n18187), .ZN(P3_U3045) );
  AOI22_X1 U20307 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n18194), .B1(
        P3_ADDRESS_REG_14__SCAN_IN), .B2(n21724), .ZN(n18188) );
  OAI21_X1 U20308 ( .B1(n21159), .B2(n18199), .A(n18188), .ZN(P3_U3046) );
  AOI22_X1 U20309 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n18194), .B1(
        P3_ADDRESS_REG_15__SCAN_IN), .B2(n21724), .ZN(n18189) );
  OAI21_X1 U20310 ( .B1(n20394), .B2(n18199), .A(n18189), .ZN(P3_U3047) );
  AOI22_X1 U20311 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n18194), .B1(
        P3_ADDRESS_REG_16__SCAN_IN), .B2(n21724), .ZN(n18190) );
  OAI21_X1 U20312 ( .B1(n21143), .B2(n18199), .A(n18190), .ZN(P3_U3048) );
  AOI22_X1 U20313 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n18194), .B1(
        P3_ADDRESS_REG_17__SCAN_IN), .B2(n21724), .ZN(n18191) );
  OAI21_X1 U20314 ( .B1(n20416), .B2(n18199), .A(n18191), .ZN(P3_U3049) );
  INV_X1 U20315 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20429) );
  AOI22_X1 U20316 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n18194), .B1(
        P3_ADDRESS_REG_18__SCAN_IN), .B2(n21724), .ZN(n18192) );
  OAI21_X1 U20317 ( .B1(n20429), .B2(n18199), .A(n18192), .ZN(P3_U3050) );
  AOI22_X1 U20318 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18194), .B1(
        P3_ADDRESS_REG_19__SCAN_IN), .B2(n21724), .ZN(n18193) );
  OAI21_X1 U20319 ( .B1(n20442), .B2(n18199), .A(n18193), .ZN(P3_U3051) );
  INV_X1 U20320 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20447) );
  AOI22_X1 U20321 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n18194), .B1(
        P3_ADDRESS_REG_20__SCAN_IN), .B2(n21724), .ZN(n18195) );
  OAI21_X1 U20322 ( .B1(n20447), .B2(n18199), .A(n18195), .ZN(P3_U3052) );
  AOI22_X1 U20323 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_21__SCAN_IN), .B2(n18214), .ZN(n18196) );
  OAI21_X1 U20324 ( .B1(n20468), .B2(n18199), .A(n18196), .ZN(P3_U3053) );
  INV_X1 U20325 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20486) );
  AOI22_X1 U20326 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_22__SCAN_IN), .B2(n18214), .ZN(n18197) );
  OAI21_X1 U20327 ( .B1(n20486), .B2(n18199), .A(n18197), .ZN(P3_U3054) );
  AOI22_X1 U20328 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_23__SCAN_IN), .B2(n21724), .ZN(n18198) );
  OAI21_X1 U20329 ( .B1(n20501), .B2(n18199), .A(n18198), .ZN(P3_U3055) );
  INV_X1 U20330 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21043) );
  AOI22_X1 U20331 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_24__SCAN_IN), .B2(n18214), .ZN(n18200) );
  OAI21_X1 U20332 ( .B1(n21043), .B2(n18209), .A(n18200), .ZN(P3_U3056) );
  AOI22_X1 U20333 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_25__SCAN_IN), .B2(n18214), .ZN(n18201) );
  OAI21_X1 U20334 ( .B1(n20539), .B2(n18209), .A(n18201), .ZN(P3_U3057) );
  INV_X1 U20335 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n20540) );
  AOI22_X1 U20336 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n18214), .ZN(n18202) );
  OAI21_X1 U20337 ( .B1(n20540), .B2(n18209), .A(n18202), .ZN(P3_U3058) );
  AOI22_X1 U20338 ( .A1(n18203), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_ADDRESS_REG_27__SCAN_IN), .B2(n18214), .ZN(n18204) );
  OAI21_X1 U20339 ( .B1(n18207), .B2(n20540), .A(n18204), .ZN(P3_U3059) );
  AOI22_X1 U20340 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n18205), .B1(
        P3_ADDRESS_REG_28__SCAN_IN), .B2(n18214), .ZN(n18206) );
  OAI21_X1 U20341 ( .B1(n20569), .B2(n18209), .A(n18206), .ZN(P3_U3060) );
  INV_X1 U20342 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19818) );
  OAI222_X1 U20343 ( .A1(n18209), .A2(n18208), .B1(n19818), .B2(n21682), .C1(
        n20569), .C2(n18207), .ZN(P3_U3061) );
  INV_X1 U20344 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18210) );
  AOI22_X1 U20345 ( .A1(n21682), .A2(n18211), .B1(n18210), .B2(n18214), .ZN(
        P3_U3277) );
  INV_X1 U20346 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18212) );
  AOI22_X1 U20347 ( .A1(n21682), .A2(n18213), .B1(n18212), .B2(n18214), .ZN(
        P3_U3276) );
  INV_X1 U20348 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18215) );
  AOI22_X1 U20349 ( .A1(n21682), .A2(n18216), .B1(n18215), .B2(n18214), .ZN(
        P3_U3275) );
  MUX2_X1 U20350 ( .A(P3_BE_N_REG_3__SCAN_IN), .B(P3_BYTEENABLE_REG_3__SCAN_IN), .S(n21682), .Z(P3_U3274) );
  NOR4_X1 U20351 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18219)
         );
  NOR4_X1 U20352 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18217), .ZN(n18218) );
  NAND3_X1 U20353 ( .A1(n18219), .A2(n18218), .A3(U215), .ZN(U213) );
  INV_X1 U20354 ( .A(n18220), .ZN(n18225) );
  INV_X1 U20355 ( .A(n18221), .ZN(n18224) );
  NAND4_X1 U20356 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n14714), .A4(n18222), .ZN(n18223) );
  OAI211_X1 U20357 ( .C1(n18619), .C2(n18225), .A(n18224), .B(n18223), .ZN(
        n18235) );
  INV_X1 U20358 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n18234) );
  NOR2_X1 U20359 ( .A1(n21699), .A2(n19214), .ZN(n18226) );
  NOR2_X1 U20360 ( .A1(n18226), .A2(n18605), .ZN(n18232) );
  INV_X1 U20361 ( .A(n18228), .ZN(n21708) );
  AND3_X1 U20362 ( .A1(n19642), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n21708), 
        .ZN(n18230) );
  AOI21_X1 U20363 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n18228), .A(n18227), 
        .ZN(n18229) );
  MUX2_X1 U20364 ( .A(n18230), .B(n18229), .S(n19585), .Z(n18231) );
  OAI21_X1 U20365 ( .B1(n18232), .B2(n18231), .A(n18235), .ZN(n18233) );
  OAI21_X1 U20366 ( .B1(n18235), .B2(n18234), .A(n18233), .ZN(P2_U3610) );
  AOI22_X1 U20367 ( .A1(n18470), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n18500), .B2(
        n18236), .ZN(n18239) );
  NAND2_X1 U20368 ( .A1(n18471), .A2(n18237), .ZN(n18238) );
  OAI211_X1 U20369 ( .C1(n18493), .C2(n18240), .A(n18239), .B(n18238), .ZN(
        n18243) );
  NOR2_X1 U20370 ( .A1(n19141), .A2(n18241), .ZN(n18242) );
  AOI211_X1 U20371 ( .C1(n18501), .C2(n18244), .A(n18243), .B(n18242), .ZN(
        n18246) );
  OAI21_X1 U20372 ( .B1(n18498), .B2(n18321), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18245) );
  OAI211_X1 U20373 ( .C1(n18247), .C2(n18505), .A(n18246), .B(n18245), .ZN(
        P2_U2855) );
  OAI21_X1 U20374 ( .B1(n18490), .B2(n18248), .A(n14141), .ZN(n18252) );
  OAI22_X1 U20375 ( .A1(n18494), .A2(n18250), .B1(n18249), .B2(n18329), .ZN(
        n18251) );
  AOI211_X1 U20376 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n18473), .A(n18252), .B(
        n18251), .ZN(n18259) );
  NAND2_X1 U20377 ( .A1(n18423), .A2(n18253), .ZN(n18254) );
  XNOR2_X1 U20378 ( .A(n18255), .B(n18254), .ZN(n18257) );
  AOI22_X1 U20379 ( .A1(n18257), .A2(n18482), .B1(n18501), .B2(n18256), .ZN(
        n18258) );
  OAI211_X1 U20380 ( .C1(n18476), .C2(n19377), .A(n18259), .B(n18258), .ZN(
        P2_U2850) );
  NAND2_X1 U20381 ( .A1(n18423), .A2(n18260), .ZN(n18262) );
  XOR2_X1 U20382 ( .A(n18262), .B(n18261), .Z(n18273) );
  NAND2_X1 U20383 ( .A1(n18470), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n18264) );
  AOI21_X1 U20384 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18498), .A(
        n18559), .ZN(n18263) );
  OAI211_X1 U20385 ( .C1(n18265), .C2(n18493), .A(n18264), .B(n18263), .ZN(
        n18266) );
  AOI21_X1 U20386 ( .B1(n18471), .B2(n18267), .A(n18266), .ZN(n18268) );
  OAI21_X1 U20387 ( .B1(n18269), .B2(n18478), .A(n18268), .ZN(n18270) );
  AOI21_X1 U20388 ( .B1(n18271), .B2(n18500), .A(n18270), .ZN(n18272) );
  OAI21_X1 U20389 ( .B1(n18273), .B2(n18602), .A(n18272), .ZN(P2_U2848) );
  NAND2_X1 U20390 ( .A1(n18470), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n18274) );
  OAI211_X1 U20391 ( .C1(n18275), .C2(n18329), .A(n18274), .B(n14141), .ZN(
        n18278) );
  NOR2_X1 U20392 ( .A1(n18276), .A2(n18494), .ZN(n18277) );
  AOI211_X1 U20393 ( .C1(n18473), .C2(P2_REIP_REG_9__SCAN_IN), .A(n18278), .B(
        n18277), .ZN(n18285) );
  NAND2_X1 U20394 ( .A1(n18423), .A2(n18279), .ZN(n18280) );
  XNOR2_X1 U20395 ( .A(n18281), .B(n18280), .ZN(n18283) );
  AOI22_X1 U20396 ( .A1(n18283), .A2(n18482), .B1(n18282), .B2(n18501), .ZN(
        n18284) );
  OAI211_X1 U20397 ( .C1(n19101), .C2(n18476), .A(n18285), .B(n18284), .ZN(
        P2_U2846) );
  AOI22_X1 U20398 ( .A1(n18470), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18474), .ZN(n18286) );
  OAI21_X1 U20399 ( .B1(n18287), .B2(n18494), .A(n18286), .ZN(n18288) );
  AOI211_X1 U20400 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n18473), .A(n18559), 
        .B(n18288), .ZN(n18295) );
  NOR2_X1 U20401 ( .A1(n18436), .A2(n18289), .ZN(n18291) );
  XNOR2_X1 U20402 ( .A(n18291), .B(n18290), .ZN(n18293) );
  AOI22_X1 U20403 ( .A1(n18293), .A2(n18482), .B1(n18292), .B2(n18501), .ZN(
        n18294) );
  OAI211_X1 U20404 ( .C1(n19098), .C2(n18476), .A(n18295), .B(n18294), .ZN(
        P2_U2845) );
  INV_X1 U20405 ( .A(n18296), .ZN(n18304) );
  OAI22_X1 U20406 ( .A1(n18297), .A2(n18329), .B1(n16457), .B2(n18493), .ZN(
        n18298) );
  INV_X1 U20407 ( .A(n18298), .ZN(n18303) );
  OAI21_X1 U20408 ( .B1(n18490), .B2(n18299), .A(n14141), .ZN(n18300) );
  AOI21_X1 U20409 ( .B1(n18301), .B2(n18501), .A(n18300), .ZN(n18302) );
  OAI211_X1 U20410 ( .C1(n18304), .C2(n18494), .A(n18303), .B(n18302), .ZN(
        n18305) );
  AOI21_X1 U20411 ( .B1(n18306), .B2(n18500), .A(n18305), .ZN(n18311) );
  INV_X1 U20412 ( .A(n18307), .ZN(n18309) );
  OAI211_X1 U20413 ( .C1(n18309), .C2(n18312), .A(n18482), .B(n18308), .ZN(
        n18310) );
  OAI211_X1 U20414 ( .C1(n18313), .C2(n18312), .A(n18311), .B(n18310), .ZN(
        P2_U2844) );
  INV_X1 U20415 ( .A(n18314), .ZN(n18317) );
  AOI21_X1 U20416 ( .B1(n18470), .B2(P2_EBX_REG_15__SCAN_IN), .A(n18559), .ZN(
        n18315) );
  OAI21_X1 U20417 ( .B1(n14969), .B2(n18493), .A(n18315), .ZN(n18316) );
  AOI21_X1 U20418 ( .B1(n18317), .B2(n18471), .A(n18316), .ZN(n18328) );
  INV_X1 U20419 ( .A(n18318), .ZN(n18325) );
  AOI21_X1 U20420 ( .B1(n18319), .B2(n18322), .A(n18505), .ZN(n18320) );
  AOI21_X1 U20421 ( .B1(n18322), .B2(n18321), .A(n18320), .ZN(n18324) );
  OAI222_X1 U20422 ( .A1(n18478), .A2(n18325), .B1(n18324), .B2(n18323), .C1(
        n19081), .C2(n18476), .ZN(n18326) );
  INV_X1 U20423 ( .A(n18326), .ZN(n18327) );
  OAI211_X1 U20424 ( .C1(n18330), .C2(n18329), .A(n18328), .B(n18327), .ZN(
        P2_U2840) );
  NAND2_X1 U20425 ( .A1(n18423), .A2(n18331), .ZN(n18332) );
  XOR2_X1 U20426 ( .A(n18333), .B(n18332), .Z(n18342) );
  AOI22_X1 U20427 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18498), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n18473), .ZN(n18334) );
  OAI211_X1 U20428 ( .C1(n18490), .C2(n18335), .A(n18334), .B(n18521), .ZN(
        n18336) );
  AOI21_X1 U20429 ( .B1(n18337), .B2(n18471), .A(n18336), .ZN(n18341) );
  AOI22_X1 U20430 ( .A1(n18339), .A2(n18501), .B1(n18338), .B2(n18500), .ZN(
        n18340) );
  OAI211_X1 U20431 ( .C1(n18602), .C2(n18342), .A(n18341), .B(n18340), .ZN(
        P2_U2838) );
  NOR2_X1 U20432 ( .A1(n18436), .A2(n18343), .ZN(n18345) );
  XOR2_X1 U20433 ( .A(n18345), .B(n18344), .Z(n18354) );
  AOI22_X1 U20434 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18498), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n18473), .ZN(n18346) );
  OAI211_X1 U20435 ( .C1(n18490), .C2(n18347), .A(n18346), .B(n18521), .ZN(
        n18348) );
  AOI21_X1 U20436 ( .B1(n18349), .B2(n18471), .A(n18348), .ZN(n18353) );
  AOI21_X1 U20437 ( .B1(n18351), .B2(n11044), .A(n18350), .ZN(n19518) );
  AOI22_X1 U20438 ( .A1(n18501), .A2(n18548), .B1(n18500), .B2(n19518), .ZN(
        n18352) );
  OAI211_X1 U20439 ( .C1(n18602), .C2(n18354), .A(n18353), .B(n18352), .ZN(
        P2_U2837) );
  NAND2_X1 U20440 ( .A1(n18423), .A2(n18355), .ZN(n18356) );
  XOR2_X1 U20441 ( .A(n18357), .B(n18356), .Z(n18366) );
  INV_X1 U20442 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n18359) );
  AOI22_X1 U20443 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18498), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n18473), .ZN(n18358) );
  OAI211_X1 U20444 ( .C1(n18490), .C2(n18359), .A(n18358), .B(n18521), .ZN(
        n18360) );
  AOI21_X1 U20445 ( .B1(n18361), .B2(n18471), .A(n18360), .ZN(n18365) );
  AOI22_X1 U20446 ( .A1(n18501), .A2(n18363), .B1(n18362), .B2(n18500), .ZN(
        n18364) );
  OAI211_X1 U20447 ( .C1(n18602), .C2(n18366), .A(n18365), .B(n18364), .ZN(
        P2_U2836) );
  NOR2_X1 U20448 ( .A1(n18436), .A2(n18367), .ZN(n18368) );
  XOR2_X1 U20449 ( .A(n18369), .B(n18368), .Z(n18380) );
  AOI21_X1 U20450 ( .B1(n18371), .B2(n11006), .A(n18370), .ZN(n19420) );
  INV_X1 U20451 ( .A(n18372), .ZN(n18377) );
  INV_X1 U20452 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n18374) );
  AOI22_X1 U20453 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18498), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18473), .ZN(n18373) );
  OAI21_X1 U20454 ( .B1(n18490), .B2(n18374), .A(n18373), .ZN(n18375) );
  AOI21_X1 U20455 ( .B1(n18533), .B2(n18501), .A(n18375), .ZN(n18376) );
  OAI21_X1 U20456 ( .B1(n18377), .B2(n18494), .A(n18376), .ZN(n18378) );
  AOI21_X1 U20457 ( .B1(n19420), .B2(n18500), .A(n18378), .ZN(n18379) );
  OAI21_X1 U20458 ( .B1(n18602), .B2(n18380), .A(n18379), .ZN(P2_U2835) );
  OAI222_X1 U20459 ( .A1(n18494), .A2(n18382), .B1(n18493), .B2(n17277), .C1(
        n18490), .C2(n18381), .ZN(n18383) );
  AOI21_X1 U20460 ( .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18498), .A(
        n18383), .ZN(n18390) );
  AOI21_X1 U20461 ( .B1(n18385), .B2(n18384), .A(n18602), .ZN(n18388) );
  AOI22_X1 U20462 ( .A1(n18388), .A2(n18387), .B1(n18386), .B2(n18501), .ZN(
        n18389) );
  OAI211_X1 U20463 ( .C1(n18391), .C2(n18476), .A(n18390), .B(n18389), .ZN(
        P2_U2834) );
  AOI22_X1 U20464 ( .A1(n18392), .A2(n18471), .B1(P2_REIP_REG_22__SCAN_IN), 
        .B2(n18473), .ZN(n18400) );
  AOI22_X1 U20465 ( .A1(n18470), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18474), .ZN(n18399) );
  AOI22_X1 U20466 ( .A1(n18501), .A2(n18393), .B1(n19322), .B2(n18500), .ZN(
        n18398) );
  OAI211_X1 U20467 ( .C1(n18396), .C2(n18395), .A(n18482), .B(n18394), .ZN(
        n18397) );
  NAND4_X1 U20468 ( .A1(n18400), .A2(n18399), .A3(n18398), .A4(n18397), .ZN(
        P2_U2833) );
  AOI22_X1 U20469 ( .A1(n18401), .A2(n18471), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n18470), .ZN(n18411) );
  AOI22_X1 U20470 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18498), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18473), .ZN(n18410) );
  INV_X1 U20471 ( .A(n18402), .ZN(n18404) );
  AOI22_X1 U20472 ( .A1(n18404), .A2(n18501), .B1(n18403), .B2(n18500), .ZN(
        n18409) );
  OAI211_X1 U20473 ( .C1(n18407), .C2(n18406), .A(n18482), .B(n18405), .ZN(
        n18408) );
  NAND4_X1 U20474 ( .A1(n18411), .A2(n18410), .A3(n18409), .A4(n18408), .ZN(
        P2_U2832) );
  AOI22_X1 U20475 ( .A1(n18412), .A2(n18471), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n18470), .ZN(n18421) );
  AOI22_X1 U20476 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18474), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18473), .ZN(n18420) );
  INV_X1 U20477 ( .A(n18413), .ZN(n18415) );
  AOI22_X1 U20478 ( .A1(n18415), .A2(n18501), .B1(n18414), .B2(n18500), .ZN(
        n18419) );
  OAI211_X1 U20479 ( .C1(n18417), .C2(n18416), .A(n18482), .B(n18422), .ZN(
        n18418) );
  NAND4_X1 U20480 ( .A1(n18421), .A2(n18420), .A3(n18419), .A4(n18418), .ZN(
        P2_U2831) );
  NAND2_X1 U20481 ( .A1(n18423), .A2(n18422), .ZN(n18425) );
  XOR2_X1 U20482 ( .A(n18425), .B(n18424), .Z(n18434) );
  AOI22_X1 U20483 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18498), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n18473), .ZN(n18426) );
  OAI21_X1 U20484 ( .B1(n18490), .B2(n16215), .A(n18426), .ZN(n18427) );
  AOI21_X1 U20485 ( .B1(n18428), .B2(n18500), .A(n18427), .ZN(n18429) );
  OAI21_X1 U20486 ( .B1(n18430), .B2(n18478), .A(n18429), .ZN(n18431) );
  AOI21_X1 U20487 ( .B1(n18432), .B2(n18471), .A(n18431), .ZN(n18433) );
  OAI21_X1 U20488 ( .B1(n18434), .B2(n18602), .A(n18433), .ZN(P2_U2830) );
  NOR2_X1 U20489 ( .A1(n18436), .A2(n18435), .ZN(n18437) );
  XOR2_X1 U20490 ( .A(n18438), .B(n18437), .Z(n18446) );
  AOI22_X1 U20491 ( .A1(n18470), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18474), .ZN(n18441) );
  AOI22_X1 U20492 ( .A1(n18473), .A2(P2_REIP_REG_26__SCAN_IN), .B1(n18500), 
        .B2(n18439), .ZN(n18440) );
  OAI211_X1 U20493 ( .C1(n18442), .C2(n18478), .A(n18441), .B(n18440), .ZN(
        n18443) );
  AOI21_X1 U20494 ( .B1(n18444), .B2(n18471), .A(n18443), .ZN(n18445) );
  OAI21_X1 U20495 ( .B1(n18602), .B2(n18446), .A(n18445), .ZN(P2_U2829) );
  INV_X1 U20496 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n18447) );
  OAI222_X1 U20497 ( .A1(n18494), .A2(n18449), .B1(n18493), .B2(n18448), .C1(
        n18490), .C2(n18447), .ZN(n18450) );
  AOI21_X1 U20498 ( .B1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18498), .A(
        n18450), .ZN(n18457) );
  AOI21_X1 U20499 ( .B1(n18452), .B2(n18451), .A(n18602), .ZN(n18455) );
  AOI22_X1 U20500 ( .A1(n18455), .A2(n18454), .B1(n18453), .B2(n18501), .ZN(
        n18456) );
  OAI211_X1 U20501 ( .C1(n18458), .C2(n18476), .A(n18457), .B(n18456), .ZN(
        P2_U2828) );
  INV_X1 U20502 ( .A(n18459), .ZN(n18460) );
  AOI22_X1 U20503 ( .A1(n18460), .A2(n18471), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n18470), .ZN(n18469) );
  AOI22_X1 U20504 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18474), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18473), .ZN(n18468) );
  AOI22_X1 U20505 ( .A1(n18462), .A2(n18501), .B1(n18461), .B2(n18500), .ZN(
        n18467) );
  OAI211_X1 U20506 ( .C1(n18465), .C2(n18464), .A(n18482), .B(n18463), .ZN(
        n18466) );
  NAND4_X1 U20507 ( .A1(n18469), .A2(n18468), .A3(n18467), .A4(n18466), .ZN(
        P2_U2827) );
  AOI22_X1 U20508 ( .A1(n18472), .A2(n18471), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n18470), .ZN(n18488) );
  AOI22_X1 U20509 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18474), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18473), .ZN(n18487) );
  INV_X1 U20510 ( .A(n18475), .ZN(n18477) );
  OAI22_X1 U20511 ( .A1(n18479), .A2(n18478), .B1(n18477), .B2(n18476), .ZN(
        n18480) );
  INV_X1 U20512 ( .A(n18480), .ZN(n18486) );
  OAI211_X1 U20513 ( .C1(n18484), .C2(n18483), .A(n18482), .B(n18481), .ZN(
        n18485) );
  NAND4_X1 U20514 ( .A1(n18488), .A2(n18487), .A3(n18486), .A4(n18485), .ZN(
        P2_U2826) );
  NOR2_X1 U20515 ( .A1(n18490), .A2(n18489), .ZN(n18497) );
  INV_X1 U20516 ( .A(n18491), .ZN(n18495) );
  OAI22_X1 U20517 ( .A1(n18495), .A2(n18494), .B1(n18493), .B2(n18492), .ZN(
        n18496) );
  AOI211_X1 U20518 ( .C1(n18498), .C2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n18497), .B(n18496), .ZN(n18504) );
  AOI22_X1 U20519 ( .A1(n18502), .A2(n18501), .B1(n18500), .B2(n18499), .ZN(
        n18503) );
  OAI211_X1 U20520 ( .C1(n18506), .C2(n18505), .A(n18504), .B(n18503), .ZN(
        P2_U2824) );
  AOI22_X1 U20521 ( .A1(n18566), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18582), .B2(n18507), .ZN(n18516) );
  OAI22_X1 U20522 ( .A1(n18576), .A2(n18509), .B1(n18579), .B2(n18508), .ZN(
        n18514) );
  OAI21_X1 U20523 ( .B1(n18512), .B2(n18511), .A(n18510), .ZN(n18513) );
  NOR2_X1 U20524 ( .A1(n18514), .A2(n18513), .ZN(n18515) );
  OAI211_X1 U20525 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18517), .A(
        n18516), .B(n18515), .ZN(P2_U3046) );
  AOI21_X1 U20526 ( .B1(n18520), .B2(n18519), .A(n18518), .ZN(n18531) );
  NOR2_X1 U20527 ( .A1(n18521), .A2(n16143), .ZN(n18522) );
  AOI211_X1 U20528 ( .C1(n18524), .C2(n18553), .A(n18523), .B(n18522), .ZN(
        n18529) );
  AOI222_X1 U20529 ( .A1(n18527), .A2(n18582), .B1(n18584), .B2(n18526), .C1(
        n18525), .C2(n18556), .ZN(n18528) );
  OAI211_X1 U20530 ( .C1(n18531), .C2(n18530), .A(n18529), .B(n18528), .ZN(
        P2_U3034) );
  AOI22_X1 U20531 ( .A1(n18532), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18553), .B2(n19420), .ZN(n18543) );
  AOI222_X1 U20532 ( .A1(n18535), .A2(n18582), .B1(n18556), .B2(n18534), .C1(
        n18584), .C2(n18533), .ZN(n18542) );
  NAND2_X1 U20533 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n18559), .ZN(n18541) );
  OAI221_X1 U20534 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C1(n18539), .C2(n18538), .A(
        n18537), .ZN(n18540) );
  NAND4_X1 U20535 ( .A1(n18543), .A2(n18542), .A3(n18541), .A4(n18540), .ZN(
        P2_U3026) );
  NAND2_X1 U20536 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n18559), .ZN(n18544) );
  OAI211_X1 U20537 ( .C1(n18546), .C2(n15407), .A(n18545), .B(n18544), .ZN(
        n18547) );
  AOI21_X1 U20538 ( .B1(n19518), .B2(n18553), .A(n18547), .ZN(n18551) );
  AOI22_X1 U20539 ( .A1(n18549), .A2(n18582), .B1(n18584), .B2(n18548), .ZN(
        n18550) );
  OAI211_X1 U20540 ( .C1(n18576), .C2(n18552), .A(n18551), .B(n18550), .ZN(
        P2_U3028) );
  AOI22_X1 U20541 ( .A1(n18554), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n18553), .B2(n19102), .ZN(n18565) );
  AOI222_X1 U20542 ( .A1(n18558), .A2(n18582), .B1(n18584), .B2(n18557), .C1(
        n18556), .C2(n18555), .ZN(n18564) );
  NAND2_X1 U20543 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18559), .ZN(n18563) );
  OAI211_X1 U20544 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n18561), .B(n18560), .ZN(n18562) );
  NAND4_X1 U20545 ( .A1(n18565), .A2(n18564), .A3(n18563), .A4(n18562), .ZN(
        P2_U3038) );
  AOI21_X1 U20546 ( .B1(n18568), .B2(n18567), .A(n18566), .ZN(n18594) );
  INV_X1 U20547 ( .A(n18569), .ZN(n18575) );
  NAND2_X1 U20548 ( .A1(n18571), .A2(n18570), .ZN(n18572) );
  NAND2_X1 U20549 ( .A1(n18573), .A2(n18572), .ZN(n18574) );
  OAI21_X1 U20550 ( .B1(n18576), .B2(n18575), .A(n18574), .ZN(n18581) );
  INV_X1 U20551 ( .A(n19523), .ZN(n18578) );
  OAI22_X1 U20552 ( .A1(n18579), .A2(n18578), .B1(n18577), .B2(n14141), .ZN(
        n18580) );
  NOR2_X1 U20553 ( .A1(n18581), .A2(n18580), .ZN(n18591) );
  NAND2_X1 U20554 ( .A1(n18583), .A2(n18582), .ZN(n18590) );
  NAND2_X1 U20555 ( .A1(n15005), .A2(n18584), .ZN(n18589) );
  INV_X1 U20556 ( .A(n18585), .ZN(n18587) );
  NAND2_X1 U20557 ( .A1(n18587), .A2(n18586), .ZN(n18588) );
  AND4_X1 U20558 ( .A1(n18591), .A2(n18590), .A3(n18589), .A4(n18588), .ZN(
        n18592) );
  OAI21_X1 U20559 ( .B1(n18594), .B2(n18593), .A(n18592), .ZN(P2_U3044) );
  AND2_X1 U20560 ( .A1(n18613), .A2(n18595), .ZN(n18608) );
  INV_X1 U20561 ( .A(n18608), .ZN(n18601) );
  OAI21_X1 U20562 ( .B1(n18597), .B2(n18596), .A(n18616), .ZN(n18600) );
  NAND2_X1 U20563 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n21699), .ZN(n18598) );
  AOI21_X1 U20564 ( .B1(n18604), .B2(n18601), .A(n18598), .ZN(n18599) );
  AOI21_X1 U20565 ( .B1(n18601), .B2(n18600), .A(n18599), .ZN(n18603) );
  NAND2_X1 U20566 ( .A1(n18603), .A2(n18602), .ZN(P2_U3177) );
  INV_X1 U20567 ( .A(n18604), .ZN(n18611) );
  AOI21_X1 U20568 ( .B1(n14714), .B2(n18606), .A(n18605), .ZN(n18607) );
  AOI21_X1 U20569 ( .B1(n18608), .B2(n21699), .A(n18607), .ZN(n18609) );
  AOI211_X1 U20570 ( .C1(n18611), .C2(n21699), .A(n18610), .B(n18609), .ZN(
        n18615) );
  OAI21_X1 U20571 ( .B1(n18613), .B2(n18612), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18614) );
  OAI211_X1 U20572 ( .C1(n18617), .C2(n18616), .A(n18615), .B(n18614), .ZN(
        P2_U3176) );
  NAND2_X1 U20573 ( .A1(n18619), .A2(n18618), .ZN(n18622) );
  NAND2_X1 U20574 ( .A1(n18622), .A2(P2_MORE_REG_SCAN_IN), .ZN(n18620) );
  OAI21_X1 U20575 ( .B1(n18622), .B2(n18621), .A(n18620), .ZN(P2_U3609) );
  INV_X1 U20576 ( .A(n18622), .ZN(n18625) );
  OAI21_X1 U20577 ( .B1(n18625), .B2(n18624), .A(n18623), .ZN(P2_U2819) );
  OAI22_X1 U20578 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n18977), .ZN(n18626) );
  INV_X1 U20579 ( .A(n18626), .ZN(U282) );
  OAI22_X1 U20580 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18977), .ZN(n18627) );
  INV_X1 U20581 ( .A(n18627), .ZN(U281) );
  OAI22_X1 U20582 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18977), .ZN(n18628) );
  INV_X1 U20583 ( .A(n18628), .ZN(U280) );
  OAI22_X1 U20584 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18977), .ZN(n18629) );
  INV_X1 U20585 ( .A(n18629), .ZN(U279) );
  OAI22_X1 U20586 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18977), .ZN(n18630) );
  INV_X1 U20587 ( .A(n18630), .ZN(U278) );
  OAI22_X1 U20588 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18977), .ZN(n18631) );
  INV_X1 U20589 ( .A(n18631), .ZN(U277) );
  OAI22_X1 U20590 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18977), .ZN(n18632) );
  INV_X1 U20591 ( .A(n18632), .ZN(U276) );
  OAI22_X1 U20592 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18977), .ZN(n18633) );
  INV_X1 U20593 ( .A(n18633), .ZN(U275) );
  INV_X1 U20594 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n18634) );
  INV_X1 U20595 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n20740) );
  AOI22_X1 U20596 ( .A1(n18977), .A2(n18634), .B1(n20740), .B2(U215), .ZN(U274) );
  OAI22_X1 U20597 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n18977), .ZN(n18635) );
  INV_X1 U20598 ( .A(n18635), .ZN(U273) );
  INV_X1 U20599 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n18636) );
  INV_X1 U20600 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n20657) );
  AOI22_X1 U20601 ( .A1(n18649), .A2(n18636), .B1(n20657), .B2(U215), .ZN(U272) );
  OAI22_X1 U20602 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18977), .ZN(n18637) );
  INV_X1 U20603 ( .A(n18637), .ZN(U271) );
  OAI22_X1 U20604 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18649), .ZN(n18638) );
  INV_X1 U20605 ( .A(n18638), .ZN(U270) );
  OAI22_X1 U20606 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18649), .ZN(n18639) );
  INV_X1 U20607 ( .A(n18639), .ZN(U269) );
  OAI22_X1 U20608 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18649), .ZN(n18640) );
  INV_X1 U20609 ( .A(n18640), .ZN(U268) );
  OAI22_X1 U20610 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18649), .ZN(n18641) );
  INV_X1 U20611 ( .A(n18641), .ZN(U267) );
  OAI22_X1 U20612 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18649), .ZN(n18642) );
  INV_X1 U20613 ( .A(n18642), .ZN(U266) );
  OAI22_X1 U20614 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n18649), .ZN(n18643) );
  INV_X1 U20615 ( .A(n18643), .ZN(U265) );
  OAI22_X1 U20616 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n18649), .ZN(n18644) );
  INV_X1 U20617 ( .A(n18644), .ZN(U264) );
  INV_X1 U20618 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n18645) );
  INV_X1 U20619 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n20609) );
  AOI22_X1 U20620 ( .A1(n18977), .A2(n18645), .B1(n20609), .B2(U215), .ZN(U263) );
  INV_X1 U20621 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n18646) );
  INV_X1 U20622 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n20614) );
  AOI22_X1 U20623 ( .A1(n18649), .A2(n18646), .B1(n20614), .B2(U215), .ZN(U262) );
  OAI22_X1 U20624 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n18977), .ZN(n18647) );
  INV_X1 U20625 ( .A(n18647), .ZN(U261) );
  INV_X1 U20626 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n18648) );
  INV_X1 U20627 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n20623) );
  AOI22_X1 U20628 ( .A1(n18649), .A2(n18648), .B1(n20623), .B2(U215), .ZN(U260) );
  OAI22_X1 U20629 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n18977), .ZN(n18650) );
  INV_X1 U20630 ( .A(n18650), .ZN(U259) );
  INV_X1 U20631 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n18651) );
  INV_X1 U20632 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20629) );
  AOI22_X1 U20633 ( .A1(n18977), .A2(n18651), .B1(n20629), .B2(U215), .ZN(U258) );
  NOR3_X1 U20634 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18652), .A3(
        n21228), .ZN(n18661) );
  NAND2_X1 U20635 ( .A1(n18661), .A2(n21216), .ZN(n18896) );
  NAND2_X1 U20636 ( .A1(n18978), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18710) );
  INV_X1 U20637 ( .A(n18661), .ZN(n18660) );
  NOR2_X2 U20638 ( .A1(n21216), .A2(n18660), .ZN(n18990) );
  NOR2_X1 U20639 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21252), .ZN(n20154) );
  INV_X1 U20640 ( .A(n20154), .ZN(n21241) );
  NOR2_X1 U20641 ( .A1(n21228), .A2(n18672), .ZN(n18718) );
  AND2_X1 U20642 ( .A1(n21241), .A2(n18718), .ZN(n18980) );
  NOR2_X2 U20643 ( .A1(n20629), .A2(n18979), .ZN(n18723) );
  AOI22_X1 U20644 ( .A1(n18990), .A2(n18724), .B1(n18980), .B2(n18723), .ZN(
        n18657) );
  NOR2_X1 U20645 ( .A1(n18653), .A2(n18979), .ZN(n18669) );
  AOI22_X1 U20646 ( .A1(n18978), .A2(n18661), .B1(n18718), .B2(n18669), .ZN(
        n18982) );
  NAND2_X1 U20647 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18718), .ZN(
        n18967) );
  INV_X1 U20648 ( .A(n18967), .ZN(n19060) );
  INV_X1 U20649 ( .A(n18654), .ZN(n18655) );
  NAND2_X1 U20650 ( .A1(n21248), .A2(n18655), .ZN(n18981) );
  NOR2_X2 U20651 ( .A1(n20667), .A2(n18981), .ZN(n18722) );
  AOI22_X1 U20652 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18982), .B1(
        n19060), .B2(n18722), .ZN(n18656) );
  OAI211_X1 U20653 ( .C1(n18896), .C2(n18710), .A(n18657), .B(n18656), .ZN(
        P3_U2995) );
  INV_X1 U20654 ( .A(n18724), .ZN(n18721) );
  INV_X1 U20655 ( .A(n18710), .ZN(n18728) );
  NAND2_X1 U20656 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18681), .ZN(
        n18668) );
  NOR2_X2 U20657 ( .A1(n21216), .A2(n18668), .ZN(n19002) );
  INV_X1 U20658 ( .A(n18990), .ZN(n19076) );
  NAND2_X1 U20659 ( .A1(n21216), .A2(n18718), .ZN(n19065) );
  NAND2_X1 U20660 ( .A1(n19076), .A2(n19065), .ZN(n18727) );
  AND2_X1 U20661 ( .A1(n21241), .A2(n18727), .ZN(n18985) );
  AOI22_X1 U20662 ( .A1(n18728), .A2(n19002), .B1(n18723), .B2(n18985), .ZN(
        n18659) );
  INV_X1 U20663 ( .A(n19002), .ZN(n18994) );
  NAND2_X1 U20664 ( .A1(n18896), .A2(n18994), .ZN(n18665) );
  AOI21_X1 U20665 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18979), .ZN(n18726) );
  OAI221_X1 U20666 ( .B1(n18727), .B2(n18693), .C1(n18727), .C2(n18665), .A(
        n18726), .ZN(n18986) );
  INV_X1 U20667 ( .A(n19065), .ZN(n19069) );
  AOI22_X1 U20668 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18986), .B1(
        n18722), .B2(n19069), .ZN(n18658) );
  OAI211_X1 U20669 ( .C1(n18896), .C2(n18721), .A(n18659), .B(n18658), .ZN(
        P3_U2987) );
  INV_X1 U20670 ( .A(n18668), .ZN(n18662) );
  NAND2_X1 U20671 ( .A1(n18662), .A2(n21216), .ZN(n19000) );
  NOR2_X1 U20672 ( .A1(n20154), .A2(n18660), .ZN(n18989) );
  AOI22_X1 U20673 ( .A1(n18724), .A2(n19002), .B1(n18723), .B2(n18989), .ZN(
        n18664) );
  AOI22_X1 U20674 ( .A1(n18978), .A2(n18662), .B1(n18669), .B2(n18661), .ZN(
        n18991) );
  AOI22_X1 U20675 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18991), .B1(
        n18722), .B2(n18990), .ZN(n18663) );
  OAI211_X1 U20676 ( .C1(n18710), .C2(n19000), .A(n18664), .B(n18663), .ZN(
        P3_U2979) );
  NOR2_X1 U20677 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21216), .ZN(
        n18702) );
  NAND2_X1 U20678 ( .A1(n18681), .A2(n18702), .ZN(n18943) );
  INV_X1 U20679 ( .A(n19000), .ZN(n19007) );
  AND2_X1 U20680 ( .A1(n21241), .A2(n18665), .ZN(n18995) );
  AOI22_X1 U20681 ( .A1(n18724), .A2(n19007), .B1(n18723), .B2(n18995), .ZN(
        n18667) );
  NAND2_X1 U20682 ( .A1(n19000), .A2(n18943), .ZN(n18673) );
  AOI22_X1 U20683 ( .A1(n18978), .A2(n18673), .B1(n18726), .B2(n18665), .ZN(
        n18997) );
  INV_X1 U20684 ( .A(n18896), .ZN(n18996) );
  AOI22_X1 U20685 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18997), .B1(
        n18996), .B2(n18722), .ZN(n18666) );
  OAI211_X1 U20686 ( .C1(n18710), .C2(n18943), .A(n18667), .B(n18666), .ZN(
        P3_U2971) );
  NOR2_X1 U20687 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21221) );
  NAND2_X1 U20688 ( .A1(n21221), .A2(n18681), .ZN(n19011) );
  INV_X1 U20689 ( .A(n18943), .ZN(n19013) );
  NOR2_X1 U20690 ( .A1(n20154), .A2(n18668), .ZN(n19001) );
  AOI22_X1 U20691 ( .A1(n18724), .A2(n19013), .B1(n18723), .B2(n19001), .ZN(
        n18671) );
  INV_X1 U20692 ( .A(n18693), .ZN(n18675) );
  INV_X1 U20693 ( .A(n18669), .ZN(n18680) );
  AOI21_X1 U20694 ( .B1(n21217), .B2(n18675), .A(n18680), .ZN(n18707) );
  NAND2_X1 U20695 ( .A1(n18681), .A2(n18707), .ZN(n19003) );
  AOI22_X1 U20696 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19003), .B1(
        n18722), .B2(n19002), .ZN(n18670) );
  OAI211_X1 U20697 ( .C1(n18710), .C2(n19011), .A(n18671), .B(n18670), .ZN(
        P3_U2963) );
  NOR2_X1 U20698 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18672), .ZN(
        n18689) );
  NAND2_X1 U20699 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18689), .ZN(
        n18948) );
  INV_X1 U20700 ( .A(n19011), .ZN(n19018) );
  INV_X1 U20701 ( .A(n18673), .ZN(n18674) );
  NOR2_X1 U20702 ( .A1(n20154), .A2(n18674), .ZN(n19006) );
  AOI22_X1 U20703 ( .A1(n18724), .A2(n19018), .B1(n18723), .B2(n19006), .ZN(
        n18678) );
  INV_X1 U20704 ( .A(n18948), .ZN(n19024) );
  NOR2_X1 U20705 ( .A1(n19018), .A2(n19024), .ZN(n18684) );
  OAI21_X1 U20706 ( .B1(n18684), .B2(n18675), .A(n18674), .ZN(n18676) );
  OAI211_X1 U20707 ( .C1(n19007), .C2(n21252), .A(n18932), .B(n18676), .ZN(
        n19008) );
  AOI22_X1 U20708 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19008), .B1(
        n18722), .B2(n19007), .ZN(n18677) );
  OAI211_X1 U20709 ( .C1(n18710), .C2(n18948), .A(n18678), .B(n18677), .ZN(
        P3_U2955) );
  NAND2_X1 U20710 ( .A1(n18689), .A2(n21216), .ZN(n19022) );
  INV_X1 U20711 ( .A(n18681), .ZN(n18679) );
  NAND2_X1 U20712 ( .A1(n21217), .A2(n21241), .ZN(n18715) );
  NOR2_X1 U20713 ( .A1(n18679), .A2(n18715), .ZN(n19012) );
  AOI22_X1 U20714 ( .A1(n18724), .A2(n19024), .B1(n18723), .B2(n19012), .ZN(
        n18683) );
  NOR2_X1 U20715 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18680), .ZN(
        n18717) );
  AOI22_X1 U20716 ( .A1(n18978), .A2(n18689), .B1(n18681), .B2(n18717), .ZN(
        n19014) );
  AOI22_X1 U20717 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19014), .B1(
        n18722), .B2(n19013), .ZN(n18682) );
  OAI211_X1 U20718 ( .C1(n18710), .C2(n19022), .A(n18683), .B(n18682), .ZN(
        P3_U2947) );
  NAND2_X1 U20719 ( .A1(n18698), .A2(n18702), .ZN(n18951) );
  INV_X1 U20720 ( .A(n19022), .ZN(n19030) );
  NOR2_X1 U20721 ( .A1(n20154), .A2(n18684), .ZN(n19017) );
  AOI22_X1 U20722 ( .A1(n18724), .A2(n19030), .B1(n18723), .B2(n19017), .ZN(
        n18687) );
  NAND2_X1 U20723 ( .A1(n19022), .A2(n18951), .ZN(n18694) );
  INV_X1 U20724 ( .A(n18684), .ZN(n18685) );
  AOI22_X1 U20725 ( .A1(n18978), .A2(n18694), .B1(n18726), .B2(n18685), .ZN(
        n19019) );
  AOI22_X1 U20726 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19019), .B1(
        n18722), .B2(n19018), .ZN(n18686) );
  OAI211_X1 U20727 ( .C1(n18710), .C2(n18951), .A(n18687), .B(n18686), .ZN(
        P3_U2939) );
  INV_X1 U20728 ( .A(n21221), .ZN(n18688) );
  INV_X1 U20729 ( .A(n18698), .ZN(n18697) );
  NOR2_X2 U20730 ( .A1(n18688), .A2(n18697), .ZN(n19041) );
  INV_X1 U20731 ( .A(n18689), .ZN(n18690) );
  NOR2_X1 U20732 ( .A1(n20154), .A2(n18690), .ZN(n19023) );
  AOI22_X1 U20733 ( .A1(n18728), .A2(n19041), .B1(n18723), .B2(n19023), .ZN(
        n18692) );
  NAND2_X1 U20734 ( .A1(n18698), .A2(n18707), .ZN(n19025) );
  AOI22_X1 U20735 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19025), .B1(
        n18722), .B2(n19024), .ZN(n18691) );
  OAI211_X1 U20736 ( .C1(n18721), .C2(n18951), .A(n18692), .B(n18691), .ZN(
        P3_U2931) );
  INV_X1 U20737 ( .A(n19041), .ZN(n19028) );
  NOR2_X1 U20738 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18716) );
  NAND2_X1 U20739 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18716), .ZN(
        n18706) );
  NOR2_X2 U20740 ( .A1(n21216), .A2(n18706), .ZN(n19047) );
  AND2_X1 U20741 ( .A1(n21241), .A2(n18694), .ZN(n19029) );
  AOI22_X1 U20742 ( .A1(n18728), .A2(n19047), .B1(n18723), .B2(n19029), .ZN(
        n18696) );
  INV_X1 U20743 ( .A(n19047), .ZN(n19034) );
  NAND2_X1 U20744 ( .A1(n19028), .A2(n19034), .ZN(n18703) );
  OAI221_X1 U20745 ( .B1(n18694), .B2(n18693), .C1(n18694), .C2(n18703), .A(
        n18726), .ZN(n19031) );
  AOI22_X1 U20746 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19031), .B1(
        n18722), .B2(n19030), .ZN(n18695) );
  OAI211_X1 U20747 ( .C1(n18721), .C2(n19028), .A(n18696), .B(n18695), .ZN(
        P3_U2923) );
  INV_X1 U20748 ( .A(n18706), .ZN(n18699) );
  NAND2_X1 U20749 ( .A1(n18699), .A2(n21216), .ZN(n19045) );
  NOR2_X1 U20750 ( .A1(n18697), .A2(n18715), .ZN(n19035) );
  AOI22_X1 U20751 ( .A1(n18724), .A2(n19047), .B1(n18723), .B2(n19035), .ZN(
        n18701) );
  AOI22_X1 U20752 ( .A1(n18978), .A2(n18699), .B1(n18698), .B2(n18717), .ZN(
        n19037) );
  INV_X1 U20753 ( .A(n18951), .ZN(n19036) );
  AOI22_X1 U20754 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19037), .B1(
        n18722), .B2(n19036), .ZN(n18700) );
  OAI211_X1 U20755 ( .C1(n18710), .C2(n19045), .A(n18701), .B(n18700), .ZN(
        P3_U2915) );
  NAND2_X1 U20756 ( .A1(n18702), .A2(n18716), .ZN(n18964) );
  INV_X1 U20757 ( .A(n19045), .ZN(n19053) );
  AND2_X1 U20758 ( .A1(n21241), .A2(n18703), .ZN(n19040) );
  AOI22_X1 U20759 ( .A1(n18724), .A2(n19053), .B1(n18723), .B2(n19040), .ZN(
        n18705) );
  NAND2_X1 U20760 ( .A1(n19045), .A2(n18964), .ZN(n18711) );
  AOI22_X1 U20761 ( .A1(n18978), .A2(n18711), .B1(n18726), .B2(n18703), .ZN(
        n19042) );
  AOI22_X1 U20762 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19042), .B1(
        n18722), .B2(n19041), .ZN(n18704) );
  OAI211_X1 U20763 ( .C1(n18710), .C2(n18964), .A(n18705), .B(n18704), .ZN(
        P3_U2907) );
  NAND2_X1 U20764 ( .A1(n21221), .A2(n18716), .ZN(n19058) );
  INV_X1 U20765 ( .A(n18964), .ZN(n19061) );
  NOR2_X1 U20766 ( .A1(n20154), .A2(n18706), .ZN(n19046) );
  AOI22_X1 U20767 ( .A1(n18724), .A2(n19061), .B1(n18723), .B2(n19046), .ZN(
        n18709) );
  NAND2_X1 U20768 ( .A1(n18707), .A2(n18716), .ZN(n19048) );
  AOI22_X1 U20769 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19048), .B1(
        n18722), .B2(n19047), .ZN(n18708) );
  OAI211_X1 U20770 ( .C1(n18710), .C2(n19058), .A(n18709), .B(n18708), .ZN(
        P3_U2899) );
  AND2_X1 U20771 ( .A1(n21241), .A2(n18711), .ZN(n19051) );
  AOI22_X1 U20772 ( .A1(n18728), .A2(n19060), .B1(n18723), .B2(n19051), .ZN(
        n18713) );
  NAND2_X1 U20773 ( .A1(n18967), .A2(n19058), .ZN(n18725) );
  AOI22_X1 U20774 ( .A1(n18978), .A2(n18725), .B1(n18726), .B2(n18711), .ZN(
        n19054) );
  AOI22_X1 U20775 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19054), .B1(
        n18722), .B2(n19053), .ZN(n18712) );
  OAI211_X1 U20776 ( .C1(n18721), .C2(n19058), .A(n18713), .B(n18712), .ZN(
        P3_U2891) );
  INV_X1 U20777 ( .A(n18716), .ZN(n18714) );
  NOR2_X1 U20778 ( .A1(n18715), .A2(n18714), .ZN(n19059) );
  AOI22_X1 U20779 ( .A1(n18728), .A2(n19069), .B1(n18723), .B2(n19059), .ZN(
        n18720) );
  AOI22_X1 U20780 ( .A1(n18978), .A2(n18718), .B1(n18717), .B2(n18716), .ZN(
        n19062) );
  AOI22_X1 U20781 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19062), .B1(
        n18722), .B2(n19061), .ZN(n18719) );
  OAI211_X1 U20782 ( .C1(n18967), .C2(n18721), .A(n18720), .B(n18719), .ZN(
        P3_U2883) );
  INV_X1 U20783 ( .A(n18722), .ZN(n18731) );
  AND2_X1 U20784 ( .A1(n21241), .A2(n18725), .ZN(n19067) );
  AOI22_X1 U20785 ( .A1(n18724), .A2(n19069), .B1(n18723), .B2(n19067), .ZN(
        n18730) );
  AOI22_X1 U20786 ( .A1(n18978), .A2(n18727), .B1(n18726), .B2(n18725), .ZN(
        n19072) );
  AOI22_X1 U20787 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19072), .B1(
        n18728), .B2(n18990), .ZN(n18729) );
  OAI211_X1 U20788 ( .C1(n18731), .C2(n19058), .A(n18730), .B(n18729), .ZN(
        P3_U2875) );
  INV_X1 U20789 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n18732) );
  INV_X1 U20790 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20674) );
  AOI22_X1 U20791 ( .A1(n18977), .A2(n18732), .B1(n20674), .B2(U215), .ZN(U257) );
  NAND2_X1 U20792 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18978), .ZN(n18764) );
  NAND2_X1 U20793 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18978), .ZN(n18770) );
  INV_X1 U20794 ( .A(n18770), .ZN(n18761) );
  NOR2_X2 U20795 ( .A1(n20674), .A2(n18979), .ZN(n18765) );
  AOI22_X1 U20796 ( .A1(n18990), .A2(n18761), .B1(n18980), .B2(n18765), .ZN(
        n18734) );
  NOR2_X2 U20797 ( .A1(n20656), .A2(n18981), .ZN(n18767) );
  AOI22_X1 U20798 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18982), .B1(
        n19060), .B2(n18767), .ZN(n18733) );
  OAI211_X1 U20799 ( .C1(n18896), .C2(n18764), .A(n18734), .B(n18733), .ZN(
        P3_U2994) );
  AOI22_X1 U20800 ( .A1(n18996), .A2(n18761), .B1(n18985), .B2(n18765), .ZN(
        n18736) );
  AOI22_X1 U20801 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18986), .B1(
        n19069), .B2(n18767), .ZN(n18735) );
  OAI211_X1 U20802 ( .C1(n18994), .C2(n18764), .A(n18736), .B(n18735), .ZN(
        P3_U2986) );
  AOI22_X1 U20803 ( .A1(n19002), .A2(n18761), .B1(n18989), .B2(n18765), .ZN(
        n18738) );
  AOI22_X1 U20804 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18991), .B1(
        n18990), .B2(n18767), .ZN(n18737) );
  OAI211_X1 U20805 ( .C1(n19000), .C2(n18764), .A(n18738), .B(n18737), .ZN(
        P3_U2978) );
  AOI22_X1 U20806 ( .A1(n19007), .A2(n18761), .B1(n18995), .B2(n18765), .ZN(
        n18740) );
  AOI22_X1 U20807 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18997), .B1(
        n18996), .B2(n18767), .ZN(n18739) );
  OAI211_X1 U20808 ( .C1(n18943), .C2(n18764), .A(n18740), .B(n18739), .ZN(
        P3_U2970) );
  AOI22_X1 U20809 ( .A1(n19013), .A2(n18761), .B1(n19001), .B2(n18765), .ZN(
        n18742) );
  AOI22_X1 U20810 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19003), .B1(
        n19002), .B2(n18767), .ZN(n18741) );
  OAI211_X1 U20811 ( .C1(n19011), .C2(n18764), .A(n18742), .B(n18741), .ZN(
        P3_U2962) );
  AOI22_X1 U20812 ( .A1(n19018), .A2(n18761), .B1(n19006), .B2(n18765), .ZN(
        n18744) );
  AOI22_X1 U20813 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19008), .B1(
        n19007), .B2(n18767), .ZN(n18743) );
  OAI211_X1 U20814 ( .C1(n18948), .C2(n18764), .A(n18744), .B(n18743), .ZN(
        P3_U2954) );
  AOI22_X1 U20815 ( .A1(n19024), .A2(n18761), .B1(n19012), .B2(n18765), .ZN(
        n18746) );
  AOI22_X1 U20816 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19014), .B1(
        n19013), .B2(n18767), .ZN(n18745) );
  OAI211_X1 U20817 ( .C1(n19022), .C2(n18764), .A(n18746), .B(n18745), .ZN(
        P3_U2946) );
  INV_X1 U20818 ( .A(n18764), .ZN(n18766) );
  AOI22_X1 U20819 ( .A1(n19036), .A2(n18766), .B1(n19017), .B2(n18765), .ZN(
        n18748) );
  AOI22_X1 U20820 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19019), .B1(
        n19018), .B2(n18767), .ZN(n18747) );
  OAI211_X1 U20821 ( .C1(n19022), .C2(n18770), .A(n18748), .B(n18747), .ZN(
        P3_U2938) );
  AOI22_X1 U20822 ( .A1(n19036), .A2(n18761), .B1(n19023), .B2(n18765), .ZN(
        n18750) );
  AOI22_X1 U20823 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19025), .B1(
        n19024), .B2(n18767), .ZN(n18749) );
  OAI211_X1 U20824 ( .C1(n19028), .C2(n18764), .A(n18750), .B(n18749), .ZN(
        P3_U2930) );
  AOI22_X1 U20825 ( .A1(n19047), .A2(n18766), .B1(n19029), .B2(n18765), .ZN(
        n18752) );
  AOI22_X1 U20826 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19031), .B1(
        n19030), .B2(n18767), .ZN(n18751) );
  OAI211_X1 U20827 ( .C1(n19028), .C2(n18770), .A(n18752), .B(n18751), .ZN(
        P3_U2922) );
  AOI22_X1 U20828 ( .A1(n19047), .A2(n18761), .B1(n19035), .B2(n18765), .ZN(
        n18754) );
  AOI22_X1 U20829 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19037), .B1(
        n19036), .B2(n18767), .ZN(n18753) );
  OAI211_X1 U20830 ( .C1(n19045), .C2(n18764), .A(n18754), .B(n18753), .ZN(
        P3_U2914) );
  AOI22_X1 U20831 ( .A1(n19061), .A2(n18766), .B1(n19040), .B2(n18765), .ZN(
        n18756) );
  AOI22_X1 U20832 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n18767), .ZN(n18755) );
  OAI211_X1 U20833 ( .C1(n19045), .C2(n18770), .A(n18756), .B(n18755), .ZN(
        P3_U2906) );
  INV_X1 U20834 ( .A(n19058), .ZN(n19071) );
  AOI22_X1 U20835 ( .A1(n19071), .A2(n18766), .B1(n19046), .B2(n18765), .ZN(
        n18758) );
  AOI22_X1 U20836 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n18767), .ZN(n18757) );
  OAI211_X1 U20837 ( .C1(n18964), .C2(n18770), .A(n18758), .B(n18757), .ZN(
        P3_U2898) );
  AOI22_X1 U20838 ( .A1(n19060), .A2(n18766), .B1(n19051), .B2(n18765), .ZN(
        n18760) );
  AOI22_X1 U20839 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n18767), .ZN(n18759) );
  OAI211_X1 U20840 ( .C1(n19058), .C2(n18770), .A(n18760), .B(n18759), .ZN(
        P3_U2890) );
  AOI22_X1 U20841 ( .A1(n19060), .A2(n18761), .B1(n19059), .B2(n18765), .ZN(
        n18763) );
  AOI22_X1 U20842 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19062), .B1(
        n19061), .B2(n18767), .ZN(n18762) );
  OAI211_X1 U20843 ( .C1(n19065), .C2(n18764), .A(n18763), .B(n18762), .ZN(
        P3_U2882) );
  AOI22_X1 U20844 ( .A1(n18990), .A2(n18766), .B1(n19067), .B2(n18765), .ZN(
        n18769) );
  AOI22_X1 U20845 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n18767), .ZN(n18768) );
  OAI211_X1 U20846 ( .C1(n19065), .C2(n18770), .A(n18769), .B(n18768), .ZN(
        P3_U2874) );
  INV_X1 U20847 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n18771) );
  INV_X1 U20848 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n20637) );
  AOI22_X1 U20849 ( .A1(n18977), .A2(n18771), .B1(n20637), .B2(U215), .ZN(U256) );
  OR2_X1 U20850 ( .A1(n18981), .A2(n18772), .ZN(n18809) );
  AND2_X1 U20851 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18978), .ZN(n18806) );
  NOR2_X2 U20852 ( .A1(n18979), .A2(n20637), .ZN(n18804) );
  AOI22_X1 U20853 ( .A1(n18996), .A2(n18806), .B1(n18980), .B2(n18804), .ZN(
        n18775) );
  NOR2_X2 U20854 ( .A1(n18773), .A2(n20657), .ZN(n18805) );
  AOI22_X1 U20855 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18982), .B1(
        n18990), .B2(n18805), .ZN(n18774) );
  OAI211_X1 U20856 ( .C1(n18967), .C2(n18809), .A(n18775), .B(n18774), .ZN(
        P3_U2993) );
  AOI22_X1 U20857 ( .A1(n19002), .A2(n18806), .B1(n18985), .B2(n18804), .ZN(
        n18777) );
  AOI22_X1 U20858 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18986), .B1(
        n18996), .B2(n18805), .ZN(n18776) );
  OAI211_X1 U20859 ( .C1(n19065), .C2(n18809), .A(n18777), .B(n18776), .ZN(
        P3_U2985) );
  AOI22_X1 U20860 ( .A1(n19007), .A2(n18806), .B1(n18989), .B2(n18804), .ZN(
        n18779) );
  AOI22_X1 U20861 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18991), .B1(
        n19002), .B2(n18805), .ZN(n18778) );
  OAI211_X1 U20862 ( .C1(n19076), .C2(n18809), .A(n18779), .B(n18778), .ZN(
        P3_U2977) );
  AOI22_X1 U20863 ( .A1(n19013), .A2(n18806), .B1(n18995), .B2(n18804), .ZN(
        n18781) );
  AOI22_X1 U20864 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18997), .B1(
        n19007), .B2(n18805), .ZN(n18780) );
  OAI211_X1 U20865 ( .C1(n18896), .C2(n18809), .A(n18781), .B(n18780), .ZN(
        P3_U2969) );
  AOI22_X1 U20866 ( .A1(n19018), .A2(n18806), .B1(n19001), .B2(n18804), .ZN(
        n18783) );
  AOI22_X1 U20867 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19003), .B1(
        n19013), .B2(n18805), .ZN(n18782) );
  OAI211_X1 U20868 ( .C1(n18994), .C2(n18809), .A(n18783), .B(n18782), .ZN(
        P3_U2961) );
  AOI22_X1 U20869 ( .A1(n19024), .A2(n18806), .B1(n19006), .B2(n18804), .ZN(
        n18785) );
  AOI22_X1 U20870 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19008), .B1(
        n19018), .B2(n18805), .ZN(n18784) );
  OAI211_X1 U20871 ( .C1(n19000), .C2(n18809), .A(n18785), .B(n18784), .ZN(
        P3_U2953) );
  AOI22_X1 U20872 ( .A1(n19024), .A2(n18805), .B1(n19012), .B2(n18804), .ZN(
        n18787) );
  AOI22_X1 U20873 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19014), .B1(
        n19030), .B2(n18806), .ZN(n18786) );
  OAI211_X1 U20874 ( .C1(n18943), .C2(n18809), .A(n18787), .B(n18786), .ZN(
        P3_U2945) );
  AOI22_X1 U20875 ( .A1(n19030), .A2(n18805), .B1(n19017), .B2(n18804), .ZN(
        n18789) );
  AOI22_X1 U20876 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19019), .B1(
        n19036), .B2(n18806), .ZN(n18788) );
  OAI211_X1 U20877 ( .C1(n19011), .C2(n18809), .A(n18789), .B(n18788), .ZN(
        P3_U2937) );
  AOI22_X1 U20878 ( .A1(n19041), .A2(n18806), .B1(n19023), .B2(n18804), .ZN(
        n18791) );
  AOI22_X1 U20879 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19025), .B1(
        n19036), .B2(n18805), .ZN(n18790) );
  OAI211_X1 U20880 ( .C1(n18948), .C2(n18809), .A(n18791), .B(n18790), .ZN(
        P3_U2929) );
  AOI22_X1 U20881 ( .A1(n19047), .A2(n18806), .B1(n19029), .B2(n18804), .ZN(
        n18793) );
  AOI22_X1 U20882 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19031), .B1(
        n19041), .B2(n18805), .ZN(n18792) );
  OAI211_X1 U20883 ( .C1(n19022), .C2(n18809), .A(n18793), .B(n18792), .ZN(
        P3_U2921) );
  AOI22_X1 U20884 ( .A1(n19047), .A2(n18805), .B1(n19035), .B2(n18804), .ZN(
        n18795) );
  AOI22_X1 U20885 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19037), .B1(
        n19053), .B2(n18806), .ZN(n18794) );
  OAI211_X1 U20886 ( .C1(n18951), .C2(n18809), .A(n18795), .B(n18794), .ZN(
        P3_U2913) );
  AOI22_X1 U20887 ( .A1(n19061), .A2(n18806), .B1(n19040), .B2(n18804), .ZN(
        n18797) );
  AOI22_X1 U20888 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19042), .B1(
        n19053), .B2(n18805), .ZN(n18796) );
  OAI211_X1 U20889 ( .C1(n19028), .C2(n18809), .A(n18797), .B(n18796), .ZN(
        P3_U2905) );
  AOI22_X1 U20890 ( .A1(n19061), .A2(n18805), .B1(n19046), .B2(n18804), .ZN(
        n18799) );
  AOI22_X1 U20891 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19048), .B1(
        n19071), .B2(n18806), .ZN(n18798) );
  OAI211_X1 U20892 ( .C1(n19034), .C2(n18809), .A(n18799), .B(n18798), .ZN(
        P3_U2897) );
  AOI22_X1 U20893 ( .A1(n19060), .A2(n18806), .B1(n19051), .B2(n18804), .ZN(
        n18801) );
  AOI22_X1 U20894 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19054), .B1(
        n19071), .B2(n18805), .ZN(n18800) );
  OAI211_X1 U20895 ( .C1(n19045), .C2(n18809), .A(n18801), .B(n18800), .ZN(
        P3_U2889) );
  AOI22_X1 U20896 ( .A1(n19069), .A2(n18806), .B1(n19059), .B2(n18804), .ZN(
        n18803) );
  AOI22_X1 U20897 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19062), .B1(
        n19060), .B2(n18805), .ZN(n18802) );
  OAI211_X1 U20898 ( .C1(n18964), .C2(n18809), .A(n18803), .B(n18802), .ZN(
        P3_U2881) );
  AOI22_X1 U20899 ( .A1(n19069), .A2(n18805), .B1(n19067), .B2(n18804), .ZN(
        n18808) );
  AOI22_X1 U20900 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19072), .B1(
        n18990), .B2(n18806), .ZN(n18807) );
  OAI211_X1 U20901 ( .C1(n19058), .C2(n18809), .A(n18808), .B(n18807), .ZN(
        P3_U2873) );
  INV_X1 U20902 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n18810) );
  AOI22_X1 U20903 ( .A1(n18977), .A2(n18810), .B1(n20643), .B2(U215), .ZN(U255) );
  NAND2_X1 U20904 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18978), .ZN(n18833) );
  NAND2_X1 U20905 ( .A1(n18978), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18849) );
  INV_X1 U20906 ( .A(n18849), .ZN(n18830) );
  NOR2_X2 U20907 ( .A1(n18979), .A2(n20643), .ZN(n18844) );
  AOI22_X1 U20908 ( .A1(n18990), .A2(n18830), .B1(n18980), .B2(n18844), .ZN(
        n18813) );
  NOR2_X2 U20909 ( .A1(n18811), .A2(n18981), .ZN(n18846) );
  AOI22_X1 U20910 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18982), .B1(
        n19060), .B2(n18846), .ZN(n18812) );
  OAI211_X1 U20911 ( .C1(n18896), .C2(n18833), .A(n18813), .B(n18812), .ZN(
        P3_U2992) );
  AOI22_X1 U20912 ( .A1(n18996), .A2(n18830), .B1(n18985), .B2(n18844), .ZN(
        n18815) );
  AOI22_X1 U20913 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18986), .B1(
        n19069), .B2(n18846), .ZN(n18814) );
  OAI211_X1 U20914 ( .C1(n18994), .C2(n18833), .A(n18815), .B(n18814), .ZN(
        P3_U2984) );
  AOI22_X1 U20915 ( .A1(n19002), .A2(n18830), .B1(n18989), .B2(n18844), .ZN(
        n18817) );
  AOI22_X1 U20916 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18991), .B1(
        n18990), .B2(n18846), .ZN(n18816) );
  OAI211_X1 U20917 ( .C1(n19000), .C2(n18833), .A(n18817), .B(n18816), .ZN(
        P3_U2976) );
  AOI22_X1 U20918 ( .A1(n19007), .A2(n18830), .B1(n18995), .B2(n18844), .ZN(
        n18819) );
  AOI22_X1 U20919 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18997), .B1(
        n18996), .B2(n18846), .ZN(n18818) );
  OAI211_X1 U20920 ( .C1(n18943), .C2(n18833), .A(n18819), .B(n18818), .ZN(
        P3_U2968) );
  AOI22_X1 U20921 ( .A1(n19013), .A2(n18830), .B1(n19001), .B2(n18844), .ZN(
        n18821) );
  AOI22_X1 U20922 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19003), .B1(
        n19002), .B2(n18846), .ZN(n18820) );
  OAI211_X1 U20923 ( .C1(n19011), .C2(n18833), .A(n18821), .B(n18820), .ZN(
        P3_U2960) );
  INV_X1 U20924 ( .A(n18833), .ZN(n18845) );
  AOI22_X1 U20925 ( .A1(n19024), .A2(n18845), .B1(n19006), .B2(n18844), .ZN(
        n18823) );
  AOI22_X1 U20926 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19008), .B1(
        n19007), .B2(n18846), .ZN(n18822) );
  OAI211_X1 U20927 ( .C1(n19011), .C2(n18849), .A(n18823), .B(n18822), .ZN(
        P3_U2952) );
  AOI22_X1 U20928 ( .A1(n19030), .A2(n18845), .B1(n19012), .B2(n18844), .ZN(
        n18825) );
  AOI22_X1 U20929 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19014), .B1(
        n19013), .B2(n18846), .ZN(n18824) );
  OAI211_X1 U20930 ( .C1(n18948), .C2(n18849), .A(n18825), .B(n18824), .ZN(
        P3_U2944) );
  AOI22_X1 U20931 ( .A1(n19030), .A2(n18830), .B1(n19017), .B2(n18844), .ZN(
        n18827) );
  AOI22_X1 U20932 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19019), .B1(
        n19018), .B2(n18846), .ZN(n18826) );
  OAI211_X1 U20933 ( .C1(n18951), .C2(n18833), .A(n18827), .B(n18826), .ZN(
        P3_U2936) );
  AOI22_X1 U20934 ( .A1(n19036), .A2(n18830), .B1(n19023), .B2(n18844), .ZN(
        n18829) );
  AOI22_X1 U20935 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19025), .B1(
        n19024), .B2(n18846), .ZN(n18828) );
  OAI211_X1 U20936 ( .C1(n19028), .C2(n18833), .A(n18829), .B(n18828), .ZN(
        P3_U2928) );
  AOI22_X1 U20937 ( .A1(n19041), .A2(n18830), .B1(n19029), .B2(n18844), .ZN(
        n18832) );
  AOI22_X1 U20938 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19031), .B1(
        n19030), .B2(n18846), .ZN(n18831) );
  OAI211_X1 U20939 ( .C1(n19034), .C2(n18833), .A(n18832), .B(n18831), .ZN(
        P3_U2920) );
  AOI22_X1 U20940 ( .A1(n19053), .A2(n18845), .B1(n19035), .B2(n18844), .ZN(
        n18835) );
  AOI22_X1 U20941 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19037), .B1(
        n19036), .B2(n18846), .ZN(n18834) );
  OAI211_X1 U20942 ( .C1(n19034), .C2(n18849), .A(n18835), .B(n18834), .ZN(
        P3_U2912) );
  AOI22_X1 U20943 ( .A1(n19061), .A2(n18845), .B1(n19040), .B2(n18844), .ZN(
        n18837) );
  AOI22_X1 U20944 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n18846), .ZN(n18836) );
  OAI211_X1 U20945 ( .C1(n19045), .C2(n18849), .A(n18837), .B(n18836), .ZN(
        P3_U2904) );
  AOI22_X1 U20946 ( .A1(n19071), .A2(n18845), .B1(n19046), .B2(n18844), .ZN(
        n18839) );
  AOI22_X1 U20947 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n18846), .ZN(n18838) );
  OAI211_X1 U20948 ( .C1(n18964), .C2(n18849), .A(n18839), .B(n18838), .ZN(
        P3_U2896) );
  AOI22_X1 U20949 ( .A1(n19060), .A2(n18845), .B1(n19051), .B2(n18844), .ZN(
        n18841) );
  AOI22_X1 U20950 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n18846), .ZN(n18840) );
  OAI211_X1 U20951 ( .C1(n19058), .C2(n18849), .A(n18841), .B(n18840), .ZN(
        P3_U2888) );
  AOI22_X1 U20952 ( .A1(n19069), .A2(n18845), .B1(n19059), .B2(n18844), .ZN(
        n18843) );
  AOI22_X1 U20953 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19062), .B1(
        n19061), .B2(n18846), .ZN(n18842) );
  OAI211_X1 U20954 ( .C1(n18967), .C2(n18849), .A(n18843), .B(n18842), .ZN(
        P3_U2880) );
  AOI22_X1 U20955 ( .A1(n18990), .A2(n18845), .B1(n19067), .B2(n18844), .ZN(
        n18848) );
  AOI22_X1 U20956 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n18846), .ZN(n18847) );
  OAI211_X1 U20957 ( .C1(n19065), .C2(n18849), .A(n18848), .B(n18847), .ZN(
        P3_U2872) );
  OAI22_X1 U20958 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n18977), .ZN(n18850) );
  INV_X1 U20959 ( .A(n18850), .ZN(U254) );
  NAND2_X1 U20960 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18978), .ZN(n18883) );
  NAND2_X1 U20961 ( .A1(n18978), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18889) );
  INV_X1 U20962 ( .A(n18889), .ZN(n18880) );
  AND2_X1 U20963 ( .A1(n18932), .A2(BUF2_REG_3__SCAN_IN), .ZN(n18884) );
  AOI22_X1 U20964 ( .A1(n18990), .A2(n18880), .B1(n18980), .B2(n18884), .ZN(
        n18853) );
  NOR2_X2 U20965 ( .A1(n18851), .A2(n18981), .ZN(n18886) );
  AOI22_X1 U20966 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18982), .B1(
        n19060), .B2(n18886), .ZN(n18852) );
  OAI211_X1 U20967 ( .C1(n18896), .C2(n18883), .A(n18853), .B(n18852), .ZN(
        P3_U2991) );
  AOI22_X1 U20968 ( .A1(n18996), .A2(n18880), .B1(n18985), .B2(n18884), .ZN(
        n18855) );
  AOI22_X1 U20969 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18986), .B1(
        n19069), .B2(n18886), .ZN(n18854) );
  OAI211_X1 U20970 ( .C1(n18994), .C2(n18883), .A(n18855), .B(n18854), .ZN(
        P3_U2983) );
  AOI22_X1 U20971 ( .A1(n19002), .A2(n18880), .B1(n18989), .B2(n18884), .ZN(
        n18857) );
  AOI22_X1 U20972 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18991), .B1(
        n18990), .B2(n18886), .ZN(n18856) );
  OAI211_X1 U20973 ( .C1(n19000), .C2(n18883), .A(n18857), .B(n18856), .ZN(
        P3_U2975) );
  INV_X1 U20974 ( .A(n18883), .ZN(n18885) );
  AOI22_X1 U20975 ( .A1(n19013), .A2(n18885), .B1(n18995), .B2(n18884), .ZN(
        n18859) );
  AOI22_X1 U20976 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18997), .B1(
        n18996), .B2(n18886), .ZN(n18858) );
  OAI211_X1 U20977 ( .C1(n19000), .C2(n18889), .A(n18859), .B(n18858), .ZN(
        P3_U2967) );
  AOI22_X1 U20978 ( .A1(n19018), .A2(n18885), .B1(n19001), .B2(n18884), .ZN(
        n18861) );
  AOI22_X1 U20979 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19003), .B1(
        n19002), .B2(n18886), .ZN(n18860) );
  OAI211_X1 U20980 ( .C1(n18943), .C2(n18889), .A(n18861), .B(n18860), .ZN(
        P3_U2959) );
  AOI22_X1 U20981 ( .A1(n19018), .A2(n18880), .B1(n19006), .B2(n18884), .ZN(
        n18863) );
  AOI22_X1 U20982 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19008), .B1(
        n19007), .B2(n18886), .ZN(n18862) );
  OAI211_X1 U20983 ( .C1(n18948), .C2(n18883), .A(n18863), .B(n18862), .ZN(
        P3_U2951) );
  AOI22_X1 U20984 ( .A1(n19024), .A2(n18880), .B1(n19012), .B2(n18884), .ZN(
        n18865) );
  AOI22_X1 U20985 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19014), .B1(
        n19013), .B2(n18886), .ZN(n18864) );
  OAI211_X1 U20986 ( .C1(n19022), .C2(n18883), .A(n18865), .B(n18864), .ZN(
        P3_U2943) );
  AOI22_X1 U20987 ( .A1(n19030), .A2(n18880), .B1(n19017), .B2(n18884), .ZN(
        n18867) );
  AOI22_X1 U20988 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19019), .B1(
        n19018), .B2(n18886), .ZN(n18866) );
  OAI211_X1 U20989 ( .C1(n18951), .C2(n18883), .A(n18867), .B(n18866), .ZN(
        P3_U2935) );
  AOI22_X1 U20990 ( .A1(n19036), .A2(n18880), .B1(n19023), .B2(n18884), .ZN(
        n18869) );
  AOI22_X1 U20991 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19025), .B1(
        n19024), .B2(n18886), .ZN(n18868) );
  OAI211_X1 U20992 ( .C1(n19028), .C2(n18883), .A(n18869), .B(n18868), .ZN(
        P3_U2927) );
  AOI22_X1 U20993 ( .A1(n19041), .A2(n18880), .B1(n19029), .B2(n18884), .ZN(
        n18871) );
  AOI22_X1 U20994 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19031), .B1(
        n19030), .B2(n18886), .ZN(n18870) );
  OAI211_X1 U20995 ( .C1(n19034), .C2(n18883), .A(n18871), .B(n18870), .ZN(
        P3_U2919) );
  AOI22_X1 U20996 ( .A1(n19053), .A2(n18885), .B1(n19035), .B2(n18884), .ZN(
        n18873) );
  AOI22_X1 U20997 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19037), .B1(
        n19036), .B2(n18886), .ZN(n18872) );
  OAI211_X1 U20998 ( .C1(n19034), .C2(n18889), .A(n18873), .B(n18872), .ZN(
        P3_U2911) );
  AOI22_X1 U20999 ( .A1(n19053), .A2(n18880), .B1(n19040), .B2(n18884), .ZN(
        n18875) );
  AOI22_X1 U21000 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n18886), .ZN(n18874) );
  OAI211_X1 U21001 ( .C1(n18964), .C2(n18883), .A(n18875), .B(n18874), .ZN(
        P3_U2903) );
  AOI22_X1 U21002 ( .A1(n19071), .A2(n18885), .B1(n19046), .B2(n18884), .ZN(
        n18877) );
  AOI22_X1 U21003 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n18886), .ZN(n18876) );
  OAI211_X1 U21004 ( .C1(n18964), .C2(n18889), .A(n18877), .B(n18876), .ZN(
        P3_U2895) );
  AOI22_X1 U21005 ( .A1(n19060), .A2(n18885), .B1(n19051), .B2(n18884), .ZN(
        n18879) );
  AOI22_X1 U21006 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n18886), .ZN(n18878) );
  OAI211_X1 U21007 ( .C1(n19058), .C2(n18889), .A(n18879), .B(n18878), .ZN(
        P3_U2887) );
  AOI22_X1 U21008 ( .A1(n19060), .A2(n18880), .B1(n19059), .B2(n18884), .ZN(
        n18882) );
  AOI22_X1 U21009 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19062), .B1(
        n19061), .B2(n18886), .ZN(n18881) );
  OAI211_X1 U21010 ( .C1(n19065), .C2(n18883), .A(n18882), .B(n18881), .ZN(
        P3_U2879) );
  AOI22_X1 U21011 ( .A1(n18990), .A2(n18885), .B1(n19067), .B2(n18884), .ZN(
        n18888) );
  AOI22_X1 U21012 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n18886), .ZN(n18887) );
  OAI211_X1 U21013 ( .C1(n19065), .C2(n18889), .A(n18888), .B(n18887), .ZN(
        P3_U2871) );
  INV_X1 U21014 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n18890) );
  AOI22_X1 U21015 ( .A1(n18977), .A2(n18890), .B1(n20130), .B2(U215), .ZN(U253) );
  NAND2_X1 U21016 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18978), .ZN(n18930) );
  NAND2_X1 U21017 ( .A1(n18978), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18912) );
  INV_X1 U21018 ( .A(n18912), .ZN(n18926) );
  NOR2_X2 U21019 ( .A1(n18979), .A2(n20130), .ZN(n18925) );
  AOI22_X1 U21020 ( .A1(n18990), .A2(n18926), .B1(n18980), .B2(n18925), .ZN(
        n18893) );
  NOR2_X2 U21021 ( .A1(n18891), .A2(n18981), .ZN(n18927) );
  AOI22_X1 U21022 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18982), .B1(
        n19060), .B2(n18927), .ZN(n18892) );
  OAI211_X1 U21023 ( .C1(n18896), .C2(n18930), .A(n18893), .B(n18892), .ZN(
        P3_U2990) );
  INV_X1 U21024 ( .A(n18930), .ZN(n18909) );
  AOI22_X1 U21025 ( .A1(n19002), .A2(n18909), .B1(n18985), .B2(n18925), .ZN(
        n18895) );
  AOI22_X1 U21026 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18986), .B1(
        n19069), .B2(n18927), .ZN(n18894) );
  OAI211_X1 U21027 ( .C1(n18896), .C2(n18912), .A(n18895), .B(n18894), .ZN(
        P3_U2982) );
  AOI22_X1 U21028 ( .A1(n19002), .A2(n18926), .B1(n18989), .B2(n18925), .ZN(
        n18898) );
  AOI22_X1 U21029 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18991), .B1(
        n18990), .B2(n18927), .ZN(n18897) );
  OAI211_X1 U21030 ( .C1(n19000), .C2(n18930), .A(n18898), .B(n18897), .ZN(
        P3_U2974) );
  AOI22_X1 U21031 ( .A1(n19007), .A2(n18926), .B1(n18995), .B2(n18925), .ZN(
        n18900) );
  AOI22_X1 U21032 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18997), .B1(
        n18996), .B2(n18927), .ZN(n18899) );
  OAI211_X1 U21033 ( .C1(n18943), .C2(n18930), .A(n18900), .B(n18899), .ZN(
        P3_U2966) );
  AOI22_X1 U21034 ( .A1(n19018), .A2(n18909), .B1(n19001), .B2(n18925), .ZN(
        n18902) );
  AOI22_X1 U21035 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19003), .B1(
        n19002), .B2(n18927), .ZN(n18901) );
  OAI211_X1 U21036 ( .C1(n18943), .C2(n18912), .A(n18902), .B(n18901), .ZN(
        P3_U2958) );
  AOI22_X1 U21037 ( .A1(n19018), .A2(n18926), .B1(n19006), .B2(n18925), .ZN(
        n18904) );
  AOI22_X1 U21038 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19008), .B1(
        n19007), .B2(n18927), .ZN(n18903) );
  OAI211_X1 U21039 ( .C1(n18948), .C2(n18930), .A(n18904), .B(n18903), .ZN(
        P3_U2950) );
  AOI22_X1 U21040 ( .A1(n19030), .A2(n18909), .B1(n19012), .B2(n18925), .ZN(
        n18906) );
  AOI22_X1 U21041 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19014), .B1(
        n19013), .B2(n18927), .ZN(n18905) );
  OAI211_X1 U21042 ( .C1(n18948), .C2(n18912), .A(n18906), .B(n18905), .ZN(
        P3_U2942) );
  AOI22_X1 U21043 ( .A1(n19036), .A2(n18909), .B1(n19017), .B2(n18925), .ZN(
        n18908) );
  AOI22_X1 U21044 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19019), .B1(
        n19018), .B2(n18927), .ZN(n18907) );
  OAI211_X1 U21045 ( .C1(n19022), .C2(n18912), .A(n18908), .B(n18907), .ZN(
        P3_U2934) );
  AOI22_X1 U21046 ( .A1(n19041), .A2(n18909), .B1(n19023), .B2(n18925), .ZN(
        n18911) );
  AOI22_X1 U21047 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19025), .B1(
        n19024), .B2(n18927), .ZN(n18910) );
  OAI211_X1 U21048 ( .C1(n18951), .C2(n18912), .A(n18911), .B(n18910), .ZN(
        P3_U2926) );
  AOI22_X1 U21049 ( .A1(n19041), .A2(n18926), .B1(n19029), .B2(n18925), .ZN(
        n18914) );
  AOI22_X1 U21050 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19031), .B1(
        n19030), .B2(n18927), .ZN(n18913) );
  OAI211_X1 U21051 ( .C1(n19034), .C2(n18930), .A(n18914), .B(n18913), .ZN(
        P3_U2918) );
  AOI22_X1 U21052 ( .A1(n19047), .A2(n18926), .B1(n19035), .B2(n18925), .ZN(
        n18916) );
  AOI22_X1 U21053 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19037), .B1(
        n19036), .B2(n18927), .ZN(n18915) );
  OAI211_X1 U21054 ( .C1(n19045), .C2(n18930), .A(n18916), .B(n18915), .ZN(
        P3_U2910) );
  AOI22_X1 U21055 ( .A1(n19053), .A2(n18926), .B1(n19040), .B2(n18925), .ZN(
        n18918) );
  AOI22_X1 U21056 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n18927), .ZN(n18917) );
  OAI211_X1 U21057 ( .C1(n18964), .C2(n18930), .A(n18918), .B(n18917), .ZN(
        P3_U2902) );
  AOI22_X1 U21058 ( .A1(n19061), .A2(n18926), .B1(n19046), .B2(n18925), .ZN(
        n18920) );
  AOI22_X1 U21059 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n18927), .ZN(n18919) );
  OAI211_X1 U21060 ( .C1(n19058), .C2(n18930), .A(n18920), .B(n18919), .ZN(
        P3_U2894) );
  AOI22_X1 U21061 ( .A1(n19071), .A2(n18926), .B1(n19051), .B2(n18925), .ZN(
        n18922) );
  AOI22_X1 U21062 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n18927), .ZN(n18921) );
  OAI211_X1 U21063 ( .C1(n18967), .C2(n18930), .A(n18922), .B(n18921), .ZN(
        P3_U2886) );
  AOI22_X1 U21064 ( .A1(n19060), .A2(n18926), .B1(n19059), .B2(n18925), .ZN(
        n18924) );
  AOI22_X1 U21065 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19062), .B1(
        n19061), .B2(n18927), .ZN(n18923) );
  OAI211_X1 U21066 ( .C1(n19065), .C2(n18930), .A(n18924), .B(n18923), .ZN(
        P3_U2878) );
  AOI22_X1 U21067 ( .A1(n19069), .A2(n18926), .B1(n19067), .B2(n18925), .ZN(
        n18929) );
  AOI22_X1 U21068 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n18927), .ZN(n18928) );
  OAI211_X1 U21069 ( .C1(n19076), .C2(n18930), .A(n18929), .B(n18928), .ZN(
        P3_U2870) );
  OAI22_X1 U21070 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n18977), .ZN(n18931) );
  INV_X1 U21071 ( .A(n18931), .ZN(U252) );
  NAND2_X1 U21072 ( .A1(n18978), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18963) );
  NAND2_X1 U21073 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18978), .ZN(n18975) );
  INV_X1 U21074 ( .A(n18975), .ZN(n18960) );
  AND2_X1 U21075 ( .A1(n18932), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18970) );
  AOI22_X1 U21076 ( .A1(n18996), .A2(n18960), .B1(n18980), .B2(n18970), .ZN(
        n18934) );
  NOR2_X2 U21077 ( .A1(n20158), .A2(n18981), .ZN(n18972) );
  AOI22_X1 U21078 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18982), .B1(
        n19060), .B2(n18972), .ZN(n18933) );
  OAI211_X1 U21079 ( .C1(n19076), .C2(n18963), .A(n18934), .B(n18933), .ZN(
        P3_U2989) );
  INV_X1 U21080 ( .A(n18963), .ZN(n18971) );
  AOI22_X1 U21081 ( .A1(n18996), .A2(n18971), .B1(n18985), .B2(n18970), .ZN(
        n18936) );
  AOI22_X1 U21082 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18986), .B1(
        n19069), .B2(n18972), .ZN(n18935) );
  OAI211_X1 U21083 ( .C1(n18994), .C2(n18975), .A(n18936), .B(n18935), .ZN(
        P3_U2981) );
  AOI22_X1 U21084 ( .A1(n19002), .A2(n18971), .B1(n18989), .B2(n18970), .ZN(
        n18938) );
  AOI22_X1 U21085 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18991), .B1(
        n18990), .B2(n18972), .ZN(n18937) );
  OAI211_X1 U21086 ( .C1(n19000), .C2(n18975), .A(n18938), .B(n18937), .ZN(
        P3_U2973) );
  AOI22_X1 U21087 ( .A1(n19013), .A2(n18960), .B1(n18995), .B2(n18970), .ZN(
        n18940) );
  AOI22_X1 U21088 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18997), .B1(
        n18996), .B2(n18972), .ZN(n18939) );
  OAI211_X1 U21089 ( .C1(n19000), .C2(n18963), .A(n18940), .B(n18939), .ZN(
        P3_U2965) );
  AOI22_X1 U21090 ( .A1(n19018), .A2(n18960), .B1(n19001), .B2(n18970), .ZN(
        n18942) );
  AOI22_X1 U21091 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19003), .B1(
        n19002), .B2(n18972), .ZN(n18941) );
  OAI211_X1 U21092 ( .C1(n18943), .C2(n18963), .A(n18942), .B(n18941), .ZN(
        P3_U2957) );
  AOI22_X1 U21093 ( .A1(n19024), .A2(n18960), .B1(n19006), .B2(n18970), .ZN(
        n18945) );
  AOI22_X1 U21094 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19008), .B1(
        n19007), .B2(n18972), .ZN(n18944) );
  OAI211_X1 U21095 ( .C1(n19011), .C2(n18963), .A(n18945), .B(n18944), .ZN(
        P3_U2949) );
  AOI22_X1 U21096 ( .A1(n19030), .A2(n18960), .B1(n19012), .B2(n18970), .ZN(
        n18947) );
  AOI22_X1 U21097 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19014), .B1(
        n19013), .B2(n18972), .ZN(n18946) );
  OAI211_X1 U21098 ( .C1(n18948), .C2(n18963), .A(n18947), .B(n18946), .ZN(
        P3_U2941) );
  AOI22_X1 U21099 ( .A1(n19030), .A2(n18971), .B1(n19017), .B2(n18970), .ZN(
        n18950) );
  AOI22_X1 U21100 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19019), .B1(
        n19018), .B2(n18972), .ZN(n18949) );
  OAI211_X1 U21101 ( .C1(n18951), .C2(n18975), .A(n18950), .B(n18949), .ZN(
        P3_U2933) );
  AOI22_X1 U21102 ( .A1(n19036), .A2(n18971), .B1(n19023), .B2(n18970), .ZN(
        n18953) );
  AOI22_X1 U21103 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19025), .B1(
        n19024), .B2(n18972), .ZN(n18952) );
  OAI211_X1 U21104 ( .C1(n19028), .C2(n18975), .A(n18953), .B(n18952), .ZN(
        P3_U2925) );
  AOI22_X1 U21105 ( .A1(n19041), .A2(n18971), .B1(n19029), .B2(n18970), .ZN(
        n18955) );
  AOI22_X1 U21106 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19031), .B1(
        n19030), .B2(n18972), .ZN(n18954) );
  OAI211_X1 U21107 ( .C1(n19034), .C2(n18975), .A(n18955), .B(n18954), .ZN(
        P3_U2917) );
  AOI22_X1 U21108 ( .A1(n19053), .A2(n18960), .B1(n19035), .B2(n18970), .ZN(
        n18957) );
  AOI22_X1 U21109 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19037), .B1(
        n19036), .B2(n18972), .ZN(n18956) );
  OAI211_X1 U21110 ( .C1(n19034), .C2(n18963), .A(n18957), .B(n18956), .ZN(
        P3_U2909) );
  AOI22_X1 U21111 ( .A1(n19053), .A2(n18971), .B1(n19040), .B2(n18970), .ZN(
        n18959) );
  AOI22_X1 U21112 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n18972), .ZN(n18958) );
  OAI211_X1 U21113 ( .C1(n18964), .C2(n18975), .A(n18959), .B(n18958), .ZN(
        P3_U2901) );
  AOI22_X1 U21114 ( .A1(n19071), .A2(n18960), .B1(n19046), .B2(n18970), .ZN(
        n18962) );
  AOI22_X1 U21115 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n18972), .ZN(n18961) );
  OAI211_X1 U21116 ( .C1(n18964), .C2(n18963), .A(n18962), .B(n18961), .ZN(
        P3_U2893) );
  AOI22_X1 U21117 ( .A1(n19071), .A2(n18971), .B1(n19051), .B2(n18970), .ZN(
        n18966) );
  AOI22_X1 U21118 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n18972), .ZN(n18965) );
  OAI211_X1 U21119 ( .C1(n18967), .C2(n18975), .A(n18966), .B(n18965), .ZN(
        P3_U2885) );
  AOI22_X1 U21120 ( .A1(n19060), .A2(n18971), .B1(n19059), .B2(n18970), .ZN(
        n18969) );
  AOI22_X1 U21121 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19062), .B1(
        n19061), .B2(n18972), .ZN(n18968) );
  OAI211_X1 U21122 ( .C1(n19065), .C2(n18975), .A(n18969), .B(n18968), .ZN(
        P3_U2877) );
  AOI22_X1 U21123 ( .A1(n19069), .A2(n18971), .B1(n19067), .B2(n18970), .ZN(
        n18974) );
  AOI22_X1 U21124 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n18972), .ZN(n18973) );
  OAI211_X1 U21125 ( .C1(n19076), .C2(n18975), .A(n18974), .B(n18973), .ZN(
        P3_U2869) );
  INV_X1 U21126 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n18976) );
  AOI22_X1 U21127 ( .A1(n18977), .A2(n18976), .B1(n20747), .B2(U215), .ZN(U251) );
  NAND2_X1 U21128 ( .A1(n18978), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19057) );
  NAND2_X1 U21129 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18978), .ZN(n19075) );
  INV_X1 U21130 ( .A(n19075), .ZN(n19052) );
  NOR2_X2 U21131 ( .A1(n18979), .A2(n20747), .ZN(n19066) );
  AOI22_X1 U21132 ( .A1(n18996), .A2(n19052), .B1(n18980), .B2(n19066), .ZN(
        n18984) );
  NOR2_X2 U21133 ( .A1(n20156), .A2(n18981), .ZN(n19070) );
  AOI22_X1 U21134 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18982), .B1(
        n19060), .B2(n19070), .ZN(n18983) );
  OAI211_X1 U21135 ( .C1(n19076), .C2(n19057), .A(n18984), .B(n18983), .ZN(
        P3_U2988) );
  INV_X1 U21136 ( .A(n19057), .ZN(n19068) );
  AOI22_X1 U21137 ( .A1(n18996), .A2(n19068), .B1(n18985), .B2(n19066), .ZN(
        n18988) );
  AOI22_X1 U21138 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18986), .B1(
        n19069), .B2(n19070), .ZN(n18987) );
  OAI211_X1 U21139 ( .C1(n18994), .C2(n19075), .A(n18988), .B(n18987), .ZN(
        P3_U2980) );
  AOI22_X1 U21140 ( .A1(n19007), .A2(n19052), .B1(n18989), .B2(n19066), .ZN(
        n18993) );
  AOI22_X1 U21141 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18991), .B1(
        n18990), .B2(n19070), .ZN(n18992) );
  OAI211_X1 U21142 ( .C1(n18994), .C2(n19057), .A(n18993), .B(n18992), .ZN(
        P3_U2972) );
  AOI22_X1 U21143 ( .A1(n19013), .A2(n19052), .B1(n18995), .B2(n19066), .ZN(
        n18999) );
  AOI22_X1 U21144 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18997), .B1(
        n18996), .B2(n19070), .ZN(n18998) );
  OAI211_X1 U21145 ( .C1(n19000), .C2(n19057), .A(n18999), .B(n18998), .ZN(
        P3_U2964) );
  AOI22_X1 U21146 ( .A1(n19013), .A2(n19068), .B1(n19001), .B2(n19066), .ZN(
        n19005) );
  AOI22_X1 U21147 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19003), .B1(
        n19002), .B2(n19070), .ZN(n19004) );
  OAI211_X1 U21148 ( .C1(n19011), .C2(n19075), .A(n19005), .B(n19004), .ZN(
        P3_U2956) );
  AOI22_X1 U21149 ( .A1(n19024), .A2(n19052), .B1(n19006), .B2(n19066), .ZN(
        n19010) );
  AOI22_X1 U21150 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19008), .B1(
        n19007), .B2(n19070), .ZN(n19009) );
  OAI211_X1 U21151 ( .C1(n19011), .C2(n19057), .A(n19010), .B(n19009), .ZN(
        P3_U2948) );
  AOI22_X1 U21152 ( .A1(n19024), .A2(n19068), .B1(n19012), .B2(n19066), .ZN(
        n19016) );
  AOI22_X1 U21153 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19014), .B1(
        n19013), .B2(n19070), .ZN(n19015) );
  OAI211_X1 U21154 ( .C1(n19022), .C2(n19075), .A(n19016), .B(n19015), .ZN(
        P3_U2940) );
  AOI22_X1 U21155 ( .A1(n19036), .A2(n19052), .B1(n19017), .B2(n19066), .ZN(
        n19021) );
  AOI22_X1 U21156 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19019), .B1(
        n19018), .B2(n19070), .ZN(n19020) );
  OAI211_X1 U21157 ( .C1(n19022), .C2(n19057), .A(n19021), .B(n19020), .ZN(
        P3_U2932) );
  AOI22_X1 U21158 ( .A1(n19036), .A2(n19068), .B1(n19023), .B2(n19066), .ZN(
        n19027) );
  AOI22_X1 U21159 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19025), .B1(
        n19024), .B2(n19070), .ZN(n19026) );
  OAI211_X1 U21160 ( .C1(n19028), .C2(n19075), .A(n19027), .B(n19026), .ZN(
        P3_U2924) );
  AOI22_X1 U21161 ( .A1(n19041), .A2(n19068), .B1(n19029), .B2(n19066), .ZN(
        n19033) );
  AOI22_X1 U21162 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19031), .B1(
        n19030), .B2(n19070), .ZN(n19032) );
  OAI211_X1 U21163 ( .C1(n19034), .C2(n19075), .A(n19033), .B(n19032), .ZN(
        P3_U2916) );
  AOI22_X1 U21164 ( .A1(n19047), .A2(n19068), .B1(n19035), .B2(n19066), .ZN(
        n19039) );
  AOI22_X1 U21165 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19037), .B1(
        n19036), .B2(n19070), .ZN(n19038) );
  OAI211_X1 U21166 ( .C1(n19045), .C2(n19075), .A(n19039), .B(n19038), .ZN(
        P3_U2908) );
  AOI22_X1 U21167 ( .A1(n19061), .A2(n19052), .B1(n19040), .B2(n19066), .ZN(
        n19044) );
  AOI22_X1 U21168 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19042), .B1(
        n19041), .B2(n19070), .ZN(n19043) );
  OAI211_X1 U21169 ( .C1(n19045), .C2(n19057), .A(n19044), .B(n19043), .ZN(
        P3_U2900) );
  AOI22_X1 U21170 ( .A1(n19061), .A2(n19068), .B1(n19046), .B2(n19066), .ZN(
        n19050) );
  AOI22_X1 U21171 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19048), .B1(
        n19047), .B2(n19070), .ZN(n19049) );
  OAI211_X1 U21172 ( .C1(n19058), .C2(n19075), .A(n19050), .B(n19049), .ZN(
        P3_U2892) );
  AOI22_X1 U21173 ( .A1(n19060), .A2(n19052), .B1(n19051), .B2(n19066), .ZN(
        n19056) );
  AOI22_X1 U21174 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19054), .B1(
        n19053), .B2(n19070), .ZN(n19055) );
  OAI211_X1 U21175 ( .C1(n19058), .C2(n19057), .A(n19056), .B(n19055), .ZN(
        P3_U2884) );
  AOI22_X1 U21176 ( .A1(n19060), .A2(n19068), .B1(n19059), .B2(n19066), .ZN(
        n19064) );
  AOI22_X1 U21177 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19062), .B1(
        n19061), .B2(n19070), .ZN(n19063) );
  OAI211_X1 U21178 ( .C1(n19065), .C2(n19075), .A(n19064), .B(n19063), .ZN(
        P3_U2876) );
  AOI22_X1 U21179 ( .A1(n19069), .A2(n19068), .B1(n19067), .B2(n19066), .ZN(
        n19074) );
  AOI22_X1 U21180 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19072), .B1(
        n19071), .B2(n19070), .ZN(n19073) );
  OAI211_X1 U21181 ( .C1(n19076), .C2(n19075), .A(n19074), .B(n19073), .ZN(
        P3_U2868) );
  AOI22_X1 U21182 ( .A1(n19630), .A2(BUF2_REG_31__SCAN_IN), .B1(n19633), .B2(
        n18499), .ZN(n19078) );
  AOI22_X1 U21183 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19627), .B1(n19631), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19077) );
  NAND2_X1 U21184 ( .A1(n19078), .A2(n19077), .ZN(P2_U2888) );
  OAI222_X1 U21185 ( .A1(n19081), .A2(n19378), .B1(n19080), .B2(n19531), .C1(
        n19079), .C2(n19583), .ZN(P2_U2904) );
  INV_X1 U21186 ( .A(n19082), .ZN(n19085) );
  AOI22_X1 U21187 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19627), .B1(n19083), 
        .B2(n19524), .ZN(n19084) );
  OAI21_X1 U21188 ( .B1(n19378), .B2(n19085), .A(n19084), .ZN(P2_U2905) );
  INV_X1 U21189 ( .A(n19086), .ZN(n19089) );
  OAI222_X1 U21190 ( .A1(n19089), .A2(n19378), .B1(n19088), .B2(n19531), .C1(
        n19583), .C2(n19087), .ZN(P2_U2906) );
  AOI22_X1 U21191 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19627), .B1(n19090), 
        .B2(n19524), .ZN(n19091) );
  OAI21_X1 U21192 ( .B1(n19378), .B2(n19092), .A(n19091), .ZN(P2_U2907) );
  OAI222_X1 U21193 ( .A1(n19095), .A2(n19378), .B1(n19094), .B2(n19531), .C1(
        n19583), .C2(n19093), .ZN(P2_U2908) );
  OAI222_X1 U21194 ( .A1(n19098), .A2(n19378), .B1(n19097), .B2(n19531), .C1(
        n19583), .C2(n19096), .ZN(P2_U2909) );
  OAI222_X1 U21195 ( .A1(n19101), .A2(n19378), .B1(n19100), .B2(n19531), .C1(
        n19583), .C2(n19099), .ZN(P2_U2910) );
  INV_X1 U21196 ( .A(n19102), .ZN(n19105) );
  OAI222_X1 U21197 ( .A1(n19105), .A2(n19378), .B1(n19104), .B2(n19531), .C1(
        n19583), .C2(n19103), .ZN(P2_U2911) );
  OAI222_X1 U21198 ( .A1(n19107), .A2(n19378), .B1(n19106), .B2(n19531), .C1(
        n19583), .C2(n19113), .ZN(P2_U2912) );
  NOR3_X4 U21199 ( .A1(n13854), .A2(n19108), .A3(n19306), .ZN(n19645) );
  NOR3_X4 U21200 ( .A1(n19109), .A2(n13854), .A3(n19306), .ZN(n19646) );
  AOI22_X1 U21201 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19645), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19646), .ZN(n19301) );
  NAND3_X1 U21202 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19124) );
  INV_X1 U21203 ( .A(n19111), .ZN(n19643) );
  OAI21_X1 U21204 ( .B1(n19115), .B2(n19643), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19112) );
  OAI21_X1 U21205 ( .B1(n19124), .B2(n19290), .A(n19112), .ZN(n19644) );
  NOR2_X2 U21206 ( .A1(n11083), .A2(n19641), .ZN(n19312) );
  AOI22_X1 U21207 ( .A1(n19644), .A2(n19114), .B1(n19643), .B2(n19312), .ZN(
        n19122) );
  OAI21_X1 U21208 ( .B1(n19143), .B2(n19259), .A(n19124), .ZN(n19120) );
  INV_X1 U21209 ( .A(n19115), .ZN(n19118) );
  NOR2_X1 U21210 ( .A1(n19116), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19294) );
  INV_X1 U21211 ( .A(n19294), .ZN(n19307) );
  INV_X1 U21212 ( .A(n19306), .ZN(n19220) );
  AOI21_X1 U21213 ( .B1(n19643), .B2(n19281), .A(n19220), .ZN(n19117) );
  OAI21_X1 U21214 ( .B1(n19118), .B2(n19307), .A(n19117), .ZN(n19119) );
  NAND2_X1 U21215 ( .A1(n19120), .A2(n19119), .ZN(n19647) );
  AOI22_X1 U21216 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19646), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19645), .ZN(n19286) );
  AOI22_X1 U21217 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19647), .B1(
        n19745), .B2(n19317), .ZN(n19121) );
  OAI211_X1 U21218 ( .C1(n19301), .C2(n19650), .A(n19122), .B(n19121), .ZN(
        P2_U3175) );
  INV_X1 U21219 ( .A(n19221), .ZN(n19283) );
  NOR2_X1 U21220 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19124), .ZN(
        n19651) );
  AOI22_X1 U21221 ( .A1(n19317), .A2(n19652), .B1(n19312), .B2(n19651), .ZN(
        n19134) );
  OAI21_X1 U21222 ( .B1(n19221), .B2(n19254), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19278) );
  OR2_X1 U21223 ( .A1(n19143), .A2(n19278), .ZN(n19126) );
  NAND3_X1 U21224 ( .A1(n19260), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19149) );
  NOR2_X1 U21225 ( .A1(n19288), .A2(n19149), .ZN(n19658) );
  INV_X1 U21226 ( .A(n19658), .ZN(n19128) );
  AOI21_X1 U21227 ( .B1(n15026), .B2(n19294), .A(n19220), .ZN(n19127) );
  AOI21_X1 U21228 ( .B1(n19130), .B2(n19128), .A(n19127), .ZN(n19129) );
  AOI21_X1 U21229 ( .B1(n19651), .B2(n19281), .A(n19129), .ZN(n19654) );
  OAI21_X1 U21230 ( .B1(n19651), .B2(n19658), .A(n19130), .ZN(n19132) );
  OAI21_X1 U21231 ( .B1(n15026), .B2(n19651), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19131) );
  NAND2_X1 U21232 ( .A1(n19132), .A2(n19131), .ZN(n19653) );
  AOI22_X1 U21233 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19654), .B1(
        n19114), .B2(n19653), .ZN(n19133) );
  OAI211_X1 U21234 ( .C1(n19301), .C2(n19657), .A(n19134), .B(n19133), .ZN(
        P2_U3167) );
  NAND2_X1 U21235 ( .A1(n19142), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19292) );
  OAI21_X1 U21236 ( .B1(n19143), .B2(n19292), .A(n19149), .ZN(n19138) );
  NAND2_X1 U21237 ( .A1(n19139), .A2(n19294), .ZN(n19136) );
  OAI21_X1 U21238 ( .B1(n19304), .B2(n19658), .A(n19281), .ZN(n19135) );
  NAND2_X1 U21239 ( .A1(n19136), .A2(n19135), .ZN(n19137) );
  INV_X1 U21240 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n19146) );
  OAI21_X1 U21241 ( .B1(n19139), .B2(n19658), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19140) );
  OAI21_X1 U21242 ( .B1(n19149), .B2(n19290), .A(n19140), .ZN(n19659) );
  AOI22_X1 U21243 ( .A1(n19659), .A2(n19114), .B1(n19312), .B2(n19658), .ZN(
        n19145) );
  NOR2_X2 U21244 ( .A1(n19287), .A2(n19143), .ZN(n19667) );
  INV_X1 U21245 ( .A(n19301), .ZN(n19313) );
  AOI22_X1 U21246 ( .A1(n19660), .A2(n19317), .B1(n19667), .B2(n19313), .ZN(
        n19144) );
  OAI211_X1 U21247 ( .C1(n19435), .C2(n19146), .A(n19145), .B(n19144), .ZN(
        P2_U3159) );
  NAND2_X1 U21248 ( .A1(n19148), .A2(n19217), .ZN(n19243) );
  NOR2_X1 U21249 ( .A1(n19255), .A2(n19243), .ZN(n19156) );
  INV_X1 U21250 ( .A(n19156), .ZN(n19152) );
  NOR2_X1 U21251 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19149), .ZN(
        n19665) );
  OAI21_X1 U21252 ( .B1(n19150), .B2(n19665), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19151) );
  OAI21_X1 U21253 ( .B1(n19152), .B2(n19290), .A(n19151), .ZN(n19666) );
  AOI22_X1 U21254 ( .A1(n19666), .A2(n19114), .B1(n19312), .B2(n19665), .ZN(
        n19159) );
  INV_X1 U21255 ( .A(n19667), .ZN(n19664) );
  AOI21_X1 U21256 ( .B1(n19664), .B2(n19676), .A(n13854), .ZN(n19157) );
  OAI21_X1 U21257 ( .B1(n19304), .B2(n19665), .A(n19281), .ZN(n19153) );
  OAI21_X1 U21258 ( .B1(n19154), .B2(n19307), .A(n19153), .ZN(n19155) );
  AOI22_X1 U21259 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19668), .B1(
        n19667), .B2(n19317), .ZN(n19158) );
  OAI211_X1 U21260 ( .C1(n19301), .C2(n19676), .A(n19159), .B(n19158), .ZN(
        P2_U3151) );
  NAND3_X1 U21261 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19256), .ZN(n19168) );
  NOR2_X1 U21262 ( .A1(n19288), .A2(n19168), .ZN(n19671) );
  OAI21_X1 U21263 ( .B1(n15096), .B2(n19671), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19160) );
  OAI21_X1 U21264 ( .B1(n19168), .B2(n19290), .A(n19160), .ZN(n19672) );
  AOI22_X1 U21265 ( .A1(n19672), .A2(n19114), .B1(n19312), .B2(n19671), .ZN(
        n19167) );
  NAND2_X1 U21266 ( .A1(n19178), .A2(n19254), .ZN(n19600) );
  INV_X1 U21267 ( .A(n15096), .ZN(n19161) );
  NOR2_X1 U21268 ( .A1(n19161), .A2(n19307), .ZN(n19165) );
  INV_X1 U21269 ( .A(n19671), .ZN(n19162) );
  AOI21_X1 U21270 ( .B1(n19162), .B2(n19290), .A(n19639), .ZN(n19164) );
  OAI21_X1 U21271 ( .B1(n19179), .B2(n19259), .A(n19168), .ZN(n19163) );
  OAI21_X1 U21272 ( .B1(n19165), .B2(n19164), .A(n19163), .ZN(n19673) );
  AOI22_X1 U21273 ( .A1(n19313), .A2(n19678), .B1(n19673), .B2(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n19166) );
  OAI211_X1 U21274 ( .C1(n19286), .C2(n19676), .A(n19167), .B(n19166), .ZN(
        P2_U3143) );
  NOR2_X1 U21275 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19168), .ZN(
        n19677) );
  AOI22_X1 U21276 ( .A1(n19317), .A2(n19678), .B1(n19312), .B2(n19677), .ZN(
        n19177) );
  OAI21_X1 U21277 ( .B1(n19179), .B2(n19278), .A(n19304), .ZN(n19175) );
  NAND3_X1 U21278 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19260), .A3(
        n19256), .ZN(n19190) );
  INV_X1 U21279 ( .A(n19190), .ZN(n19184) );
  NAND2_X1 U21280 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19184), .ZN(
        n19181) );
  INV_X1 U21281 ( .A(n19181), .ZN(n19683) );
  NOR2_X1 U21282 ( .A1(n19677), .A2(n19683), .ZN(n19174) );
  INV_X1 U21283 ( .A(n19174), .ZN(n19172) );
  INV_X1 U21284 ( .A(n19677), .ZN(n19169) );
  OAI211_X1 U21285 ( .C1(n19170), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19169), 
        .B(n19290), .ZN(n19171) );
  OAI211_X1 U21286 ( .C1(n19175), .C2(n19172), .A(n19281), .B(n19171), .ZN(
        n19680) );
  OAI21_X1 U21287 ( .B1(n15110), .B2(n19677), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19173) );
  OAI21_X1 U21288 ( .B1(n19175), .B2(n19174), .A(n19173), .ZN(n19679) );
  AOI22_X1 U21289 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19680), .B1(
        n19114), .B2(n19679), .ZN(n19176) );
  OAI211_X1 U21290 ( .C1(n19301), .C2(n19688), .A(n19177), .B(n19176), .ZN(
        P2_U3135) );
  AOI22_X1 U21291 ( .A1(n19313), .A2(n19690), .B1(n19312), .B2(n19683), .ZN(
        n19189) );
  OAI21_X1 U21292 ( .B1(n19179), .B2(n19292), .A(n19304), .ZN(n19187) );
  INV_X1 U21293 ( .A(n19185), .ZN(n19180) );
  NOR2_X1 U21294 ( .A1(n19180), .A2(n19307), .ZN(n19183) );
  AOI21_X1 U21295 ( .B1(n19181), .B2(n19290), .A(n19639), .ZN(n19182) );
  OAI22_X1 U21296 ( .A1(n19187), .A2(n19184), .B1(n19183), .B2(n19182), .ZN(
        n19685) );
  OAI21_X1 U21297 ( .B1(n19185), .B2(n19683), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19186) );
  OAI21_X1 U21298 ( .B1(n19187), .B2(n19190), .A(n19186), .ZN(n19684) );
  AOI22_X1 U21299 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19685), .B1(
        n19114), .B2(n19684), .ZN(n19188) );
  OAI211_X1 U21300 ( .C1(n19286), .C2(n19688), .A(n19189), .B(n19188), .ZN(
        P2_U3127) );
  NOR2_X1 U21301 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19190), .ZN(
        n19689) );
  AOI22_X1 U21302 ( .A1(n19317), .A2(n19690), .B1(n19312), .B2(n19689), .ZN(
        n19201) );
  INV_X1 U21303 ( .A(n19196), .ZN(n19194) );
  OAI21_X1 U21304 ( .B1(n19690), .B2(n19698), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19191) );
  NAND2_X1 U21305 ( .A1(n19191), .A2(n19304), .ZN(n19199) );
  NOR2_X1 U21306 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19256), .ZN(
        n19226) );
  AND2_X1 U21307 ( .A1(n19192), .A2(n19226), .ZN(n19696) );
  NOR2_X1 U21308 ( .A1(n19199), .A2(n19696), .ZN(n19193) );
  AOI211_X1 U21309 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19194), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19193), .ZN(n19195) );
  OAI21_X1 U21310 ( .B1(n19689), .B2(n19195), .A(n19281), .ZN(n19692) );
  NOR2_X1 U21311 ( .A1(n19696), .A2(n19689), .ZN(n19198) );
  OAI21_X1 U21312 ( .B1(n19196), .B2(n19689), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19197) );
  AOI22_X1 U21313 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19692), .B1(
        n19691), .B2(n19114), .ZN(n19200) );
  OAI211_X1 U21314 ( .C1(n19301), .C2(n19695), .A(n19201), .B(n19200), .ZN(
        P2_U3119) );
  NAND2_X1 U21315 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19226), .ZN(
        n19211) );
  OAI21_X1 U21316 ( .B1(n19204), .B2(n19696), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19202) );
  OAI21_X1 U21317 ( .B1(n19211), .B2(n19290), .A(n19202), .ZN(n19697) );
  AOI22_X1 U21318 ( .A1(n19697), .A2(n19114), .B1(n19696), .B2(n19312), .ZN(
        n19210) );
  INV_X1 U21319 ( .A(n19203), .ZN(n19208) );
  INV_X1 U21320 ( .A(n19211), .ZN(n19207) );
  AOI21_X1 U21321 ( .B1(n19204), .B2(n19294), .A(n19696), .ZN(n19205) );
  OAI21_X1 U21322 ( .B1(n19205), .B2(n19639), .A(n19306), .ZN(n19206) );
  OAI21_X1 U21323 ( .B1(n19208), .B2(n19207), .A(n19206), .ZN(n19699) );
  AOI22_X1 U21324 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19317), .ZN(n19209) );
  OAI211_X1 U21325 ( .C1(n19301), .C2(n19708), .A(n19210), .B(n19209), .ZN(
        P2_U3111) );
  NOR2_X1 U21326 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19211), .ZN(
        n19702) );
  NOR2_X1 U21327 ( .A1(n19212), .A2(n19702), .ZN(n19216) );
  INV_X1 U21328 ( .A(n19272), .ZN(n19213) );
  INV_X1 U21329 ( .A(n19226), .ZN(n19241) );
  OAI22_X1 U21330 ( .A1(n19216), .A2(n19214), .B1(n19213), .B2(n19241), .ZN(
        n19703) );
  AOI22_X1 U21331 ( .A1(n19703), .A2(n19114), .B1(n19312), .B2(n19702), .ZN(
        n19223) );
  INV_X1 U21332 ( .A(n19702), .ZN(n19215) );
  OAI22_X1 U21333 ( .A1(n19216), .A2(n19307), .B1(n19639), .B2(n19215), .ZN(
        n19219) );
  INV_X1 U21334 ( .A(n19225), .ZN(n19227) );
  OAI22_X1 U21335 ( .A1(n19217), .A2(n19241), .B1(n19227), .B2(n19278), .ZN(
        n19218) );
  OAI21_X1 U21336 ( .B1(n19220), .B2(n19219), .A(n19218), .ZN(n19705) );
  NAND2_X1 U21337 ( .A1(n19225), .A2(n19221), .ZN(n19714) );
  AOI22_X1 U21338 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19313), .ZN(n19222) );
  OAI211_X1 U21339 ( .C1(n19286), .C2(n19708), .A(n19223), .B(n19222), .ZN(
        P2_U3103) );
  NAND2_X1 U21340 ( .A1(n19226), .A2(n19260), .ZN(n19234) );
  NOR2_X1 U21341 ( .A1(n19288), .A2(n19234), .ZN(n19709) );
  AOI22_X1 U21342 ( .A1(n19313), .A2(n19716), .B1(n19312), .B2(n19709), .ZN(
        n19237) );
  OAI21_X1 U21343 ( .B1(n19227), .B2(n19292), .A(n19304), .ZN(n19235) );
  INV_X1 U21344 ( .A(n19234), .ZN(n19231) );
  INV_X1 U21345 ( .A(n19232), .ZN(n19229) );
  OAI21_X1 U21346 ( .B1(n19304), .B2(n19709), .A(n19281), .ZN(n19228) );
  OAI21_X1 U21347 ( .B1(n19229), .B2(n19307), .A(n19228), .ZN(n19230) );
  OAI21_X1 U21348 ( .B1(n19235), .B2(n19231), .A(n19230), .ZN(n19711) );
  OAI21_X1 U21349 ( .B1(n19232), .B2(n19709), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19233) );
  OAI21_X1 U21350 ( .B1(n19235), .B2(n19234), .A(n19233), .ZN(n19710) );
  AOI22_X1 U21351 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19711), .B1(
        n19114), .B2(n19710), .ZN(n19236) );
  OAI211_X1 U21352 ( .C1(n19286), .C2(n19714), .A(n19237), .B(n19236), .ZN(
        P2_U3095) );
  NOR2_X1 U21353 ( .A1(n19303), .A2(n19241), .ZN(n19715) );
  AOI22_X1 U21354 ( .A1(n19317), .A2(n19716), .B1(n19312), .B2(n19715), .ZN(
        n19253) );
  OAI21_X1 U21355 ( .B1(n19723), .B2(n19716), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19242) );
  NAND2_X1 U21356 ( .A1(n19242), .A2(n19304), .ZN(n19251) );
  NOR2_X1 U21357 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19243), .ZN(
        n19247) );
  NOR2_X1 U21358 ( .A1(n15103), .A2(n19307), .ZN(n19246) );
  INV_X1 U21359 ( .A(n19715), .ZN(n19244) );
  AOI21_X1 U21360 ( .B1(n19244), .B2(n19290), .A(n19639), .ZN(n19245) );
  INV_X1 U21361 ( .A(n19247), .ZN(n19250) );
  OAI21_X1 U21362 ( .B1(n19248), .B2(n19715), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19249) );
  AOI22_X1 U21363 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19718), .B1(
        n19114), .B2(n19717), .ZN(n19252) );
  OAI211_X1 U21364 ( .C1(n19301), .C2(n19721), .A(n19253), .B(n19252), .ZN(
        P2_U3087) );
  NAND2_X1 U21365 ( .A1(n19256), .A2(n19255), .ZN(n19302) );
  NOR2_X1 U21366 ( .A1(n19257), .A2(n19302), .ZN(n19722) );
  AOI22_X1 U21367 ( .A1(n19317), .A2(n19723), .B1(n19722), .B2(n19312), .ZN(
        n19269) );
  OAI21_X1 U21368 ( .B1(n19293), .B2(n19259), .A(n19304), .ZN(n19267) );
  NOR2_X1 U21369 ( .A1(n19260), .A2(n19302), .ZN(n19264) );
  INV_X1 U21370 ( .A(n19265), .ZN(n19262) );
  OAI21_X1 U21371 ( .B1(n19304), .B2(n19722), .A(n19281), .ZN(n19261) );
  OAI21_X1 U21372 ( .B1(n19262), .B2(n19307), .A(n19261), .ZN(n19263) );
  OAI21_X1 U21373 ( .B1(n19267), .B2(n19264), .A(n19263), .ZN(n19725) );
  INV_X1 U21374 ( .A(n19264), .ZN(n19270) );
  OAI21_X1 U21375 ( .B1(n19265), .B2(n19722), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19266) );
  OAI21_X1 U21376 ( .B1(n19267), .B2(n19270), .A(n19266), .ZN(n19724) );
  AOI22_X1 U21377 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19725), .B1(
        n19114), .B2(n19724), .ZN(n19268) );
  OAI211_X1 U21378 ( .C1(n19301), .C2(n19733), .A(n19269), .B(n19268), .ZN(
        P2_U3079) );
  NOR2_X1 U21379 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19270), .ZN(
        n19728) );
  OAI21_X1 U21380 ( .B1(n19274), .B2(n19728), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19273) );
  INV_X1 U21381 ( .A(n19302), .ZN(n19271) );
  NAND2_X1 U21382 ( .A1(n19272), .A2(n19271), .ZN(n19277) );
  NAND2_X1 U21383 ( .A1(n19273), .A2(n19277), .ZN(n19729) );
  AOI22_X1 U21384 ( .A1(n19729), .A2(n19114), .B1(n19312), .B2(n19728), .ZN(
        n19285) );
  INV_X1 U21385 ( .A(n19274), .ZN(n19276) );
  INV_X1 U21386 ( .A(n19728), .ZN(n19275) );
  OAI21_X1 U21387 ( .B1(n19276), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19275), 
        .ZN(n19280) );
  OAI21_X1 U21388 ( .B1(n19293), .B2(n19278), .A(n19277), .ZN(n19279) );
  MUX2_X1 U21389 ( .A(n19280), .B(n19279), .S(n19304), .Z(n19282) );
  NAND2_X1 U21390 ( .A1(n19282), .A2(n19281), .ZN(n19730) );
  NOR2_X2 U21391 ( .A1(n19293), .A2(n19283), .ZN(n19737) );
  AOI22_X1 U21392 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19730), .B1(
        n19737), .B2(n19313), .ZN(n19284) );
  OAI211_X1 U21393 ( .C1(n19286), .C2(n19733), .A(n19285), .B(n19284), .ZN(
        P2_U3071) );
  OR2_X1 U21394 ( .A1(n19302), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19291) );
  NOR2_X1 U21395 ( .A1(n19288), .A2(n19291), .ZN(n19735) );
  OAI21_X1 U21396 ( .B1(n15095), .B2(n19735), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19289) );
  OAI21_X1 U21397 ( .B1(n19291), .B2(n19290), .A(n19289), .ZN(n19736) );
  AOI22_X1 U21398 ( .A1(n19736), .A2(n19114), .B1(n19312), .B2(n19735), .ZN(
        n19300) );
  OAI21_X1 U21399 ( .B1(n19293), .B2(n19292), .A(n19291), .ZN(n19298) );
  INV_X1 U21400 ( .A(n19735), .ZN(n19296) );
  NAND2_X1 U21401 ( .A1(n15095), .A2(n19294), .ZN(n19295) );
  OAI211_X1 U21402 ( .C1(n19639), .C2(n19296), .A(n19295), .B(n19306), .ZN(
        n19297) );
  NAND2_X1 U21403 ( .A1(n19298), .A2(n19297), .ZN(n19738) );
  AOI22_X1 U21404 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19738), .B1(
        n19737), .B2(n19317), .ZN(n19299) );
  OAI211_X1 U21405 ( .C1(n19301), .C2(n19741), .A(n19300), .B(n19299), .ZN(
        P2_U3063) );
  NOR2_X1 U21406 ( .A1(n19303), .A2(n19302), .ZN(n19743) );
  INV_X1 U21407 ( .A(n19743), .ZN(n19311) );
  NOR2_X1 U21408 ( .A1(n19745), .A2(n19750), .ZN(n19305) );
  OAI21_X1 U21409 ( .B1(n19305), .B2(n13854), .A(n19304), .ZN(n19316) );
  OAI21_X1 U21410 ( .B1(n19308), .B2(n19307), .A(n19306), .ZN(n19309) );
  OAI21_X1 U21411 ( .B1(n19316), .B2(n19643), .A(n19309), .ZN(n19310) );
  AOI22_X1 U21412 ( .A1(n19313), .A2(n19745), .B1(n19312), .B2(n19743), .ZN(
        n19319) );
  NOR2_X1 U21413 ( .A1(n19643), .A2(n19743), .ZN(n19315) );
  OAI21_X1 U21414 ( .B1(n15109), .B2(n19743), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19314) );
  AOI22_X1 U21415 ( .A1(n19114), .A2(n19748), .B1(n19750), .B2(n19317), .ZN(
        n19318) );
  OAI211_X1 U21416 ( .C1(n19754), .C2(n19320), .A(n19319), .B(n19318), .ZN(
        P2_U3055) );
  AOI22_X1 U21417 ( .A1(n19629), .A2(n19321), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19627), .ZN(n19326) );
  AOI22_X1 U21418 ( .A1(n19631), .A2(BUF1_REG_22__SCAN_IN), .B1(n19630), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n19325) );
  AOI22_X1 U21419 ( .A1(n19323), .A2(n19634), .B1(n19633), .B2(n19322), .ZN(
        n19324) );
  NAND3_X1 U21420 ( .A1(n19326), .A2(n19325), .A3(n19324), .ZN(P2_U2897) );
  OAI222_X1 U21421 ( .A1(n19328), .A2(n19378), .B1(n19327), .B2(n19531), .C1(
        n19583), .C2(n19329), .ZN(P2_U2913) );
  AOI22_X1 U21422 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19645), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19646), .ZN(n19363) );
  NOR2_X2 U21423 ( .A1(n13035), .A2(n19641), .ZN(n19364) );
  AOI22_X1 U21424 ( .A1(n19644), .A2(n19330), .B1(n19643), .B2(n19364), .ZN(
        n19332) );
  AOI22_X1 U21425 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19645), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19646), .ZN(n19360) );
  AOI22_X1 U21426 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19647), .B1(
        n19745), .B2(n19366), .ZN(n19331) );
  OAI211_X1 U21427 ( .C1(n19363), .C2(n19650), .A(n19332), .B(n19331), .ZN(
        P2_U3174) );
  AOI22_X1 U21428 ( .A1(n19365), .A2(n19660), .B1(n19364), .B2(n19651), .ZN(
        n19334) );
  AOI22_X1 U21429 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19654), .B1(
        n19330), .B2(n19653), .ZN(n19333) );
  OAI211_X1 U21430 ( .C1(n19360), .C2(n19650), .A(n19334), .B(n19333), .ZN(
        P2_U3166) );
  INV_X1 U21431 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n19337) );
  AOI22_X1 U21432 ( .A1(n19659), .A2(n19330), .B1(n19364), .B2(n19658), .ZN(
        n19336) );
  AOI22_X1 U21433 ( .A1(n19660), .A2(n19366), .B1(n19667), .B2(n19365), .ZN(
        n19335) );
  OAI211_X1 U21434 ( .C1(n19435), .C2(n19337), .A(n19336), .B(n19335), .ZN(
        P2_U3158) );
  AOI22_X1 U21435 ( .A1(n19666), .A2(n19330), .B1(n19364), .B2(n19665), .ZN(
        n19339) );
  AOI22_X1 U21436 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19668), .B1(
        n19667), .B2(n19366), .ZN(n19338) );
  OAI211_X1 U21437 ( .C1(n19363), .C2(n19676), .A(n19339), .B(n19338), .ZN(
        P2_U3150) );
  AOI22_X1 U21438 ( .A1(n19672), .A2(n19330), .B1(n19364), .B2(n19671), .ZN(
        n19341) );
  AOI22_X1 U21439 ( .A1(n19365), .A2(n19678), .B1(n19673), .B2(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n19340) );
  OAI211_X1 U21440 ( .C1(n19360), .C2(n19676), .A(n19341), .B(n19340), .ZN(
        P2_U3142) );
  INV_X1 U21441 ( .A(n19688), .ZN(n19597) );
  AOI22_X1 U21442 ( .A1(n19365), .A2(n19597), .B1(n19364), .B2(n19677), .ZN(
        n19343) );
  AOI22_X1 U21443 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19680), .B1(
        n19330), .B2(n19679), .ZN(n19342) );
  OAI211_X1 U21444 ( .C1(n19360), .C2(n19600), .A(n19343), .B(n19342), .ZN(
        P2_U3134) );
  AOI22_X1 U21445 ( .A1(n19365), .A2(n19690), .B1(n19364), .B2(n19683), .ZN(
        n19345) );
  AOI22_X1 U21446 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19685), .B1(
        n19330), .B2(n19684), .ZN(n19344) );
  OAI211_X1 U21447 ( .C1(n19360), .C2(n19688), .A(n19345), .B(n19344), .ZN(
        P2_U3126) );
  AOI22_X1 U21448 ( .A1(n19366), .A2(n19690), .B1(n19364), .B2(n19689), .ZN(
        n19347) );
  AOI22_X1 U21449 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19692), .B1(
        n19691), .B2(n19330), .ZN(n19346) );
  OAI211_X1 U21450 ( .C1(n19363), .C2(n19695), .A(n19347), .B(n19346), .ZN(
        P2_U3118) );
  AOI22_X1 U21451 ( .A1(n19697), .A2(n19330), .B1(n19696), .B2(n19364), .ZN(
        n19349) );
  AOI22_X1 U21452 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19366), .ZN(n19348) );
  OAI211_X1 U21453 ( .C1(n19363), .C2(n19708), .A(n19349), .B(n19348), .ZN(
        P2_U3110) );
  AOI22_X1 U21454 ( .A1(n19703), .A2(n19330), .B1(n19364), .B2(n19702), .ZN(
        n19351) );
  AOI22_X1 U21455 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19365), .ZN(n19350) );
  OAI211_X1 U21456 ( .C1(n19360), .C2(n19708), .A(n19351), .B(n19350), .ZN(
        P2_U3102) );
  AOI22_X1 U21457 ( .A1(n19365), .A2(n19716), .B1(n19364), .B2(n19709), .ZN(
        n19353) );
  AOI22_X1 U21458 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19711), .B1(
        n19330), .B2(n19710), .ZN(n19352) );
  OAI211_X1 U21459 ( .C1(n19360), .C2(n19714), .A(n19353), .B(n19352), .ZN(
        P2_U3094) );
  AOI22_X1 U21460 ( .A1(n19366), .A2(n19716), .B1(n19364), .B2(n19715), .ZN(
        n19355) );
  AOI22_X1 U21461 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19718), .B1(
        n19330), .B2(n19717), .ZN(n19354) );
  OAI211_X1 U21462 ( .C1(n19363), .C2(n19721), .A(n19355), .B(n19354), .ZN(
        P2_U3086) );
  AOI22_X1 U21463 ( .A1(n19366), .A2(n19723), .B1(n19722), .B2(n19364), .ZN(
        n19357) );
  AOI22_X1 U21464 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19725), .B1(
        n19330), .B2(n19724), .ZN(n19356) );
  OAI211_X1 U21465 ( .C1(n19363), .C2(n19733), .A(n19357), .B(n19356), .ZN(
        P2_U3078) );
  AOI22_X1 U21466 ( .A1(n19729), .A2(n19330), .B1(n19364), .B2(n19728), .ZN(
        n19359) );
  AOI22_X1 U21467 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19730), .B1(
        n19737), .B2(n19365), .ZN(n19358) );
  OAI211_X1 U21468 ( .C1(n19360), .C2(n19733), .A(n19359), .B(n19358), .ZN(
        P2_U3070) );
  AOI22_X1 U21469 ( .A1(n19736), .A2(n19330), .B1(n19364), .B2(n19735), .ZN(
        n19362) );
  AOI22_X1 U21470 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19738), .B1(
        n19737), .B2(n19366), .ZN(n19361) );
  OAI211_X1 U21471 ( .C1(n19363), .C2(n19741), .A(n19362), .B(n19361), .ZN(
        P2_U3062) );
  AOI22_X1 U21472 ( .A1(n19365), .A2(n19745), .B1(n19364), .B2(n19743), .ZN(
        n19368) );
  AOI22_X1 U21473 ( .A1(n19750), .A2(n19366), .B1(n19748), .B2(n19330), .ZN(
        n19367) );
  OAI211_X1 U21474 ( .C1(n19754), .C2(n19369), .A(n19368), .B(n19367), .ZN(
        P2_U3054) );
  OAI22_X1 U21475 ( .A1(n19370), .A2(n19531), .B1(n19379), .B2(n19583), .ZN(
        n19371) );
  INV_X1 U21476 ( .A(n19371), .ZN(n19376) );
  INV_X1 U21477 ( .A(n19372), .ZN(n19373) );
  NAND3_X1 U21478 ( .A1(n19374), .A2(n19373), .A3(n19634), .ZN(n19375) );
  OAI211_X1 U21479 ( .C1(n19378), .C2(n19377), .A(n19376), .B(n19375), .ZN(
        P2_U2914) );
  AOI22_X1 U21480 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19645), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19646), .ZN(n19411) );
  AOI22_X1 U21481 ( .A1(n19644), .A2(n19380), .B1(n19643), .B2(n19382), .ZN(
        n19384) );
  AOI22_X1 U21482 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19645), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19646), .ZN(n19414) );
  AOI22_X1 U21483 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19647), .B1(
        n19652), .B2(n19415), .ZN(n19383) );
  OAI211_X1 U21484 ( .C1(n19411), .C2(n19537), .A(n19384), .B(n19383), .ZN(
        P2_U3173) );
  AOI22_X1 U21485 ( .A1(n19415), .A2(n19660), .B1(n19382), .B2(n19651), .ZN(
        n19386) );
  AOI22_X1 U21486 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19654), .B1(
        n19380), .B2(n19653), .ZN(n19385) );
  OAI211_X1 U21487 ( .C1(n19411), .C2(n19650), .A(n19386), .B(n19385), .ZN(
        P2_U3165) );
  AOI22_X1 U21488 ( .A1(n19659), .A2(n19380), .B1(n19382), .B2(n19658), .ZN(
        n19388) );
  AOI22_X1 U21489 ( .A1(n19660), .A2(n19416), .B1(n19667), .B2(n19415), .ZN(
        n19387) );
  OAI211_X1 U21490 ( .C1(n19435), .C2(n13453), .A(n19388), .B(n19387), .ZN(
        P2_U3157) );
  AOI22_X1 U21491 ( .A1(n19666), .A2(n19380), .B1(n19382), .B2(n19665), .ZN(
        n19390) );
  AOI22_X1 U21492 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19668), .B1(
        n19667), .B2(n19416), .ZN(n19389) );
  OAI211_X1 U21493 ( .C1(n19414), .C2(n19676), .A(n19390), .B(n19389), .ZN(
        P2_U3149) );
  AOI22_X1 U21494 ( .A1(n19672), .A2(n19380), .B1(n19382), .B2(n19671), .ZN(
        n19392) );
  AOI22_X1 U21495 ( .A1(n19415), .A2(n19678), .B1(n19673), .B2(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n19391) );
  OAI211_X1 U21496 ( .C1(n19411), .C2(n19676), .A(n19392), .B(n19391), .ZN(
        P2_U3141) );
  AOI22_X1 U21497 ( .A1(n19416), .A2(n19678), .B1(n19382), .B2(n19677), .ZN(
        n19394) );
  AOI22_X1 U21498 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19680), .B1(
        n19380), .B2(n19679), .ZN(n19393) );
  OAI211_X1 U21499 ( .C1(n19414), .C2(n19688), .A(n19394), .B(n19393), .ZN(
        P2_U3133) );
  AOI22_X1 U21500 ( .A1(n19415), .A2(n19690), .B1(n19382), .B2(n19683), .ZN(
        n19396) );
  AOI22_X1 U21501 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19685), .B1(
        n19380), .B2(n19684), .ZN(n19395) );
  OAI211_X1 U21502 ( .C1(n19411), .C2(n19688), .A(n19396), .B(n19395), .ZN(
        P2_U3125) );
  AOI22_X1 U21503 ( .A1(n19416), .A2(n19690), .B1(n19382), .B2(n19689), .ZN(
        n19398) );
  AOI22_X1 U21504 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19692), .B1(
        n19691), .B2(n19380), .ZN(n19397) );
  OAI211_X1 U21505 ( .C1(n19414), .C2(n19695), .A(n19398), .B(n19397), .ZN(
        P2_U3117) );
  AOI22_X1 U21506 ( .A1(n19697), .A2(n19380), .B1(n19696), .B2(n19382), .ZN(
        n19400) );
  AOI22_X1 U21507 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19416), .ZN(n19399) );
  OAI211_X1 U21508 ( .C1(n19414), .C2(n19708), .A(n19400), .B(n19399), .ZN(
        P2_U3109) );
  AOI22_X1 U21509 ( .A1(n19703), .A2(n19380), .B1(n19382), .B2(n19702), .ZN(
        n19402) );
  AOI22_X1 U21510 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19415), .ZN(n19401) );
  OAI211_X1 U21511 ( .C1(n19411), .C2(n19708), .A(n19402), .B(n19401), .ZN(
        P2_U3101) );
  AOI22_X1 U21512 ( .A1(n19415), .A2(n19716), .B1(n19382), .B2(n19709), .ZN(
        n19404) );
  AOI22_X1 U21513 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19711), .B1(
        n19380), .B2(n19710), .ZN(n19403) );
  OAI211_X1 U21514 ( .C1(n19411), .C2(n19714), .A(n19404), .B(n19403), .ZN(
        P2_U3093) );
  AOI22_X1 U21515 ( .A1(n19416), .A2(n19716), .B1(n19382), .B2(n19715), .ZN(
        n19406) );
  AOI22_X1 U21516 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19718), .B1(
        n19380), .B2(n19717), .ZN(n19405) );
  OAI211_X1 U21517 ( .C1(n19414), .C2(n19721), .A(n19406), .B(n19405), .ZN(
        P2_U3085) );
  AOI22_X1 U21518 ( .A1(n19416), .A2(n19723), .B1(n19722), .B2(n19382), .ZN(
        n19408) );
  AOI22_X1 U21519 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19725), .B1(
        n19380), .B2(n19724), .ZN(n19407) );
  OAI211_X1 U21520 ( .C1(n19414), .C2(n19733), .A(n19408), .B(n19407), .ZN(
        P2_U3077) );
  AOI22_X1 U21521 ( .A1(n19729), .A2(n19380), .B1(n19382), .B2(n19728), .ZN(
        n19410) );
  AOI22_X1 U21522 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19730), .B1(
        n19737), .B2(n19415), .ZN(n19409) );
  OAI211_X1 U21523 ( .C1(n19411), .C2(n19733), .A(n19410), .B(n19409), .ZN(
        P2_U3069) );
  AOI22_X1 U21524 ( .A1(n19736), .A2(n19380), .B1(n19382), .B2(n19735), .ZN(
        n19413) );
  AOI22_X1 U21525 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19738), .B1(
        n19737), .B2(n19416), .ZN(n19412) );
  OAI211_X1 U21526 ( .C1(n19414), .C2(n19741), .A(n19413), .B(n19412), .ZN(
        P2_U3061) );
  AOI22_X1 U21527 ( .A1(n19415), .A2(n19745), .B1(n19382), .B2(n19743), .ZN(
        n19418) );
  AOI22_X1 U21528 ( .A1(n19750), .A2(n19416), .B1(n19748), .B2(n19380), .ZN(
        n19417) );
  OAI211_X1 U21529 ( .C1(n19754), .C2(n19419), .A(n19418), .B(n19417), .ZN(
        P2_U3053) );
  AOI22_X1 U21530 ( .A1(n19629), .A2(n19428), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19627), .ZN(n19427) );
  AOI22_X1 U21531 ( .A1(n19631), .A2(BUF1_REG_20__SCAN_IN), .B1(n19630), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n19426) );
  INV_X1 U21532 ( .A(n19633), .ZN(n19422) );
  INV_X1 U21533 ( .A(n19420), .ZN(n19421) );
  OAI22_X1 U21534 ( .A1(n19423), .A2(n19579), .B1(n19422), .B2(n19421), .ZN(
        n19424) );
  INV_X1 U21535 ( .A(n19424), .ZN(n19425) );
  NAND3_X1 U21536 ( .A1(n19427), .A2(n19426), .A3(n19425), .ZN(P2_U2899) );
  AOI22_X1 U21537 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19646), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19645), .ZN(n19463) );
  INV_X1 U21538 ( .A(n19428), .ZN(n19429) );
  NOR2_X2 U21539 ( .A1(n12992), .A2(n19641), .ZN(n19464) );
  AOI22_X1 U21540 ( .A1(n19644), .A2(n19430), .B1(n19643), .B2(n19464), .ZN(
        n19432) );
  AOI22_X1 U21541 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19645), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19646), .ZN(n19460) );
  AOI22_X1 U21542 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19647), .B1(
        n19745), .B2(n19466), .ZN(n19431) );
  OAI211_X1 U21543 ( .C1(n19463), .C2(n19650), .A(n19432), .B(n19431), .ZN(
        P2_U3172) );
  AOI22_X1 U21544 ( .A1(n19466), .A2(n19652), .B1(n19464), .B2(n19651), .ZN(
        n19434) );
  AOI22_X1 U21545 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19654), .B1(
        n19430), .B2(n19653), .ZN(n19433) );
  OAI211_X1 U21546 ( .C1(n19463), .C2(n19657), .A(n19434), .B(n19433), .ZN(
        P2_U3164) );
  AOI22_X1 U21547 ( .A1(n19659), .A2(n19430), .B1(n19464), .B2(n19658), .ZN(
        n19437) );
  INV_X1 U21548 ( .A(n19435), .ZN(n19661) );
  AOI22_X1 U21549 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19661), .B1(
        n19660), .B2(n19466), .ZN(n19436) );
  OAI211_X1 U21550 ( .C1(n19463), .C2(n19664), .A(n19437), .B(n19436), .ZN(
        P2_U3156) );
  AOI22_X1 U21551 ( .A1(n19666), .A2(n19430), .B1(n19464), .B2(n19665), .ZN(
        n19439) );
  AOI22_X1 U21552 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19668), .B1(
        n19667), .B2(n19466), .ZN(n19438) );
  OAI211_X1 U21553 ( .C1(n19463), .C2(n19676), .A(n19439), .B(n19438), .ZN(
        P2_U3148) );
  AOI22_X1 U21554 ( .A1(n19672), .A2(n19430), .B1(n19464), .B2(n19671), .ZN(
        n19441) );
  INV_X1 U21555 ( .A(n19463), .ZN(n19465) );
  AOI22_X1 U21556 ( .A1(n19465), .A2(n19678), .B1(n19673), .B2(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n19440) );
  OAI211_X1 U21557 ( .C1(n19460), .C2(n19676), .A(n19441), .B(n19440), .ZN(
        P2_U3140) );
  AOI22_X1 U21558 ( .A1(n19466), .A2(n19678), .B1(n19464), .B2(n19677), .ZN(
        n19443) );
  AOI22_X1 U21559 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19680), .B1(
        n19430), .B2(n19679), .ZN(n19442) );
  OAI211_X1 U21560 ( .C1(n19463), .C2(n19688), .A(n19443), .B(n19442), .ZN(
        P2_U3132) );
  AOI22_X1 U21561 ( .A1(n19465), .A2(n19690), .B1(n19464), .B2(n19683), .ZN(
        n19445) );
  AOI22_X1 U21562 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19685), .B1(
        n19430), .B2(n19684), .ZN(n19444) );
  OAI211_X1 U21563 ( .C1(n19460), .C2(n19688), .A(n19445), .B(n19444), .ZN(
        P2_U3124) );
  AOI22_X1 U21564 ( .A1(n19466), .A2(n19690), .B1(n19464), .B2(n19689), .ZN(
        n19447) );
  AOI22_X1 U21565 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19692), .B1(
        n19691), .B2(n19430), .ZN(n19446) );
  OAI211_X1 U21566 ( .C1(n19463), .C2(n19695), .A(n19447), .B(n19446), .ZN(
        P2_U3116) );
  AOI22_X1 U21567 ( .A1(n19697), .A2(n19430), .B1(n19696), .B2(n19464), .ZN(
        n19449) );
  AOI22_X1 U21568 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19466), .ZN(n19448) );
  OAI211_X1 U21569 ( .C1(n19463), .C2(n19708), .A(n19449), .B(n19448), .ZN(
        P2_U3108) );
  AOI22_X1 U21570 ( .A1(n19703), .A2(n19430), .B1(n19464), .B2(n19702), .ZN(
        n19451) );
  AOI22_X1 U21571 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19465), .ZN(n19450) );
  OAI211_X1 U21572 ( .C1(n19460), .C2(n19708), .A(n19451), .B(n19450), .ZN(
        P2_U3100) );
  AOI22_X1 U21573 ( .A1(n19465), .A2(n19716), .B1(n19464), .B2(n19709), .ZN(
        n19453) );
  AOI22_X1 U21574 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19711), .B1(
        n19430), .B2(n19710), .ZN(n19452) );
  OAI211_X1 U21575 ( .C1(n19460), .C2(n19714), .A(n19453), .B(n19452), .ZN(
        P2_U3092) );
  AOI22_X1 U21576 ( .A1(n19466), .A2(n19716), .B1(n19464), .B2(n19715), .ZN(
        n19455) );
  AOI22_X1 U21577 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19718), .B1(
        n19430), .B2(n19717), .ZN(n19454) );
  OAI211_X1 U21578 ( .C1(n19463), .C2(n19721), .A(n19455), .B(n19454), .ZN(
        P2_U3084) );
  AOI22_X1 U21579 ( .A1(n19466), .A2(n19723), .B1(n19722), .B2(n19464), .ZN(
        n19457) );
  AOI22_X1 U21580 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19725), .B1(
        n19430), .B2(n19724), .ZN(n19456) );
  OAI211_X1 U21581 ( .C1(n19463), .C2(n19733), .A(n19457), .B(n19456), .ZN(
        P2_U3076) );
  AOI22_X1 U21582 ( .A1(n19729), .A2(n19430), .B1(n19464), .B2(n19728), .ZN(
        n19459) );
  AOI22_X1 U21583 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19730), .B1(
        n19737), .B2(n19465), .ZN(n19458) );
  OAI211_X1 U21584 ( .C1(n19460), .C2(n19733), .A(n19459), .B(n19458), .ZN(
        P2_U3068) );
  AOI22_X1 U21585 ( .A1(n19736), .A2(n19430), .B1(n19464), .B2(n19735), .ZN(
        n19462) );
  AOI22_X1 U21586 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19738), .B1(
        n19737), .B2(n19466), .ZN(n19461) );
  OAI211_X1 U21587 ( .C1(n19463), .C2(n19741), .A(n19462), .B(n19461), .ZN(
        P2_U3060) );
  AOI22_X1 U21588 ( .A1(n19465), .A2(n19745), .B1(n19464), .B2(n19743), .ZN(
        n19468) );
  AOI22_X1 U21589 ( .A1(n19750), .A2(n19466), .B1(n19748), .B2(n19430), .ZN(
        n19467) );
  OAI211_X1 U21590 ( .C1(n19754), .C2(n19469), .A(n19468), .B(n19467), .ZN(
        P2_U3052) );
  AOI22_X1 U21591 ( .A1(n19470), .A2(n19633), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19627), .ZN(n19476) );
  AOI21_X1 U21592 ( .B1(n19473), .B2(n19472), .A(n19471), .ZN(n19474) );
  OR2_X1 U21593 ( .A1(n19474), .A2(n19579), .ZN(n19475) );
  OAI211_X1 U21594 ( .C1(n19477), .C2(n19583), .A(n19476), .B(n19475), .ZN(
        P2_U2916) );
  AOI22_X1 U21595 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19645), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19646), .ZN(n19510) );
  NOR2_X2 U21596 ( .A1(n19477), .A2(n19639), .ZN(n19513) );
  NOR2_X2 U21597 ( .A1(n19478), .A2(n19641), .ZN(n19511) );
  AOI22_X1 U21598 ( .A1(n19644), .A2(n19513), .B1(n19643), .B2(n19511), .ZN(
        n19480) );
  AOI22_X1 U21599 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n19646), .B1(
        BUF1_REG_19__SCAN_IN), .B2(n19645), .ZN(n19507) );
  AOI22_X1 U21600 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19647), .B1(
        n19745), .B2(n19514), .ZN(n19479) );
  OAI211_X1 U21601 ( .C1(n19510), .C2(n19650), .A(n19480), .B(n19479), .ZN(
        P2_U3171) );
  AOI22_X1 U21602 ( .A1(n19514), .A2(n19652), .B1(n19511), .B2(n19651), .ZN(
        n19482) );
  AOI22_X1 U21603 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19654), .B1(
        n19513), .B2(n19653), .ZN(n19481) );
  OAI211_X1 U21604 ( .C1(n19510), .C2(n19657), .A(n19482), .B(n19481), .ZN(
        P2_U3163) );
  AOI22_X1 U21605 ( .A1(n19659), .A2(n19513), .B1(n19511), .B2(n19658), .ZN(
        n19484) );
  INV_X1 U21606 ( .A(n19510), .ZN(n19512) );
  AOI22_X1 U21607 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19661), .B1(
        n19667), .B2(n19512), .ZN(n19483) );
  OAI211_X1 U21608 ( .C1(n19507), .C2(n19657), .A(n19484), .B(n19483), .ZN(
        P2_U3155) );
  AOI22_X1 U21609 ( .A1(n19666), .A2(n19513), .B1(n19511), .B2(n19665), .ZN(
        n19486) );
  AOI22_X1 U21610 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19668), .B1(
        n19667), .B2(n19514), .ZN(n19485) );
  OAI211_X1 U21611 ( .C1(n19510), .C2(n19676), .A(n19486), .B(n19485), .ZN(
        P2_U3147) );
  AOI22_X1 U21612 ( .A1(n19672), .A2(n19513), .B1(n19511), .B2(n19671), .ZN(
        n19488) );
  AOI22_X1 U21613 ( .A1(n19512), .A2(n19678), .B1(n19673), .B2(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n19487) );
  OAI211_X1 U21614 ( .C1(n19507), .C2(n19676), .A(n19488), .B(n19487), .ZN(
        P2_U3139) );
  AOI22_X1 U21615 ( .A1(n19512), .A2(n19597), .B1(n19511), .B2(n19677), .ZN(
        n19490) );
  AOI22_X1 U21616 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19680), .B1(
        n19513), .B2(n19679), .ZN(n19489) );
  OAI211_X1 U21617 ( .C1(n19507), .C2(n19600), .A(n19490), .B(n19489), .ZN(
        P2_U3131) );
  AOI22_X1 U21618 ( .A1(n19512), .A2(n19690), .B1(n19511), .B2(n19683), .ZN(
        n19492) );
  AOI22_X1 U21619 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19685), .B1(
        n19513), .B2(n19684), .ZN(n19491) );
  OAI211_X1 U21620 ( .C1(n19507), .C2(n19688), .A(n19492), .B(n19491), .ZN(
        P2_U3123) );
  AOI22_X1 U21621 ( .A1(n19514), .A2(n19690), .B1(n19511), .B2(n19689), .ZN(
        n19494) );
  AOI22_X1 U21622 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19692), .B1(
        n19691), .B2(n19513), .ZN(n19493) );
  OAI211_X1 U21623 ( .C1(n19510), .C2(n19695), .A(n19494), .B(n19493), .ZN(
        P2_U3115) );
  AOI22_X1 U21624 ( .A1(n19697), .A2(n19513), .B1(n19696), .B2(n19511), .ZN(
        n19496) );
  AOI22_X1 U21625 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19514), .ZN(n19495) );
  OAI211_X1 U21626 ( .C1(n19510), .C2(n19708), .A(n19496), .B(n19495), .ZN(
        P2_U3107) );
  AOI22_X1 U21627 ( .A1(n19703), .A2(n19513), .B1(n19511), .B2(n19702), .ZN(
        n19498) );
  AOI22_X1 U21628 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19512), .ZN(n19497) );
  OAI211_X1 U21629 ( .C1(n19507), .C2(n19708), .A(n19498), .B(n19497), .ZN(
        P2_U3099) );
  AOI22_X1 U21630 ( .A1(n19512), .A2(n19716), .B1(n19511), .B2(n19709), .ZN(
        n19500) );
  AOI22_X1 U21631 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19711), .B1(
        n19513), .B2(n19710), .ZN(n19499) );
  OAI211_X1 U21632 ( .C1(n19507), .C2(n19714), .A(n19500), .B(n19499), .ZN(
        P2_U3091) );
  AOI22_X1 U21633 ( .A1(n19514), .A2(n19716), .B1(n19511), .B2(n19715), .ZN(
        n19502) );
  AOI22_X1 U21634 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19718), .B1(
        n19513), .B2(n19717), .ZN(n19501) );
  OAI211_X1 U21635 ( .C1(n19510), .C2(n19721), .A(n19502), .B(n19501), .ZN(
        P2_U3083) );
  AOI22_X1 U21636 ( .A1(n19514), .A2(n19723), .B1(n19722), .B2(n19511), .ZN(
        n19504) );
  AOI22_X1 U21637 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19725), .B1(
        n19513), .B2(n19724), .ZN(n19503) );
  OAI211_X1 U21638 ( .C1(n19510), .C2(n19733), .A(n19504), .B(n19503), .ZN(
        P2_U3075) );
  AOI22_X1 U21639 ( .A1(n19729), .A2(n19513), .B1(n19511), .B2(n19728), .ZN(
        n19506) );
  AOI22_X1 U21640 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19730), .B1(
        n19737), .B2(n19512), .ZN(n19505) );
  OAI211_X1 U21641 ( .C1(n19507), .C2(n19733), .A(n19506), .B(n19505), .ZN(
        P2_U3067) );
  AOI22_X1 U21642 ( .A1(n19736), .A2(n19513), .B1(n19511), .B2(n19735), .ZN(
        n19509) );
  AOI22_X1 U21643 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19738), .B1(
        n19737), .B2(n19514), .ZN(n19508) );
  OAI211_X1 U21644 ( .C1(n19510), .C2(n19741), .A(n19509), .B(n19508), .ZN(
        P2_U3059) );
  AOI22_X1 U21645 ( .A1(n19512), .A2(n19745), .B1(n19511), .B2(n19743), .ZN(
        n19516) );
  AOI22_X1 U21646 ( .A1(n19750), .A2(n19514), .B1(n19748), .B2(n19513), .ZN(
        n19515) );
  OAI211_X1 U21647 ( .C1(n19754), .C2(n19517), .A(n19516), .B(n19515), .ZN(
        P2_U3051) );
  AOI22_X1 U21648 ( .A1(n19629), .A2(n19532), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19627), .ZN(n19522) );
  AOI22_X1 U21649 ( .A1(n19631), .A2(BUF1_REG_18__SCAN_IN), .B1(n19630), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n19521) );
  AOI22_X1 U21650 ( .A1(n19519), .A2(n19634), .B1(n19633), .B2(n19518), .ZN(
        n19520) );
  NAND3_X1 U21651 ( .A1(n19522), .A2(n19521), .A3(n19520), .ZN(P2_U2901) );
  AOI22_X1 U21652 ( .A1(n19524), .A2(n19532), .B1(n19633), .B2(n19523), .ZN(
        n19529) );
  XNOR2_X1 U21653 ( .A(n19526), .B(n19525), .ZN(n19527) );
  NAND2_X1 U21654 ( .A1(n19527), .A2(n19634), .ZN(n19528) );
  OAI211_X1 U21655 ( .C1(n19531), .C2(n19530), .A(n19529), .B(n19528), .ZN(
        P2_U2917) );
  AOI22_X1 U21656 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19645), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19646), .ZN(n19564) );
  INV_X1 U21657 ( .A(n19532), .ZN(n19533) );
  NOR2_X2 U21658 ( .A1(n19533), .A2(n19639), .ZN(n19570) );
  NOR2_X2 U21659 ( .A1(n19534), .A2(n19641), .ZN(n19568) );
  AOI22_X1 U21660 ( .A1(n19644), .A2(n19570), .B1(n19643), .B2(n19568), .ZN(
        n19536) );
  AOI22_X1 U21661 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19645), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19646), .ZN(n19567) );
  AOI22_X1 U21662 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19647), .B1(
        n19652), .B2(n19569), .ZN(n19535) );
  OAI211_X1 U21663 ( .C1(n19564), .C2(n19537), .A(n19536), .B(n19535), .ZN(
        P2_U3170) );
  INV_X1 U21664 ( .A(n19564), .ZN(n19571) );
  AOI22_X1 U21665 ( .A1(n19571), .A2(n19652), .B1(n19568), .B2(n19651), .ZN(
        n19539) );
  AOI22_X1 U21666 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19654), .B1(
        n19570), .B2(n19653), .ZN(n19538) );
  OAI211_X1 U21667 ( .C1(n19567), .C2(n19657), .A(n19539), .B(n19538), .ZN(
        P2_U3162) );
  AOI22_X1 U21668 ( .A1(n19659), .A2(n19570), .B1(n19568), .B2(n19658), .ZN(
        n19541) );
  AOI22_X1 U21669 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19661), .B1(
        n19667), .B2(n19569), .ZN(n19540) );
  OAI211_X1 U21670 ( .C1(n19564), .C2(n19657), .A(n19541), .B(n19540), .ZN(
        P2_U3154) );
  AOI22_X1 U21671 ( .A1(n19666), .A2(n19570), .B1(n19568), .B2(n19665), .ZN(
        n19543) );
  AOI22_X1 U21672 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19668), .B1(
        n19667), .B2(n19571), .ZN(n19542) );
  OAI211_X1 U21673 ( .C1(n19567), .C2(n19676), .A(n19543), .B(n19542), .ZN(
        P2_U3146) );
  AOI22_X1 U21674 ( .A1(n19672), .A2(n19570), .B1(n19568), .B2(n19671), .ZN(
        n19545) );
  AOI22_X1 U21675 ( .A1(n19569), .A2(n19678), .B1(n19673), .B2(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n19544) );
  OAI211_X1 U21676 ( .C1(n19564), .C2(n19676), .A(n19545), .B(n19544), .ZN(
        P2_U3138) );
  AOI22_X1 U21677 ( .A1(n19569), .A2(n19597), .B1(n19568), .B2(n19677), .ZN(
        n19547) );
  AOI22_X1 U21678 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19680), .B1(
        n19570), .B2(n19679), .ZN(n19546) );
  OAI211_X1 U21679 ( .C1(n19564), .C2(n19600), .A(n19547), .B(n19546), .ZN(
        P2_U3130) );
  AOI22_X1 U21680 ( .A1(n19569), .A2(n19690), .B1(n19568), .B2(n19683), .ZN(
        n19549) );
  AOI22_X1 U21681 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19685), .B1(
        n19570), .B2(n19684), .ZN(n19548) );
  OAI211_X1 U21682 ( .C1(n19564), .C2(n19688), .A(n19549), .B(n19548), .ZN(
        P2_U3122) );
  AOI22_X1 U21683 ( .A1(n19571), .A2(n19690), .B1(n19568), .B2(n19689), .ZN(
        n19551) );
  AOI22_X1 U21684 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19692), .B1(
        n19691), .B2(n19570), .ZN(n19550) );
  OAI211_X1 U21685 ( .C1(n19567), .C2(n19695), .A(n19551), .B(n19550), .ZN(
        P2_U3114) );
  AOI22_X1 U21686 ( .A1(n19697), .A2(n19570), .B1(n19696), .B2(n19568), .ZN(
        n19553) );
  AOI22_X1 U21687 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19571), .ZN(n19552) );
  OAI211_X1 U21688 ( .C1(n19567), .C2(n19708), .A(n19553), .B(n19552), .ZN(
        P2_U3106) );
  AOI22_X1 U21689 ( .A1(n19703), .A2(n19570), .B1(n19568), .B2(n19702), .ZN(
        n19555) );
  AOI22_X1 U21690 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19569), .ZN(n19554) );
  OAI211_X1 U21691 ( .C1(n19564), .C2(n19708), .A(n19555), .B(n19554), .ZN(
        P2_U3098) );
  AOI22_X1 U21692 ( .A1(n19569), .A2(n19716), .B1(n19568), .B2(n19709), .ZN(
        n19557) );
  AOI22_X1 U21693 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19711), .B1(
        n19570), .B2(n19710), .ZN(n19556) );
  OAI211_X1 U21694 ( .C1(n19564), .C2(n19714), .A(n19557), .B(n19556), .ZN(
        P2_U3090) );
  AOI22_X1 U21695 ( .A1(n19571), .A2(n19716), .B1(n19568), .B2(n19715), .ZN(
        n19559) );
  AOI22_X1 U21696 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19718), .B1(
        n19570), .B2(n19717), .ZN(n19558) );
  OAI211_X1 U21697 ( .C1(n19567), .C2(n19721), .A(n19559), .B(n19558), .ZN(
        P2_U3082) );
  AOI22_X1 U21698 ( .A1(n19571), .A2(n19723), .B1(n19722), .B2(n19568), .ZN(
        n19561) );
  AOI22_X1 U21699 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19725), .B1(
        n19570), .B2(n19724), .ZN(n19560) );
  OAI211_X1 U21700 ( .C1(n19567), .C2(n19733), .A(n19561), .B(n19560), .ZN(
        P2_U3074) );
  AOI22_X1 U21701 ( .A1(n19729), .A2(n19570), .B1(n19568), .B2(n19728), .ZN(
        n19563) );
  AOI22_X1 U21702 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19730), .B1(
        n19737), .B2(n19569), .ZN(n19562) );
  OAI211_X1 U21703 ( .C1(n19564), .C2(n19733), .A(n19563), .B(n19562), .ZN(
        P2_U3066) );
  AOI22_X1 U21704 ( .A1(n19736), .A2(n19570), .B1(n19568), .B2(n19735), .ZN(
        n19566) );
  AOI22_X1 U21705 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19738), .B1(
        n19737), .B2(n19571), .ZN(n19565) );
  OAI211_X1 U21706 ( .C1(n19567), .C2(n19741), .A(n19566), .B(n19565), .ZN(
        P2_U3058) );
  AOI22_X1 U21707 ( .A1(n19569), .A2(n19745), .B1(n19568), .B2(n19743), .ZN(
        n19573) );
  AOI22_X1 U21708 ( .A1(n19750), .A2(n19571), .B1(n19748), .B2(n19570), .ZN(
        n19572) );
  OAI211_X1 U21709 ( .C1(n19754), .C2(n19574), .A(n19573), .B(n19572), .ZN(
        P2_U3050) );
  AOI22_X1 U21710 ( .A1(n19633), .A2(n19575), .B1(n19627), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19582) );
  AOI21_X1 U21711 ( .B1(n19578), .B2(n19577), .A(n19576), .ZN(n19580) );
  OR2_X1 U21712 ( .A1(n19580), .A2(n19579), .ZN(n19581) );
  OAI211_X1 U21713 ( .C1(n19584), .C2(n19583), .A(n19582), .B(n19581), .ZN(
        P2_U2918) );
  AOI22_X1 U21714 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19646), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19645), .ZN(n19620) );
  NOR2_X2 U21715 ( .A1(n19584), .A2(n19639), .ZN(n19622) );
  AOI22_X1 U21716 ( .A1(n19644), .A2(n19622), .B1(n19643), .B2(n19586), .ZN(
        n19588) );
  AOI22_X1 U21717 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n19646), .B1(
        BUF1_REG_17__SCAN_IN), .B2(n19645), .ZN(n19617) );
  INV_X1 U21718 ( .A(n19617), .ZN(n19623) );
  AOI22_X1 U21719 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19647), .B1(
        n19745), .B2(n19623), .ZN(n19587) );
  OAI211_X1 U21720 ( .C1(n19620), .C2(n19650), .A(n19588), .B(n19587), .ZN(
        P2_U3169) );
  AOI22_X1 U21721 ( .A1(n19621), .A2(n19660), .B1(n19586), .B2(n19651), .ZN(
        n19590) );
  AOI22_X1 U21722 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19654), .B1(
        n19622), .B2(n19653), .ZN(n19589) );
  OAI211_X1 U21723 ( .C1(n19617), .C2(n19650), .A(n19590), .B(n19589), .ZN(
        P2_U3161) );
  AOI22_X1 U21724 ( .A1(n19659), .A2(n19622), .B1(n19586), .B2(n19658), .ZN(
        n19592) );
  AOI22_X1 U21725 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19661), .B1(
        n19667), .B2(n19621), .ZN(n19591) );
  OAI211_X1 U21726 ( .C1(n19617), .C2(n19657), .A(n19592), .B(n19591), .ZN(
        P2_U3153) );
  AOI22_X1 U21727 ( .A1(n19666), .A2(n19622), .B1(n19586), .B2(n19665), .ZN(
        n19594) );
  AOI22_X1 U21728 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19668), .B1(
        n19667), .B2(n19623), .ZN(n19593) );
  OAI211_X1 U21729 ( .C1(n19620), .C2(n19676), .A(n19594), .B(n19593), .ZN(
        P2_U3145) );
  AOI22_X1 U21730 ( .A1(n19672), .A2(n19622), .B1(n19586), .B2(n19671), .ZN(
        n19596) );
  AOI22_X1 U21731 ( .A1(n19621), .A2(n19678), .B1(n19673), .B2(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n19595) );
  OAI211_X1 U21732 ( .C1(n19617), .C2(n19676), .A(n19596), .B(n19595), .ZN(
        P2_U3137) );
  AOI22_X1 U21733 ( .A1(n19621), .A2(n19597), .B1(n19586), .B2(n19677), .ZN(
        n19599) );
  AOI22_X1 U21734 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19680), .B1(
        n19622), .B2(n19679), .ZN(n19598) );
  OAI211_X1 U21735 ( .C1(n19617), .C2(n19600), .A(n19599), .B(n19598), .ZN(
        P2_U3129) );
  AOI22_X1 U21736 ( .A1(n19621), .A2(n19690), .B1(n19586), .B2(n19683), .ZN(
        n19602) );
  AOI22_X1 U21737 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19685), .B1(
        n19622), .B2(n19684), .ZN(n19601) );
  OAI211_X1 U21738 ( .C1(n19617), .C2(n19688), .A(n19602), .B(n19601), .ZN(
        P2_U3121) );
  AOI22_X1 U21739 ( .A1(n19623), .A2(n19690), .B1(n19586), .B2(n19689), .ZN(
        n19604) );
  AOI22_X1 U21740 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19692), .B1(
        n19691), .B2(n19622), .ZN(n19603) );
  OAI211_X1 U21741 ( .C1(n19620), .C2(n19695), .A(n19604), .B(n19603), .ZN(
        P2_U3113) );
  AOI22_X1 U21742 ( .A1(n19697), .A2(n19622), .B1(n19696), .B2(n19586), .ZN(
        n19606) );
  AOI22_X1 U21743 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19623), .ZN(n19605) );
  OAI211_X1 U21744 ( .C1(n19620), .C2(n19708), .A(n19606), .B(n19605), .ZN(
        P2_U3105) );
  AOI22_X1 U21745 ( .A1(n19703), .A2(n19622), .B1(n19586), .B2(n19702), .ZN(
        n19608) );
  AOI22_X1 U21746 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19621), .ZN(n19607) );
  OAI211_X1 U21747 ( .C1(n19617), .C2(n19708), .A(n19608), .B(n19607), .ZN(
        P2_U3097) );
  AOI22_X1 U21748 ( .A1(n19621), .A2(n19716), .B1(n19586), .B2(n19709), .ZN(
        n19610) );
  AOI22_X1 U21749 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19711), .B1(
        n19622), .B2(n19710), .ZN(n19609) );
  OAI211_X1 U21750 ( .C1(n19617), .C2(n19714), .A(n19610), .B(n19609), .ZN(
        P2_U3089) );
  AOI22_X1 U21751 ( .A1(n19623), .A2(n19716), .B1(n19586), .B2(n19715), .ZN(
        n19612) );
  AOI22_X1 U21752 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19718), .B1(
        n19622), .B2(n19717), .ZN(n19611) );
  OAI211_X1 U21753 ( .C1(n19620), .C2(n19721), .A(n19612), .B(n19611), .ZN(
        P2_U3081) );
  AOI22_X1 U21754 ( .A1(n19623), .A2(n19723), .B1(n19722), .B2(n19586), .ZN(
        n19614) );
  AOI22_X1 U21755 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19725), .B1(
        n19622), .B2(n19724), .ZN(n19613) );
  OAI211_X1 U21756 ( .C1(n19620), .C2(n19733), .A(n19614), .B(n19613), .ZN(
        P2_U3073) );
  AOI22_X1 U21757 ( .A1(n19729), .A2(n19622), .B1(n19586), .B2(n19728), .ZN(
        n19616) );
  AOI22_X1 U21758 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19730), .B1(
        n19737), .B2(n19621), .ZN(n19615) );
  OAI211_X1 U21759 ( .C1(n19617), .C2(n19733), .A(n19616), .B(n19615), .ZN(
        P2_U3065) );
  AOI22_X1 U21760 ( .A1(n19736), .A2(n19622), .B1(n19586), .B2(n19735), .ZN(
        n19619) );
  AOI22_X1 U21761 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19738), .B1(
        n19737), .B2(n19623), .ZN(n19618) );
  OAI211_X1 U21762 ( .C1(n19620), .C2(n19741), .A(n19619), .B(n19618), .ZN(
        P2_U3057) );
  AOI22_X1 U21763 ( .A1(n19621), .A2(n19745), .B1(n19586), .B2(n19743), .ZN(
        n19625) );
  AOI22_X1 U21764 ( .A1(n19750), .A2(n19623), .B1(n19748), .B2(n19622), .ZN(
        n19624) );
  OAI211_X1 U21765 ( .C1(n19754), .C2(n19626), .A(n19625), .B(n19624), .ZN(
        P2_U3049) );
  AOI22_X1 U21766 ( .A1(n19629), .A2(n19628), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19627), .ZN(n19638) );
  AOI22_X1 U21767 ( .A1(n19631), .A2(BUF1_REG_16__SCAN_IN), .B1(n19630), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19637) );
  AOI22_X1 U21768 ( .A1(n19635), .A2(n19634), .B1(n19633), .B2(n19632), .ZN(
        n19636) );
  NAND3_X1 U21769 ( .A1(n19638), .A2(n19637), .A3(n19636), .ZN(P2_U2903) );
  AOI22_X1 U21770 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19646), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19645), .ZN(n19742) );
  NOR2_X2 U21771 ( .A1(n19640), .A2(n19639), .ZN(n19747) );
  NOR2_X2 U21772 ( .A1(n19642), .A2(n19641), .ZN(n19744) );
  AOI22_X1 U21773 ( .A1(n19644), .A2(n19747), .B1(n19643), .B2(n19744), .ZN(
        n19649) );
  AOI22_X1 U21774 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n19646), .B1(
        BUF1_REG_16__SCAN_IN), .B2(n19645), .ZN(n19734) );
  AOI22_X1 U21775 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19647), .B1(
        n19745), .B2(n19749), .ZN(n19648) );
  OAI211_X1 U21776 ( .C1(n19742), .C2(n19650), .A(n19649), .B(n19648), .ZN(
        P2_U3168) );
  AOI22_X1 U21777 ( .A1(n19749), .A2(n19652), .B1(n19744), .B2(n19651), .ZN(
        n19656) );
  AOI22_X1 U21778 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19654), .B1(
        n19747), .B2(n19653), .ZN(n19655) );
  OAI211_X1 U21779 ( .C1(n19742), .C2(n19657), .A(n19656), .B(n19655), .ZN(
        P2_U3160) );
  AOI22_X1 U21780 ( .A1(n19659), .A2(n19747), .B1(n19744), .B2(n19658), .ZN(
        n19663) );
  AOI22_X1 U21781 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19661), .B1(
        n19660), .B2(n19749), .ZN(n19662) );
  OAI211_X1 U21782 ( .C1(n19742), .C2(n19664), .A(n19663), .B(n19662), .ZN(
        P2_U3152) );
  AOI22_X1 U21783 ( .A1(n19666), .A2(n19747), .B1(n19744), .B2(n19665), .ZN(
        n19670) );
  AOI22_X1 U21784 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19668), .B1(
        n19667), .B2(n19749), .ZN(n19669) );
  OAI211_X1 U21785 ( .C1(n19742), .C2(n19676), .A(n19670), .B(n19669), .ZN(
        P2_U3144) );
  AOI22_X1 U21786 ( .A1(n19672), .A2(n19747), .B1(n19744), .B2(n19671), .ZN(
        n19675) );
  INV_X1 U21787 ( .A(n19742), .ZN(n19746) );
  AOI22_X1 U21788 ( .A1(n19746), .A2(n19678), .B1(n19673), .B2(
        P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n19674) );
  OAI211_X1 U21789 ( .C1(n19734), .C2(n19676), .A(n19675), .B(n19674), .ZN(
        P2_U3136) );
  AOI22_X1 U21790 ( .A1(n19749), .A2(n19678), .B1(n19744), .B2(n19677), .ZN(
        n19682) );
  AOI22_X1 U21791 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19680), .B1(
        n19747), .B2(n19679), .ZN(n19681) );
  OAI211_X1 U21792 ( .C1(n19742), .C2(n19688), .A(n19682), .B(n19681), .ZN(
        P2_U3128) );
  AOI22_X1 U21793 ( .A1(n19746), .A2(n19690), .B1(n19744), .B2(n19683), .ZN(
        n19687) );
  AOI22_X1 U21794 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19685), .B1(
        n19747), .B2(n19684), .ZN(n19686) );
  OAI211_X1 U21795 ( .C1(n19734), .C2(n19688), .A(n19687), .B(n19686), .ZN(
        P2_U3120) );
  AOI22_X1 U21796 ( .A1(n19749), .A2(n19690), .B1(n19744), .B2(n19689), .ZN(
        n19694) );
  AOI22_X1 U21797 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19692), .B1(
        n19691), .B2(n19747), .ZN(n19693) );
  OAI211_X1 U21798 ( .C1(n19742), .C2(n19695), .A(n19694), .B(n19693), .ZN(
        P2_U3112) );
  AOI22_X1 U21799 ( .A1(n19697), .A2(n19747), .B1(n19696), .B2(n19744), .ZN(
        n19701) );
  AOI22_X1 U21800 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19699), .B1(
        n19698), .B2(n19749), .ZN(n19700) );
  OAI211_X1 U21801 ( .C1(n19742), .C2(n19708), .A(n19701), .B(n19700), .ZN(
        P2_U3104) );
  AOI22_X1 U21802 ( .A1(n19703), .A2(n19747), .B1(n19744), .B2(n19702), .ZN(
        n19707) );
  AOI22_X1 U21803 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19705), .B1(
        n19704), .B2(n19746), .ZN(n19706) );
  OAI211_X1 U21804 ( .C1(n19734), .C2(n19708), .A(n19707), .B(n19706), .ZN(
        P2_U3096) );
  AOI22_X1 U21805 ( .A1(n19746), .A2(n19716), .B1(n19744), .B2(n19709), .ZN(
        n19713) );
  AOI22_X1 U21806 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19711), .B1(
        n19747), .B2(n19710), .ZN(n19712) );
  OAI211_X1 U21807 ( .C1(n19734), .C2(n19714), .A(n19713), .B(n19712), .ZN(
        P2_U3088) );
  AOI22_X1 U21808 ( .A1(n19749), .A2(n19716), .B1(n19744), .B2(n19715), .ZN(
        n19720) );
  AOI22_X1 U21809 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19718), .B1(
        n19747), .B2(n19717), .ZN(n19719) );
  OAI211_X1 U21810 ( .C1(n19742), .C2(n19721), .A(n19720), .B(n19719), .ZN(
        P2_U3080) );
  AOI22_X1 U21811 ( .A1(n19749), .A2(n19723), .B1(n19722), .B2(n19744), .ZN(
        n19727) );
  AOI22_X1 U21812 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19725), .B1(
        n19747), .B2(n19724), .ZN(n19726) );
  OAI211_X1 U21813 ( .C1(n19742), .C2(n19733), .A(n19727), .B(n19726), .ZN(
        P2_U3072) );
  AOI22_X1 U21814 ( .A1(n19729), .A2(n19747), .B1(n19744), .B2(n19728), .ZN(
        n19732) );
  AOI22_X1 U21815 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19730), .B1(
        n19737), .B2(n19746), .ZN(n19731) );
  OAI211_X1 U21816 ( .C1(n19734), .C2(n19733), .A(n19732), .B(n19731), .ZN(
        P2_U3064) );
  AOI22_X1 U21817 ( .A1(n19736), .A2(n19747), .B1(n19744), .B2(n19735), .ZN(
        n19740) );
  AOI22_X1 U21818 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19738), .B1(
        n19737), .B2(n19749), .ZN(n19739) );
  OAI211_X1 U21819 ( .C1(n19742), .C2(n19741), .A(n19740), .B(n19739), .ZN(
        P2_U3056) );
  AOI22_X1 U21820 ( .A1(n19746), .A2(n19745), .B1(n19744), .B2(n19743), .ZN(
        n19752) );
  AOI22_X1 U21821 ( .A1(n19750), .A2(n19749), .B1(n19748), .B2(n19747), .ZN(
        n19751) );
  OAI211_X1 U21822 ( .C1(n19754), .C2(n19753), .A(n19752), .B(n19751), .ZN(
        P2_U3048) );
  INV_X1 U21823 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20092) );
  INV_X1 U21824 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20094) );
  INV_X1 U21825 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n19755) );
  AOI222_X1 U21826 ( .A1(n20092), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n20094), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n19755), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n19756) );
  INV_X1 U21827 ( .A(n19816), .ZN(n19805) );
  INV_X1 U21828 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19758) );
  AOI22_X1 U21829 ( .A1(n19805), .A2(n19758), .B1(n19757), .B2(n19816), .ZN(
        U376) );
  INV_X1 U21830 ( .A(n19816), .ZN(n19819) );
  INV_X1 U21831 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19760) );
  AOI22_X1 U21832 ( .A1(n19819), .A2(n19760), .B1(n19759), .B2(n19816), .ZN(
        U365) );
  INV_X1 U21833 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19762) );
  AOI22_X1 U21834 ( .A1(n19805), .A2(n19762), .B1(n19761), .B2(n19816), .ZN(
        U354) );
  INV_X1 U21835 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19764) );
  AOI22_X1 U21836 ( .A1(n19805), .A2(n19764), .B1(n19763), .B2(n19816), .ZN(
        U353) );
  INV_X1 U21837 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19766) );
  AOI22_X1 U21838 ( .A1(n19805), .A2(n19766), .B1(n19765), .B2(n19816), .ZN(
        U352) );
  INV_X1 U21839 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19768) );
  AOI22_X1 U21840 ( .A1(n19805), .A2(n19768), .B1(n19767), .B2(n19816), .ZN(
        U351) );
  INV_X1 U21841 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19770) );
  AOI22_X1 U21842 ( .A1(n19819), .A2(n19770), .B1(n19769), .B2(n19816), .ZN(
        U350) );
  INV_X1 U21843 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19772) );
  AOI22_X1 U21844 ( .A1(n19805), .A2(n19772), .B1(n19771), .B2(n19816), .ZN(
        U349) );
  INV_X1 U21845 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19774) );
  AOI22_X1 U21846 ( .A1(n19805), .A2(n19774), .B1(n19773), .B2(n19816), .ZN(
        U348) );
  INV_X1 U21847 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19776) );
  AOI22_X1 U21848 ( .A1(n19805), .A2(n19776), .B1(n19775), .B2(n19816), .ZN(
        U347) );
  INV_X1 U21849 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19778) );
  AOI22_X1 U21850 ( .A1(n19805), .A2(n19778), .B1(n19777), .B2(n19816), .ZN(
        U375) );
  INV_X1 U21851 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19780) );
  AOI22_X1 U21852 ( .A1(n19805), .A2(n19780), .B1(n19779), .B2(n19816), .ZN(
        U374) );
  INV_X1 U21853 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19782) );
  AOI22_X1 U21854 ( .A1(n19805), .A2(n19782), .B1(n19781), .B2(n19816), .ZN(
        U373) );
  INV_X1 U21855 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19784) );
  AOI22_X1 U21856 ( .A1(n19805), .A2(n19784), .B1(n19783), .B2(n19816), .ZN(
        U372) );
  INV_X1 U21857 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19786) );
  AOI22_X1 U21858 ( .A1(n19805), .A2(n19786), .B1(n19785), .B2(n19816), .ZN(
        U371) );
  INV_X1 U21859 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U21860 ( .A1(n19805), .A2(n19788), .B1(n19787), .B2(n19816), .ZN(
        U370) );
  INV_X1 U21861 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19790) );
  AOI22_X1 U21862 ( .A1(n19805), .A2(n19790), .B1(n19789), .B2(n19816), .ZN(
        U369) );
  INV_X1 U21863 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19792) );
  AOI22_X1 U21864 ( .A1(n19805), .A2(n19792), .B1(n19791), .B2(n19816), .ZN(
        U368) );
  INV_X1 U21865 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19794) );
  AOI22_X1 U21866 ( .A1(n19805), .A2(n19794), .B1(n19793), .B2(n19816), .ZN(
        U367) );
  INV_X1 U21867 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19796) );
  AOI22_X1 U21868 ( .A1(n19805), .A2(n19796), .B1(n19795), .B2(n19816), .ZN(
        U366) );
  INV_X1 U21869 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19798) );
  AOI22_X1 U21870 ( .A1(n19805), .A2(n19798), .B1(n19797), .B2(n19816), .ZN(
        U364) );
  INV_X1 U21871 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19800) );
  AOI22_X1 U21872 ( .A1(n19805), .A2(n19800), .B1(n19799), .B2(n19816), .ZN(
        U363) );
  INV_X1 U21873 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19802) );
  AOI22_X1 U21874 ( .A1(n19805), .A2(n19802), .B1(n19801), .B2(n19816), .ZN(
        U362) );
  INV_X1 U21875 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19804) );
  AOI22_X1 U21876 ( .A1(n19805), .A2(n19804), .B1(n19803), .B2(n19816), .ZN(
        U361) );
  INV_X1 U21877 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19807) );
  AOI22_X1 U21878 ( .A1(n19819), .A2(n19807), .B1(n19806), .B2(n19816), .ZN(
        U360) );
  INV_X1 U21879 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19809) );
  AOI22_X1 U21880 ( .A1(n19819), .A2(n19809), .B1(n19808), .B2(n19816), .ZN(
        U359) );
  INV_X1 U21881 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19811) );
  AOI22_X1 U21882 ( .A1(n19819), .A2(n19811), .B1(n19810), .B2(n19816), .ZN(
        U358) );
  INV_X1 U21883 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19813) );
  AOI22_X1 U21884 ( .A1(n19819), .A2(n19813), .B1(n19812), .B2(n19816), .ZN(
        U357) );
  INV_X1 U21885 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19815) );
  AOI22_X1 U21886 ( .A1(n19819), .A2(n19815), .B1(n19814), .B2(n19816), .ZN(
        U356) );
  AOI22_X1 U21887 ( .A1(n19819), .A2(n19818), .B1(n19817), .B2(n19816), .ZN(
        U355) );
  AOI22_X1 U21888 ( .A1(n21278), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19821) );
  OAI21_X1 U21889 ( .B1(n19822), .B2(n19843), .A(n19821), .ZN(P1_U2936) );
  AOI22_X1 U21890 ( .A1(n21278), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19823) );
  OAI21_X1 U21891 ( .B1(n19824), .B2(n19843), .A(n19823), .ZN(P1_U2935) );
  AOI22_X1 U21892 ( .A1(n21278), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19825) );
  OAI21_X1 U21893 ( .B1(n19826), .B2(n19843), .A(n19825), .ZN(P1_U2934) );
  AOI22_X1 U21894 ( .A1(n21278), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19827) );
  OAI21_X1 U21895 ( .B1(n19828), .B2(n19843), .A(n19827), .ZN(P1_U2933) );
  AOI22_X1 U21896 ( .A1(n21278), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19829) );
  OAI21_X1 U21897 ( .B1(n19830), .B2(n19843), .A(n19829), .ZN(P1_U2932) );
  AOI22_X1 U21898 ( .A1(n21278), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19831) );
  OAI21_X1 U21899 ( .B1(n19832), .B2(n19843), .A(n19831), .ZN(P1_U2931) );
  AOI22_X1 U21900 ( .A1(n21278), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19833) );
  OAI21_X1 U21901 ( .B1(n11934), .B2(n19843), .A(n19833), .ZN(P1_U2930) );
  AOI22_X1 U21902 ( .A1(n21278), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19834) );
  OAI21_X1 U21903 ( .B1(n11948), .B2(n19843), .A(n19834), .ZN(P1_U2929) );
  AOI22_X1 U21904 ( .A1(n21278), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19835) );
  OAI21_X1 U21905 ( .B1(n14805), .B2(n19843), .A(n19835), .ZN(P1_U2928) );
  AOI22_X1 U21906 ( .A1(n21278), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19836) );
  OAI21_X1 U21907 ( .B1(n14939), .B2(n19843), .A(n19836), .ZN(P1_U2926) );
  AOI22_X1 U21908 ( .A1(n21278), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19837) );
  OAI21_X1 U21909 ( .B1(n15168), .B2(n19843), .A(n19837), .ZN(P1_U2925) );
  INV_X1 U21910 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n21762) );
  AOI22_X1 U21911 ( .A1(n21278), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19838) );
  OAI21_X1 U21912 ( .B1(n21762), .B2(n19843), .A(n19838), .ZN(P1_U2924) );
  INV_X1 U21913 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n21769) );
  AOI22_X1 U21914 ( .A1(n21278), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19839) );
  OAI21_X1 U21915 ( .B1(n21769), .B2(n19843), .A(n19839), .ZN(P1_U2923) );
  INV_X1 U21916 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n21778) );
  AOI22_X1 U21917 ( .A1(n21278), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19840) );
  OAI21_X1 U21918 ( .B1(n21778), .B2(n19843), .A(n19840), .ZN(P1_U2922) );
  AOI22_X1 U21919 ( .A1(n21278), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n19841), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19842) );
  OAI21_X1 U21920 ( .B1(n19844), .B2(n19843), .A(n19842), .ZN(P1_U2921) );
  AND2_X1 U21921 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22279), .ZN(n19882) );
  INV_X1 U21922 ( .A(n19882), .ZN(n19893) );
  AND2_X1 U21923 ( .A1(n22279), .A2(n21690), .ZN(n19879) );
  INV_X1 U21924 ( .A(n19879), .ZN(n19890) );
  OAI222_X1 U21925 ( .A1(n19893), .A2(n14210), .B1(n19845), .B2(n22279), .C1(
        n21443), .C2(n19890), .ZN(P1_U3197) );
  INV_X1 U21926 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n19846) );
  OAI222_X1 U21927 ( .A1(n19890), .A2(n19847), .B1(n19846), .B2(n22279), .C1(
        n21443), .C2(n19893), .ZN(P1_U3198) );
  INV_X1 U21928 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n19848) );
  OAI222_X1 U21929 ( .A1(n19890), .A2(n21460), .B1(n19848), .B2(n22279), .C1(
        n19847), .C2(n19893), .ZN(P1_U3199) );
  AOI22_X1 U21930 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19879), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n22276), .ZN(n19849) );
  OAI21_X1 U21931 ( .B1(n21460), .B2(n19893), .A(n19849), .ZN(P1_U3200) );
  AOI22_X1 U21932 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19882), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n22276), .ZN(n19850) );
  OAI21_X1 U21933 ( .B1(n19852), .B2(n19890), .A(n19850), .ZN(P1_U3201) );
  AOI22_X1 U21934 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19879), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n22276), .ZN(n19851) );
  OAI21_X1 U21935 ( .B1(n19852), .B2(n19893), .A(n19851), .ZN(P1_U3202) );
  AOI22_X1 U21936 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19882), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n22276), .ZN(n19853) );
  OAI21_X1 U21937 ( .B1(n19855), .B2(n19890), .A(n19853), .ZN(P1_U3203) );
  AOI22_X1 U21938 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19879), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n22276), .ZN(n19854) );
  OAI21_X1 U21939 ( .B1(n19855), .B2(n19893), .A(n19854), .ZN(P1_U3204) );
  AOI22_X1 U21940 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19882), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n22276), .ZN(n19856) );
  OAI21_X1 U21941 ( .B1(n19857), .B2(n19890), .A(n19856), .ZN(P1_U3205) );
  INV_X1 U21942 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n19858) );
  OAI222_X1 U21943 ( .A1(n19890), .A2(n19969), .B1(n19858), .B2(n22279), .C1(
        n19857), .C2(n19893), .ZN(P1_U3206) );
  INV_X1 U21944 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21516) );
  INV_X1 U21945 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n19859) );
  OAI222_X1 U21946 ( .A1(n19890), .A2(n21516), .B1(n19859), .B2(n22279), .C1(
        n19969), .C2(n19893), .ZN(P1_U3207) );
  INV_X1 U21947 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n19860) );
  OAI222_X1 U21948 ( .A1(n19890), .A2(n19861), .B1(n19860), .B2(n22279), .C1(
        n21516), .C2(n19893), .ZN(P1_U3208) );
  INV_X1 U21949 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n19863) );
  INV_X1 U21950 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n19862) );
  OAI222_X1 U21951 ( .A1(n19890), .A2(n19863), .B1(n19862), .B2(n22279), .C1(
        n19861), .C2(n19893), .ZN(P1_U3209) );
  INV_X1 U21952 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n19864) );
  OAI222_X1 U21953 ( .A1(n19890), .A2(n19866), .B1(n19864), .B2(n22279), .C1(
        n19863), .C2(n19893), .ZN(P1_U3210) );
  AOI22_X1 U21954 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n19879), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n22276), .ZN(n19865) );
  OAI21_X1 U21955 ( .B1(n19866), .B2(n19893), .A(n19865), .ZN(P1_U3211) );
  AOI22_X1 U21956 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n19882), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n22276), .ZN(n19867) );
  OAI21_X1 U21957 ( .B1(n21539), .B2(n19890), .A(n19867), .ZN(P1_U3212) );
  AOI22_X1 U21958 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n19879), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n22276), .ZN(n19868) );
  OAI21_X1 U21959 ( .B1(n21539), .B2(n19893), .A(n19868), .ZN(P1_U3213) );
  AOI22_X1 U21960 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n19882), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n22276), .ZN(n19869) );
  OAI21_X1 U21961 ( .B1(n19870), .B2(n19890), .A(n19869), .ZN(P1_U3214) );
  INV_X1 U21962 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n19871) );
  OAI222_X1 U21963 ( .A1(n19890), .A2(n19872), .B1(n19871), .B2(n22279), .C1(
        n19870), .C2(n19893), .ZN(P1_U3215) );
  INV_X1 U21964 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n19873) );
  OAI222_X1 U21965 ( .A1(n19890), .A2(n21592), .B1(n19873), .B2(n22279), .C1(
        n19872), .C2(n19893), .ZN(P1_U3216) );
  INV_X1 U21966 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21587) );
  INV_X1 U21967 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n19874) );
  OAI222_X1 U21968 ( .A1(n19890), .A2(n21587), .B1(n19874), .B2(n22279), .C1(
        n21592), .C2(n19893), .ZN(P1_U3217) );
  INV_X1 U21969 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n19875) );
  OAI222_X1 U21970 ( .A1(n19890), .A2(n21600), .B1(n19875), .B2(n22279), .C1(
        n21587), .C2(n19893), .ZN(P1_U3218) );
  INV_X1 U21971 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n19876) );
  OAI222_X1 U21972 ( .A1(n19890), .A2(n19877), .B1(n19876), .B2(n22279), .C1(
        n21600), .C2(n19893), .ZN(P1_U3219) );
  INV_X1 U21973 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n19878) );
  OAI222_X1 U21974 ( .A1(n19890), .A2(n19881), .B1(n19878), .B2(n22279), .C1(
        n19877), .C2(n19893), .ZN(P1_U3220) );
  AOI22_X1 U21975 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n19879), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n22276), .ZN(n19880) );
  OAI21_X1 U21976 ( .B1(n19881), .B2(n19893), .A(n19880), .ZN(P1_U3221) );
  AOI22_X1 U21977 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n19882), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n22276), .ZN(n19883) );
  OAI21_X1 U21978 ( .B1(n19884), .B2(n19890), .A(n19883), .ZN(P1_U3222) );
  INV_X1 U21979 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n19885) );
  OAI222_X1 U21980 ( .A1(n19890), .A2(n19887), .B1(n19885), .B2(n22279), .C1(
        n19884), .C2(n19893), .ZN(P1_U3223) );
  INV_X1 U21981 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n19886) );
  OAI222_X1 U21982 ( .A1(n19893), .A2(n19887), .B1(n19886), .B2(n22279), .C1(
        n19888), .C2(n19890), .ZN(P1_U3224) );
  INV_X1 U21983 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n19889) );
  OAI222_X1 U21984 ( .A1(n19890), .A2(n15807), .B1(n19889), .B2(n22279), .C1(
        n19888), .C2(n19893), .ZN(P1_U3225) );
  INV_X1 U21985 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n19892) );
  OAI222_X1 U21986 ( .A1(n19893), .A2(n15807), .B1(n19892), .B2(n22279), .C1(
        n19891), .C2(n19890), .ZN(P1_U3226) );
  INV_X1 U21987 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n19894) );
  AOI22_X1 U21988 ( .A1(n22279), .A2(n19895), .B1(n19894), .B2(n22276), .ZN(
        P1_U3458) );
  AOI221_X1 U21989 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19906) );
  NOR4_X1 U21990 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19899) );
  NOR4_X1 U21991 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19898) );
  NOR4_X1 U21992 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19897) );
  NOR4_X1 U21993 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19896) );
  NAND4_X1 U21994 ( .A1(n19899), .A2(n19898), .A3(n19897), .A4(n19896), .ZN(
        n19905) );
  NOR4_X1 U21995 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19903) );
  AOI211_X1 U21996 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19902) );
  NOR4_X1 U21997 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19901) );
  NOR4_X1 U21998 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19900) );
  NAND4_X1 U21999 ( .A1(n19903), .A2(n19902), .A3(n19901), .A4(n19900), .ZN(
        n19904) );
  NOR2_X1 U22000 ( .A1(n19905), .A2(n19904), .ZN(n19918) );
  MUX2_X1 U22001 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(n19906), .S(n19918), 
        .Z(P1_U2808) );
  INV_X1 U22002 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n19907) );
  AOI22_X1 U22003 ( .A1(n22279), .A2(n19910), .B1(n19907), .B2(n22276), .ZN(
        P1_U3459) );
  AOI21_X1 U22004 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19908) );
  OAI221_X1 U22005 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19908), .C1(n14210), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n19918), .ZN(n19909) );
  OAI21_X1 U22006 ( .B1(n19918), .B2(n19910), .A(n19909), .ZN(P1_U3481) );
  INV_X1 U22007 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n19911) );
  AOI22_X1 U22008 ( .A1(n22279), .A2(n19914), .B1(n19911), .B2(n22276), .ZN(
        P1_U3460) );
  NOR3_X1 U22009 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19912) );
  OAI21_X1 U22010 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19912), .A(n19918), .ZN(
        n19913) );
  OAI21_X1 U22011 ( .B1(n19918), .B2(n19914), .A(n19913), .ZN(P1_U2807) );
  INV_X1 U22012 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n19915) );
  AOI22_X1 U22013 ( .A1(n22279), .A2(n19917), .B1(n19915), .B2(n22276), .ZN(
        P1_U3461) );
  OAI21_X1 U22014 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n19918), .ZN(n19916) );
  OAI21_X1 U22015 ( .B1(n19918), .B2(n19917), .A(n19916), .ZN(P1_U3482) );
  INV_X1 U22016 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n19927) );
  INV_X1 U22017 ( .A(n19919), .ZN(n21520) );
  OAI21_X1 U22018 ( .B1(n19922), .B2(n19921), .A(n19920), .ZN(n19924) );
  AND2_X1 U22019 ( .A1(n19924), .A2(n19923), .ZN(n21519) );
  AOI22_X1 U22020 ( .A1(n21520), .A2(n19932), .B1(n19925), .B2(n21519), .ZN(
        n19926) );
  OAI21_X1 U22021 ( .B1(n19946), .B2(n19927), .A(n19926), .ZN(P1_U2860) );
  NOR2_X1 U22022 ( .A1(n19929), .A2(n19928), .ZN(n19930) );
  OR2_X1 U22023 ( .A1(n15671), .A2(n19930), .ZN(n21616) );
  NOR2_X1 U22024 ( .A1(n21616), .A2(n19942), .ZN(n19931) );
  AOI21_X1 U22025 ( .B1(n21619), .B2(n19932), .A(n19931), .ZN(n19933) );
  OAI21_X1 U22026 ( .B1(n19946), .B2(n21611), .A(n19933), .ZN(P1_U2848) );
  NOR2_X1 U22027 ( .A1(n15705), .A2(n19934), .ZN(n19935) );
  OR2_X1 U22028 ( .A1(n19936), .A2(n19935), .ZN(n21568) );
  OAI22_X1 U22029 ( .A1(n21569), .A2(n15726), .B1(n21568), .B2(n19942), .ZN(
        n19937) );
  INV_X1 U22030 ( .A(n19937), .ZN(n19938) );
  OAI21_X1 U22031 ( .B1(n19946), .B2(n21565), .A(n19938), .ZN(P1_U2852) );
  INV_X1 U22032 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19945) );
  INV_X1 U22033 ( .A(n19939), .ZN(n19940) );
  XNOR2_X1 U22034 ( .A(n19941), .B(n19940), .ZN(n21495) );
  OAI22_X1 U22035 ( .A1(n21500), .A2(n15726), .B1(n21495), .B2(n19942), .ZN(
        n19943) );
  INV_X1 U22036 ( .A(n19943), .ZN(n19944) );
  OAI21_X1 U22037 ( .B1(n19946), .B2(n19945), .A(n19944), .ZN(P1_U2865) );
  AOI22_X1 U22038 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20014), .B1(
        n14073), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19952) );
  OAI21_X1 U22039 ( .B1(n19949), .B2(n19948), .A(n19947), .ZN(n19950) );
  INV_X1 U22040 ( .A(n19950), .ZN(n21307) );
  AOI22_X1 U22041 ( .A1(n21307), .A2(n20020), .B1(n21463), .B2(n20021), .ZN(
        n19951) );
  OAI211_X1 U22042 ( .C1(n20024), .C2(n21466), .A(n19952), .B(n19951), .ZN(
        P1_U2995) );
  AOI22_X1 U22043 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20014), .B1(
        n14073), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n19956) );
  INV_X1 U22044 ( .A(n19953), .ZN(n21475) );
  AOI22_X1 U22045 ( .A1(n19954), .A2(n20020), .B1(n21475), .B2(n20021), .ZN(
        n19955) );
  OAI211_X1 U22046 ( .C1(n20024), .C2(n21478), .A(n19956), .B(n19955), .ZN(
        P1_U2994) );
  AOI22_X1 U22047 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20014), .B1(
        n14073), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n19962) );
  INV_X1 U22048 ( .A(n19957), .ZN(n19958) );
  AOI21_X1 U22049 ( .B1(n19960), .B2(n19959), .A(n19958), .ZN(n21318) );
  AOI22_X1 U22050 ( .A1(n21318), .A2(n20020), .B1(n20021), .B2(n21489), .ZN(
        n19961) );
  OAI211_X1 U22051 ( .C1(n20024), .C2(n21492), .A(n19962), .B(n19961), .ZN(
        P1_U2993) );
  AOI22_X1 U22052 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20014), .B1(
        n14073), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n19968) );
  OAI21_X1 U22053 ( .B1(n19965), .B2(n19964), .A(n19963), .ZN(n21328) );
  OAI22_X1 U22054 ( .A1(n21328), .A2(n21639), .B1(n19975), .B2(n21500), .ZN(
        n19966) );
  INV_X1 U22055 ( .A(n19966), .ZN(n19967) );
  OAI211_X1 U22056 ( .C1(n20024), .C2(n21505), .A(n19968), .B(n19967), .ZN(
        P1_U2992) );
  NOR2_X1 U22057 ( .A1(n21419), .A2(n19969), .ZN(n21376) );
  OAI21_X1 U22058 ( .B1(n19975), .B2(n19974), .A(n19973), .ZN(P1_U2988) );
  OAI21_X1 U22059 ( .B1(n19978), .B2(n19977), .A(n19976), .ZN(n19979) );
  INV_X1 U22060 ( .A(n19979), .ZN(n21375) );
  AOI22_X1 U22061 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20014), .B1(
        n14073), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U22062 ( .A1(n19989), .A2(n21521), .B1(n20021), .B2(n21520), .ZN(
        n19980) );
  OAI211_X1 U22063 ( .C1(n21375), .C2(n21639), .A(n19981), .B(n19980), .ZN(
        P1_U2987) );
  INV_X1 U22064 ( .A(n19982), .ZN(n19985) );
  OAI21_X1 U22065 ( .B1(n19985), .B2(n19984), .A(n19983), .ZN(n19987) );
  XNOR2_X1 U22066 ( .A(n12852), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n19986) );
  XNOR2_X1 U22067 ( .A(n19987), .B(n19986), .ZN(n21292) );
  AOI22_X1 U22068 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20014), .B1(
        n14073), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n19991) );
  INV_X1 U22069 ( .A(n19988), .ZN(n21528) );
  AOI22_X1 U22070 ( .A1(n21528), .A2(n20021), .B1(n19989), .B2(n21527), .ZN(
        n19990) );
  OAI211_X1 U22071 ( .C1(n21292), .C2(n21639), .A(n19991), .B(n19990), .ZN(
        P1_U2985) );
  AOI22_X1 U22072 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n20014), .B1(
        n14073), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n19999) );
  MUX2_X1 U22073 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n19993), .S(
        n19992), .Z(n19995) );
  NAND2_X1 U22074 ( .A1(n19995), .A2(n19994), .ZN(n19996) );
  XNOR2_X1 U22075 ( .A(n19996), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n21388) );
  AOI22_X1 U22076 ( .A1(n21388), .A2(n20020), .B1(n20021), .B2(n19997), .ZN(
        n19998) );
  OAI211_X1 U22077 ( .C1(n20024), .C2(n20000), .A(n19999), .B(n19998), .ZN(
        P1_U2983) );
  AOI22_X1 U22078 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n20014), .B1(
        n14073), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n20007) );
  INV_X1 U22079 ( .A(n20001), .ZN(n20003) );
  AOI21_X1 U22080 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n20003), .A(
        n20002), .ZN(n20004) );
  XOR2_X1 U22081 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n20004), .Z(
        n21394) );
  INV_X1 U22082 ( .A(n21569), .ZN(n20005) );
  AOI22_X1 U22083 ( .A1(n21394), .A2(n20020), .B1(n20021), .B2(n20005), .ZN(
        n20006) );
  OAI211_X1 U22084 ( .C1(n20024), .C2(n21566), .A(n20007), .B(n20006), .ZN(
        P1_U2979) );
  AOI22_X1 U22085 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20014), .B1(
        n14073), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n20012) );
  NAND2_X1 U22086 ( .A1(n20009), .A2(n20008), .ZN(n20010) );
  XNOR2_X1 U22087 ( .A(n20010), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n21399) );
  AOI22_X1 U22088 ( .A1(n21591), .A2(n20021), .B1(n20020), .B2(n21399), .ZN(
        n20011) );
  OAI211_X1 U22089 ( .C1(n20024), .C2(n20013), .A(n20012), .B(n20011), .ZN(
        P1_U2977) );
  AOI22_X1 U22090 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20014), .B1(
        n14073), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n20023) );
  OR2_X1 U22091 ( .A1(n20015), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n20017) );
  NAND3_X1 U22092 ( .A1(n20018), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n20015), .ZN(n20016) );
  OAI21_X1 U22093 ( .B1(n20018), .B2(n20017), .A(n20016), .ZN(n20019) );
  XNOR2_X1 U22094 ( .A(n20019), .B(n21429), .ZN(n21423) );
  AOI22_X1 U22095 ( .A1(n21619), .A2(n20021), .B1(n20020), .B2(n21423), .ZN(
        n20022) );
  OAI211_X1 U22096 ( .C1(n20024), .C2(n21612), .A(n20023), .B(n20022), .ZN(
        P1_U2975) );
  OAI21_X1 U22097 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21690), .A(n21696), 
        .ZN(n20025) );
  AOI22_X1 U22098 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n22279), .B1(n20026), 
        .B2(n20025), .ZN(P1_U2804) );
  INV_X2 U22099 ( .A(U212), .ZN(n20089) );
  AOI22_X1 U22100 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n20088), .ZN(n20028) );
  OAI21_X1 U22101 ( .B1(n20029), .B2(n20074), .A(n20028), .ZN(U247) );
  AOI22_X1 U22102 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n20088), .ZN(n20030) );
  OAI21_X1 U22103 ( .B1(n20031), .B2(n20074), .A(n20030), .ZN(U246) );
  AOI22_X1 U22104 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n20088), .ZN(n20032) );
  OAI21_X1 U22105 ( .B1(n20033), .B2(n20074), .A(n20032), .ZN(U245) );
  AOI22_X1 U22106 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n20088), .ZN(n20034) );
  OAI21_X1 U22107 ( .B1(n20035), .B2(n20074), .A(n20034), .ZN(U244) );
  AOI22_X1 U22108 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n20088), .ZN(n20036) );
  OAI21_X1 U22109 ( .B1(n20037), .B2(n20074), .A(n20036), .ZN(U243) );
  AOI22_X1 U22110 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n20088), .ZN(n20038) );
  OAI21_X1 U22111 ( .B1(n20039), .B2(n20074), .A(n20038), .ZN(U242) );
  AOI22_X1 U22112 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n20088), .ZN(n20040) );
  OAI21_X1 U22113 ( .B1(n20041), .B2(n20074), .A(n20040), .ZN(U241) );
  AOI22_X1 U22114 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n20088), .ZN(n20042) );
  OAI21_X1 U22115 ( .B1(n20043), .B2(n20074), .A(n20042), .ZN(U240) );
  INV_X1 U22116 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20045) );
  AOI22_X1 U22117 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n20088), .ZN(n20044) );
  OAI21_X1 U22118 ( .B1(n20045), .B2(n20074), .A(n20044), .ZN(U239) );
  INV_X1 U22119 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20047) );
  AOI22_X1 U22120 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20088), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n20089), .ZN(n20046) );
  OAI21_X1 U22121 ( .B1(n20047), .B2(n20074), .A(n20046), .ZN(U238) );
  INV_X1 U22122 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20049) );
  AOI22_X1 U22123 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n20088), .ZN(n20048) );
  OAI21_X1 U22124 ( .B1(n20049), .B2(n20074), .A(n20048), .ZN(U237) );
  INV_X1 U22125 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20051) );
  AOI22_X1 U22126 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n20088), .ZN(n20050) );
  OAI21_X1 U22127 ( .B1(n20051), .B2(n20074), .A(n20050), .ZN(U236) );
  AOI22_X1 U22128 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n20088), .ZN(n20052) );
  OAI21_X1 U22129 ( .B1(n20053), .B2(n20074), .A(n20052), .ZN(U235) );
  INV_X1 U22130 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20055) );
  AOI22_X1 U22131 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n20088), .ZN(n20054) );
  OAI21_X1 U22132 ( .B1(n20055), .B2(n20074), .A(n20054), .ZN(U234) );
  AOI22_X1 U22133 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n20088), .ZN(n20056) );
  OAI21_X1 U22134 ( .B1(n20057), .B2(n20074), .A(n20056), .ZN(U233) );
  AOI22_X1 U22135 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n20088), .ZN(n20058) );
  OAI21_X1 U22136 ( .B1(n14260), .B2(n20074), .A(n20058), .ZN(U232) );
  AOI22_X1 U22137 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20088), .ZN(n20059) );
  OAI21_X1 U22138 ( .B1(n20060), .B2(n20074), .A(n20059), .ZN(U231) );
  AOI22_X1 U22139 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n20088), .ZN(n20061) );
  OAI21_X1 U22140 ( .B1(n20062), .B2(n20074), .A(n20061), .ZN(U230) );
  AOI22_X1 U22141 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n20088), .ZN(n20063) );
  OAI21_X1 U22142 ( .B1(n20064), .B2(n20074), .A(n20063), .ZN(U229) );
  AOI22_X1 U22143 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n20088), .ZN(n20065) );
  OAI21_X1 U22144 ( .B1(n20066), .B2(n20074), .A(n20065), .ZN(U228) );
  AOI22_X1 U22145 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n20088), .ZN(n20067) );
  OAI21_X1 U22146 ( .B1(n20068), .B2(n20074), .A(n20067), .ZN(U227) );
  AOI22_X1 U22147 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n20088), .ZN(n20069) );
  OAI21_X1 U22148 ( .B1(n20070), .B2(n20074), .A(n20069), .ZN(U226) );
  AOI22_X1 U22149 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n20088), .ZN(n20071) );
  OAI21_X1 U22150 ( .B1(n20072), .B2(n20074), .A(n20071), .ZN(U225) );
  AOI22_X1 U22151 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n20088), .ZN(n20073) );
  OAI21_X1 U22152 ( .B1(n20075), .B2(n20074), .A(n20073), .ZN(U224) );
  AOI22_X1 U22153 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n20088), .ZN(n20076) );
  OAI21_X1 U22154 ( .B1(n20077), .B2(n20074), .A(n20076), .ZN(U223) );
  AOI22_X1 U22155 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n20088), .ZN(n20078) );
  OAI21_X1 U22156 ( .B1(n20079), .B2(n20074), .A(n20078), .ZN(U222) );
  AOI22_X1 U22157 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n20088), .ZN(n20080) );
  OAI21_X1 U22158 ( .B1(n20081), .B2(n20074), .A(n20080), .ZN(U221) );
  AOI22_X1 U22159 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n20088), .ZN(n20082) );
  OAI21_X1 U22160 ( .B1(n20083), .B2(n20074), .A(n20082), .ZN(U220) );
  AOI22_X1 U22161 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n20088), .ZN(n20084) );
  OAI21_X1 U22162 ( .B1(n20085), .B2(n20074), .A(n20084), .ZN(U219) );
  AOI22_X1 U22163 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n20088), .ZN(n20086) );
  OAI21_X1 U22164 ( .B1(n20087), .B2(n20074), .A(n20086), .ZN(U218) );
  AOI22_X1 U22165 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n20089), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20088), .ZN(n20090) );
  OAI21_X1 U22166 ( .B1(n20091), .B2(n20074), .A(n20090), .ZN(U217) );
  OAI222_X1 U22167 ( .A1(U214), .A2(n20094), .B1(n20074), .B2(n20093), .C1(
        U212), .C2(n20092), .ZN(U216) );
  AOI22_X1 U22168 ( .A1(n22279), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20095), 
        .B2(n22276), .ZN(P1_U3483) );
  INV_X1 U22169 ( .A(n20096), .ZN(n20099) );
  OAI21_X1 U22170 ( .B1(n21679), .B2(n20097), .A(n20157), .ZN(n20098) );
  AOI21_X1 U22171 ( .B1(n20099), .B2(n21263), .A(n20098), .ZN(n20106) );
  AOI21_X1 U22172 ( .B1(n20158), .B2(n21672), .A(n20100), .ZN(n20101) );
  OAI211_X1 U22173 ( .C1(n20102), .C2(n20101), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n21723), .ZN(n20103) );
  AOI21_X1 U22174 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20103), .A(n21255), 
        .ZN(n20105) );
  NAND2_X1 U22175 ( .A1(n20106), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20104) );
  OAI21_X1 U22176 ( .B1(n20106), .B2(n20105), .A(n20104), .ZN(P3_U3296) );
  INV_X1 U22177 ( .A(n20594), .ZN(n20107) );
  NOR2_X2 U22178 ( .A1(n21205), .A2(n20107), .ZN(n20151) );
  NOR2_X2 U22179 ( .A1(n21239), .A2(n20108), .ZN(n20143) );
  AOI22_X1 U22180 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20150), .ZN(n20109) );
  OAI21_X1 U22181 ( .B1(n20747), .B2(n20145), .A(n20109), .ZN(P3_U2768) );
  INV_X1 U22182 ( .A(n20143), .ZN(n20153) );
  AOI22_X1 U22183 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20151), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20150), .ZN(n20110) );
  OAI21_X1 U22184 ( .B1(n20654), .B2(n20153), .A(n20110), .ZN(P3_U2769) );
  AOI22_X1 U22185 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20150), .ZN(n20111) );
  OAI21_X1 U22186 ( .B1(n20130), .B2(n20145), .A(n20111), .ZN(P3_U2770) );
  AOI22_X1 U22187 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20151), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20150), .ZN(n20112) );
  OAI21_X1 U22188 ( .B1(n20676), .B2(n20153), .A(n20112), .ZN(P3_U2771) );
  AOI22_X1 U22189 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20150), .ZN(n20113) );
  OAI21_X1 U22190 ( .B1(n20643), .B2(n20145), .A(n20113), .ZN(P3_U2772) );
  AOI22_X1 U22191 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20142), .ZN(n20114) );
  OAI21_X1 U22192 ( .B1(n20637), .B2(n20145), .A(n20114), .ZN(P3_U2773) );
  AOI22_X1 U22193 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20142), .ZN(n20115) );
  OAI21_X1 U22194 ( .B1(n20674), .B2(n20145), .A(n20115), .ZN(P3_U2774) );
  AOI22_X1 U22195 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20142), .ZN(n20116) );
  OAI21_X1 U22196 ( .B1(n20629), .B2(n20145), .A(n20116), .ZN(P3_U2775) );
  AOI22_X1 U22197 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20151), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20142), .ZN(n20117) );
  OAI21_X1 U22198 ( .B1(n20118), .B2(n20153), .A(n20117), .ZN(P3_U2776) );
  AOI22_X1 U22199 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20142), .ZN(n20119) );
  OAI21_X1 U22200 ( .B1(n20623), .B2(n20145), .A(n20119), .ZN(P3_U2777) );
  AOI22_X1 U22201 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20151), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20142), .ZN(n20120) );
  OAI21_X1 U22202 ( .B1(n20121), .B2(n20153), .A(n20120), .ZN(P3_U2778) );
  AOI22_X1 U22203 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20142), .ZN(n20122) );
  OAI21_X1 U22204 ( .B1(n20614), .B2(n20145), .A(n20122), .ZN(P3_U2779) );
  AOI22_X1 U22205 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20150), .ZN(n20123) );
  OAI21_X1 U22206 ( .B1(n20609), .B2(n20145), .A(n20123), .ZN(P3_U2780) );
  AOI22_X1 U22207 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20151), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20150), .ZN(n20124) );
  OAI21_X1 U22208 ( .B1(n20711), .B2(n20153), .A(n20124), .ZN(P3_U2781) );
  AOI22_X1 U22209 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20151), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20150), .ZN(n20125) );
  OAI21_X1 U22210 ( .B1(n20126), .B2(n20153), .A(n20125), .ZN(P3_U2782) );
  AOI22_X1 U22211 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20150), .ZN(n20127) );
  OAI21_X1 U22212 ( .B1(n20747), .B2(n20145), .A(n20127), .ZN(P3_U2783) );
  AOI22_X1 U22213 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20151), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20150), .ZN(n20128) );
  OAI21_X1 U22214 ( .B1(n20769), .B2(n20153), .A(n20128), .ZN(P3_U2784) );
  AOI22_X1 U22215 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20150), .ZN(n20129) );
  OAI21_X1 U22216 ( .B1(n20130), .B2(n20145), .A(n20129), .ZN(P3_U2785) );
  AOI22_X1 U22217 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20151), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20150), .ZN(n20131) );
  OAI21_X1 U22218 ( .B1(n20132), .B2(n20153), .A(n20131), .ZN(P3_U2786) );
  AOI22_X1 U22219 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20150), .ZN(n20133) );
  OAI21_X1 U22220 ( .B1(n20643), .B2(n20145), .A(n20133), .ZN(P3_U2787) );
  AOI22_X1 U22221 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20150), .ZN(n20134) );
  OAI21_X1 U22222 ( .B1(n20637), .B2(n20145), .A(n20134), .ZN(P3_U2788) );
  AOI22_X1 U22223 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20150), .ZN(n20135) );
  OAI21_X1 U22224 ( .B1(n20674), .B2(n20145), .A(n20135), .ZN(P3_U2789) );
  AOI22_X1 U22225 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20150), .ZN(n20136) );
  OAI21_X1 U22226 ( .B1(n20629), .B2(n20145), .A(n20136), .ZN(P3_U2790) );
  AOI22_X1 U22227 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20151), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20150), .ZN(n20137) );
  OAI21_X1 U22228 ( .B1(n20762), .B2(n20153), .A(n20137), .ZN(P3_U2791) );
  AOI22_X1 U22229 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20142), .ZN(n20138) );
  OAI21_X1 U22230 ( .B1(n20623), .B2(n20145), .A(n20138), .ZN(P3_U2792) );
  AOI22_X1 U22231 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20151), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20142), .ZN(n20139) );
  OAI21_X1 U22232 ( .B1(n20140), .B2(n20153), .A(n20139), .ZN(P3_U2793) );
  AOI22_X1 U22233 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20142), .ZN(n20141) );
  OAI21_X1 U22234 ( .B1(n20614), .B2(n20145), .A(n20141), .ZN(P3_U2794) );
  AOI22_X1 U22235 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20142), .ZN(n20144) );
  OAI21_X1 U22236 ( .B1(n20609), .B2(n20145), .A(n20144), .ZN(P3_U2795) );
  AOI22_X1 U22237 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20151), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20150), .ZN(n20146) );
  OAI21_X1 U22238 ( .B1(n20147), .B2(n20153), .A(n20146), .ZN(P3_U2796) );
  AOI22_X1 U22239 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20151), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20150), .ZN(n20148) );
  OAI21_X1 U22240 ( .B1(n20149), .B2(n20153), .A(n20148), .ZN(P3_U2797) );
  AOI22_X1 U22241 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20151), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20150), .ZN(n20152) );
  OAI21_X1 U22242 ( .B1(n20756), .B2(n20153), .A(n20152), .ZN(P3_U2798) );
  NAND2_X1 U22243 ( .A1(n21243), .A2(n20154), .ZN(n21261) );
  NAND4_X1 U22244 ( .A1(n10961), .A2(n20157), .A3(n21247), .A4(n21261), .ZN(
        n20588) );
  INV_X1 U22245 ( .A(n20588), .ZN(n20505) );
  NOR2_X1 U22246 ( .A1(n20789), .A2(n10962), .ZN(n20788) );
  AOI22_X1 U22247 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20505), .B1(n20788), 
        .B2(n20584), .ZN(n20168) );
  INV_X1 U22248 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n20571) );
  OAI211_X1 U22249 ( .C1(n12661), .C2(n20155), .A(n21723), .B(n21672), .ZN(
        n21240) );
  OAI211_X2 U22250 ( .C1(n20571), .C2(n20158), .A(n21240), .B(n20159), .ZN(
        n20570) );
  AOI21_X1 U22251 ( .B1(n20396), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21247), .ZN(n20265) );
  AOI22_X1 U22252 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n20587), .B1(n20163), .B2(
        n20265), .ZN(n20167) );
  NAND2_X1 U22253 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n12661), .ZN(n20160) );
  AOI211_X4 U22254 ( .C1(n21723), .C2(n21672), .A(n20161), .B(n20160), .ZN(
        n20586) );
  AOI22_X1 U22255 ( .A1(n20586), .A2(n20162), .B1(n20502), .B2(n20859), .ZN(
        n20166) );
  NAND2_X1 U22256 ( .A1(n20396), .A2(n20560), .ZN(n20582) );
  INV_X1 U22257 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20350) );
  AOI221_X1 U22258 ( .B1(n20572), .B2(n20582), .C1(n20572), .C2(n20350), .A(
        n20163), .ZN(n20164) );
  INV_X1 U22259 ( .A(n20164), .ZN(n20165) );
  NAND4_X1 U22260 ( .A1(n20168), .A2(n20167), .A3(n20166), .A4(n20165), .ZN(
        P3_U2670) );
  AOI22_X1 U22261 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n10962), .B1(
        n20809), .B2(n20808), .ZN(n20801) );
  AOI22_X1 U22262 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n20505), .B1(n20584), 
        .B2(n20801), .ZN(n20182) );
  AOI221_X1 U22263 ( .B1(P3_REIP_REG_2__SCAN_IN), .B2(P3_REIP_REG_1__SCAN_IN), 
        .C1(n20169), .C2(n20859), .A(n20517), .ZN(n20180) );
  NOR2_X1 U22264 ( .A1(n20396), .A2(n21247), .ZN(n20353) );
  INV_X1 U22265 ( .A(n20353), .ZN(n20178) );
  NAND2_X1 U22266 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n20350), .ZN(
        n20197) );
  INV_X1 U22267 ( .A(n20197), .ZN(n20311) );
  AOI21_X1 U22268 ( .B1(n20350), .B2(n20171), .A(n11194), .ZN(n20186) );
  OAI211_X1 U22269 ( .C1(n20311), .C2(n20177), .A(n20560), .B(n20186), .ZN(
        n20176) );
  NOR3_X1 U22270 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20191) );
  INV_X1 U22271 ( .A(n20191), .ZN(n20172) );
  OAI211_X1 U22272 ( .C1(n20174), .C2(n20173), .A(n20586), .B(n20172), .ZN(
        n20175) );
  OAI211_X1 U22273 ( .C1(n20178), .C2(n20177), .A(n20176), .B(n20175), .ZN(
        n20179) );
  AOI211_X1 U22274 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20587), .A(n20180), .B(
        n20179), .ZN(n20181) );
  OAI211_X1 U22275 ( .C1(n20183), .C2(n20572), .A(n20182), .B(n20181), .ZN(
        P3_U2669) );
  NAND2_X1 U22276 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20811) );
  OAI21_X1 U22277 ( .B1(n20784), .B2(n20811), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20816) );
  NAND2_X1 U22278 ( .A1(n20816), .A2(n20184), .ZN(n20825) );
  AOI22_X1 U22279 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n20528), .B1(
        n20584), .B2(n20825), .ZN(n20195) );
  NAND3_X1 U22280 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n20210) );
  AOI21_X1 U22281 ( .B1(n20210), .B2(n20502), .A(n20505), .ZN(n20185) );
  INV_X1 U22282 ( .A(n20185), .ZN(n20204) );
  XOR2_X1 U22283 ( .A(n20187), .B(n20186), .Z(n20188) );
  OAI22_X1 U22284 ( .A1(n20570), .A2(n20190), .B1(n21247), .B2(n20188), .ZN(
        n20189) );
  AOI21_X1 U22285 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n20204), .A(n20189), .ZN(
        n20194) );
  NAND2_X1 U22286 ( .A1(n20191), .A2(n20190), .ZN(n20201) );
  OAI211_X1 U22287 ( .C1(n20191), .C2(n20190), .A(n20586), .B(n20201), .ZN(
        n20193) );
  NAND4_X1 U22288 ( .A1(n20502), .A2(P3_REIP_REG_2__SCAN_IN), .A3(
        P3_REIP_REG_1__SCAN_IN), .A4(n20879), .ZN(n20192) );
  NAND4_X1 U22289 ( .A1(n20195), .A2(n20194), .A3(n20193), .A4(n20192), .ZN(
        P3_U2668) );
  AOI22_X1 U22290 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20528), .B1(
        n20587), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n20209) );
  NAND2_X1 U22291 ( .A1(n20196), .A2(n21234), .ZN(n20200) );
  NOR2_X1 U22292 ( .A1(n20198), .A2(n20197), .ZN(n20212) );
  NOR3_X1 U22293 ( .A1(n20205), .A2(n20212), .A3(n20582), .ZN(n20199) );
  AOI211_X1 U22294 ( .C1(n20584), .C2(n20200), .A(n21189), .B(n20199), .ZN(
        n20208) );
  NOR2_X1 U22295 ( .A1(n20517), .A2(n20210), .ZN(n20203) );
  NOR2_X1 U22296 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20201), .ZN(n20218) );
  AOI211_X1 U22297 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20201), .A(n20218), .B(
        n20562), .ZN(n20202) );
  AOI221_X1 U22298 ( .B1(n20204), .B2(P3_REIP_REG_4__SCAN_IN), .C1(n20203), 
        .C2(n20211), .A(n20202), .ZN(n20207) );
  OAI211_X1 U22299 ( .C1(n20353), .C2(n11185), .A(n20205), .B(n20265), .ZN(
        n20206) );
  NAND4_X1 U22300 ( .A1(n20209), .A2(n20208), .A3(n20207), .A4(n20206), .ZN(
        P3_U2667) );
  INV_X1 U22301 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20225) );
  NOR2_X1 U22302 ( .A1(n20211), .A2(n20210), .ZN(n20216) );
  NAND2_X1 U22303 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n20216), .ZN(n20240) );
  INV_X1 U22304 ( .A(n20240), .ZN(n20235) );
  NOR2_X1 U22305 ( .A1(n20517), .A2(n20235), .ZN(n20215) );
  NOR2_X1 U22306 ( .A1(n20505), .A2(n20215), .ZN(n20251) );
  INV_X1 U22307 ( .A(n20251), .ZN(n20223) );
  NOR2_X1 U22308 ( .A1(n20212), .A2(n11194), .ZN(n20213) );
  XOR2_X1 U22309 ( .A(n20214), .B(n20213), .Z(n20217) );
  AOI22_X1 U22310 ( .A1(n20560), .A2(n20217), .B1(n20216), .B2(n20215), .ZN(
        n20220) );
  NAND2_X1 U22311 ( .A1(n20218), .A2(n20225), .ZN(n20226) );
  OAI211_X1 U22312 ( .C1(n20218), .C2(n20225), .A(n20586), .B(n20226), .ZN(
        n20219) );
  OAI211_X1 U22313 ( .C1(n20572), .C2(n20221), .A(n20220), .B(n20219), .ZN(
        n20222) );
  AOI21_X1 U22314 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n20223), .A(n20222), .ZN(
        n20224) );
  OAI211_X1 U22315 ( .C1(n20570), .C2(n20225), .A(n20224), .B(n10961), .ZN(
        P3_U2666) );
  NOR2_X1 U22316 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20226), .ZN(n20244) );
  AOI211_X1 U22317 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20226), .A(n20244), .B(
        n20562), .ZN(n20234) );
  AOI211_X1 U22318 ( .C1(n20286), .C2(n20350), .A(n20229), .B(n20582), .ZN(
        n20227) );
  NOR2_X1 U22319 ( .A1(n21189), .A2(n20227), .ZN(n20232) );
  INV_X1 U22320 ( .A(n20228), .ZN(n20230) );
  OAI211_X1 U22321 ( .C1(n20230), .C2(n11194), .A(n20229), .B(n20265), .ZN(
        n20231) );
  OAI211_X1 U22322 ( .C1(n20251), .C2(n20908), .A(n20232), .B(n20231), .ZN(
        n20233) );
  AOI211_X1 U22323 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20587), .A(n20234), .B(
        n20233), .ZN(n20236) );
  NAND3_X1 U22324 ( .A1(n20502), .A2(n20235), .A3(n20908), .ZN(n20250) );
  OAI211_X1 U22325 ( .C1(n20572), .C2(n20237), .A(n20236), .B(n20250), .ZN(
        P3_U2665) );
  AOI21_X1 U22326 ( .B1(n20286), .B2(n20350), .A(n11194), .ZN(n20239) );
  XNOR2_X1 U22327 ( .A(n20239), .B(n20238), .ZN(n20242) );
  NOR2_X1 U22328 ( .A1(n20908), .A2(n20240), .ZN(n20256) );
  NOR2_X1 U22329 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20517), .ZN(n20241) );
  AOI22_X1 U22330 ( .A1(n20560), .A2(n20242), .B1(n20256), .B2(n20241), .ZN(
        n20246) );
  INV_X1 U22331 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20243) );
  NAND2_X1 U22332 ( .A1(n20244), .A2(n20243), .ZN(n20259) );
  OAI211_X1 U22333 ( .C1(n20244), .C2(n20243), .A(n20586), .B(n20259), .ZN(
        n20245) );
  OAI211_X1 U22334 ( .C1(n20572), .C2(n20247), .A(n20246), .B(n20245), .ZN(
        n20248) );
  AOI211_X1 U22335 ( .C1(n20587), .C2(P3_EBX_REG_7__SCAN_IN), .A(n21189), .B(
        n20248), .ZN(n20249) );
  OAI221_X1 U22336 ( .B1(n20252), .B2(n20251), .C1(n20252), .C2(n20250), .A(
        n20249), .ZN(P3_U2664) );
  OAI21_X1 U22337 ( .B1(n20253), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n10956), .ZN(n20254) );
  XOR2_X1 U22338 ( .A(n20255), .B(n20254), .Z(n20264) );
  AOI21_X1 U22339 ( .B1(n20587), .B2(P3_EBX_REG_8__SCAN_IN), .A(n21189), .ZN(
        n20263) );
  NAND2_X1 U22340 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20256), .ZN(n20257) );
  NOR2_X1 U22341 ( .A1(n20258), .A2(n20257), .ZN(n20283) );
  OAI21_X1 U22342 ( .B1(n20517), .B2(n20283), .A(n20588), .ZN(n20273) );
  INV_X1 U22343 ( .A(n20273), .ZN(n20282) );
  AOI221_X1 U22344 ( .B1(n20517), .B2(n20258), .C1(n20257), .C2(n20258), .A(
        n20282), .ZN(n20261) );
  NOR2_X1 U22345 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20259), .ZN(n20275) );
  AOI211_X1 U22346 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n20259), .A(n20275), .B(
        n20562), .ZN(n20260) );
  AOI211_X1 U22347 ( .C1(n20528), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20261), .B(n20260), .ZN(n20262) );
  OAI211_X1 U22348 ( .C1(n21247), .C2(n20264), .A(n20263), .B(n20262), .ZN(
        P3_U2663) );
  INV_X1 U22349 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20274) );
  OAI21_X1 U22350 ( .B1(n20266), .B2(n20353), .A(n20265), .ZN(n20267) );
  OAI22_X1 U22351 ( .A1(n20570), .A2(n20274), .B1(n20268), .B2(n20267), .ZN(
        n20272) );
  OAI21_X1 U22352 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20289), .A(
        n20268), .ZN(n20270) );
  NAND3_X1 U22353 ( .A1(n20502), .A2(n20283), .A3(n20269), .ZN(n20281) );
  OAI211_X1 U22354 ( .C1(n20582), .C2(n20270), .A(n10961), .B(n20281), .ZN(
        n20271) );
  AOI211_X1 U22355 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n20273), .A(n20272), .B(
        n20271), .ZN(n20277) );
  NAND2_X1 U22356 ( .A1(n20275), .A2(n20274), .ZN(n20279) );
  OAI211_X1 U22357 ( .C1(n20275), .C2(n20274), .A(n20586), .B(n20279), .ZN(
        n20276) );
  OAI211_X1 U22358 ( .C1(n20572), .C2(n20278), .A(n20277), .B(n20276), .ZN(
        P3_U2662) );
  NOR2_X1 U22359 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20279), .ZN(n20305) );
  AOI211_X1 U22360 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20279), .A(n20305), .B(
        n20562), .ZN(n20280) );
  AOI21_X1 U22361 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n20587), .A(n20280), .ZN(
        n20295) );
  AOI21_X1 U22362 ( .B1(n20282), .B2(n20281), .A(n20297), .ZN(n20285) );
  NAND2_X1 U22363 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20283), .ZN(n20296) );
  NOR3_X1 U22364 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n20517), .A3(n20296), 
        .ZN(n20284) );
  AOI211_X1 U22365 ( .C1(n20528), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20285), .B(n20284), .ZN(n20294) );
  AND2_X1 U22366 ( .A1(n20350), .A2(n20286), .ZN(n20287) );
  AOI21_X1 U22367 ( .B1(n20288), .B2(n20287), .A(n11194), .ZN(n20300) );
  OR2_X1 U22368 ( .A1(n20289), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20290) );
  AOI21_X1 U22369 ( .B1(n20292), .B2(n20290), .A(n21247), .ZN(n20291) );
  OAI22_X1 U22370 ( .A1(n20292), .A2(n20300), .B1(n20353), .B2(n20291), .ZN(
        n20293) );
  NAND4_X1 U22371 ( .A1(n20295), .A2(n20294), .A3(n10961), .A4(n20293), .ZN(
        P3_U2661) );
  AOI22_X1 U22372 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n20528), .B1(
        n20587), .B2(P3_EBX_REG_11__SCAN_IN), .ZN(n20308) );
  NOR2_X1 U22373 ( .A1(n20297), .A2(n20296), .ZN(n20309) );
  NAND2_X1 U22374 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n20309), .ZN(n20460) );
  AOI21_X1 U22375 ( .B1(n20502), .B2(n20460), .A(n20505), .ZN(n20378) );
  INV_X1 U22376 ( .A(n20378), .ZN(n20339) );
  AND2_X1 U22377 ( .A1(n20502), .A2(n20309), .ZN(n20303) );
  INV_X1 U22378 ( .A(n20299), .ZN(n20301) );
  INV_X1 U22379 ( .A(n20300), .ZN(n20298) );
  AOI221_X1 U22380 ( .B1(n20301), .B2(n20300), .C1(n20299), .C2(n20298), .A(
        n21247), .ZN(n20302) );
  AOI221_X1 U22381 ( .B1(P3_REIP_REG_11__SCAN_IN), .B2(n20339), .C1(n20303), 
        .C2(n20339), .A(n20302), .ZN(n20307) );
  NAND2_X1 U22382 ( .A1(n20305), .A2(n20304), .ZN(n20310) );
  OAI211_X1 U22383 ( .C1(n20305), .C2(n20304), .A(n20586), .B(n20310), .ZN(
        n20306) );
  NAND4_X1 U22384 ( .A1(n20308), .A2(n20307), .A3(n10961), .A4(n20306), .ZN(
        P3_U2660) );
  NAND3_X1 U22385 ( .A1(n20502), .A2(P3_REIP_REG_11__SCAN_IN), .A3(n20309), 
        .ZN(n20461) );
  NOR2_X1 U22386 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20310), .ZN(n20333) );
  AOI211_X1 U22387 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20310), .A(n20333), .B(
        n20562), .ZN(n20318) );
  AOI21_X1 U22388 ( .B1(n17743), .B2(n20311), .A(n11194), .ZN(n20313) );
  INV_X1 U22389 ( .A(n20314), .ZN(n20312) );
  INV_X1 U22390 ( .A(n20313), .ZN(n20321) );
  OAI221_X1 U22391 ( .B1(n20314), .B2(n20313), .C1(n20312), .C2(n20321), .A(
        n20560), .ZN(n20315) );
  OAI211_X1 U22392 ( .C1(n20316), .C2(n20572), .A(n10961), .B(n20315), .ZN(
        n20317) );
  AOI211_X1 U22393 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20587), .A(n20318), .B(
        n20317), .ZN(n20319) );
  OAI221_X1 U22394 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n20461), .C1(n20320), 
        .C2(n20378), .A(n20319), .ZN(P3_U2659) );
  OAI21_X1 U22395 ( .B1(n20322), .B2(n11194), .A(n20321), .ZN(n20337) );
  NAND2_X1 U22396 ( .A1(n20560), .A2(n20337), .ZN(n20327) );
  INV_X1 U22397 ( .A(n20328), .ZN(n20326) );
  NOR2_X1 U22398 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21247), .ZN(
        n20324) );
  AOI21_X1 U22399 ( .B1(n20324), .B2(n20323), .A(n20353), .ZN(n20325) );
  OAI221_X1 U22400 ( .B1(n20328), .B2(n20327), .C1(n20326), .C2(n20325), .A(
        n10961), .ZN(n20332) );
  NAND2_X1 U22401 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_12__SCAN_IN), 
        .ZN(n20341) );
  OAI21_X1 U22402 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(P3_REIP_REG_12__SCAN_IN), 
        .A(n20341), .ZN(n20329) );
  OAI22_X1 U22403 ( .A1(n20378), .A2(n20330), .B1(n20461), .B2(n20329), .ZN(
        n20331) );
  AOI211_X1 U22404 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n20528), .A(
        n20332), .B(n20331), .ZN(n20335) );
  NAND2_X1 U22405 ( .A1(n20333), .A2(n20336), .ZN(n20342) );
  OAI211_X1 U22406 ( .C1(n20333), .C2(n20336), .A(n20586), .B(n20342), .ZN(
        n20334) );
  OAI211_X1 U22407 ( .C1(n20336), .C2(n20570), .A(n20335), .B(n20334), .ZN(
        P3_U2658) );
  XNOR2_X1 U22408 ( .A(n20338), .B(n20337), .ZN(n20347) );
  AOI21_X1 U22409 ( .B1(n20587), .B2(P3_EBX_REG_14__SCAN_IN), .A(n21189), .ZN(
        n20346) );
  OR2_X1 U22410 ( .A1(n20340), .A2(n20341), .ZN(n20377) );
  NAND2_X1 U22411 ( .A1(n20517), .A2(n20588), .ZN(n20585) );
  AOI21_X1 U22412 ( .B1(n20377), .B2(n20585), .A(n20339), .ZN(n20374) );
  AOI221_X1 U22413 ( .B1(n20341), .B2(n20340), .C1(n20461), .C2(n20340), .A(
        n20374), .ZN(n20344) );
  NOR2_X1 U22414 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20342), .ZN(n20359) );
  AOI211_X1 U22415 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20342), .A(n20359), .B(
        n20562), .ZN(n20343) );
  AOI211_X1 U22416 ( .C1(n20528), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20344), .B(n20343), .ZN(n20345) );
  OAI211_X1 U22417 ( .C1(n21247), .C2(n20347), .A(n20346), .B(n20345), .ZN(
        P3_U2657) );
  NOR2_X1 U22418 ( .A1(n20377), .A2(n20461), .ZN(n20375) );
  INV_X1 U22419 ( .A(n20374), .ZN(n20357) );
  INV_X1 U22420 ( .A(n20348), .ZN(n20354) );
  NAND2_X1 U22421 ( .A1(n20350), .A2(n20349), .ZN(n20351) );
  OAI21_X1 U22422 ( .B1(n20362), .B2(n20351), .A(n20396), .ZN(n20364) );
  INV_X1 U22423 ( .A(n20364), .ZN(n20366) );
  AOI21_X1 U22424 ( .B1(n20354), .B2(n20351), .A(n21247), .ZN(n20352) );
  OAI22_X1 U22425 ( .A1(n20354), .A2(n20366), .B1(n20353), .B2(n20352), .ZN(
        n20355) );
  OAI211_X1 U22426 ( .C1(n20570), .C2(n20358), .A(n10961), .B(n20355), .ZN(
        n20356) );
  AOI221_X1 U22427 ( .B1(n20375), .B2(n20376), .C1(n20357), .C2(
        P3_REIP_REG_15__SCAN_IN), .A(n20356), .ZN(n20361) );
  NAND2_X1 U22428 ( .A1(n20359), .A2(n20358), .ZN(n20363) );
  OAI211_X1 U22429 ( .C1(n20359), .C2(n20358), .A(n20586), .B(n20363), .ZN(
        n20360) );
  OAI211_X1 U22430 ( .C1(n20572), .C2(n20362), .A(n20361), .B(n20360), .ZN(
        P3_U2656) );
  NOR2_X1 U22431 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20363), .ZN(n20387) );
  AOI211_X1 U22432 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20363), .A(n20387), .B(
        n20562), .ZN(n20371) );
  INV_X1 U22433 ( .A(n20367), .ZN(n20365) );
  OAI221_X1 U22434 ( .B1(n20367), .B2(n20366), .C1(n20365), .C2(n20364), .A(
        n20560), .ZN(n20368) );
  OAI211_X1 U22435 ( .C1(n20369), .C2(n20572), .A(n10961), .B(n20368), .ZN(
        n20370) );
  AOI211_X1 U22436 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20587), .A(n20371), .B(
        n20370), .ZN(n20373) );
  OAI221_X1 U22437 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n21159), .C2(n20376), .A(n20375), .ZN(n20372) );
  OAI211_X1 U22438 ( .C1(n20374), .C2(n21159), .A(n20373), .B(n20372), .ZN(
        P3_U2655) );
  NAND3_X1 U22439 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n20375), .ZN(n20393) );
  INV_X1 U22440 ( .A(n20393), .ZN(n20386) );
  NOR4_X1 U22441 ( .A1(n20394), .A2(n20377), .A3(n21159), .A4(n20376), .ZN(
        n20446) );
  INV_X1 U22442 ( .A(n20585), .ZN(n20379) );
  OAI21_X1 U22443 ( .B1(n20446), .B2(n20379), .A(n20378), .ZN(n20417) );
  INV_X1 U22444 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n20384) );
  NAND2_X1 U22445 ( .A1(n20382), .A2(n20381), .ZN(n20395) );
  OAI211_X1 U22446 ( .C1(n20382), .C2(n20381), .A(n20560), .B(n20395), .ZN(
        n20383) );
  OAI211_X1 U22447 ( .C1(n20384), .C2(n20572), .A(n10961), .B(n20383), .ZN(
        n20385) );
  AOI221_X1 U22448 ( .B1(n20386), .B2(n20394), .C1(n20417), .C2(
        P3_REIP_REG_17__SCAN_IN), .A(n20385), .ZN(n20389) );
  NAND2_X1 U22449 ( .A1(n20387), .A2(n20390), .ZN(n20391) );
  OAI211_X1 U22450 ( .C1(n20387), .C2(n20390), .A(n20586), .B(n20391), .ZN(
        n20388) );
  OAI211_X1 U22451 ( .C1(n20390), .C2(n20570), .A(n20389), .B(n20388), .ZN(
        P3_U2654) );
  NOR2_X1 U22452 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20391), .ZN(n20408) );
  AOI211_X1 U22453 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20391), .A(n20408), .B(
        n20562), .ZN(n20392) );
  AOI211_X1 U22454 ( .C1(n20587), .C2(P3_EBX_REG_18__SCAN_IN), .A(n21189), .B(
        n20392), .ZN(n20401) );
  NOR2_X1 U22455 ( .A1(n20394), .A2(n20393), .ZN(n20440) );
  NAND2_X1 U22456 ( .A1(n20396), .A2(n20395), .ZN(n20404) );
  INV_X1 U22457 ( .A(n20404), .ZN(n20398) );
  INV_X1 U22458 ( .A(n20405), .ZN(n20397) );
  AOI221_X1 U22459 ( .B1(n20398), .B2(n20397), .C1(n20404), .C2(n20405), .A(
        n21247), .ZN(n20399) );
  AOI221_X1 U22460 ( .B1(n20440), .B2(n21143), .C1(n20417), .C2(
        P3_REIP_REG_18__SCAN_IN), .A(n20399), .ZN(n20400) );
  OAI211_X1 U22461 ( .C1(n20402), .C2(n20572), .A(n20401), .B(n20400), .ZN(
        P3_U2653) );
  INV_X1 U22462 ( .A(n20417), .ZN(n20415) );
  INV_X1 U22463 ( .A(n20403), .ZN(n20407) );
  OAI21_X1 U22464 ( .B1(n11194), .B2(n20405), .A(n20404), .ZN(n20406) );
  AOI211_X1 U22465 ( .C1(n20407), .C2(n20406), .A(n20419), .B(n21247), .ZN(
        n20412) );
  INV_X1 U22466 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20410) );
  NAND2_X1 U22467 ( .A1(n20408), .A2(n20410), .ZN(n20422) );
  OAI211_X1 U22468 ( .C1(n20408), .C2(n20410), .A(n20586), .B(n20422), .ZN(
        n20409) );
  OAI211_X1 U22469 ( .C1(n20570), .C2(n20410), .A(n10961), .B(n20409), .ZN(
        n20411) );
  AOI211_X1 U22470 ( .C1(n20528), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20412), .B(n20411), .ZN(n20414) );
  OAI221_X1 U22471 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n21143), .C2(n20416), .A(n20440), .ZN(n20413) );
  OAI211_X1 U22472 ( .C1(n20415), .C2(n20416), .A(n20414), .B(n20413), .ZN(
        P3_U2652) );
  NAND3_X1 U22473 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(n20440), .ZN(n20430) );
  NOR3_X1 U22474 ( .A1(n20429), .A2(n21143), .A3(n20416), .ZN(n20445) );
  INV_X1 U22475 ( .A(n20445), .ZN(n20418) );
  AOI21_X1 U22476 ( .B1(n20502), .B2(n20418), .A(n20417), .ZN(n20449) );
  AOI211_X1 U22477 ( .C1(n20421), .C2(n20420), .A(n20432), .B(n21247), .ZN(
        n20427) );
  NOR2_X1 U22478 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n20422), .ZN(n20435) );
  AOI211_X1 U22479 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n20422), .A(n20435), .B(
        n20562), .ZN(n20426) );
  OAI22_X1 U22480 ( .A1(n20424), .A2(n20572), .B1(n20570), .B2(n20423), .ZN(
        n20425) );
  NOR3_X1 U22481 ( .A1(n20427), .A2(n20426), .A3(n20425), .ZN(n20428) );
  OAI221_X1 U22482 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n20430), .C1(n20429), 
        .C2(n20449), .A(n20428), .ZN(P3_U2651) );
  INV_X1 U22483 ( .A(n20431), .ZN(n20434) );
  NOR2_X1 U22484 ( .A1(n20434), .A2(n20433), .ZN(n20450) );
  AOI211_X1 U22485 ( .C1(n20434), .C2(n20433), .A(n20450), .B(n21247), .ZN(
        n20439) );
  NAND2_X1 U22486 ( .A1(n20435), .A2(n20437), .ZN(n20443) );
  OAI211_X1 U22487 ( .C1(n20435), .C2(n20437), .A(n20586), .B(n20443), .ZN(
        n20436) );
  OAI21_X1 U22488 ( .B1(n20437), .B2(n20570), .A(n20436), .ZN(n20438) );
  AOI211_X1 U22489 ( .C1(n20528), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n20439), .B(n20438), .ZN(n20441) );
  NAND3_X1 U22490 ( .A1(n20445), .A2(n20440), .A3(n20442), .ZN(n20448) );
  OAI211_X1 U22491 ( .C1(n20449), .C2(n20442), .A(n20441), .B(n20448), .ZN(
        P3_U2650) );
  NOR2_X1 U22492 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n20443), .ZN(n20471) );
  AOI211_X1 U22493 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n20443), .A(n20471), .B(
        n20562), .ZN(n20444) );
  AOI21_X1 U22494 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n20587), .A(n20444), .ZN(
        n20457) );
  AND3_X1 U22495 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n20446), .A3(n20445), 
        .ZN(n20459) );
  NOR2_X1 U22496 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n20461), .ZN(n20455) );
  AOI21_X1 U22497 ( .B1(n20449), .B2(n20448), .A(n20447), .ZN(n20454) );
  NOR2_X1 U22498 ( .A1(n20450), .A2(n11194), .ZN(n20451) );
  NOR2_X1 U22499 ( .A1(n20452), .A2(n20451), .ZN(n20464) );
  AOI211_X1 U22500 ( .C1(n20452), .C2(n20451), .A(n20464), .B(n21247), .ZN(
        n20453) );
  AOI211_X1 U22501 ( .C1(n20459), .C2(n20455), .A(n20454), .B(n20453), .ZN(
        n20456) );
  OAI211_X1 U22502 ( .C1(n20458), .C2(n20572), .A(n20457), .B(n20456), .ZN(
        P3_U2649) );
  AOI22_X1 U22503 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20528), .B1(
        n20587), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n20474) );
  NAND2_X1 U22504 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n20459), .ZN(n20462) );
  NOR3_X1 U22505 ( .A1(n20468), .A2(n20460), .A3(n20462), .ZN(n20490) );
  OAI21_X1 U22506 ( .B1(n20490), .B2(n20517), .A(n20588), .ZN(n20485) );
  NOR2_X1 U22507 ( .A1(n20462), .A2(n20461), .ZN(n20469) );
  INV_X1 U22508 ( .A(n20463), .ZN(n20466) );
  NOR2_X1 U22509 ( .A1(n20464), .A2(n11194), .ZN(n20465) );
  NOR2_X1 U22510 ( .A1(n20466), .A2(n20465), .ZN(n20475) );
  AOI211_X1 U22511 ( .C1(n20466), .C2(n20465), .A(n20475), .B(n21247), .ZN(
        n20467) );
  AOI221_X1 U22512 ( .B1(n20485), .B2(P3_REIP_REG_23__SCAN_IN), .C1(n20469), 
        .C2(n20468), .A(n20467), .ZN(n20473) );
  INV_X1 U22513 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20470) );
  NAND2_X1 U22514 ( .A1(n20471), .A2(n20470), .ZN(n20478) );
  OAI211_X1 U22515 ( .C1(n20471), .C2(n20470), .A(n20586), .B(n20478), .ZN(
        n20472) );
  NAND3_X1 U22516 ( .A1(n20474), .A2(n20473), .A3(n20472), .ZN(P3_U2648) );
  INV_X1 U22517 ( .A(n20485), .ZN(n20484) );
  AOI22_X1 U22518 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20528), .B1(
        n20587), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n20483) );
  NOR2_X1 U22519 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20517), .ZN(n20481) );
  NOR2_X1 U22520 ( .A1(n20475), .A2(n11194), .ZN(n20476) );
  NOR2_X1 U22521 ( .A1(n20477), .A2(n20476), .ZN(n20487) );
  AOI211_X1 U22522 ( .C1(n20477), .C2(n20476), .A(n20487), .B(n21247), .ZN(
        n20480) );
  NOR2_X1 U22523 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n20478), .ZN(n20496) );
  AOI211_X1 U22524 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n20478), .A(n20496), .B(
        n20562), .ZN(n20479) );
  AOI211_X1 U22525 ( .C1(n20481), .C2(n20490), .A(n20480), .B(n20479), .ZN(
        n20482) );
  OAI211_X1 U22526 ( .C1(n20486), .C2(n20484), .A(n20483), .B(n20482), .ZN(
        P3_U2647) );
  AOI21_X1 U22527 ( .B1(n20502), .B2(n20486), .A(n20485), .ZN(n20499) );
  NOR2_X1 U22528 ( .A1(n20487), .A2(n11194), .ZN(n20488) );
  NOR2_X1 U22529 ( .A1(n20489), .A2(n20488), .ZN(n20508) );
  AOI211_X1 U22530 ( .C1(n20489), .C2(n20488), .A(n20508), .B(n21247), .ZN(
        n20494) );
  NAND2_X1 U22531 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20490), .ZN(n20500) );
  NOR3_X1 U22532 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n20517), .A3(n20500), 
        .ZN(n20493) );
  OAI22_X1 U22533 ( .A1(n20491), .A2(n20572), .B1(n20570), .B2(n20495), .ZN(
        n20492) );
  NOR3_X1 U22534 ( .A1(n20494), .A2(n20493), .A3(n20492), .ZN(n20498) );
  NAND2_X1 U22535 ( .A1(n20496), .A2(n20495), .ZN(n20506) );
  OAI211_X1 U22536 ( .C1(n20496), .C2(n20495), .A(n20586), .B(n20506), .ZN(
        n20497) );
  OAI211_X1 U22537 ( .C1(n20499), .C2(n20501), .A(n20498), .B(n20497), .ZN(
        P3_U2646) );
  NOR2_X1 U22538 ( .A1(n20501), .A2(n20500), .ZN(n20503) );
  NAND2_X1 U22539 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n20503), .ZN(n20516) );
  AND2_X1 U22540 ( .A1(n20502), .A2(n20516), .ZN(n20504) );
  AOI22_X1 U22541 ( .A1(n20587), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n20503), 
        .B2(n20504), .ZN(n20514) );
  NOR2_X1 U22542 ( .A1(n20505), .A2(n20504), .ZN(n20527) );
  INV_X1 U22543 ( .A(n20527), .ZN(n20542) );
  NOR2_X1 U22544 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n20506), .ZN(n20524) );
  AOI211_X1 U22545 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20506), .A(n20524), .B(
        n20562), .ZN(n20512) );
  INV_X1 U22546 ( .A(n20507), .ZN(n20510) );
  NOR2_X1 U22547 ( .A1(n20510), .A2(n20509), .ZN(n20518) );
  AOI211_X1 U22548 ( .C1(n20510), .C2(n20509), .A(n20518), .B(n21247), .ZN(
        n20511) );
  AOI211_X1 U22549 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n20542), .A(n20512), 
        .B(n20511), .ZN(n20513) );
  OAI211_X1 U22550 ( .C1(n20515), .C2(n20572), .A(n20514), .B(n20513), .ZN(
        P3_U2645) );
  NOR2_X1 U22551 ( .A1(n20517), .A2(n20516), .ZN(n20556) );
  AND2_X1 U22552 ( .A1(n20539), .A2(n20556), .ZN(n20531) );
  AOI211_X1 U22553 ( .C1(n20520), .C2(n20519), .A(n10988), .B(n21247), .ZN(
        n20522) );
  INV_X1 U22554 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n20523) );
  OAI22_X1 U22555 ( .A1(n11201), .A2(n20572), .B1(n20570), .B2(n20523), .ZN(
        n20521) );
  NOR3_X1 U22556 ( .A1(n20531), .A2(n20522), .A3(n20521), .ZN(n20526) );
  NAND2_X1 U22557 ( .A1(n20524), .A2(n20523), .ZN(n20529) );
  OAI211_X1 U22558 ( .C1(n20524), .C2(n20523), .A(n20586), .B(n20529), .ZN(
        n20525) );
  OAI211_X1 U22559 ( .C1(n20527), .C2(n20539), .A(n20526), .B(n20525), .ZN(
        P3_U2644) );
  AOI22_X1 U22560 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20528), .B1(
        n20587), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n20538) );
  NOR2_X1 U22561 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n20529), .ZN(n20545) );
  AOI211_X1 U22562 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n20529), .A(n20545), .B(
        n20562), .ZN(n20530) );
  AOI221_X1 U22563 ( .B1(n20531), .B2(P3_REIP_REG_28__SCAN_IN), .C1(n20542), 
        .C2(P3_REIP_REG_28__SCAN_IN), .A(n20530), .ZN(n20537) );
  NOR2_X1 U22564 ( .A1(n10988), .A2(n11194), .ZN(n20533) );
  INV_X1 U22565 ( .A(n20533), .ZN(n20532) );
  OAI221_X1 U22566 ( .B1(n20534), .B2(n20533), .C1(n20547), .C2(n20532), .A(
        n20560), .ZN(n20536) );
  NAND3_X1 U22567 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n20556), .A3(n20540), 
        .ZN(n20535) );
  NAND4_X1 U22568 ( .A1(n20538), .A2(n20537), .A3(n20536), .A4(n20535), .ZN(
        P3_U2643) );
  NOR3_X1 U22569 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n20540), .A3(n20539), 
        .ZN(n20541) );
  AOI22_X1 U22570 ( .A1(n20587), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n20556), 
        .B2(n20541), .ZN(n20553) );
  NAND3_X1 U22571 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n20543) );
  AOI21_X1 U22572 ( .B1(n20543), .B2(n20585), .A(n20542), .ZN(n20558) );
  INV_X1 U22573 ( .A(n20558), .ZN(n20578) );
  INV_X1 U22574 ( .A(n20545), .ZN(n20546) );
  NAND2_X1 U22575 ( .A1(n20545), .A2(n20544), .ZN(n20561) );
  NAND2_X1 U22576 ( .A1(n20586), .A2(n20561), .ZN(n20565) );
  AOI21_X1 U22577 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n20546), .A(n20565), .ZN(
        n20551) );
  AOI211_X1 U22578 ( .C1(n20549), .C2(n20548), .A(n20555), .B(n21247), .ZN(
        n20550) );
  AOI211_X1 U22579 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n20578), .A(n20551), 
        .B(n20550), .ZN(n20552) );
  OAI211_X1 U22580 ( .C1(n20554), .C2(n20572), .A(n20553), .B(n20552), .ZN(
        P3_U2642) );
  NAND4_X1 U22582 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n20556), .ZN(n20568) );
  NOR2_X1 U22583 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n20568), .ZN(n20579) );
  OAI22_X1 U22584 ( .A1(n20558), .A2(n20569), .B1(n20557), .B2(n20572), .ZN(
        n20559) );
  NOR2_X1 U22585 ( .A1(n20562), .A2(n20561), .ZN(n20577) );
  OAI21_X1 U22586 ( .B1(n20587), .B2(n20577), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n20563) );
  OAI211_X1 U22587 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n20565), .A(n20564), .B(
        n20563), .ZN(P3_U2641) );
  NAND2_X1 U22588 ( .A1(n20567), .A2(n20566), .ZN(n20583) );
  NOR3_X1 U22589 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n20569), .A3(n20568), 
        .ZN(n20575) );
  OAI22_X1 U22590 ( .A1(n20573), .A2(n20572), .B1(n20571), .B2(n20570), .ZN(
        n20574) );
  AOI211_X1 U22591 ( .C1(n20577), .C2(n20576), .A(n20575), .B(n20574), .ZN(
        n20581) );
  OAI21_X1 U22592 ( .B1(n20579), .B2(n20578), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n20580) );
  OAI211_X1 U22593 ( .C1(n20583), .C2(n20582), .A(n20581), .B(n20580), .ZN(
        P3_U2640) );
  AOI22_X1 U22594 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n20585), .B1(n20584), 
        .B2(n20784), .ZN(n20591) );
  OAI21_X1 U22595 ( .B1(n20587), .B2(n20586), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n20590) );
  NAND3_X1 U22596 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20588), .A3(
        n20790), .ZN(n20589) );
  NAND3_X1 U22597 ( .A1(n20591), .A2(n20590), .A3(n20589), .ZN(P3_U2671) );
  NOR2_X1 U22598 ( .A1(n12661), .A2(n20592), .ZN(n20596) );
  NAND2_X1 U22599 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .ZN(n20624) );
  NAND4_X1 U22600 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .A4(P3_EAX_REG_7__SCAN_IN), .ZN(n20597) );
  NOR2_X1 U22601 ( .A1(n20624), .A2(n20597), .ZN(n20651) );
  NAND4_X1 U22602 ( .A1(n20667), .A2(n20767), .A3(n20651), .A4(
        P3_EAX_REG_8__SCAN_IN), .ZN(n20619) );
  NOR2_X1 U22603 ( .A1(n20598), .A2(n20619), .ZN(n20622) );
  NAND2_X1 U22604 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20622), .ZN(n20616) );
  NOR2_X1 U22605 ( .A1(n20599), .A2(n20616), .ZN(n20613) );
  NAND2_X1 U22606 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n20613), .ZN(n20606) );
  NAND2_X1 U22607 ( .A1(n20606), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n20605) );
  NOR2_X1 U22608 ( .A1(n20601), .A2(n20600), .ZN(n20777) );
  AOI22_X1 U22609 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20777), .B1(n20776), .B2(
        n20603), .ZN(n20604) );
  OAI221_X1 U22610 ( .B1(n20606), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n20605), 
        .C2(n20768), .A(n20604), .ZN(P3_U2722) );
  INV_X1 U22611 ( .A(n20777), .ZN(n20642) );
  INV_X1 U22612 ( .A(n20606), .ZN(n20749) );
  AOI21_X1 U22613 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n20751), .A(n20613), .ZN(
        n20608) );
  OAI222_X1 U22614 ( .A1(n20642), .A2(n20609), .B1(n20749), .B2(n20608), .C1(
        n20773), .C2(n20607), .ZN(P3_U2723) );
  INV_X1 U22615 ( .A(n20616), .ZN(n20610) );
  AOI21_X1 U22616 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n20751), .A(n20610), .ZN(
        n20612) );
  OAI222_X1 U22617 ( .A1(n20642), .A2(n20614), .B1(n20613), .B2(n20612), .C1(
        n20773), .C2(n20611), .ZN(P3_U2724) );
  AOI22_X1 U22618 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20777), .B1(n20776), .B2(
        n20615), .ZN(n20618) );
  OAI211_X1 U22619 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n20622), .A(n20751), .B(
        n20616), .ZN(n20617) );
  NAND2_X1 U22620 ( .A1(n20618), .A2(n20617), .ZN(P3_U2725) );
  INV_X1 U22621 ( .A(n20619), .ZN(n20761) );
  AOI21_X1 U22622 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n20751), .A(n20761), .ZN(
        n20621) );
  OAI222_X1 U22623 ( .A1(n20642), .A2(n20623), .B1(n20622), .B2(n20621), .C1(
        n20773), .C2(n20620), .ZN(P3_U2726) );
  AND2_X1 U22624 ( .A1(n20651), .A2(n20767), .ZN(n20628) );
  NAND3_X1 U22625 ( .A1(n20667), .A2(n20767), .A3(P3_EAX_REG_2__SCAN_IN), .ZN(
        n20648) );
  NOR2_X1 U22626 ( .A1(n20624), .A2(n20648), .ZN(n20641) );
  NAND2_X1 U22627 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n20641), .ZN(n20630) );
  NOR2_X1 U22628 ( .A1(n20625), .A2(n20630), .ZN(n20633) );
  AOI21_X1 U22629 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n20751), .A(n20633), .ZN(
        n20627) );
  OAI222_X1 U22630 ( .A1(n20629), .A2(n20642), .B1(n20628), .B2(n20627), .C1(
        n20773), .C2(n20626), .ZN(P3_U2728) );
  INV_X1 U22631 ( .A(n20630), .ZN(n20636) );
  AOI21_X1 U22632 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n20751), .A(n20636), .ZN(
        n20632) );
  OAI222_X1 U22633 ( .A1(n20674), .A2(n20642), .B1(n20633), .B2(n20632), .C1(
        n20773), .C2(n20631), .ZN(P3_U2729) );
  AOI21_X1 U22634 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n20751), .A(n20641), .ZN(
        n20635) );
  OAI222_X1 U22635 ( .A1(n20637), .A2(n20642), .B1(n20636), .B2(n20635), .C1(
        n20773), .C2(n20634), .ZN(P3_U2730) );
  INV_X1 U22636 ( .A(n20648), .ZN(n20638) );
  AOI22_X1 U22637 ( .A1(n20638), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n20751), .ZN(n20640) );
  OAI222_X1 U22638 ( .A1(n20643), .A2(n20642), .B1(n20641), .B2(n20640), .C1(
        n20773), .C2(n20639), .ZN(P3_U2731) );
  NAND2_X1 U22639 ( .A1(n20648), .A2(P3_EAX_REG_3__SCAN_IN), .ZN(n20646) );
  AOI22_X1 U22640 ( .A1(n20777), .A2(BUF2_REG_3__SCAN_IN), .B1(n20776), .B2(
        n20644), .ZN(n20645) );
  OAI221_X1 U22641 ( .B1(n20648), .B2(P3_EAX_REG_3__SCAN_IN), .C1(n20646), 
        .C2(n20768), .A(n20645), .ZN(P3_U2732) );
  AOI22_X1 U22642 ( .A1(n20777), .A2(BUF2_REG_2__SCAN_IN), .B1(n20776), .B2(
        n20647), .ZN(n20650) );
  OAI211_X1 U22643 ( .C1(n20767), .C2(P3_EAX_REG_2__SCAN_IN), .A(n20751), .B(
        n20648), .ZN(n20649) );
  NAND2_X1 U22644 ( .A1(n20650), .A2(n20649), .ZN(P3_U2733) );
  NAND2_X1 U22645 ( .A1(n20767), .A2(n20651), .ZN(n20763) );
  NAND4_X1 U22646 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(P3_EAX_REG_13__SCAN_IN), .ZN(n20652)
         );
  NOR2_X1 U22647 ( .A1(n20763), .A2(n20652), .ZN(n20653) );
  NAND4_X1 U22648 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(n20653), .ZN(n20757) );
  NAND2_X1 U22649 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n20685), .ZN(n20681) );
  NAND2_X1 U22650 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20675), .ZN(n20662) );
  NAND2_X1 U22651 ( .A1(n20751), .A2(n20662), .ZN(n20668) );
  NOR2_X2 U22652 ( .A1(n20655), .A2(n20751), .ZN(n20735) );
  NOR2_X2 U22653 ( .A1(n20656), .A2(n20751), .ZN(n20743) );
  INV_X1 U22654 ( .A(n20743), .ZN(n20741) );
  OAI22_X1 U22655 ( .A1(n20658), .A2(n20773), .B1(n20657), .B2(n20741), .ZN(
        n20659) );
  AOI21_X1 U22656 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n20735), .A(n20659), .ZN(
        n20660) );
  OAI221_X1 U22657 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n20662), .C1(n20661), 
        .C2(n20668), .A(n20660), .ZN(P3_U2714) );
  AOI22_X1 U22658 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20735), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20743), .ZN(n20664) );
  OAI211_X1 U22659 ( .C1(n20675), .C2(P3_EAX_REG_20__SCAN_IN), .A(n20751), .B(
        n20662), .ZN(n20663) );
  OAI211_X1 U22660 ( .C1(n20665), .C2(n20773), .A(n20664), .B(n20663), .ZN(
        P3_U2715) );
  INV_X1 U22661 ( .A(n20735), .ZN(n20748) );
  AOI22_X1 U22662 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n20743), .B1(n20776), .B2(
        n20666), .ZN(n20673) );
  NAND2_X1 U22663 ( .A1(n20667), .A2(n20779), .ZN(n20781) );
  OAI21_X1 U22664 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n20781), .A(n20668), .ZN(
        n20671) );
  NAND2_X1 U22665 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .ZN(n20692) );
  INV_X1 U22666 ( .A(n20675), .ZN(n20669) );
  NOR3_X1 U22667 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n20692), .A3(n20669), .ZN(
        n20670) );
  AOI21_X1 U22668 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(n20671), .A(n20670), .ZN(
        n20672) );
  OAI211_X1 U22669 ( .C1(n20674), .C2(n20748), .A(n20673), .B(n20672), .ZN(
        P3_U2713) );
  AOI22_X1 U22670 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20735), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20743), .ZN(n20679) );
  AOI211_X1 U22671 ( .C1(n20676), .C2(n20681), .A(n20675), .B(n20768), .ZN(
        n20677) );
  INV_X1 U22672 ( .A(n20677), .ZN(n20678) );
  OAI211_X1 U22673 ( .C1(n20680), .C2(n20773), .A(n20679), .B(n20678), .ZN(
        P3_U2716) );
  AOI22_X1 U22674 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20735), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20743), .ZN(n20683) );
  OAI211_X1 U22675 ( .C1(n20685), .C2(P3_EAX_REG_18__SCAN_IN), .A(n20751), .B(
        n20681), .ZN(n20682) );
  OAI211_X1 U22676 ( .C1(n20684), .C2(n20773), .A(n20683), .B(n20682), .ZN(
        P3_U2717) );
  AOI22_X1 U22677 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20735), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20743), .ZN(n20689) );
  INV_X1 U22678 ( .A(n20744), .ZN(n20687) );
  INV_X1 U22679 ( .A(n20685), .ZN(n20686) );
  OAI211_X1 U22680 ( .C1(n20687), .C2(P3_EAX_REG_17__SCAN_IN), .A(n20751), .B(
        n20686), .ZN(n20688) );
  OAI211_X1 U22681 ( .C1(n20690), .C2(n20773), .A(n20689), .B(n20688), .ZN(
        P3_U2718) );
  NAND4_X1 U22682 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n20691)
         );
  NAND2_X1 U22683 ( .A1(n20737), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n20736) );
  INV_X1 U22684 ( .A(n20700), .ZN(n20696) );
  OAI21_X1 U22685 ( .B1(n20768), .B2(n20694), .A(n20729), .ZN(n20695) );
  AOI22_X1 U22686 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n20743), .B1(n20696), .B2(
        n20695), .ZN(n20699) );
  AOI22_X1 U22687 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20735), .B1(n20776), .B2(
        n20697), .ZN(n20698) );
  NAND2_X1 U22688 ( .A1(n20699), .A2(n20698), .ZN(P3_U2710) );
  AOI22_X1 U22689 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20735), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20743), .ZN(n20702) );
  NAND2_X1 U22690 ( .A1(n20700), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n20722) );
  OAI211_X1 U22691 ( .C1(n20700), .C2(P3_EAX_REG_26__SCAN_IN), .A(n20751), .B(
        n20722), .ZN(n20701) );
  OAI211_X1 U22692 ( .C1(n20703), .C2(n20773), .A(n20702), .B(n20701), .ZN(
        P3_U2709) );
  NAND2_X1 U22693 ( .A1(n20721), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n20717) );
  NAND2_X1 U22694 ( .A1(n20710), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n20706) );
  NAND2_X1 U22695 ( .A1(n20706), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n20705) );
  NAND2_X1 U22696 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n20743), .ZN(n20704) );
  OAI221_X1 U22697 ( .B1(n20706), .B2(P3_EAX_REG_31__SCAN_IN), .C1(n20705), 
        .C2(n20768), .A(n20704), .ZN(P3_U2704) );
  AOI22_X1 U22698 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20735), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20743), .ZN(n20708) );
  OAI211_X1 U22699 ( .C1(n20710), .C2(P3_EAX_REG_30__SCAN_IN), .A(n20751), .B(
        n20706), .ZN(n20707) );
  OAI211_X1 U22700 ( .C1(n20709), .C2(n20773), .A(n20708), .B(n20707), .ZN(
        P3_U2705) );
  INV_X1 U22701 ( .A(n20710), .ZN(n20713) );
  OAI21_X1 U22702 ( .B1(n20768), .B2(n20711), .A(n20717), .ZN(n20712) );
  AOI22_X1 U22703 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20743), .B1(n20713), .B2(
        n20712), .ZN(n20716) );
  AOI22_X1 U22704 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20735), .B1(n20776), .B2(
        n20714), .ZN(n20715) );
  NAND2_X1 U22705 ( .A1(n20716), .A2(n20715), .ZN(P3_U2706) );
  AOI22_X1 U22706 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20735), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20743), .ZN(n20719) );
  OAI211_X1 U22707 ( .C1(n20721), .C2(P3_EAX_REG_28__SCAN_IN), .A(n20751), .B(
        n20717), .ZN(n20718) );
  OAI211_X1 U22708 ( .C1(n20720), .C2(n20773), .A(n20719), .B(n20718), .ZN(
        P3_U2707) );
  INV_X1 U22709 ( .A(n20721), .ZN(n20725) );
  OAI21_X1 U22710 ( .B1(n20768), .B2(n20723), .A(n20722), .ZN(n20724) );
  AOI22_X1 U22711 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20743), .B1(n20725), .B2(
        n20724), .ZN(n20728) );
  AOI22_X1 U22712 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20735), .B1(n20776), .B2(
        n20726), .ZN(n20727) );
  NAND2_X1 U22713 ( .A1(n20728), .A2(n20727), .ZN(P3_U2708) );
  AOI22_X1 U22714 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20735), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20743), .ZN(n20732) );
  OAI211_X1 U22715 ( .C1(n20730), .C2(P3_EAX_REG_24__SCAN_IN), .A(n20751), .B(
        n20729), .ZN(n20731) );
  OAI211_X1 U22716 ( .C1(n20733), .C2(n20773), .A(n20732), .B(n20731), .ZN(
        P3_U2711) );
  AOI22_X1 U22717 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20735), .B1(n20776), .B2(
        n20734), .ZN(n20739) );
  OAI211_X1 U22718 ( .C1(n20737), .C2(P3_EAX_REG_23__SCAN_IN), .A(n20751), .B(
        n20736), .ZN(n20738) );
  OAI211_X1 U22719 ( .C1(n20741), .C2(n20740), .A(n20739), .B(n20738), .ZN(
        P3_U2712) );
  AOI22_X1 U22720 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n20743), .B1(n20776), .B2(
        n20742), .ZN(n20746) );
  OAI211_X1 U22721 ( .C1(n20755), .C2(P3_EAX_REG_16__SCAN_IN), .A(n20751), .B(
        n20744), .ZN(n20745) );
  OAI211_X1 U22722 ( .C1(n20748), .C2(n20747), .A(n20746), .B(n20745), .ZN(
        P3_U2719) );
  NAND2_X1 U22723 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n20749), .ZN(n20754) );
  AOI22_X1 U22724 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20777), .B1(n20776), .B2(
        n20750), .ZN(n20753) );
  NAND3_X1 U22725 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n20751), .A3(n20757), 
        .ZN(n20752) );
  OAI211_X1 U22726 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n20754), .A(n20753), .B(
        n20752), .ZN(P3_U2721) );
  AOI211_X1 U22727 ( .C1(n20757), .C2(n20756), .A(n20768), .B(n20755), .ZN(
        n20758) );
  AOI21_X1 U22728 ( .B1(n20777), .B2(BUF2_REG_15__SCAN_IN), .A(n20758), .ZN(
        n20759) );
  OAI21_X1 U22729 ( .B1(n20760), .B2(n20773), .A(n20759), .ZN(P3_U2720) );
  AOI211_X1 U22730 ( .C1(n20763), .C2(n20762), .A(n20768), .B(n20761), .ZN(
        n20764) );
  AOI21_X1 U22731 ( .B1(n20777), .B2(BUF2_REG_8__SCAN_IN), .A(n20764), .ZN(
        n20765) );
  OAI21_X1 U22732 ( .B1(n20766), .B2(n20773), .A(n20765), .ZN(P3_U2727) );
  AOI211_X1 U22733 ( .C1(n20770), .C2(n20769), .A(n20768), .B(n20767), .ZN(
        n20771) );
  AOI21_X1 U22734 ( .B1(n20777), .B2(BUF2_REG_1__SCAN_IN), .A(n20771), .ZN(
        n20772) );
  OAI21_X1 U22735 ( .B1(n20774), .B2(n20773), .A(n20772), .ZN(P3_U2734) );
  AOI22_X1 U22736 ( .A1(n20777), .A2(BUF2_REG_0__SCAN_IN), .B1(n20776), .B2(
        n20775), .ZN(n20778) );
  OAI221_X1 U22737 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n20781), .C1(n20780), 
        .C2(n20779), .A(n20778), .ZN(P3_U2735) );
  NAND2_X1 U22738 ( .A1(n21004), .A2(n20782), .ZN(n20787) );
  AOI22_X1 U22739 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20955), .B1(
        n20787), .B2(n20784), .ZN(n21218) );
  INV_X1 U22740 ( .A(n21218), .ZN(n21215) );
  AOI222_X1 U22741 ( .A1(n20860), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21215), 
        .B2(n20824), .C1(n20784), .C2(n21254), .ZN(n20783) );
  AOI22_X1 U22742 ( .A1(n20828), .A2(n20784), .B1(n20783), .B2(n20826), .ZN(
        P3_U3290) );
  NOR2_X1 U22743 ( .A1(n20785), .A2(n20860), .ZN(n20804) );
  AOI22_X1 U22744 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12891), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n12489), .ZN(n20802) );
  AOI21_X1 U22745 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20954), .A(
        n20786), .ZN(n20818) );
  NAND2_X1 U22746 ( .A1(n20818), .A2(n21204), .ZN(n20793) );
  AOI22_X1 U22747 ( .A1(n20788), .A2(n20787), .B1(n20794), .B2(n20793), .ZN(
        n21220) );
  NAND2_X1 U22748 ( .A1(n21254), .A2(n20809), .ZN(n20807) );
  OAI22_X1 U22749 ( .A1(n21220), .A2(n20790), .B1(n20789), .B2(n20807), .ZN(
        n20791) );
  AOI21_X1 U22750 ( .B1(n20804), .B2(n20802), .A(n20791), .ZN(n20792) );
  AOI22_X1 U22751 ( .A1(n20828), .A2(n20794), .B1(n20792), .B2(n20826), .ZN(
        P3_U3289) );
  OAI221_X1 U22752 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C1(n20794), .C2(n20808), .A(
        n20793), .ZN(n20800) );
  NOR2_X1 U22753 ( .A1(n20796), .A2(n20795), .ZN(n20797) );
  NOR2_X1 U22754 ( .A1(n20798), .A2(n20797), .ZN(n20815) );
  OR3_X1 U22755 ( .A1(n20808), .A2(n10962), .A3(n20815), .ZN(n20799) );
  OAI211_X1 U22756 ( .C1(n21203), .C2(n20801), .A(n20800), .B(n20799), .ZN(
        n21223) );
  INV_X1 U22757 ( .A(n20802), .ZN(n20805) );
  NOR2_X1 U22758 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20809), .ZN(
        n20803) );
  AOI222_X1 U22759 ( .A1(n21223), .A2(n20824), .B1(n20805), .B2(n20804), .C1(
        n21254), .C2(n20803), .ZN(n20806) );
  OAI222_X1 U22760 ( .A1(n20808), .A2(n20807), .B1(n20808), .B2(n20826), .C1(
        n20828), .C2(n20806), .ZN(P3_U3288) );
  AOI211_X1 U22761 ( .C1(n20810), .C2(n20809), .A(n17642), .B(n21203), .ZN(
        n20822) );
  NAND2_X1 U22762 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20811), .ZN(
        n20813) );
  AOI221_X1 U22763 ( .B1(n20814), .B2(n20813), .C1(n20817), .C2(n20813), .A(
        n20812), .ZN(n20820) );
  OAI22_X1 U22764 ( .A1(n20818), .A2(n20817), .B1(n20816), .B2(n20815), .ZN(
        n20819) );
  AOI211_X1 U22765 ( .C1(n20822), .C2(n20821), .A(n20820), .B(n20819), .ZN(
        n21213) );
  INV_X1 U22766 ( .A(n21213), .ZN(n20823) );
  AOI22_X1 U22767 ( .A1(n21254), .A2(n20825), .B1(n20824), .B2(n20823), .ZN(
        n20827) );
  AOI22_X1 U22768 ( .A1(n20828), .A2(n21214), .B1(n20827), .B2(n20826), .ZN(
        P3_U3285) );
  NAND2_X1 U22769 ( .A1(n21078), .A2(n20829), .ZN(n21127) );
  AOI21_X1 U22770 ( .B1(n21194), .B2(n20831), .A(n20830), .ZN(n20844) );
  NAND3_X1 U22771 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20832), .A3(
        n21184), .ZN(n20986) );
  AOI221_X1 U22772 ( .B1(n20986), .B2(n20954), .C1(n20833), .C2(n20954), .A(
        n21068), .ZN(n21113) );
  INV_X1 U22773 ( .A(n20841), .ZN(n20840) );
  NAND2_X1 U22774 ( .A1(n21162), .A2(n21203), .ZN(n21006) );
  OAI21_X1 U22775 ( .B1(n21134), .B2(n20834), .A(n20955), .ZN(n20835) );
  OAI21_X1 U22776 ( .B1(n20836), .B2(n21203), .A(n20835), .ZN(n21115) );
  OAI22_X1 U22777 ( .A1(n20838), .A2(n21202), .B1(n20837), .B2(n21063), .ZN(
        n20839) );
  AOI211_X1 U22778 ( .C1(n20840), .C2(n21006), .A(n21115), .B(n20839), .ZN(
        n21003) );
  OAI211_X1 U22779 ( .C1(n20841), .C2(n21004), .A(n21113), .B(n21003), .ZN(
        n20842) );
  NAND3_X1 U22780 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n10961), .A3(
        n20842), .ZN(n20843) );
  OAI211_X1 U22781 ( .C1(n21127), .C2(n20845), .A(n20844), .B(n20843), .ZN(
        P3_U2841) );
  INV_X1 U22782 ( .A(n20921), .ZN(n21033) );
  INV_X1 U22783 ( .A(n20923), .ZN(n20911) );
  NAND2_X1 U22784 ( .A1(n21004), .A2(n21203), .ZN(n21119) );
  NAND2_X1 U22785 ( .A1(n20860), .A2(n21119), .ZN(n20853) );
  AOI221_X1 U22786 ( .B1(n21162), .B2(n20853), .C1(n20860), .C2(n20853), .A(
        n21068), .ZN(n20846) );
  AOI221_X1 U22787 ( .B1(n21033), .B2(n20848), .C1(n20911), .C2(n20847), .A(
        n20846), .ZN(n20850) );
  NAND2_X1 U22788 ( .A1(n21189), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n20849) );
  OAI211_X1 U22789 ( .C1(n21086), .C2(n20860), .A(n20850), .B(n20849), .ZN(
        P3_U2862) );
  AOI22_X1 U22790 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21092), .B1(
        n20911), .B2(n20851), .ZN(n20858) );
  NOR3_X1 U22791 ( .A1(n21103), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n20852), .ZN(n20856) );
  OAI22_X1 U22792 ( .A1(n20854), .A2(n21202), .B1(n12489), .B2(n20853), .ZN(
        n20855) );
  OAI21_X1 U22793 ( .B1(n20856), .B2(n20855), .A(n21078), .ZN(n20857) );
  OAI211_X1 U22794 ( .C1(n20859), .C2(n10961), .A(n20858), .B(n20857), .ZN(
        P3_U2861) );
  INV_X1 U22795 ( .A(n20873), .ZN(n20877) );
  NOR2_X1 U22796 ( .A1(n12489), .A2(n20860), .ZN(n20861) );
  OAI221_X1 U22797 ( .B1(n20877), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n20877), .C2(n20861), .A(n21133), .ZN(n20866) );
  AOI211_X1 U22798 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n21049), .A(
        n20874), .B(n20871), .ZN(n20863) );
  AND3_X1 U22799 ( .A1(n20871), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n20872), .ZN(n20862) );
  AOI211_X1 U22800 ( .C1(n20864), .C2(n21209), .A(n20863), .B(n20862), .ZN(
        n20865) );
  AOI21_X1 U22801 ( .B1(n20866), .B2(n20865), .A(n21068), .ZN(n20867) );
  AOI211_X1 U22802 ( .C1(n21092), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n20868), .B(n20867), .ZN(n20869) );
  OAI21_X1 U22803 ( .B1(n20921), .B2(n20870), .A(n20869), .ZN(P3_U2860) );
  NOR2_X1 U22804 ( .A1(n20871), .A2(n12489), .ZN(n20875) );
  AOI22_X1 U22805 ( .A1(n20873), .A2(n21133), .B1(n20872), .B2(n20875), .ZN(
        n20886) );
  AOI21_X1 U22806 ( .B1(n20875), .B2(n21049), .A(n20874), .ZN(n20876) );
  AOI211_X1 U22807 ( .C1(n21133), .C2(n20877), .A(n20876), .B(n20878), .ZN(
        n20887) );
  AOI211_X1 U22808 ( .C1(n20886), .C2(n20878), .A(n20887), .B(n21068), .ZN(
        n20881) );
  OAI22_X1 U22809 ( .A1(n10961), .A2(n20879), .B1(n20878), .B2(n21086), .ZN(
        n20880) );
  AOI211_X1 U22810 ( .C1(n20882), .C2(n20911), .A(n20881), .B(n20880), .ZN(
        n20883) );
  OAI21_X1 U22811 ( .B1(n20921), .B2(n20884), .A(n20883), .ZN(P3_U2859) );
  AOI21_X1 U22812 ( .B1(n21092), .B2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n20885), .ZN(n20893) );
  INV_X1 U22813 ( .A(n20886), .ZN(n20905) );
  AND2_X1 U22814 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n20905), .ZN(
        n20889) );
  NOR2_X1 U22815 ( .A1(n21103), .A2(n20887), .ZN(n20888) );
  MUX2_X1 U22816 ( .A(n20889), .B(n20888), .S(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n20891) );
  AOI22_X1 U22817 ( .A1(n21078), .A2(n20891), .B1(n20911), .B2(n20890), .ZN(
        n20892) );
  OAI211_X1 U22818 ( .C1(n20921), .C2(n20894), .A(n20893), .B(n20892), .ZN(
        P3_U2858) );
  NAND4_X1 U22819 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n21078), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A4(n20905), .ZN(n20904) );
  INV_X1 U22820 ( .A(n21049), .ZN(n21187) );
  AOI21_X1 U22821 ( .B1(n21185), .B2(n20895), .A(n21187), .ZN(n20896) );
  OAI21_X1 U22822 ( .B1(n20897), .B2(n21203), .A(n20896), .ZN(n20915) );
  OAI21_X1 U22823 ( .B1(n21068), .B2(n20915), .A(n10961), .ZN(n20907) );
  OAI22_X1 U22824 ( .A1(n10961), .A2(n20899), .B1(n20921), .B2(n20898), .ZN(
        n20900) );
  AOI21_X1 U22825 ( .B1(n20911), .B2(n20901), .A(n20900), .ZN(n20902) );
  OAI221_X1 U22826 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n20904), .C1(
        n20903), .C2(n20907), .A(n20902), .ZN(P3_U2857) );
  NAND2_X1 U22827 ( .A1(n20906), .A2(n20905), .ZN(n20917) );
  NOR3_X1 U22828 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21068), .A3(
        n20917), .ZN(n20910) );
  INV_X1 U22829 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n20918) );
  OAI22_X1 U22830 ( .A1(n10961), .A2(n20908), .B1(n20918), .B2(n20907), .ZN(
        n20909) );
  AOI211_X1 U22831 ( .C1(n20912), .C2(n20911), .A(n20910), .B(n20909), .ZN(
        n20913) );
  OAI21_X1 U22832 ( .B1(n20921), .B2(n20914), .A(n20913), .ZN(P3_U2856) );
  AOI211_X1 U22833 ( .C1(n21153), .C2(n20918), .A(n20927), .B(n20915), .ZN(
        n20916) );
  NOR2_X1 U22834 ( .A1(n20916), .A2(n21068), .ZN(n20928) );
  NOR2_X1 U22835 ( .A1(n20918), .A2(n20917), .ZN(n20929) );
  INV_X1 U22836 ( .A(n20919), .ZN(n20922) );
  OAI22_X1 U22837 ( .A1(n20923), .A2(n20922), .B1(n20921), .B2(n20920), .ZN(
        n20924) );
  AOI221_X1 U22838 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n20928), .C1(
        n20929), .C2(n20928), .A(n20924), .ZN(n20926) );
  NAND2_X1 U22839 ( .A1(n21161), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n20925) );
  OAI211_X1 U22840 ( .C1(n21086), .C2(n20927), .A(n20926), .B(n20925), .ZN(
        P3_U2855) );
  AOI21_X1 U22841 ( .B1(n20928), .B2(n21153), .A(n21092), .ZN(n20935) );
  NAND2_X1 U22842 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n20929), .ZN(
        n20942) );
  OAI222_X1 U22843 ( .A1(n20930), .A2(n21202), .B1(n21063), .B2(n20931), .C1(
        n20942), .C2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20932) );
  AOI22_X1 U22844 ( .A1(n21078), .A2(n20932), .B1(n21194), .B2(n20931), .ZN(
        n20934) );
  OAI211_X1 U22845 ( .C1(n20935), .C2(n20943), .A(n20934), .B(n20933), .ZN(
        P3_U2854) );
  NAND2_X1 U22846 ( .A1(n21133), .A2(n20951), .ZN(n20972) );
  OAI221_X1 U22847 ( .B1(n21162), .B2(n20940), .C1(n21162), .C2(n21184), .A(
        n20972), .ZN(n20959) );
  NOR2_X1 U22848 ( .A1(n21111), .A2(n21131), .ZN(n21138) );
  NOR2_X1 U22849 ( .A1(n20958), .A2(n21063), .ZN(n20937) );
  NAND2_X1 U22850 ( .A1(n21133), .A2(n20936), .ZN(n20983) );
  NAND2_X1 U22851 ( .A1(n21078), .A2(n20983), .ZN(n21164) );
  AOI211_X1 U22852 ( .C1(n20938), .C2(n21111), .A(n20937), .B(n21164), .ZN(
        n21191) );
  NAND2_X1 U22853 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21184), .ZN(
        n20952) );
  OAI21_X1 U22854 ( .B1(n21188), .B2(n20952), .A(n20954), .ZN(n20939) );
  OAI211_X1 U22855 ( .C1(n20940), .C2(n21138), .A(n21191), .B(n20939), .ZN(
        n21179) );
  AOI211_X1 U22856 ( .C1(n21174), .C2(n20954), .A(n20959), .B(n21179), .ZN(
        n20941) );
  NOR2_X1 U22857 ( .A1(n20941), .A2(n20956), .ZN(n20948) );
  NOR2_X1 U22858 ( .A1(n20943), .A2(n20942), .ZN(n20987) );
  INV_X1 U22859 ( .A(n20944), .ZN(n20945) );
  NOR3_X1 U22860 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n20946), .A3(
        n21197), .ZN(n20947) );
  AOI221_X1 U22861 ( .B1(P3_REIP_REG_11__SCAN_IN), .B2(n21189), .C1(n20948), 
        .C2(n10961), .A(n20947), .ZN(n20949) );
  OAI21_X1 U22862 ( .B1(n20950), .B2(n21150), .A(n20949), .ZN(P3_U2851) );
  OAI22_X1 U22863 ( .A1(n21068), .A2(n20968), .B1(n21197), .B2(n20951), .ZN(
        n20964) );
  INV_X1 U22864 ( .A(n20957), .ZN(n20953) );
  NOR2_X1 U22865 ( .A1(n20953), .A2(n20952), .ZN(n20970) );
  AOI211_X1 U22866 ( .C1(n20956), .C2(n20955), .A(n20968), .B(n20954), .ZN(
        n20962) );
  AOI21_X1 U22867 ( .B1(n20958), .B2(n20957), .A(n21063), .ZN(n20960) );
  AOI211_X1 U22868 ( .C1(n21111), .C2(n20961), .A(n20960), .B(n20959), .ZN(
        n21168) );
  OAI211_X1 U22869 ( .C1(n20970), .C2(n20962), .A(n21168), .B(n20983), .ZN(
        n20963) );
  AOI22_X1 U22870 ( .A1(n21194), .A2(n20965), .B1(n20964), .B2(n20963), .ZN(
        n20967) );
  OAI211_X1 U22871 ( .C1(n21086), .C2(n20968), .A(n20967), .B(n20966), .ZN(
        P3_U2850) );
  AOI22_X1 U22872 ( .A1(n21161), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21092), .ZN(n20981) );
  NAND2_X1 U22873 ( .A1(n20969), .A2(n20987), .ZN(n20977) );
  AOI21_X1 U22874 ( .B1(n20969), .B2(n21184), .A(n21162), .ZN(n20971) );
  OAI22_X1 U22875 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21203), .B1(
        n21004), .B2(n20970), .ZN(n21163) );
  AOI211_X1 U22876 ( .C1(n21166), .C2(n21119), .A(n20971), .B(n21163), .ZN(
        n20973) );
  NAND3_X1 U22877 ( .A1(n20973), .A2(n20983), .A3(n20972), .ZN(n20974) );
  AOI22_X1 U22878 ( .A1(n21131), .A2(n20975), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n20974), .ZN(n20976) );
  OAI21_X1 U22879 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n20977), .A(
        n20976), .ZN(n20979) );
  AOI22_X1 U22880 ( .A1(n21078), .A2(n20979), .B1(n21033), .B2(n20978), .ZN(
        n20980) );
  OAI211_X1 U22881 ( .C1(n20982), .C2(n21150), .A(n20981), .B(n20980), .ZN(
        P3_U2848) );
  NAND2_X1 U22882 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21004), .ZN(
        n20985) );
  NOR2_X1 U22883 ( .A1(n21162), .A2(n21184), .ZN(n21176) );
  INV_X1 U22884 ( .A(n20983), .ZN(n20984) );
  AOI211_X1 U22885 ( .C1(n20986), .C2(n20985), .A(n21176), .B(n20984), .ZN(
        n20994) );
  NAND2_X1 U22886 ( .A1(n20995), .A2(n20987), .ZN(n20991) );
  INV_X1 U22887 ( .A(n20988), .ZN(n20990) );
  NAND2_X1 U22888 ( .A1(n21131), .A2(n20989), .ZN(n20996) );
  OAI22_X1 U22889 ( .A1(n20994), .A2(n20991), .B1(n20990), .B2(n20996), .ZN(
        n20993) );
  AOI22_X1 U22890 ( .A1(n21078), .A2(n20993), .B1(n21194), .B2(n20992), .ZN(
        n21002) );
  INV_X1 U22891 ( .A(n21006), .ZN(n21177) );
  OAI21_X1 U22892 ( .B1(n20995), .B2(n21177), .A(n20994), .ZN(n21152) );
  INV_X1 U22893 ( .A(n21129), .ZN(n20997) );
  OAI211_X1 U22894 ( .C1(n20997), .C2(n21202), .A(n21078), .B(n20996), .ZN(
        n21154) );
  OAI211_X1 U22895 ( .C1(n21152), .C2(n21154), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n10961), .ZN(n21001) );
  NAND3_X1 U22896 ( .A1(n20998), .A2(n21033), .A3(n12545), .ZN(n20999) );
  NAND4_X1 U22897 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        P3_U2847) );
  OAI211_X1 U22898 ( .C1(n21004), .C2(n21013), .A(n21003), .B(n21049), .ZN(
        n21005) );
  AOI21_X1 U22899 ( .B1(n21007), .B2(n21006), .A(n21005), .ZN(n21008) );
  AOI221_X1 U22900 ( .B1(n21008), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), 
        .C1(n21093), .C2(n21094), .A(n21068), .ZN(n21009) );
  AOI21_X1 U22901 ( .B1(n21092), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n21009), .ZN(n21011) );
  NAND2_X1 U22902 ( .A1(n21189), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n21010) );
  OAI211_X1 U22903 ( .C1(n21012), .C2(n21150), .A(n21011), .B(n21010), .ZN(
        P3_U2840) );
  AOI22_X1 U22904 ( .A1(n21161), .A2(P3_REIP_REG_25__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21092), .ZN(n21029) );
  NAND3_X1 U22905 ( .A1(n21049), .A2(n21013), .A3(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21014) );
  NAND2_X1 U22906 ( .A1(n21014), .A2(n21185), .ZN(n21085) );
  OAI21_X1 U22907 ( .B1(n21094), .B2(n21015), .A(n21133), .ZN(n21090) );
  NAND4_X1 U22908 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n21085), .A4(n21090), .ZN(
        n21017) );
  AOI21_X1 U22909 ( .B1(n21153), .B2(n21017), .A(n21016), .ZN(n21035) );
  NAND2_X1 U22910 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21018) );
  NOR2_X1 U22911 ( .A1(n21094), .A2(n21018), .ZN(n21022) );
  NOR2_X1 U22912 ( .A1(n21020), .A2(n21019), .ZN(n21021) );
  AOI21_X1 U22913 ( .B1(n21022), .B2(n21021), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21025) );
  INV_X1 U22914 ( .A(n21023), .ZN(n21024) );
  OAI22_X1 U22915 ( .A1(n21035), .A2(n21025), .B1(n21063), .B2(n21024), .ZN(
        n21027) );
  AOI22_X1 U22916 ( .A1(n21078), .A2(n21027), .B1(n21033), .B2(n21026), .ZN(
        n21028) );
  OAI211_X1 U22917 ( .C1(n21150), .C2(n21030), .A(n21029), .B(n21028), .ZN(
        P3_U2837) );
  OAI21_X1 U22918 ( .B1(n21093), .B2(n21031), .A(n21038), .ZN(n21040) );
  NAND2_X1 U22919 ( .A1(n21033), .A2(n21032), .ZN(n21048) );
  AND2_X1 U22920 ( .A1(n21034), .A2(n21131), .ZN(n21046) );
  OAI21_X1 U22921 ( .B1(n21103), .B2(n21035), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21036) );
  OAI21_X1 U22922 ( .B1(n21046), .B2(n21036), .A(n21078), .ZN(n21037) );
  OAI211_X1 U22923 ( .C1(n21086), .C2(n21038), .A(n21048), .B(n21037), .ZN(
        n21039) );
  AOI22_X1 U22924 ( .A1(n21194), .A2(n21041), .B1(n21040), .B2(n21039), .ZN(
        n21042) );
  OAI21_X1 U22925 ( .B1(n10961), .B2(n21043), .A(n21042), .ZN(P3_U2836) );
  OAI21_X1 U22926 ( .B1(n21044), .B2(n21093), .A(n21057), .ZN(n21052) );
  AOI211_X1 U22927 ( .C1(n21185), .C2(n21047), .A(n21046), .B(n21045), .ZN(
        n21050) );
  OAI221_X1 U22928 ( .B1(n21068), .B2(n21050), .C1(n21068), .C2(n21049), .A(
        n21048), .ZN(n21051) );
  AOI22_X1 U22929 ( .A1(n21194), .A2(n21053), .B1(n21052), .B2(n21051), .ZN(
        n21056) );
  INV_X1 U22930 ( .A(n21054), .ZN(n21055) );
  OAI211_X1 U22931 ( .C1(n21086), .C2(n21057), .A(n21056), .B(n21055), .ZN(
        P3_U2835) );
  AND2_X1 U22932 ( .A1(n21131), .A2(n21058), .ZN(n21059) );
  AOI211_X1 U22933 ( .C1(n21061), .C2(n21111), .A(n21060), .B(n21059), .ZN(
        n21076) );
  NAND2_X1 U22934 ( .A1(n21078), .A2(n21075), .ZN(n21073) );
  OAI221_X1 U22935 ( .B1(n21068), .B2(n21067), .C1(n21068), .C2(n21066), .A(
        n21086), .ZN(n21069) );
  AOI22_X1 U22936 ( .A1(n21194), .A2(n21070), .B1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n21069), .ZN(n21072) );
  NAND2_X1 U22937 ( .A1(n21161), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n21071) );
  OAI211_X1 U22938 ( .C1(n21076), .C2(n21073), .A(n21072), .B(n21071), .ZN(
        P3_U2833) );
  AOI22_X1 U22939 ( .A1(n21161), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n21092), 
        .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21082) );
  OAI21_X1 U22940 ( .B1(n21076), .B2(n21075), .A(n21074), .ZN(n21077) );
  OAI211_X1 U22941 ( .C1(n21080), .C2(n21079), .A(n21078), .B(n21077), .ZN(
        n21081) );
  OAI211_X1 U22942 ( .C1(n21083), .C2(n21150), .A(n21082), .B(n21081), .ZN(
        P3_U2832) );
  INV_X1 U22943 ( .A(n21084), .ZN(n21089) );
  OAI211_X1 U22944 ( .C1(n21087), .C2(n21202), .A(n21086), .B(n21085), .ZN(
        n21088) );
  AOI21_X1 U22945 ( .B1(n21131), .B2(n21089), .A(n21088), .ZN(n21102) );
  NAND3_X1 U22946 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21102), .A3(
        n21090), .ZN(n21091) );
  NAND2_X1 U22947 ( .A1(n10961), .A2(n21091), .ZN(n21100) );
  INV_X1 U22948 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21099) );
  OR3_X1 U22949 ( .A1(n21094), .A2(n21093), .A3(n21092), .ZN(n21098) );
  AOI21_X1 U22950 ( .B1(n21096), .B2(n21194), .A(n21095), .ZN(n21097) );
  OAI221_X1 U22951 ( .B1(n21100), .B2(n21099), .C1(n21100), .C2(n21098), .A(
        n21097), .ZN(P3_U2839) );
  AOI211_X1 U22952 ( .C1(n21103), .C2(n21102), .A(n21101), .B(n21100), .ZN(
        n21104) );
  AOI21_X1 U22953 ( .B1(n21194), .B2(n21105), .A(n21104), .ZN(n21107) );
  OAI211_X1 U22954 ( .C1(n21108), .C2(n21127), .A(n21107), .B(n21106), .ZN(
        P3_U2838) );
  AOI22_X1 U22955 ( .A1(n21111), .A2(n21110), .B1(n21131), .B2(n21109), .ZN(
        n21112) );
  NAND2_X1 U22956 ( .A1(n21113), .A2(n21112), .ZN(n21114) );
  OAI21_X1 U22957 ( .B1(n21115), .B2(n21114), .A(n10961), .ZN(n21121) );
  AOI21_X1 U22958 ( .B1(n21194), .B2(n21117), .A(n21116), .ZN(n21118) );
  OAI221_X1 U22959 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21127), 
        .C1(n21120), .C2(n21121), .A(n21118), .ZN(P3_U2843) );
  NAND3_X1 U22960 ( .A1(n21120), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n21119), 
        .ZN(n21122) );
  NAND2_X1 U22961 ( .A1(n21122), .A2(n21121), .ZN(n21124) );
  AOI22_X1 U22962 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21124), .B1(
        n21194), .B2(n21123), .ZN(n21126) );
  OAI211_X1 U22963 ( .C1(n21128), .C2(n21127), .A(n21126), .B(n21125), .ZN(
        P3_U2842) );
  AOI211_X1 U22964 ( .C1(n21131), .C2(n21130), .A(n21132), .B(n21129), .ZN(
        n21137) );
  AOI221_X1 U22965 ( .B1(n21139), .B2(n21133), .C1(n21132), .C2(n21133), .A(
        n21164), .ZN(n21136) );
  AOI221_X1 U22966 ( .B1(n21155), .B2(n21185), .C1(n21134), .C2(n21185), .A(
        n21187), .ZN(n21135) );
  OAI211_X1 U22967 ( .C1(n21138), .C2(n21137), .A(n21136), .B(n21135), .ZN(
        n21147) );
  OAI221_X1 U22968 ( .B1(n21147), .B2(n21185), .C1(n21147), .C2(n11246), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21144) );
  NOR2_X1 U22969 ( .A1(n21139), .A2(n21197), .ZN(n21156) );
  AOI22_X1 U22970 ( .A1(n21194), .A2(n21141), .B1(n21140), .B2(n21156), .ZN(
        n21142) );
  OAI221_X1 U22971 ( .B1(n21189), .B2(n21144), .C1(n10961), .C2(n21143), .A(
        n21142), .ZN(P3_U2844) );
  NOR2_X1 U22972 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21155), .ZN(
        n21146) );
  AOI21_X1 U22973 ( .B1(n21156), .B2(n21146), .A(n21145), .ZN(n21149) );
  NAND3_X1 U22974 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n10961), .A3(
        n21147), .ZN(n21148) );
  OAI211_X1 U22975 ( .C1(n21151), .C2(n21150), .A(n21149), .B(n21148), .ZN(
        P3_U2845) );
  OAI221_X1 U22976 ( .B1(n21154), .B2(n21153), .C1(n21154), .C2(n21152), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21160) );
  AOI22_X1 U22977 ( .A1(n21157), .A2(n21194), .B1(n21156), .B2(n21155), .ZN(
        n21158) );
  OAI221_X1 U22978 ( .B1(n21161), .B2(n21160), .C1(n10961), .C2(n21159), .A(
        n21158), .ZN(P3_U2846) );
  AOI21_X1 U22979 ( .B1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n21162), .ZN(n21165) );
  NOR3_X1 U22980 ( .A1(n21165), .A2(n21164), .A3(n21163), .ZN(n21167) );
  AOI211_X1 U22981 ( .C1(n21168), .C2(n21167), .A(n21189), .B(n21166), .ZN(
        n21169) );
  AOI21_X1 U22982 ( .B1(n21194), .B2(n21170), .A(n21169), .ZN(n21172) );
  OAI211_X1 U22983 ( .C1(n21197), .C2(n21173), .A(n21172), .B(n21171), .ZN(
        P3_U2849) );
  NAND2_X1 U22984 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21174), .ZN(
        n21183) );
  AOI22_X1 U22985 ( .A1(n21161), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21194), 
        .B2(n21175), .ZN(n21182) );
  INV_X1 U22986 ( .A(n21176), .ZN(n21178) );
  AOI21_X1 U22987 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21178), .A(
        n21177), .ZN(n21180) );
  OAI211_X1 U22988 ( .C1(n21180), .C2(n21179), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n10961), .ZN(n21181) );
  OAI211_X1 U22989 ( .C1(n21183), .C2(n21197), .A(n21182), .B(n21181), .ZN(
        P3_U2852) );
  INV_X1 U22990 ( .A(n21184), .ZN(n21186) );
  OAI21_X1 U22991 ( .B1(n21187), .B2(n21186), .A(n21185), .ZN(n21190) );
  AOI211_X1 U22992 ( .C1(n21191), .C2(n21190), .A(n21189), .B(n21188), .ZN(
        n21192) );
  AOI21_X1 U22993 ( .B1(n21194), .B2(n21193), .A(n21192), .ZN(n21196) );
  OAI211_X1 U22994 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n21197), .A(
        n21196), .B(n21195), .ZN(P3_U2853) );
  NAND2_X1 U22995 ( .A1(n21679), .A2(n21253), .ZN(n21246) );
  INV_X1 U22996 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n21268) );
  INV_X1 U22997 ( .A(n21198), .ZN(n21199) );
  NAND3_X1 U22998 ( .A1(n21201), .A2(n21200), .A3(n21199), .ZN(n21265) );
  AOI21_X1 U22999 ( .B1(n21271), .B2(n21268), .A(n21265), .ZN(n21237) );
  NAND2_X1 U23000 ( .A1(n21203), .A2(n21202), .ZN(n21212) );
  NAND3_X1 U23001 ( .A1(n21206), .A2(n21205), .A3(n21204), .ZN(n21208) );
  AOI222_X1 U23002 ( .A1(n21212), .A2(n21211), .B1(n21210), .B2(n21209), .C1(
        n21208), .C2(n21207), .ZN(n21269) );
  AOI22_X1 U23003 ( .A1(n21224), .A2(n21214), .B1(n21213), .B2(n21233), .ZN(
        n21231) );
  NOR3_X1 U23004 ( .A1(n21217), .A2(n21216), .A3(n21215), .ZN(n21219) );
  OAI22_X1 U23005 ( .A1(n21220), .A2(n21219), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n21218), .ZN(n21222) );
  AOI21_X1 U23006 ( .B1(n21222), .B2(n21233), .A(n21221), .ZN(n21226) );
  AOI22_X1 U23007 ( .A1(n21224), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n21223), .B2(n21233), .ZN(n21227) );
  OR2_X1 U23008 ( .A1(n21227), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21225) );
  AOI221_X1 U23009 ( .B1(n21226), .B2(n21225), .C1(n21227), .C2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21230) );
  OAI21_X1 U23010 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n21227), .ZN(n21229) );
  AOI222_X1 U23011 ( .A1(n21231), .A2(n21230), .B1(n21231), .B2(n21229), .C1(
        n21230), .C2(n21228), .ZN(n21232) );
  OAI211_X1 U23012 ( .C1(n21234), .C2(n21233), .A(n21269), .B(n21232), .ZN(
        n21235) );
  NOR4_X1 U23013 ( .A1(n21238), .A2(n21237), .A3(n21236), .A4(n21235), .ZN(
        n21264) );
  OAI211_X1 U23014 ( .C1(n21240), .C2(n21239), .A(n21266), .B(n21264), .ZN(
        n21251) );
  OAI21_X1 U23015 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n21723), .A(n21251), 
        .ZN(n21257) );
  INV_X1 U23016 ( .A(n21257), .ZN(n21242) );
  NAND3_X1 U23017 ( .A1(n21243), .A2(n21242), .A3(n21241), .ZN(n21244) );
  NAND4_X1 U23018 ( .A1(n21247), .A2(n21246), .A3(n21245), .A4(n21244), .ZN(
        P3_U2997) );
  NOR2_X1 U23019 ( .A1(n21249), .A2(n21248), .ZN(n21250) );
  OAI21_X1 U23020 ( .B1(n21252), .B2(n21251), .A(n21250), .ZN(P3_U3282) );
  AOI22_X1 U23021 ( .A1(n21255), .A2(n21254), .B1(n21679), .B2(n21253), .ZN(
        n21256) );
  INV_X1 U23022 ( .A(n21256), .ZN(n21260) );
  NOR2_X1 U23023 ( .A1(n21258), .A2(n21257), .ZN(n21259) );
  MUX2_X1 U23024 ( .A(n21260), .B(n21259), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n21262) );
  OAI211_X1 U23025 ( .C1(n21264), .C2(n21263), .A(n21262), .B(n21261), .ZN(
        P3_U2996) );
  NAND2_X1 U23026 ( .A1(n21266), .A2(n21265), .ZN(n21267) );
  INV_X1 U23027 ( .A(n21267), .ZN(n21272) );
  AOI22_X1 U23028 ( .A1(n21272), .A2(n21269), .B1(n21268), .B2(n21267), .ZN(
        P3_U3295) );
  OAI21_X1 U23029 ( .B1(n21272), .B2(n21271), .A(n21270), .ZN(P3_U2637) );
  AOI211_X1 U23030 ( .C1(n21274), .C2(n14439), .A(n21922), .B(n21273), .ZN(
        n21276) );
  OAI21_X1 U23031 ( .B1(n21276), .B2(n21655), .A(n21275), .ZN(n21280) );
  AOI211_X1 U23032 ( .C1(n21278), .C2(n21683), .A(n21277), .B(n13858), .ZN(
        n21279) );
  MUX2_X1 U23033 ( .A(n21280), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21279), 
        .Z(P1_U3485) );
  NOR3_X1 U23034 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21282), .A3(
        n21281), .ZN(n21290) );
  NOR3_X1 U23035 ( .A1(n21285), .A2(n21284), .A3(n21283), .ZN(n21288) );
  AOI22_X1 U23036 ( .A1(n21526), .A2(n21421), .B1(n14073), .B2(
        P1_REIP_REG_14__SCAN_IN), .ZN(n21286) );
  OAI21_X1 U23037 ( .B1(n21288), .B2(n21287), .A(n21286), .ZN(n21289) );
  NOR2_X1 U23038 ( .A1(n21290), .A2(n21289), .ZN(n21291) );
  OAI21_X1 U23039 ( .B1(n21292), .B2(n21382), .A(n21291), .ZN(P1_U3017) );
  INV_X1 U23040 ( .A(n21293), .ZN(n21439) );
  AOI21_X1 U23041 ( .B1(n21421), .B2(n21439), .A(n21294), .ZN(n21305) );
  NAND2_X1 U23042 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21296) );
  OAI21_X1 U23043 ( .B1(n21296), .B2(n21368), .A(n21295), .ZN(n21299) );
  INV_X1 U23044 ( .A(n21297), .ZN(n21298) );
  AOI22_X1 U23045 ( .A1(n21299), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21298), .B2(n21422), .ZN(n21304) );
  NAND3_X1 U23046 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21301), .A3(
        n21300), .ZN(n21302) );
  NAND4_X1 U23047 ( .A1(n21305), .A2(n21304), .A3(n21303), .A4(n21302), .ZN(
        P1_U3029) );
  AOI22_X1 U23048 ( .A1(n21421), .A2(n21455), .B1(n14073), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n21311) );
  AOI22_X1 U23049 ( .A1(n21307), .A2(n21422), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n21306), .ZN(n21310) );
  OAI211_X1 U23050 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n21312), .B(n21308), .ZN(n21309) );
  NAND3_X1 U23051 ( .A1(n21311), .A2(n21310), .A3(n21309), .ZN(P1_U3027) );
  NAND3_X1 U23052 ( .A1(n21313), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n21312), .ZN(n21325) );
  AOI22_X1 U23053 ( .A1(n21421), .A2(n21480), .B1(n14073), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n21320) );
  OAI21_X1 U23054 ( .B1(n21316), .B2(n21315), .A(n21314), .ZN(n21317) );
  AOI22_X1 U23055 ( .A1(n21318), .A2(n21422), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n21317), .ZN(n21319) );
  OAI211_X1 U23056 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n21325), .A(
        n21320), .B(n21319), .ZN(P1_U3025) );
  OAI22_X1 U23057 ( .A1(n21400), .A2(n21401), .B1(n21322), .B2(n21321), .ZN(
        n21339) );
  INV_X1 U23058 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21323) );
  OAI22_X1 U23059 ( .A1(n21414), .A2(n21495), .B1(n21419), .B2(n21323), .ZN(
        n21324) );
  INV_X1 U23060 ( .A(n21324), .ZN(n21331) );
  INV_X1 U23061 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21326) );
  NOR2_X1 U23062 ( .A1(n21326), .A2(n21325), .ZN(n21341) );
  INV_X1 U23063 ( .A(n21341), .ZN(n21327) );
  OAI22_X1 U23064 ( .A1(n21328), .A2(n21382), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21327), .ZN(n21329) );
  INV_X1 U23065 ( .A(n21329), .ZN(n21330) );
  OAI211_X1 U23066 ( .C1(n21334), .C2(n21339), .A(n21331), .B(n21330), .ZN(
        P1_U3024) );
  AOI21_X1 U23067 ( .B1(n21421), .B2(n21333), .A(n21332), .ZN(n21338) );
  AOI21_X1 U23068 ( .B1(n21340), .B2(n21334), .A(n21342), .ZN(n21335) );
  AOI22_X1 U23069 ( .A1(n21336), .A2(n21422), .B1(n21341), .B2(n21335), .ZN(
        n21337) );
  OAI211_X1 U23070 ( .C1(n21340), .C2(n21339), .A(n21338), .B(n21337), .ZN(
        P1_U3023) );
  NAND2_X1 U23071 ( .A1(n21342), .A2(n21341), .ZN(n21362) );
  INV_X1 U23072 ( .A(n21343), .ZN(n21344) );
  AOI21_X1 U23073 ( .B1(n21421), .B2(n21345), .A(n21344), .ZN(n21352) );
  NAND2_X1 U23074 ( .A1(n21366), .A2(n21346), .ZN(n21347) );
  OAI211_X1 U23075 ( .C1(n21349), .C2(n21368), .A(n21348), .B(n21347), .ZN(
        n21358) );
  AOI22_X1 U23076 ( .A1(n21350), .A2(n21422), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21358), .ZN(n21351) );
  OAI211_X1 U23077 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n21362), .A(
        n21352), .B(n21351), .ZN(P1_U3022) );
  OAI21_X1 U23078 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n21353), .ZN(n21361) );
  INV_X1 U23079 ( .A(n21354), .ZN(n21356) );
  AOI21_X1 U23080 ( .B1(n21421), .B2(n21356), .A(n21355), .ZN(n21360) );
  AOI22_X1 U23081 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n21358), .B1(
        n21422), .B2(n21357), .ZN(n21359) );
  OAI211_X1 U23082 ( .C1(n21362), .C2(n21361), .A(n21360), .B(n21359), .ZN(
        P1_U3021) );
  NOR2_X1 U23083 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n11614), .ZN(
        n21363) );
  AOI22_X1 U23084 ( .A1(n14073), .A2(P1_REIP_REG_12__SCAN_IN), .B1(n21363), 
        .B2(n21378), .ZN(n21374) );
  INV_X1 U23085 ( .A(n21364), .ZN(n21365) );
  AOI21_X1 U23086 ( .B1(n21366), .B2(n21365), .A(n21401), .ZN(n21367) );
  OAI21_X1 U23087 ( .B1(n21369), .B2(n21368), .A(n21367), .ZN(n21379) );
  INV_X1 U23088 ( .A(n21379), .ZN(n21370) );
  OAI21_X1 U23089 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n21371), .A(
        n21370), .ZN(n21372) );
  AOI22_X1 U23090 ( .A1(n21372), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n21421), .B2(n21519), .ZN(n21373) );
  OAI211_X1 U23091 ( .C1(n21375), .C2(n21382), .A(n21374), .B(n21373), .ZN(
        P1_U3019) );
  INV_X1 U23092 ( .A(n21509), .ZN(n21377) );
  AOI21_X1 U23093 ( .B1(n21421), .B2(n21377), .A(n21376), .ZN(n21381) );
  AOI22_X1 U23094 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21379), .B1(
        n21378), .B2(n11614), .ZN(n21380) );
  OAI211_X1 U23095 ( .C1(n21383), .C2(n21382), .A(n21381), .B(n21380), .ZN(
        P1_U3020) );
  NAND2_X1 U23096 ( .A1(n21385), .A2(n21384), .ZN(n21391) );
  AOI22_X1 U23097 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21386), .B1(
        n14073), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n21390) );
  AOI22_X1 U23098 ( .A1(n21388), .A2(n21422), .B1(n21421), .B2(n21387), .ZN(
        n21389) );
  OAI211_X1 U23099 ( .C1(n21392), .C2(n21391), .A(n21390), .B(n21389), .ZN(
        P1_U3015) );
  INV_X1 U23100 ( .A(n21405), .ZN(n21402) );
  NAND2_X1 U23101 ( .A1(n21404), .A2(n21402), .ZN(n21397) );
  AOI22_X1 U23102 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21403), .B1(
        n14073), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n21396) );
  INV_X1 U23103 ( .A(n21568), .ZN(n21393) );
  AOI22_X1 U23104 ( .A1(n21394), .A2(n21422), .B1(n21421), .B2(n21393), .ZN(
        n21395) );
  OAI211_X1 U23105 ( .C1(n21398), .C2(n21397), .A(n21396), .B(n21395), .ZN(
        P1_U3011) );
  AOI22_X1 U23106 ( .A1(n21399), .A2(n21422), .B1(n21421), .B2(n21589), .ZN(
        n21412) );
  OAI22_X1 U23107 ( .A1(n21403), .A2(n21402), .B1(n21401), .B2(n21400), .ZN(
        n21413) );
  NAND3_X1 U23108 ( .A1(n21405), .A2(n21404), .A3(n12869), .ZN(n21417) );
  AOI21_X1 U23109 ( .B1(n21413), .B2(n21417), .A(n21406), .ZN(n21410) );
  NOR3_X1 U23110 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21408), .A3(
        n21407), .ZN(n21409) );
  AOI211_X1 U23111 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14073), .A(n21410), 
        .B(n21409), .ZN(n21411) );
  NAND2_X1 U23112 ( .A1(n21412), .A2(n21411), .ZN(P1_U3009) );
  OAI22_X1 U23113 ( .A1(n21585), .A2(n21414), .B1(n21413), .B2(n12869), .ZN(
        n21415) );
  AOI21_X1 U23114 ( .B1(n21422), .B2(n21416), .A(n21415), .ZN(n21418) );
  OAI211_X1 U23115 ( .C1(n21592), .C2(n21419), .A(n21418), .B(n21417), .ZN(
        P1_U3010) );
  INV_X1 U23116 ( .A(n21616), .ZN(n21420) );
  AOI22_X1 U23117 ( .A1(n21423), .A2(n21422), .B1(n21421), .B2(n21420), .ZN(
        n21433) );
  NAND2_X1 U23118 ( .A1(n14073), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n21432) );
  NOR2_X1 U23119 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21425), .ZN(
        n21427) );
  OAI21_X1 U23120 ( .B1(n21427), .B2(n21426), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21431) );
  NAND3_X1 U23121 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21429), .A3(
        n21428), .ZN(n21430) );
  NAND4_X1 U23122 ( .A1(n21433), .A2(n21432), .A3(n21431), .A4(n21430), .ZN(
        P1_U3007) );
  AOI22_X1 U23123 ( .A1(n21627), .A2(P1_REIP_REG_0__SCAN_IN), .B1(
        P1_EBX_REG_0__SCAN_IN), .B2(n21597), .ZN(n21437) );
  NAND2_X1 U23124 ( .A1(n21626), .A2(n21613), .ZN(n21435) );
  OAI211_X1 U23125 ( .C1(n21440), .C2(n21438), .A(n21437), .B(n21436), .ZN(
        P1_U2840) );
  AOI21_X1 U23126 ( .B1(n21493), .B2(n14210), .A(n14660), .ZN(n21454) );
  AOI22_X1 U23127 ( .A1(n21439), .A2(n21590), .B1(n21597), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n21453) );
  INV_X1 U23128 ( .A(n21440), .ZN(n21474) );
  NAND2_X1 U23129 ( .A1(n21615), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n21449) );
  INV_X1 U23130 ( .A(n21441), .ZN(n21442) );
  NAND2_X1 U23131 ( .A1(n21634), .A2(n21442), .ZN(n21448) );
  INV_X1 U23132 ( .A(n21456), .ZN(n21445) );
  NAND2_X1 U23133 ( .A1(n21443), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21444) );
  OAI22_X1 U23134 ( .A1(n21877), .A2(n21445), .B1(n21484), .B2(n21444), .ZN(
        n21446) );
  INV_X1 U23135 ( .A(n21446), .ZN(n21447) );
  NAND3_X1 U23136 ( .A1(n21449), .A2(n21448), .A3(n21447), .ZN(n21450) );
  AOI21_X1 U23137 ( .B1(n21451), .B2(n21474), .A(n21450), .ZN(n21452) );
  OAI211_X1 U23138 ( .C1(n21454), .C2(n21443), .A(n21453), .B(n21452), .ZN(
        P1_U2838) );
  AOI222_X1 U23139 ( .A1(n21457), .A2(n21456), .B1(n21590), .B2(n21455), .C1(
        n21597), .C2(P1_EBX_REG_4__SCAN_IN), .ZN(n21458) );
  INV_X1 U23140 ( .A(n21458), .ZN(n21459) );
  AOI211_X1 U23141 ( .C1(n21615), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21557), .B(n21459), .ZN(n21465) );
  OAI21_X1 U23142 ( .B1(n21467), .B2(n21484), .A(n21483), .ZN(n21473) );
  OAI21_X1 U23143 ( .B1(n21484), .B2(n21461), .A(n21460), .ZN(n21462) );
  AOI22_X1 U23144 ( .A1(n21463), .A2(n21474), .B1(n21473), .B2(n21462), .ZN(
        n21464) );
  OAI211_X1 U23145 ( .C1(n21466), .C2(n21613), .A(n21465), .B(n21464), .ZN(
        P1_U2836) );
  INV_X1 U23146 ( .A(n21467), .ZN(n21468) );
  NOR3_X1 U23147 ( .A1(n21484), .A2(P1_REIP_REG_5__SCAN_IN), .A3(n21468), .ZN(
        n21469) );
  AOI21_X1 U23148 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(n21597), .A(n21469), .ZN(
        n21470) );
  OAI21_X1 U23149 ( .B1(n21638), .B2(n21471), .A(n21470), .ZN(n21472) );
  AOI211_X1 U23150 ( .C1(n21615), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n21557), .B(n21472), .ZN(n21477) );
  AOI22_X1 U23151 ( .A1(n21475), .A2(n21474), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n21473), .ZN(n21476) );
  OAI211_X1 U23152 ( .C1(n21478), .C2(n21613), .A(n21477), .B(n21476), .ZN(
        P1_U2835) );
  INV_X1 U23153 ( .A(n21479), .ZN(n21482) );
  NOR2_X1 U23154 ( .A1(n21494), .A2(n21484), .ZN(n21481) );
  AOI22_X1 U23155 ( .A1(n21482), .A2(n21481), .B1(n21590), .B2(n21480), .ZN(
        n21491) );
  OAI21_X1 U23156 ( .B1(n21494), .B2(n21484), .A(n21483), .ZN(n21501) );
  AOI22_X1 U23157 ( .A1(n21615), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n21501), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n21486) );
  OAI211_X1 U23158 ( .C1(n21623), .C2(n21487), .A(n21486), .B(n21485), .ZN(
        n21488) );
  AOI21_X1 U23159 ( .B1(n21489), .B2(n21618), .A(n21488), .ZN(n21490) );
  OAI211_X1 U23160 ( .C1(n21492), .C2(n21613), .A(n21491), .B(n21490), .ZN(
        P1_U2834) );
  NAND2_X1 U23161 ( .A1(n21494), .A2(n21493), .ZN(n21498) );
  INV_X1 U23162 ( .A(n21495), .ZN(n21496) );
  AOI22_X1 U23163 ( .A1(n21496), .A2(n21590), .B1(n21597), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n21497) );
  OAI21_X1 U23164 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n21498), .A(n21497), .ZN(
        n21499) );
  AOI211_X1 U23165 ( .C1(n21615), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n21557), .B(n21499), .ZN(n21504) );
  INV_X1 U23166 ( .A(n21500), .ZN(n21502) );
  AOI22_X1 U23167 ( .A1(n21502), .A2(n21618), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n21501), .ZN(n21503) );
  OAI211_X1 U23168 ( .C1(n21505), .C2(n21613), .A(n21504), .B(n21503), .ZN(
        P1_U2833) );
  OAI22_X1 U23169 ( .A1(n21626), .A2(n12000), .B1(n21506), .B2(n21623), .ZN(
        n21507) );
  AOI211_X1 U23170 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n21508), .A(n21557), 
        .B(n21507), .ZN(n21514) );
  OAI22_X1 U23171 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n21510), .B1(n21638), 
        .B2(n21509), .ZN(n21511) );
  AOI21_X1 U23172 ( .B1(n21618), .B2(n21512), .A(n21511), .ZN(n21513) );
  OAI211_X1 U23173 ( .C1(n21515), .C2(n21613), .A(n21514), .B(n21513), .ZN(
        P1_U2829) );
  AOI22_X1 U23174 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n21518), .B1(n21517), 
        .B2(n21516), .ZN(n21525) );
  AOI22_X1 U23175 ( .A1(n21615), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n21597), .B2(P1_EBX_REG_12__SCAN_IN), .ZN(n21524) );
  AOI21_X1 U23176 ( .B1(n21519), .B2(n21590), .A(n21557), .ZN(n21523) );
  AOI22_X1 U23177 ( .A1(n21521), .A2(n21634), .B1(n21618), .B2(n21520), .ZN(
        n21522) );
  NAND4_X1 U23178 ( .A1(n21525), .A2(n21524), .A3(n21523), .A4(n21522), .ZN(
        P1_U2828) );
  AOI22_X1 U23179 ( .A1(n21615), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n21597), .B2(P1_EBX_REG_14__SCAN_IN), .ZN(n21533) );
  AOI21_X1 U23180 ( .B1(n21526), .B2(n21590), .A(n21557), .ZN(n21532) );
  AOI22_X1 U23181 ( .A1(n21528), .A2(n21618), .B1(n21634), .B2(n21527), .ZN(
        n21531) );
  OAI211_X1 U23182 ( .C1(n21529), .C2(P1_REIP_REG_14__SCAN_IN), .A(n21627), 
        .B(n15235), .ZN(n21530) );
  NAND4_X1 U23183 ( .A1(n21533), .A2(n21532), .A3(n21531), .A4(n21530), .ZN(
        P1_U2826) );
  OAI22_X1 U23184 ( .A1(n21626), .A2(n21535), .B1(n21534), .B2(n21623), .ZN(
        n21536) );
  AOI211_X1 U23185 ( .C1(n21634), .C2(n21537), .A(n21557), .B(n21536), .ZN(
        n21544) );
  NAND2_X1 U23186 ( .A1(n21540), .A2(n21539), .ZN(n21541) );
  AOI22_X1 U23187 ( .A1(n21542), .A2(n21618), .B1(n11388), .B2(n21541), .ZN(
        n21543) );
  OAI211_X1 U23188 ( .C1(n21638), .C2(n21545), .A(n21544), .B(n21543), .ZN(
        P1_U2823) );
  AOI22_X1 U23189 ( .A1(n21634), .A2(n21546), .B1(n21597), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n21553) );
  INV_X1 U23190 ( .A(n21538), .ZN(n21547) );
  NOR2_X1 U23191 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n21547), .ZN(n21561) );
  AOI211_X1 U23192 ( .C1(n21615), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n21561), .B(n21557), .ZN(n21552) );
  AOI22_X1 U23193 ( .A1(n21548), .A2(n21618), .B1(P1_REIP_REG_18__SCAN_IN), 
        .B2(n11388), .ZN(n21551) );
  NAND2_X1 U23194 ( .A1(n21590), .A2(n21549), .ZN(n21550) );
  NAND4_X1 U23195 ( .A1(n21553), .A2(n21552), .A3(n21551), .A4(n21550), .ZN(
        P1_U2822) );
  OAI22_X1 U23196 ( .A1(n21555), .A2(n21638), .B1(n21554), .B2(n21623), .ZN(
        n21556) );
  AOI211_X1 U23197 ( .C1(n21615), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n21557), .B(n21556), .ZN(n21563) );
  OAI22_X1 U23198 ( .A1(n21559), .A2(n21630), .B1(P1_REIP_REG_19__SCAN_IN), 
        .B2(n21558), .ZN(n21560) );
  AOI221_X1 U23199 ( .B1(n11388), .B2(P1_REIP_REG_19__SCAN_IN), .C1(n21561), 
        .C2(P1_REIP_REG_19__SCAN_IN), .A(n21560), .ZN(n21562) );
  OAI211_X1 U23200 ( .C1(n21564), .C2(n21613), .A(n21563), .B(n21562), .ZN(
        P1_U2821) );
  OAI22_X1 U23201 ( .A1(n21613), .A2(n21566), .B1(n21565), .B2(n21623), .ZN(
        n21567) );
  AOI21_X1 U23202 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21615), .A(
        n21567), .ZN(n21575) );
  OAI22_X1 U23203 ( .A1(n21569), .A2(n21630), .B1(n21568), .B2(n21638), .ZN(
        n21570) );
  INV_X1 U23204 ( .A(n21570), .ZN(n21574) );
  INV_X1 U23205 ( .A(n21571), .ZN(n21572) );
  NOR2_X1 U23206 ( .A1(n21572), .A2(n21601), .ZN(n21581) );
  OAI21_X1 U23207 ( .B1(n11063), .B2(P1_REIP_REG_20__SCAN_IN), .A(n21581), 
        .ZN(n21573) );
  NAND3_X1 U23208 ( .A1(n21575), .A2(n21574), .A3(n21573), .ZN(P1_U2820) );
  NOR2_X1 U23209 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n21571), .ZN(n21579) );
  OAI22_X1 U23210 ( .A1(n21626), .A2(n21577), .B1(n21576), .B2(n21623), .ZN(
        n21578) );
  AOI211_X1 U23211 ( .C1(n21634), .C2(n21580), .A(n21579), .B(n21578), .ZN(
        n21584) );
  AOI22_X1 U23212 ( .A1(n21582), .A2(n21618), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n21581), .ZN(n21583) );
  OAI211_X1 U23213 ( .C1(n21638), .C2(n21585), .A(n21584), .B(n21583), .ZN(
        P1_U2819) );
  AOI22_X1 U23214 ( .A1(n21634), .A2(n21586), .B1(n21597), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n21596) );
  AOI22_X1 U23215 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n21615), .B1(
        n21588), .B2(n21587), .ZN(n21595) );
  AOI22_X1 U23216 ( .A1(n21591), .A2(n21618), .B1(n21590), .B2(n21589), .ZN(
        n21594) );
  OAI211_X1 U23217 ( .C1(n21571), .C2(n21592), .A(n21627), .B(
        P1_REIP_REG_22__SCAN_IN), .ZN(n21593) );
  NAND4_X1 U23218 ( .A1(n21596), .A2(n21595), .A3(n21594), .A4(n21593), .ZN(
        P1_U2818) );
  AOI22_X1 U23219 ( .A1(n21634), .A2(n21598), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n21597), .ZN(n21608) );
  INV_X1 U23220 ( .A(n21610), .ZN(n21606) );
  OAI21_X1 U23221 ( .B1(n21601), .B2(n21600), .A(n21599), .ZN(n21605) );
  OAI22_X1 U23222 ( .A1(n21603), .A2(n21630), .B1(n21638), .B2(n21602), .ZN(
        n21604) );
  AOI21_X1 U23223 ( .B1(n21606), .B2(n21605), .A(n21604), .ZN(n21607) );
  OAI211_X1 U23224 ( .C1(n21609), .C2(n21626), .A(n21608), .B(n21607), .ZN(
        P1_U2817) );
  AOI21_X1 U23225 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n21627), .A(n21610), 
        .ZN(n21622) );
  OAI22_X1 U23226 ( .A1(n21613), .A2(n21612), .B1(n21611), .B2(n21623), .ZN(
        n21614) );
  AOI21_X1 U23227 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n21615), .A(
        n21614), .ZN(n21621) );
  NOR2_X1 U23228 ( .A1(n21616), .A2(n21638), .ZN(n21617) );
  AOI21_X1 U23229 ( .B1(n21619), .B2(n21618), .A(n21617), .ZN(n21620) );
  OAI211_X1 U23230 ( .C1(n11390), .C2(n21622), .A(n21621), .B(n21620), .ZN(
        P1_U2816) );
  INV_X1 U23231 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n21625) );
  OAI22_X1 U23232 ( .A1(n21626), .A2(n21625), .B1(n21624), .B2(n21623), .ZN(
        n21633) );
  AOI21_X1 U23233 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n21627), .A(n11390), 
        .ZN(n21628) );
  OAI22_X1 U23234 ( .A1(n21631), .A2(n21630), .B1(n21629), .B2(n21628), .ZN(
        n21632) );
  AOI211_X1 U23235 ( .C1(n21635), .C2(n21634), .A(n21633), .B(n21632), .ZN(
        n21636) );
  OAI21_X1 U23236 ( .B1(n21638), .B2(n21637), .A(n21636), .ZN(P1_U2815) );
  OAI21_X1 U23237 ( .B1(n21641), .B2(n21640), .A(n21639), .ZN(P1_U2806) );
  INV_X1 U23238 ( .A(n21642), .ZN(n21644) );
  OAI22_X1 U23239 ( .A1(n21646), .A2(n21645), .B1(n21644), .B2(n21643), .ZN(
        n21648) );
  MUX2_X1 U23240 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21648), .S(
        n21647), .Z(P1_U3469) );
  AOI21_X1 U23241 ( .B1(n21651), .B2(n21650), .A(n21649), .ZN(n21653) );
  OAI211_X1 U23242 ( .C1(n21656), .C2(n21922), .A(n21653), .B(n21652), .ZN(
        P1_U3163) );
  OAI22_X1 U23243 ( .A1(n21656), .A2(n21837), .B1(n21655), .B2(n21654), .ZN(
        P1_U3466) );
  AOI21_X1 U23244 ( .B1(n21659), .B2(n21658), .A(n21657), .ZN(n21660) );
  OAI22_X1 U23245 ( .A1(n21662), .A2(n21661), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n21660), .ZN(n21663) );
  OAI21_X1 U23246 ( .B1(n21665), .B2(n21664), .A(n21663), .ZN(P1_U3161) );
  OAI21_X1 U23247 ( .B1(n21668), .B2(n14439), .A(n21666), .ZN(P1_U2805) );
  INV_X1 U23248 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21667) );
  OAI21_X1 U23249 ( .B1(n21668), .B2(n21667), .A(n21666), .ZN(P1_U3465) );
  OAI21_X1 U23250 ( .B1(n21671), .B2(n13854), .A(n21669), .ZN(P2_U2818) );
  OAI21_X1 U23251 ( .B1(n21671), .B2(n21670), .A(n21669), .ZN(P2_U3592) );
  OAI21_X1 U23252 ( .B1(n21675), .B2(n21672), .A(n21673), .ZN(P3_U2636) );
  INV_X1 U23253 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21674) );
  OAI21_X1 U23254 ( .B1(n21675), .B2(n21674), .A(n21673), .ZN(P3_U3281) );
  INV_X1 U23255 ( .A(HOLD), .ZN(n21725) );
  OAI21_X1 U23256 ( .B1(n21725), .B2(n21676), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21677) );
  INV_X1 U23257 ( .A(n21677), .ZN(n21681) );
  AOI21_X1 U23258 ( .B1(n21679), .B2(P3_STATE_REG_1__SCAN_IN), .A(n21678), 
        .ZN(n21731) );
  INV_X1 U23259 ( .A(NA), .ZN(n21727) );
  OAI21_X1 U23260 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n21727), .A(
        P3_STATE_REG_2__SCAN_IN), .ZN(n21730) );
  INV_X1 U23261 ( .A(n21730), .ZN(n21680) );
  OAI22_X1 U23262 ( .A1(n21682), .A2(n21681), .B1(n21731), .B2(n21680), .ZN(
        P3_U3029) );
  NAND4_X1 U23263 ( .A1(n21691), .A2(P1_STATE_REG_1__SCAN_IN), .A3(
        P1_REQUESTPENDING_REG_SCAN_IN), .A4(n21727), .ZN(n21689) );
  NOR2_X1 U23264 ( .A1(NA), .A2(n21683), .ZN(n21685) );
  OAI21_X1 U23265 ( .B1(n21690), .B2(n21725), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21694) );
  OAI211_X1 U23266 ( .C1(n21685), .C2(n21684), .A(HOLD), .B(n21694), .ZN(
        n21688) );
  AOI21_X1 U23267 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21691), .A(n21696), 
        .ZN(n21698) );
  INV_X1 U23268 ( .A(n21698), .ZN(n21686) );
  OAI211_X1 U23269 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n21727), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n21686), .ZN(n21687) );
  OAI221_X1 U23270 ( .B1(n21696), .B2(n21689), .C1(n21696), .C2(n21688), .A(
        n21687), .ZN(P1_U3196) );
  OAI221_X1 U23271 ( .B1(n21691), .B2(HOLD), .C1(n21691), .C2(n21690), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n21693) );
  OAI211_X1 U23272 ( .C1(n21696), .C2(n21694), .A(n21693), .B(n21692), .ZN(
        P1_U3195) );
  NOR2_X1 U23273 ( .A1(n11585), .A2(n21725), .ZN(n21695) );
  AOI211_X1 U23274 ( .C1(NA), .C2(n21696), .A(n21695), .B(n21694), .ZN(n21697)
         );
  OAI22_X1 U23275 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21698), .B1(n22279), 
        .B2(n21697), .ZN(P1_U3194) );
  NAND2_X1 U23276 ( .A1(n21699), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21710) );
  NAND2_X1 U23277 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21710), .ZN(n21709) );
  OAI22_X1 U23278 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21727), .B1(n21700), 
        .B2(n21725), .ZN(n21701) );
  AOI22_X1 U23279 ( .A1(n21713), .A2(n21709), .B1(n21702), .B2(n21701), .ZN(
        n21703) );
  OAI21_X1 U23280 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n21704), .A(n21703), .ZN(P2_U3209) );
  NAND2_X1 U23281 ( .A1(n21705), .A2(HOLD), .ZN(n21707) );
  OAI211_X1 U23282 ( .C1(n21713), .C2(n21725), .A(P2_STATE_REG_0__SCAN_IN), 
        .B(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21706) );
  NAND4_X1 U23283 ( .A1(n21708), .A2(n21707), .A3(n21710), .A4(n21706), .ZN(
        P2_U3210) );
  OAI22_X1 U23284 ( .A1(HOLD), .A2(n21709), .B1(P2_STATE_REG_0__SCAN_IN), .B2(
        n21727), .ZN(n21714) );
  OAI22_X1 U23285 ( .A1(NA), .A2(n21710), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21711) );
  OAI211_X1 U23286 ( .C1(HOLD), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n21711), .ZN(n21712) );
  OAI211_X1 U23287 ( .C1(n21714), .C2(n21713), .A(n21712), .B(n10969), .ZN(
        P2_U3211) );
  NOR2_X1 U23288 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21733)
         );
  OAI21_X1 U23289 ( .B1(n21726), .B2(n21725), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n21717) );
  NOR2_X1 U23290 ( .A1(n21723), .A2(n21715), .ZN(n21728) );
  INV_X1 U23291 ( .A(n21728), .ZN(n21716) );
  OAI21_X1 U23292 ( .B1(n21733), .B2(n21717), .A(n21716), .ZN(n21720) );
  OAI211_X1 U23293 ( .C1(n21726), .C2(n21725), .A(P3_STATE_REG_0__SCAN_IN), 
        .B(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21718) );
  AOI21_X1 U23294 ( .B1(n21718), .B2(n21721), .A(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n21719) );
  AOI21_X1 U23295 ( .B1(n21721), .B2(n21720), .A(n21719), .ZN(n21722) );
  OAI221_X1 U23296 ( .B1(n21724), .B2(P3_STATE_REG_2__SCAN_IN), .C1(n21724), 
        .C2(n21723), .A(n21722), .ZN(P3_U3030) );
  OAI22_X1 U23297 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n21726), .B2(n21725), .ZN(n21729)
         );
  OAI221_X1 U23298 ( .B1(n21729), .B2(n21728), .C1(n21729), .C2(n21727), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n21732) );
  OAI22_X1 U23299 ( .A1(n21733), .A2(n21732), .B1(n21731), .B2(n21730), .ZN(
        P3_U3031) );
  NOR2_X1 U23300 ( .A1(n21772), .A2(n21734), .ZN(n21737) );
  AOI21_X1 U23301 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n21775), .A(n21737), 
        .ZN(n21735) );
  OAI21_X1 U23302 ( .B1(n21736), .B2(n21777), .A(n21735), .ZN(P1_U2945) );
  AOI21_X1 U23303 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n21775), .A(n21737), 
        .ZN(n21738) );
  OAI21_X1 U23304 ( .B1(n14805), .B2(n21777), .A(n21738), .ZN(P1_U2960) );
  NAND2_X1 U23305 ( .A1(n21740), .A2(n21739), .ZN(n21745) );
  INV_X1 U23306 ( .A(n21745), .ZN(n21741) );
  AOI21_X1 U23307 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n21775), .A(n21741), 
        .ZN(n21742) );
  OAI21_X1 U23308 ( .B1(n21743), .B2(n21777), .A(n21742), .ZN(P1_U2946) );
  AOI22_X1 U23309 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21775), .B1(n21744), 
        .B2(P1_EAX_REG_9__SCAN_IN), .ZN(n21746) );
  NAND2_X1 U23310 ( .A1(n21746), .A2(n21745), .ZN(P1_U2961) );
  NOR2_X1 U23311 ( .A1(n21772), .A2(n21747), .ZN(n21750) );
  AOI21_X1 U23312 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n21775), .A(n21750), 
        .ZN(n21748) );
  OAI21_X1 U23313 ( .B1(n21749), .B2(n21777), .A(n21748), .ZN(P1_U2947) );
  AOI21_X1 U23314 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n21775), .A(n21750), 
        .ZN(n21751) );
  OAI21_X1 U23315 ( .B1(n14939), .B2(n21777), .A(n21751), .ZN(P1_U2962) );
  NOR2_X1 U23316 ( .A1(n21772), .A2(n21752), .ZN(n21755) );
  AOI21_X1 U23317 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n21775), .A(n21755), 
        .ZN(n21753) );
  OAI21_X1 U23318 ( .B1(n21754), .B2(n21777), .A(n21753), .ZN(P1_U2948) );
  AOI21_X1 U23319 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(n21775), .A(n21755), 
        .ZN(n21756) );
  OAI21_X1 U23320 ( .B1(n15168), .B2(n21777), .A(n21756), .ZN(P1_U2963) );
  INV_X1 U23321 ( .A(n21757), .ZN(n21758) );
  NOR2_X1 U23322 ( .A1(n21772), .A2(n21758), .ZN(n21760) );
  AOI21_X1 U23323 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n21775), .A(n21760), 
        .ZN(n21759) );
  OAI21_X1 U23324 ( .B1(n15730), .B2(n21777), .A(n21759), .ZN(P1_U2949) );
  AOI21_X1 U23325 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n21775), .A(n21760), 
        .ZN(n21761) );
  OAI21_X1 U23326 ( .B1(n21762), .B2(n21777), .A(n21761), .ZN(P1_U2964) );
  INV_X1 U23327 ( .A(n21763), .ZN(n21764) );
  NOR2_X1 U23328 ( .A1(n21772), .A2(n21764), .ZN(n21767) );
  AOI21_X1 U23329 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n21775), .A(n21767), 
        .ZN(n21765) );
  OAI21_X1 U23330 ( .B1(n21766), .B2(n21777), .A(n21765), .ZN(P1_U2950) );
  AOI21_X1 U23331 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n21775), .A(n21767), 
        .ZN(n21768) );
  OAI21_X1 U23332 ( .B1(n21769), .B2(n21777), .A(n21768), .ZN(P1_U2965) );
  INV_X1 U23333 ( .A(n21770), .ZN(n21771) );
  NOR2_X1 U23334 ( .A1(n21772), .A2(n21771), .ZN(n21774) );
  AOI21_X1 U23335 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n21775), .A(n21774), 
        .ZN(n21773) );
  OAI21_X1 U23336 ( .B1(n12760), .B2(n21777), .A(n21773), .ZN(P1_U2951) );
  AOI21_X1 U23337 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(n21775), .A(n21774), 
        .ZN(n21776) );
  OAI21_X1 U23338 ( .B1(n21778), .B2(n21777), .A(n21776), .ZN(P1_U2966) );
  INV_X1 U23339 ( .A(n21868), .ZN(n21779) );
  NAND2_X1 U23340 ( .A1(n22270), .A2(n21900), .ZN(n21780) );
  NAND2_X1 U23341 ( .A1(n21900), .A2(n14439), .ZN(n21847) );
  OAI21_X1 U23342 ( .B1(n22189), .B2(n21780), .A(n21847), .ZN(n21786) );
  INV_X1 U23343 ( .A(n21877), .ZN(n21781) );
  OR2_X1 U23344 ( .A1(n21829), .A2(n21781), .ZN(n21798) );
  NOR2_X1 U23345 ( .A1(n21798), .A2(n21906), .ZN(n21784) );
  AOI22_X1 U23346 ( .A1(n21786), .A2(n21784), .B1(n11386), .B2(n21850), .ZN(
        n22186) );
  NAND3_X1 U23347 ( .A1(n11834), .A2(n16851), .A3(n21880), .ZN(n21791) );
  INV_X1 U23348 ( .A(n21791), .ZN(n21794) );
  NAND2_X1 U23349 ( .A1(n21892), .A2(n21794), .ZN(n22181) );
  OAI22_X1 U23350 ( .A1(n22270), .A2(n21938), .B1(n21852), .B2(n22181), .ZN(
        n21782) );
  INV_X1 U23351 ( .A(n21782), .ZN(n21789) );
  INV_X1 U23352 ( .A(n21784), .ZN(n21785) );
  AOI22_X1 U23353 ( .A1(n21786), .A2(n21785), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22181), .ZN(n21787) );
  OAI211_X1 U23354 ( .C1(n11386), .C2(n21922), .A(n21858), .B(n21787), .ZN(
        n22183) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22183), .B1(
        n22189), .B2(n21881), .ZN(n21788) );
  OAI211_X1 U23356 ( .C1(n22186), .C2(n21889), .A(n21789), .B(n21788), .ZN(
        P1_U3033) );
  INV_X1 U23357 ( .A(n21807), .ZN(n21790) );
  INV_X1 U23358 ( .A(n21798), .ZN(n21806) );
  NOR2_X1 U23359 ( .A1(n21892), .A2(n21791), .ZN(n22187) );
  AOI21_X1 U23360 ( .B1(n21806), .B2(n21893), .A(n22187), .ZN(n21792) );
  OAI22_X1 U23361 ( .A1(n21792), .A2(n21924), .B1(n21791), .B2(n21922), .ZN(
        n22188) );
  INV_X1 U23362 ( .A(n21889), .ZN(n21926) );
  AOI22_X1 U23363 ( .A1(n22188), .A2(n21926), .B1(n21925), .B2(n22187), .ZN(
        n21796) );
  OAI211_X1 U23364 ( .C1(n21807), .C2(n14439), .A(n21900), .B(n21792), .ZN(
        n21793) );
  OAI211_X1 U23365 ( .C1(n21900), .C2(n21794), .A(n21898), .B(n21793), .ZN(
        n22190) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22190), .B1(
        n22189), .B2(n21916), .ZN(n21795) );
  OAI211_X1 U23367 ( .C1(n21934), .C2(n22193), .A(n21796), .B(n21795), .ZN(
        P1_U3041) );
  NAND2_X1 U23368 ( .A1(n22193), .A2(n21900), .ZN(n21797) );
  OAI21_X1 U23369 ( .B1(n21797), .B2(n22201), .A(n21847), .ZN(n21800) );
  NOR2_X1 U23370 ( .A1(n21798), .A2(n14662), .ZN(n21802) );
  NOR2_X1 U23371 ( .A1(n21830), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21818) );
  AOI22_X1 U23372 ( .A1(n21800), .A2(n21802), .B1(n21850), .B2(n21818), .ZN(
        n22199) );
  NAND3_X1 U23373 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n11834), .A3(
        n16851), .ZN(n21810) );
  NOR2_X1 U23374 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21810), .ZN(
        n22194) );
  INV_X1 U23375 ( .A(n22194), .ZN(n22143) );
  OAI22_X1 U23376 ( .A1(n22193), .A2(n21938), .B1(n21852), .B2(n22143), .ZN(
        n21799) );
  INV_X1 U23377 ( .A(n21799), .ZN(n21805) );
  INV_X1 U23378 ( .A(n21800), .ZN(n21803) );
  NOR2_X1 U23379 ( .A1(n21818), .A2(n21922), .ZN(n21821) );
  AOI21_X1 U23380 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22143), .A(n21821), 
        .ZN(n21801) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22196), .B1(
        n22201), .B2(n21881), .ZN(n21804) );
  OAI211_X1 U23382 ( .C1(n22199), .C2(n21889), .A(n21805), .B(n21804), .ZN(
        P1_U3049) );
  NOR2_X1 U23383 ( .A1(n21892), .A2(n21810), .ZN(n22200) );
  AOI21_X1 U23384 ( .B1(n21806), .B2(n10998), .A(n22200), .ZN(n21809) );
  AOI21_X1 U23385 ( .B1(n21807), .B2(n21900), .A(n21862), .ZN(n21813) );
  OAI22_X1 U23386 ( .A1(n21922), .A2(n21810), .B1(n21809), .B2(n21813), .ZN(
        n21808) );
  AOI22_X1 U23387 ( .A1(n22201), .A2(n21916), .B1(n21925), .B2(n22200), .ZN(
        n21815) );
  INV_X1 U23388 ( .A(n21809), .ZN(n21812) );
  AOI21_X1 U23389 ( .B1(n21924), .B2(n21810), .A(n21928), .ZN(n21811) );
  OAI21_X1 U23390 ( .B1(n21813), .B2(n21812), .A(n21811), .ZN(n22203) );
  AOI22_X1 U23391 ( .A1(n22203), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n22202), .B2(n21881), .ZN(n21814) );
  OAI211_X1 U23392 ( .C1(n22206), .C2(n21889), .A(n21815), .B(n21814), .ZN(
        P1_U3057) );
  NOR2_X1 U23393 ( .A1(n22210), .A2(n21924), .ZN(n21816) );
  INV_X1 U23394 ( .A(n21847), .ZN(n21873) );
  AOI21_X1 U23395 ( .B1(n21816), .B2(n22208), .A(n21873), .ZN(n21824) );
  INV_X1 U23396 ( .A(n21824), .ZN(n21819) );
  AND2_X1 U23397 ( .A1(n21817), .A2(n21906), .ZN(n21823) );
  OR3_X1 U23398 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n21921), .ZN(n22207) );
  OAI22_X1 U23399 ( .A1(n22067), .A2(n21934), .B1(n21852), .B2(n22207), .ZN(
        n21820) );
  INV_X1 U23400 ( .A(n21820), .ZN(n21826) );
  AOI21_X1 U23401 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22207), .A(n21821), 
        .ZN(n21822) );
  OAI211_X1 U23402 ( .C1(n21824), .C2(n21823), .A(n21914), .B(n21822), .ZN(
        n22211) );
  AOI22_X1 U23403 ( .A1(n22211), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n21916), .B2(n22069), .ZN(n21825) );
  OAI211_X1 U23404 ( .C1(n22214), .C2(n21889), .A(n21826), .B(n21825), .ZN(
        P1_U3081) );
  INV_X1 U23405 ( .A(n21869), .ZN(n21828) );
  AND2_X1 U23406 ( .A1(n21829), .A2(n21877), .ZN(n21861) );
  NAND3_X1 U23407 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16851), .A3(
        n21880), .ZN(n21840) );
  NOR2_X1 U23408 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21840), .ZN(
        n22215) );
  AOI21_X1 U23409 ( .B1(n21861), .B2(n14662), .A(n22215), .ZN(n21834) );
  NAND2_X1 U23410 ( .A1(n21831), .A2(n21830), .ZN(n21883) );
  INV_X1 U23411 ( .A(n21850), .ZN(n21832) );
  OAI22_X1 U23412 ( .A1(n21834), .A2(n21924), .B1(n21883), .B2(n21832), .ZN(
        n22216) );
  AOI22_X1 U23413 ( .A1(n22216), .A2(n21926), .B1(n21925), .B2(n22215), .ZN(
        n21839) );
  INV_X1 U23414 ( .A(n22226), .ZN(n21833) );
  OAI21_X1 U23415 ( .B1(n21833), .B2(n22217), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21835) );
  NAND2_X1 U23416 ( .A1(n21835), .A2(n21834), .ZN(n21836) );
  AOI22_X1 U23417 ( .A1(n22218), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n21916), .B2(n22217), .ZN(n21838) );
  OAI211_X1 U23418 ( .C1(n21934), .C2(n22226), .A(n21839), .B(n21838), .ZN(
        P1_U3097) );
  NOR2_X1 U23419 ( .A1(n21892), .A2(n21840), .ZN(n22221) );
  AOI21_X1 U23420 ( .B1(n21861), .B2(n21893), .A(n22221), .ZN(n21841) );
  OAI22_X1 U23421 ( .A1(n21841), .A2(n21924), .B1(n21840), .B2(n21922), .ZN(
        n22222) );
  AOI22_X1 U23422 ( .A1(n22222), .A2(n21926), .B1(n21925), .B2(n22221), .ZN(
        n21846) );
  INV_X1 U23423 ( .A(n21840), .ZN(n21843) );
  OAI211_X1 U23424 ( .C1(n21869), .C2(n14439), .A(n21900), .B(n21841), .ZN(
        n21842) );
  OAI211_X1 U23425 ( .C1(n21900), .C2(n21843), .A(n21898), .B(n21842), .ZN(
        n22223) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22223), .B1(
        n22230), .B2(n21881), .ZN(n21845) );
  OAI211_X1 U23427 ( .C1(n21938), .C2(n22226), .A(n21846), .B(n21845), .ZN(
        P1_U3105) );
  NAND3_X1 U23428 ( .A1(n22240), .A2(n22157), .A3(n21900), .ZN(n21848) );
  NAND2_X1 U23429 ( .A1(n21848), .A2(n21847), .ZN(n21856) );
  AND2_X1 U23430 ( .A1(n21861), .A2(n21906), .ZN(n21854) );
  NAND2_X1 U23431 ( .A1(n21849), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21908) );
  INV_X1 U23432 ( .A(n21908), .ZN(n21851) );
  NAND3_X1 U23433 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n16851), .ZN(n21864) );
  OR2_X1 U23434 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21864), .ZN(
        n22227) );
  OAI22_X1 U23435 ( .A1(n22240), .A2(n21934), .B1(n21852), .B2(n22227), .ZN(
        n21853) );
  INV_X1 U23436 ( .A(n21853), .ZN(n21860) );
  INV_X1 U23437 ( .A(n21854), .ZN(n21855) );
  AOI22_X1 U23438 ( .A1(n21856), .A2(n21855), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22227), .ZN(n21857) );
  NAND2_X1 U23439 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21908), .ZN(n21913) );
  NAND3_X1 U23440 ( .A1(n21858), .A2(n21857), .A3(n21913), .ZN(n22231) );
  AOI22_X1 U23441 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22231), .B1(
        n22230), .B2(n21916), .ZN(n21859) );
  OAI211_X1 U23442 ( .C1(n22234), .C2(n21889), .A(n21860), .B(n21859), .ZN(
        P1_U3113) );
  NOR2_X1 U23443 ( .A1(n21892), .A2(n21864), .ZN(n22235) );
  AOI21_X1 U23444 ( .B1(n21861), .B2(n10998), .A(n22235), .ZN(n21863) );
  OAI22_X1 U23445 ( .A1(n21863), .A2(n21924), .B1(n21864), .B2(n21922), .ZN(
        n22236) );
  AOI22_X1 U23446 ( .A1(n22236), .A2(n21926), .B1(n21925), .B2(n22235), .ZN(
        n21871) );
  AOI21_X1 U23447 ( .B1(n21869), .B2(n21900), .A(n21862), .ZN(n21867) );
  INV_X1 U23448 ( .A(n21863), .ZN(n21866) );
  AOI21_X1 U23449 ( .B1(n21924), .B2(n21864), .A(n21928), .ZN(n21865) );
  OAI21_X1 U23450 ( .B1(n21867), .B2(n21866), .A(n21865), .ZN(n22237) );
  AOI22_X1 U23451 ( .A1(n22237), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n21881), .B2(n22243), .ZN(n21870) );
  OAI211_X1 U23452 ( .C1(n21938), .C2(n22240), .A(n21871), .B(n21870), .ZN(
        P1_U3121) );
  NOR2_X1 U23453 ( .A1(n22251), .A2(n21924), .ZN(n21875) );
  AOI21_X1 U23454 ( .B1(n21875), .B2(n21874), .A(n21873), .ZN(n21886) );
  INV_X1 U23455 ( .A(n21886), .ZN(n21879) );
  OR2_X1 U23456 ( .A1(n21877), .A2(n21876), .ZN(n21891) );
  NOR2_X1 U23457 ( .A1(n21891), .A2(n21906), .ZN(n21885) );
  INV_X1 U23458 ( .A(n21883), .ZN(n21878) );
  NAND3_X1 U23459 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n21880), .ZN(n21894) );
  NOR2_X1 U23460 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21894), .ZN(
        n22241) );
  AOI22_X1 U23461 ( .A1(n22251), .A2(n21881), .B1(n21925), .B2(n22241), .ZN(
        n21888) );
  INV_X1 U23462 ( .A(n22241), .ZN(n21882) );
  AOI22_X1 U23463 ( .A1(n21883), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n21882), .ZN(n21884) );
  OAI211_X1 U23464 ( .C1(n21886), .C2(n21885), .A(n21914), .B(n21884), .ZN(
        n22244) );
  AOI22_X1 U23465 ( .A1(n22244), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n21916), .B2(n22243), .ZN(n21887) );
  OAI211_X1 U23466 ( .C1(n22248), .C2(n21889), .A(n21888), .B(n21887), .ZN(
        P1_U3129) );
  INV_X1 U23467 ( .A(n21891), .ZN(n21920) );
  NOR2_X1 U23468 ( .A1(n21892), .A2(n21894), .ZN(n22249) );
  AOI21_X1 U23469 ( .B1(n21920), .B2(n21893), .A(n22249), .ZN(n21895) );
  OAI22_X1 U23470 ( .A1(n21895), .A2(n21924), .B1(n21894), .B2(n21922), .ZN(
        n22250) );
  AOI22_X1 U23471 ( .A1(n21926), .A2(n22250), .B1(n21925), .B2(n22249), .ZN(
        n21902) );
  INV_X1 U23472 ( .A(n21894), .ZN(n21899) );
  INV_X1 U23473 ( .A(n21905), .ZN(n21896) );
  OAI211_X1 U23474 ( .C1(n21896), .C2(n14439), .A(n21900), .B(n21895), .ZN(
        n21897) );
  OAI211_X1 U23475 ( .C1(n21900), .C2(n21899), .A(n21898), .B(n21897), .ZN(
        n22252) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22252), .B1(
        n22251), .B2(n21916), .ZN(n21901) );
  OAI211_X1 U23477 ( .C1(n21934), .C2(n22255), .A(n21902), .B(n21901), .ZN(
        P1_U3137) );
  INV_X1 U23478 ( .A(n21903), .ZN(n21904) );
  NOR3_X2 U23479 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11834), .A3(
        n21921), .ZN(n22257) );
  NAND2_X1 U23480 ( .A1(n21920), .A2(n21906), .ZN(n21911) );
  INV_X1 U23481 ( .A(n21907), .ZN(n21909) );
  OAI22_X1 U23482 ( .A1(n21911), .A2(n21924), .B1(n21909), .B2(n21908), .ZN(
        n22256) );
  AOI22_X1 U23483 ( .A1(n21925), .A2(n22257), .B1(n21926), .B2(n22256), .ZN(
        n21918) );
  INV_X1 U23484 ( .A(n22274), .ZN(n21910) );
  OAI21_X1 U23485 ( .B1(n22259), .B2(n21910), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21912) );
  AOI21_X1 U23486 ( .B1(n21912), .B2(n21911), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21915) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22260), .B1(
        n22259), .B2(n21916), .ZN(n21917) );
  OAI211_X1 U23488 ( .C1(n21934), .C2(n22274), .A(n21918), .B(n21917), .ZN(
        P1_U3145) );
  NOR2_X1 U23489 ( .A1(n21919), .A2(n11834), .ZN(n22263) );
  AOI21_X1 U23490 ( .B1(n21920), .B2(n10998), .A(n22263), .ZN(n21930) );
  NOR2_X1 U23491 ( .A1(n11834), .A2(n21921), .ZN(n21927) );
  INV_X1 U23492 ( .A(n21927), .ZN(n21923) );
  OAI22_X1 U23493 ( .A1(n21930), .A2(n21924), .B1(n21923), .B2(n21922), .ZN(
        n22266) );
  AOI22_X1 U23494 ( .A1(n22266), .A2(n21926), .B1(n21925), .B2(n22263), .ZN(
        n21937) );
  OR2_X1 U23495 ( .A1(n21900), .A2(n21927), .ZN(n21932) );
  AOI21_X1 U23496 ( .B1(n21930), .B2(n21929), .A(n21928), .ZN(n21931) );
  INV_X1 U23497 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n21933) );
  OAI22_X1 U23498 ( .A1(n22270), .A2(n21934), .B1(n22268), .B2(n21933), .ZN(
        n21935) );
  INV_X1 U23499 ( .A(n21935), .ZN(n21936) );
  OAI211_X1 U23500 ( .C1(n21938), .C2(n22274), .A(n21937), .B(n21936), .ZN(
        P1_U3153) );
  OAI22_X1 U23501 ( .A1(n22270), .A2(n21978), .B1(n21956), .B2(n22181), .ZN(
        n21939) );
  INV_X1 U23502 ( .A(n21939), .ZN(n21941) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22183), .B1(
        n22189), .B2(n21962), .ZN(n21940) );
  OAI211_X1 U23504 ( .C1(n22186), .C2(n21965), .A(n21941), .B(n21940), .ZN(
        P1_U3034) );
  INV_X1 U23505 ( .A(n21962), .ZN(n21974) );
  INV_X1 U23506 ( .A(n21965), .ZN(n21972) );
  AOI22_X1 U23507 ( .A1(n22188), .A2(n21972), .B1(n21971), .B2(n22187), .ZN(
        n21943) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22190), .B1(
        n22189), .B2(n21968), .ZN(n21942) );
  OAI211_X1 U23509 ( .C1(n21974), .C2(n22193), .A(n21943), .B(n21942), .ZN(
        P1_U3042) );
  OAI22_X1 U23510 ( .A1(n22193), .A2(n21978), .B1(n21956), .B2(n22143), .ZN(
        n21944) );
  INV_X1 U23511 ( .A(n21944), .ZN(n21946) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n22196), .B1(
        n22201), .B2(n21962), .ZN(n21945) );
  OAI211_X1 U23513 ( .C1(n22199), .C2(n21965), .A(n21946), .B(n21945), .ZN(
        P1_U3050) );
  AOI22_X1 U23514 ( .A1(n22202), .A2(n21962), .B1(n21971), .B2(n22200), .ZN(
        n21948) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22203), .B1(
        n22201), .B2(n21968), .ZN(n21947) );
  OAI211_X1 U23516 ( .C1(n22206), .C2(n21965), .A(n21948), .B(n21947), .ZN(
        P1_U3058) );
  OAI22_X1 U23517 ( .A1(n22067), .A2(n21974), .B1(n21956), .B2(n22207), .ZN(
        n21949) );
  INV_X1 U23518 ( .A(n21949), .ZN(n21951) );
  AOI22_X1 U23519 ( .A1(n22211), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n21968), .B2(n22069), .ZN(n21950) );
  OAI211_X1 U23520 ( .C1(n22214), .C2(n21965), .A(n21951), .B(n21950), .ZN(
        P1_U3082) );
  AOI22_X1 U23521 ( .A1(n22216), .A2(n21972), .B1(n21971), .B2(n22215), .ZN(
        n21953) );
  AOI22_X1 U23522 ( .A1(n22218), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n21968), .B2(n22217), .ZN(n21952) );
  OAI211_X1 U23523 ( .C1(n21974), .C2(n22226), .A(n21953), .B(n21952), .ZN(
        P1_U3098) );
  AOI22_X1 U23524 ( .A1(n22222), .A2(n21972), .B1(n21971), .B2(n22221), .ZN(
        n21955) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22223), .B1(
        n22230), .B2(n21962), .ZN(n21954) );
  OAI211_X1 U23526 ( .C1(n21978), .C2(n22226), .A(n21955), .B(n21954), .ZN(
        P1_U3106) );
  OAI22_X1 U23527 ( .A1(n22157), .A2(n21978), .B1(n21956), .B2(n22227), .ZN(
        n21957) );
  INV_X1 U23528 ( .A(n21957), .ZN(n21959) );
  INV_X1 U23529 ( .A(n22240), .ZN(n22159) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22231), .B1(
        n22159), .B2(n21962), .ZN(n21958) );
  OAI211_X1 U23531 ( .C1(n22234), .C2(n21965), .A(n21959), .B(n21958), .ZN(
        P1_U3114) );
  AOI22_X1 U23532 ( .A1(n22236), .A2(n21972), .B1(n21971), .B2(n22235), .ZN(
        n21961) );
  AOI22_X1 U23533 ( .A1(n22237), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n21962), .B2(n22243), .ZN(n21960) );
  OAI211_X1 U23534 ( .C1(n21978), .C2(n22240), .A(n21961), .B(n21960), .ZN(
        P1_U3122) );
  AOI22_X1 U23535 ( .A1(n22251), .A2(n21962), .B1(n21971), .B2(n22241), .ZN(
        n21964) );
  AOI22_X1 U23536 ( .A1(n22244), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n21968), .B2(n22243), .ZN(n21963) );
  OAI211_X1 U23537 ( .C1(n22248), .C2(n21965), .A(n21964), .B(n21963), .ZN(
        P1_U3130) );
  AOI22_X1 U23538 ( .A1(n21972), .A2(n22250), .B1(n21971), .B2(n22249), .ZN(
        n21967) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22252), .B1(
        n22251), .B2(n21968), .ZN(n21966) );
  OAI211_X1 U23540 ( .C1(n21974), .C2(n22255), .A(n21967), .B(n21966), .ZN(
        P1_U3138) );
  AOI22_X1 U23541 ( .A1(n21971), .A2(n22257), .B1(n21972), .B2(n22256), .ZN(
        n21970) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22260), .B1(
        n22259), .B2(n21968), .ZN(n21969) );
  OAI211_X1 U23543 ( .C1(n21974), .C2(n22274), .A(n21970), .B(n21969), .ZN(
        P1_U3146) );
  AOI22_X1 U23544 ( .A1(n22266), .A2(n21972), .B1(n21971), .B2(n22263), .ZN(
        n21977) );
  INV_X1 U23545 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n21973) );
  OAI22_X1 U23546 ( .A1(n22270), .A2(n21974), .B1(n22268), .B2(n21973), .ZN(
        n21975) );
  INV_X1 U23547 ( .A(n21975), .ZN(n21976) );
  OAI211_X1 U23548 ( .C1(n21978), .C2(n22274), .A(n21977), .B(n21976), .ZN(
        P1_U3154) );
  OAI22_X1 U23549 ( .A1(n22270), .A2(n22017), .B1(n21995), .B2(n22181), .ZN(
        n21979) );
  INV_X1 U23550 ( .A(n21979), .ZN(n21981) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22183), .B1(
        n22189), .B2(n22001), .ZN(n21980) );
  OAI211_X1 U23552 ( .C1(n22186), .C2(n22004), .A(n21981), .B(n21980), .ZN(
        P1_U3035) );
  INV_X1 U23553 ( .A(n22001), .ZN(n22013) );
  INV_X1 U23554 ( .A(n22004), .ZN(n22011) );
  AOI22_X1 U23555 ( .A1(n22188), .A2(n22011), .B1(n22010), .B2(n22187), .ZN(
        n21983) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22190), .B1(
        n22189), .B2(n22007), .ZN(n21982) );
  OAI211_X1 U23557 ( .C1(n22013), .C2(n22193), .A(n21983), .B(n21982), .ZN(
        P1_U3043) );
  AOI22_X1 U23558 ( .A1(n22201), .A2(n22001), .B1(n22010), .B2(n22194), .ZN(
        n21985) );
  INV_X1 U23559 ( .A(n22193), .ZN(n22195) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22196), .B1(
        n22195), .B2(n22007), .ZN(n21984) );
  OAI211_X1 U23561 ( .C1(n22199), .C2(n22004), .A(n21985), .B(n21984), .ZN(
        P1_U3051) );
  AOI22_X1 U23562 ( .A1(n22201), .A2(n22007), .B1(n22010), .B2(n22200), .ZN(
        n21987) );
  AOI22_X1 U23563 ( .A1(n22203), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n22202), .B2(n22001), .ZN(n21986) );
  OAI211_X1 U23564 ( .C1(n22206), .C2(n22004), .A(n21987), .B(n21986), .ZN(
        P1_U3059) );
  OAI22_X1 U23565 ( .A1(n22208), .A2(n22017), .B1(n21995), .B2(n22207), .ZN(
        n21988) );
  INV_X1 U23566 ( .A(n21988), .ZN(n21990) );
  AOI22_X1 U23567 ( .A1(n22211), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n22001), .B2(n22210), .ZN(n21989) );
  OAI211_X1 U23568 ( .C1(n22214), .C2(n22004), .A(n21990), .B(n21989), .ZN(
        P1_U3083) );
  AOI22_X1 U23569 ( .A1(n22216), .A2(n22011), .B1(n22010), .B2(n22215), .ZN(
        n21992) );
  AOI22_X1 U23570 ( .A1(n22218), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n22007), .B2(n22217), .ZN(n21991) );
  OAI211_X1 U23571 ( .C1(n22013), .C2(n22226), .A(n21992), .B(n21991), .ZN(
        P1_U3099) );
  AOI22_X1 U23572 ( .A1(n22222), .A2(n22011), .B1(n22010), .B2(n22221), .ZN(
        n21994) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22223), .B1(
        n22230), .B2(n22001), .ZN(n21993) );
  OAI211_X1 U23574 ( .C1(n22017), .C2(n22226), .A(n21994), .B(n21993), .ZN(
        P1_U3107) );
  OAI22_X1 U23575 ( .A1(n22157), .A2(n22017), .B1(n21995), .B2(n22227), .ZN(
        n21996) );
  INV_X1 U23576 ( .A(n21996), .ZN(n21998) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22231), .B1(
        n22159), .B2(n22001), .ZN(n21997) );
  OAI211_X1 U23578 ( .C1(n22234), .C2(n22004), .A(n21998), .B(n21997), .ZN(
        P1_U3115) );
  AOI22_X1 U23579 ( .A1(n22236), .A2(n22011), .B1(n22010), .B2(n22235), .ZN(
        n22000) );
  AOI22_X1 U23580 ( .A1(n22237), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n22001), .B2(n22243), .ZN(n21999) );
  OAI211_X1 U23581 ( .C1(n22017), .C2(n22240), .A(n22000), .B(n21999), .ZN(
        P1_U3123) );
  AOI22_X1 U23582 ( .A1(n22251), .A2(n22001), .B1(n22010), .B2(n22241), .ZN(
        n22003) );
  AOI22_X1 U23583 ( .A1(n22244), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n22007), .B2(n22243), .ZN(n22002) );
  OAI211_X1 U23584 ( .C1(n22248), .C2(n22004), .A(n22003), .B(n22002), .ZN(
        P1_U3131) );
  AOI22_X1 U23585 ( .A1(n22011), .A2(n22250), .B1(n22010), .B2(n22249), .ZN(
        n22006) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22252), .B1(
        n22251), .B2(n22007), .ZN(n22005) );
  OAI211_X1 U23587 ( .C1(n22013), .C2(n22255), .A(n22006), .B(n22005), .ZN(
        P1_U3139) );
  AOI22_X1 U23588 ( .A1(n22010), .A2(n22257), .B1(n22011), .B2(n22256), .ZN(
        n22009) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22260), .B1(
        n22259), .B2(n22007), .ZN(n22008) );
  OAI211_X1 U23590 ( .C1(n22013), .C2(n22274), .A(n22009), .B(n22008), .ZN(
        P1_U3147) );
  AOI22_X1 U23591 ( .A1(n22266), .A2(n22011), .B1(n22010), .B2(n22263), .ZN(
        n22016) );
  INV_X1 U23592 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n22012) );
  OAI22_X1 U23593 ( .A1(n22270), .A2(n22013), .B1(n22268), .B2(n22012), .ZN(
        n22014) );
  INV_X1 U23594 ( .A(n22014), .ZN(n22015) );
  OAI211_X1 U23595 ( .C1(n22017), .C2(n22274), .A(n22016), .B(n22015), .ZN(
        P1_U3155) );
  OAI22_X1 U23596 ( .A1(n22270), .A2(n22056), .B1(n22034), .B2(n22181), .ZN(
        n22018) );
  INV_X1 U23597 ( .A(n22018), .ZN(n22020) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22183), .B1(
        n22189), .B2(n22040), .ZN(n22019) );
  OAI211_X1 U23599 ( .C1(n22186), .C2(n22043), .A(n22020), .B(n22019), .ZN(
        P1_U3036) );
  INV_X1 U23600 ( .A(n22040), .ZN(n22052) );
  INV_X1 U23601 ( .A(n22043), .ZN(n22050) );
  AOI22_X1 U23602 ( .A1(n22188), .A2(n22050), .B1(n22049), .B2(n22187), .ZN(
        n22022) );
  AOI22_X1 U23603 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n22190), .B1(
        n22189), .B2(n22046), .ZN(n22021) );
  OAI211_X1 U23604 ( .C1(n22052), .C2(n22193), .A(n22022), .B(n22021), .ZN(
        P1_U3044) );
  AOI22_X1 U23605 ( .A1(n22201), .A2(n22040), .B1(n22049), .B2(n22194), .ZN(
        n22024) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22196), .B1(
        n22195), .B2(n22046), .ZN(n22023) );
  OAI211_X1 U23607 ( .C1(n22199), .C2(n22043), .A(n22024), .B(n22023), .ZN(
        P1_U3052) );
  AOI22_X1 U23608 ( .A1(n22202), .A2(n22040), .B1(n22049), .B2(n22200), .ZN(
        n22026) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n22203), .B1(
        n22201), .B2(n22046), .ZN(n22025) );
  OAI211_X1 U23610 ( .C1(n22206), .C2(n22043), .A(n22026), .B(n22025), .ZN(
        P1_U3060) );
  OAI22_X1 U23611 ( .A1(n22208), .A2(n22056), .B1(n22034), .B2(n22207), .ZN(
        n22027) );
  INV_X1 U23612 ( .A(n22027), .ZN(n22029) );
  AOI22_X1 U23613 ( .A1(n22211), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22040), .B2(n22210), .ZN(n22028) );
  OAI211_X1 U23614 ( .C1(n22214), .C2(n22043), .A(n22029), .B(n22028), .ZN(
        P1_U3084) );
  AOI22_X1 U23615 ( .A1(n22216), .A2(n22050), .B1(n22049), .B2(n22215), .ZN(
        n22031) );
  AOI22_X1 U23616 ( .A1(n22218), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n22046), .B2(n22217), .ZN(n22030) );
  OAI211_X1 U23617 ( .C1(n22052), .C2(n22226), .A(n22031), .B(n22030), .ZN(
        P1_U3100) );
  AOI22_X1 U23618 ( .A1(n22222), .A2(n22050), .B1(n22049), .B2(n22221), .ZN(
        n22033) );
  AOI22_X1 U23619 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n22223), .B1(
        n22230), .B2(n22040), .ZN(n22032) );
  OAI211_X1 U23620 ( .C1(n22056), .C2(n22226), .A(n22033), .B(n22032), .ZN(
        P1_U3108) );
  OAI22_X1 U23621 ( .A1(n22240), .A2(n22052), .B1(n22034), .B2(n22227), .ZN(
        n22035) );
  INV_X1 U23622 ( .A(n22035), .ZN(n22037) );
  AOI22_X1 U23623 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n22231), .B1(
        n22230), .B2(n22046), .ZN(n22036) );
  OAI211_X1 U23624 ( .C1(n22234), .C2(n22043), .A(n22037), .B(n22036), .ZN(
        P1_U3116) );
  AOI22_X1 U23625 ( .A1(n22236), .A2(n22050), .B1(n22049), .B2(n22235), .ZN(
        n22039) );
  AOI22_X1 U23626 ( .A1(n22237), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n22040), .B2(n22243), .ZN(n22038) );
  OAI211_X1 U23627 ( .C1(n22056), .C2(n22240), .A(n22039), .B(n22038), .ZN(
        P1_U3124) );
  AOI22_X1 U23628 ( .A1(n22251), .A2(n22040), .B1(n22049), .B2(n22241), .ZN(
        n22042) );
  AOI22_X1 U23629 ( .A1(n22244), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22046), .B2(n22243), .ZN(n22041) );
  OAI211_X1 U23630 ( .C1(n22248), .C2(n22043), .A(n22042), .B(n22041), .ZN(
        P1_U3132) );
  AOI22_X1 U23631 ( .A1(n22050), .A2(n22250), .B1(n22049), .B2(n22249), .ZN(
        n22045) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n22252), .B1(
        n22251), .B2(n22046), .ZN(n22044) );
  OAI211_X1 U23633 ( .C1(n22052), .C2(n22255), .A(n22045), .B(n22044), .ZN(
        P1_U3140) );
  AOI22_X1 U23634 ( .A1(n22049), .A2(n22257), .B1(n22050), .B2(n22256), .ZN(
        n22048) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n22260), .B1(
        n22259), .B2(n22046), .ZN(n22047) );
  OAI211_X1 U23636 ( .C1(n22052), .C2(n22274), .A(n22048), .B(n22047), .ZN(
        P1_U3148) );
  AOI22_X1 U23637 ( .A1(n22266), .A2(n22050), .B1(n22049), .B2(n22263), .ZN(
        n22055) );
  INV_X1 U23638 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n22051) );
  OAI22_X1 U23639 ( .A1(n22270), .A2(n22052), .B1(n22268), .B2(n22051), .ZN(
        n22053) );
  INV_X1 U23640 ( .A(n22053), .ZN(n22054) );
  OAI211_X1 U23641 ( .C1(n22056), .C2(n22274), .A(n22055), .B(n22054), .ZN(
        P1_U3156) );
  OAI22_X1 U23642 ( .A1(n22270), .A2(n22098), .B1(n22076), .B2(n22181), .ZN(
        n22057) );
  INV_X1 U23643 ( .A(n22057), .ZN(n22059) );
  AOI22_X1 U23644 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22183), .B1(
        n22189), .B2(n22082), .ZN(n22058) );
  OAI211_X1 U23645 ( .C1(n22186), .C2(n22085), .A(n22059), .B(n22058), .ZN(
        P1_U3037) );
  INV_X1 U23646 ( .A(n22082), .ZN(n22094) );
  INV_X1 U23647 ( .A(n22085), .ZN(n22092) );
  AOI22_X1 U23648 ( .A1(n22188), .A2(n22092), .B1(n22091), .B2(n22187), .ZN(
        n22061) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22190), .B1(
        n22189), .B2(n22088), .ZN(n22060) );
  OAI211_X1 U23650 ( .C1(n22094), .C2(n22193), .A(n22061), .B(n22060), .ZN(
        P1_U3045) );
  OAI22_X1 U23651 ( .A1(n22193), .A2(n22098), .B1(n22076), .B2(n22143), .ZN(
        n22062) );
  INV_X1 U23652 ( .A(n22062), .ZN(n22064) );
  AOI22_X1 U23653 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22196), .B1(
        n22201), .B2(n22082), .ZN(n22063) );
  OAI211_X1 U23654 ( .C1(n22199), .C2(n22085), .A(n22064), .B(n22063), .ZN(
        P1_U3053) );
  AOI22_X1 U23655 ( .A1(n22201), .A2(n22088), .B1(n22091), .B2(n22200), .ZN(
        n22066) );
  AOI22_X1 U23656 ( .A1(n22203), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n22202), .B2(n22082), .ZN(n22065) );
  OAI211_X1 U23657 ( .C1(n22206), .C2(n22085), .A(n22066), .B(n22065), .ZN(
        P1_U3061) );
  OAI22_X1 U23658 ( .A1(n22067), .A2(n22094), .B1(n22076), .B2(n22207), .ZN(
        n22068) );
  INV_X1 U23659 ( .A(n22068), .ZN(n22071) );
  AOI22_X1 U23660 ( .A1(n22211), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n22088), .B2(n22069), .ZN(n22070) );
  OAI211_X1 U23661 ( .C1(n22214), .C2(n22085), .A(n22071), .B(n22070), .ZN(
        P1_U3085) );
  AOI22_X1 U23662 ( .A1(n22216), .A2(n22092), .B1(n22091), .B2(n22215), .ZN(
        n22073) );
  AOI22_X1 U23663 ( .A1(n22218), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n22088), .B2(n22217), .ZN(n22072) );
  OAI211_X1 U23664 ( .C1(n22094), .C2(n22226), .A(n22073), .B(n22072), .ZN(
        P1_U3101) );
  AOI22_X1 U23665 ( .A1(n22222), .A2(n22092), .B1(n22091), .B2(n22221), .ZN(
        n22075) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22223), .B1(
        n22230), .B2(n22082), .ZN(n22074) );
  OAI211_X1 U23667 ( .C1(n22098), .C2(n22226), .A(n22075), .B(n22074), .ZN(
        P1_U3109) );
  OAI22_X1 U23668 ( .A1(n22240), .A2(n22094), .B1(n22076), .B2(n22227), .ZN(
        n22077) );
  INV_X1 U23669 ( .A(n22077), .ZN(n22079) );
  AOI22_X1 U23670 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22231), .B1(
        n22230), .B2(n22088), .ZN(n22078) );
  OAI211_X1 U23671 ( .C1(n22234), .C2(n22085), .A(n22079), .B(n22078), .ZN(
        P1_U3117) );
  AOI22_X1 U23672 ( .A1(n22236), .A2(n22092), .B1(n22091), .B2(n22235), .ZN(
        n22081) );
  AOI22_X1 U23673 ( .A1(n22237), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n22082), .B2(n22243), .ZN(n22080) );
  OAI211_X1 U23674 ( .C1(n22098), .C2(n22240), .A(n22081), .B(n22080), .ZN(
        P1_U3125) );
  AOI22_X1 U23675 ( .A1(n22251), .A2(n22082), .B1(n22091), .B2(n22241), .ZN(
        n22084) );
  AOI22_X1 U23676 ( .A1(n22244), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n22088), .B2(n22243), .ZN(n22083) );
  OAI211_X1 U23677 ( .C1(n22248), .C2(n22085), .A(n22084), .B(n22083), .ZN(
        P1_U3133) );
  AOI22_X1 U23678 ( .A1(n22092), .A2(n22250), .B1(n22091), .B2(n22249), .ZN(
        n22087) );
  AOI22_X1 U23679 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22252), .B1(
        n22251), .B2(n22088), .ZN(n22086) );
  OAI211_X1 U23680 ( .C1(n22094), .C2(n22255), .A(n22087), .B(n22086), .ZN(
        P1_U3141) );
  AOI22_X1 U23681 ( .A1(n22091), .A2(n22257), .B1(n22092), .B2(n22256), .ZN(
        n22090) );
  AOI22_X1 U23682 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22260), .B1(
        n22259), .B2(n22088), .ZN(n22089) );
  OAI211_X1 U23683 ( .C1(n22094), .C2(n22274), .A(n22090), .B(n22089), .ZN(
        P1_U3149) );
  AOI22_X1 U23684 ( .A1(n22266), .A2(n22092), .B1(n22091), .B2(n22263), .ZN(
        n22097) );
  INV_X1 U23685 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n22093) );
  OAI22_X1 U23686 ( .A1(n22270), .A2(n22094), .B1(n22268), .B2(n22093), .ZN(
        n22095) );
  INV_X1 U23687 ( .A(n22095), .ZN(n22096) );
  OAI211_X1 U23688 ( .C1(n22098), .C2(n22274), .A(n22097), .B(n22096), .ZN(
        P1_U3157) );
  OAI22_X1 U23689 ( .A1(n22270), .A2(n22137), .B1(n22115), .B2(n22181), .ZN(
        n22099) );
  INV_X1 U23690 ( .A(n22099), .ZN(n22101) );
  AOI22_X1 U23691 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22183), .B1(
        n22189), .B2(n22121), .ZN(n22100) );
  OAI211_X1 U23692 ( .C1(n22186), .C2(n22124), .A(n22101), .B(n22100), .ZN(
        P1_U3038) );
  INV_X1 U23693 ( .A(n22121), .ZN(n22133) );
  INV_X1 U23694 ( .A(n22124), .ZN(n22131) );
  AOI22_X1 U23695 ( .A1(n22188), .A2(n22131), .B1(n22130), .B2(n22187), .ZN(
        n22103) );
  AOI22_X1 U23696 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22190), .B1(
        n22189), .B2(n22127), .ZN(n22102) );
  OAI211_X1 U23697 ( .C1(n22133), .C2(n22193), .A(n22103), .B(n22102), .ZN(
        P1_U3046) );
  AOI22_X1 U23698 ( .A1(n22201), .A2(n22121), .B1(n22130), .B2(n22194), .ZN(
        n22105) );
  AOI22_X1 U23699 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22196), .B1(
        n22195), .B2(n22127), .ZN(n22104) );
  OAI211_X1 U23700 ( .C1(n22199), .C2(n22124), .A(n22105), .B(n22104), .ZN(
        P1_U3054) );
  AOI22_X1 U23701 ( .A1(n22202), .A2(n22121), .B1(n22130), .B2(n22200), .ZN(
        n22107) );
  AOI22_X1 U23702 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n22203), .B1(
        n22201), .B2(n22127), .ZN(n22106) );
  OAI211_X1 U23703 ( .C1(n22206), .C2(n22124), .A(n22107), .B(n22106), .ZN(
        P1_U3062) );
  OAI22_X1 U23704 ( .A1(n22208), .A2(n22137), .B1(n22115), .B2(n22207), .ZN(
        n22108) );
  INV_X1 U23705 ( .A(n22108), .ZN(n22110) );
  AOI22_X1 U23706 ( .A1(n22211), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n22121), .B2(n22210), .ZN(n22109) );
  OAI211_X1 U23707 ( .C1(n22214), .C2(n22124), .A(n22110), .B(n22109), .ZN(
        P1_U3086) );
  AOI22_X1 U23708 ( .A1(n22216), .A2(n22131), .B1(n22130), .B2(n22215), .ZN(
        n22112) );
  AOI22_X1 U23709 ( .A1(n22218), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n22127), .B2(n22217), .ZN(n22111) );
  OAI211_X1 U23710 ( .C1(n22133), .C2(n22226), .A(n22112), .B(n22111), .ZN(
        P1_U3102) );
  AOI22_X1 U23711 ( .A1(n22222), .A2(n22131), .B1(n22130), .B2(n22221), .ZN(
        n22114) );
  AOI22_X1 U23712 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22223), .B1(
        n22230), .B2(n22121), .ZN(n22113) );
  OAI211_X1 U23713 ( .C1(n22137), .C2(n22226), .A(n22114), .B(n22113), .ZN(
        P1_U3110) );
  OAI22_X1 U23714 ( .A1(n22157), .A2(n22137), .B1(n22115), .B2(n22227), .ZN(
        n22116) );
  INV_X1 U23715 ( .A(n22116), .ZN(n22118) );
  AOI22_X1 U23716 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22231), .B1(
        n22159), .B2(n22121), .ZN(n22117) );
  OAI211_X1 U23717 ( .C1(n22234), .C2(n22124), .A(n22118), .B(n22117), .ZN(
        P1_U3118) );
  AOI22_X1 U23718 ( .A1(n22236), .A2(n22131), .B1(n22130), .B2(n22235), .ZN(
        n22120) );
  AOI22_X1 U23719 ( .A1(n22237), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n22121), .B2(n22243), .ZN(n22119) );
  OAI211_X1 U23720 ( .C1(n22137), .C2(n22240), .A(n22120), .B(n22119), .ZN(
        P1_U3126) );
  AOI22_X1 U23721 ( .A1(n22251), .A2(n22121), .B1(n22130), .B2(n22241), .ZN(
        n22123) );
  AOI22_X1 U23722 ( .A1(n22244), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n22127), .B2(n22243), .ZN(n22122) );
  OAI211_X1 U23723 ( .C1(n22248), .C2(n22124), .A(n22123), .B(n22122), .ZN(
        P1_U3134) );
  AOI22_X1 U23724 ( .A1(n22131), .A2(n22250), .B1(n22130), .B2(n22249), .ZN(
        n22126) );
  AOI22_X1 U23725 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22252), .B1(
        n22251), .B2(n22127), .ZN(n22125) );
  OAI211_X1 U23726 ( .C1(n22133), .C2(n22255), .A(n22126), .B(n22125), .ZN(
        P1_U3142) );
  AOI22_X1 U23727 ( .A1(n22130), .A2(n22257), .B1(n22131), .B2(n22256), .ZN(
        n22129) );
  AOI22_X1 U23728 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22260), .B1(
        n22259), .B2(n22127), .ZN(n22128) );
  OAI211_X1 U23729 ( .C1(n22133), .C2(n22274), .A(n22129), .B(n22128), .ZN(
        P1_U3150) );
  AOI22_X1 U23730 ( .A1(n22266), .A2(n22131), .B1(n22130), .B2(n22263), .ZN(
        n22136) );
  INV_X1 U23731 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n22132) );
  OAI22_X1 U23732 ( .A1(n22270), .A2(n22133), .B1(n22268), .B2(n22132), .ZN(
        n22134) );
  INV_X1 U23733 ( .A(n22134), .ZN(n22135) );
  OAI211_X1 U23734 ( .C1(n22137), .C2(n22274), .A(n22136), .B(n22135), .ZN(
        P1_U3158) );
  OAI22_X1 U23735 ( .A1(n22270), .A2(n22180), .B1(n22156), .B2(n22181), .ZN(
        n22138) );
  INV_X1 U23736 ( .A(n22138), .ZN(n22140) );
  AOI22_X1 U23737 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22183), .B1(
        n22189), .B2(n22164), .ZN(n22139) );
  OAI211_X1 U23738 ( .C1(n22186), .C2(n22167), .A(n22140), .B(n22139), .ZN(
        P1_U3039) );
  INV_X1 U23739 ( .A(n22164), .ZN(n22176) );
  INV_X1 U23740 ( .A(n22167), .ZN(n22174) );
  AOI22_X1 U23741 ( .A1(n22188), .A2(n22174), .B1(n22173), .B2(n22187), .ZN(
        n22142) );
  AOI22_X1 U23742 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n22190), .B1(
        n22189), .B2(n22170), .ZN(n22141) );
  OAI211_X1 U23743 ( .C1(n22176), .C2(n22193), .A(n22142), .B(n22141), .ZN(
        P1_U3047) );
  OAI22_X1 U23744 ( .A1(n22193), .A2(n22180), .B1(n22156), .B2(n22143), .ZN(
        n22144) );
  INV_X1 U23745 ( .A(n22144), .ZN(n22146) );
  AOI22_X1 U23746 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22196), .B1(
        n22201), .B2(n22164), .ZN(n22145) );
  OAI211_X1 U23747 ( .C1(n22199), .C2(n22167), .A(n22146), .B(n22145), .ZN(
        P1_U3055) );
  AOI22_X1 U23748 ( .A1(n22201), .A2(n22170), .B1(n22173), .B2(n22200), .ZN(
        n22148) );
  AOI22_X1 U23749 ( .A1(n22203), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22202), .B2(n22164), .ZN(n22147) );
  OAI211_X1 U23750 ( .C1(n22206), .C2(n22167), .A(n22148), .B(n22147), .ZN(
        P1_U3063) );
  OAI22_X1 U23751 ( .A1(n22208), .A2(n22180), .B1(n22156), .B2(n22207), .ZN(
        n22149) );
  INV_X1 U23752 ( .A(n22149), .ZN(n22151) );
  AOI22_X1 U23753 ( .A1(n22211), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22164), .B2(n22210), .ZN(n22150) );
  OAI211_X1 U23754 ( .C1(n22214), .C2(n22167), .A(n22151), .B(n22150), .ZN(
        P1_U3087) );
  AOI22_X1 U23755 ( .A1(n22216), .A2(n22174), .B1(n22173), .B2(n22215), .ZN(
        n22153) );
  AOI22_X1 U23756 ( .A1(n22218), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n22170), .B2(n22217), .ZN(n22152) );
  OAI211_X1 U23757 ( .C1(n22176), .C2(n22226), .A(n22153), .B(n22152), .ZN(
        P1_U3103) );
  AOI22_X1 U23758 ( .A1(n22222), .A2(n22174), .B1(n22173), .B2(n22221), .ZN(
        n22155) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n22223), .B1(
        n22230), .B2(n22164), .ZN(n22154) );
  OAI211_X1 U23760 ( .C1(n22180), .C2(n22226), .A(n22155), .B(n22154), .ZN(
        P1_U3111) );
  OAI22_X1 U23761 ( .A1(n22157), .A2(n22180), .B1(n22156), .B2(n22227), .ZN(
        n22158) );
  INV_X1 U23762 ( .A(n22158), .ZN(n22161) );
  AOI22_X1 U23763 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22231), .B1(
        n22159), .B2(n22164), .ZN(n22160) );
  OAI211_X1 U23764 ( .C1(n22234), .C2(n22167), .A(n22161), .B(n22160), .ZN(
        P1_U3119) );
  AOI22_X1 U23765 ( .A1(n22236), .A2(n22174), .B1(n22173), .B2(n22235), .ZN(
        n22163) );
  AOI22_X1 U23766 ( .A1(n22237), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n22164), .B2(n22243), .ZN(n22162) );
  OAI211_X1 U23767 ( .C1(n22180), .C2(n22240), .A(n22163), .B(n22162), .ZN(
        P1_U3127) );
  AOI22_X1 U23768 ( .A1(n22251), .A2(n22164), .B1(n22173), .B2(n22241), .ZN(
        n22166) );
  AOI22_X1 U23769 ( .A1(n22244), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n22170), .B2(n22243), .ZN(n22165) );
  OAI211_X1 U23770 ( .C1(n22248), .C2(n22167), .A(n22166), .B(n22165), .ZN(
        P1_U3135) );
  AOI22_X1 U23771 ( .A1(n22174), .A2(n22250), .B1(n22173), .B2(n22249), .ZN(
        n22169) );
  AOI22_X1 U23772 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n22252), .B1(
        n22251), .B2(n22170), .ZN(n22168) );
  OAI211_X1 U23773 ( .C1(n22176), .C2(n22255), .A(n22169), .B(n22168), .ZN(
        P1_U3143) );
  AOI22_X1 U23774 ( .A1(n22173), .A2(n22257), .B1(n22174), .B2(n22256), .ZN(
        n22172) );
  AOI22_X1 U23775 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n22260), .B1(
        n22259), .B2(n22170), .ZN(n22171) );
  OAI211_X1 U23776 ( .C1(n22176), .C2(n22274), .A(n22172), .B(n22171), .ZN(
        P1_U3151) );
  AOI22_X1 U23777 ( .A1(n22266), .A2(n22174), .B1(n22173), .B2(n22263), .ZN(
        n22179) );
  INV_X1 U23778 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n22175) );
  OAI22_X1 U23779 ( .A1(n22270), .A2(n22176), .B1(n22268), .B2(n22175), .ZN(
        n22177) );
  INV_X1 U23780 ( .A(n22177), .ZN(n22178) );
  OAI211_X1 U23781 ( .C1(n22180), .C2(n22274), .A(n22179), .B(n22178), .ZN(
        P1_U3159) );
  OAI22_X1 U23782 ( .A1(n22270), .A2(n22275), .B1(n22228), .B2(n22181), .ZN(
        n22182) );
  INV_X1 U23783 ( .A(n22182), .ZN(n22185) );
  AOI22_X1 U23784 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22183), .B1(
        n22189), .B2(n22242), .ZN(n22184) );
  OAI211_X1 U23785 ( .C1(n22186), .C2(n22247), .A(n22185), .B(n22184), .ZN(
        P1_U3040) );
  INV_X1 U23786 ( .A(n22242), .ZN(n22269) );
  INV_X1 U23787 ( .A(n22247), .ZN(n22265) );
  AOI22_X1 U23788 ( .A1(n22188), .A2(n22265), .B1(n22264), .B2(n22187), .ZN(
        n22192) );
  AOI22_X1 U23789 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22190), .B1(
        n22189), .B2(n22258), .ZN(n22191) );
  OAI211_X1 U23790 ( .C1(n22269), .C2(n22193), .A(n22192), .B(n22191), .ZN(
        P1_U3048) );
  AOI22_X1 U23791 ( .A1(n22201), .A2(n22242), .B1(n22264), .B2(n22194), .ZN(
        n22198) );
  AOI22_X1 U23792 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22196), .B1(
        n22195), .B2(n22258), .ZN(n22197) );
  OAI211_X1 U23793 ( .C1(n22199), .C2(n22247), .A(n22198), .B(n22197), .ZN(
        P1_U3056) );
  AOI22_X1 U23794 ( .A1(n22201), .A2(n22258), .B1(n22264), .B2(n22200), .ZN(
        n22205) );
  AOI22_X1 U23795 ( .A1(n22203), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n22202), .B2(n22242), .ZN(n22204) );
  OAI211_X1 U23796 ( .C1(n22206), .C2(n22247), .A(n22205), .B(n22204), .ZN(
        P1_U3064) );
  OAI22_X1 U23797 ( .A1(n22208), .A2(n22275), .B1(n22228), .B2(n22207), .ZN(
        n22209) );
  INV_X1 U23798 ( .A(n22209), .ZN(n22213) );
  AOI22_X1 U23799 ( .A1(n22211), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n22242), .B2(n22210), .ZN(n22212) );
  OAI211_X1 U23800 ( .C1(n22214), .C2(n22247), .A(n22213), .B(n22212), .ZN(
        P1_U3088) );
  AOI22_X1 U23801 ( .A1(n22216), .A2(n22265), .B1(n22264), .B2(n22215), .ZN(
        n22220) );
  AOI22_X1 U23802 ( .A1(n22218), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n22258), .B2(n22217), .ZN(n22219) );
  OAI211_X1 U23803 ( .C1(n22269), .C2(n22226), .A(n22220), .B(n22219), .ZN(
        P1_U3104) );
  AOI22_X1 U23804 ( .A1(n22222), .A2(n22265), .B1(n22264), .B2(n22221), .ZN(
        n22225) );
  AOI22_X1 U23805 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22223), .B1(
        n22230), .B2(n22242), .ZN(n22224) );
  OAI211_X1 U23806 ( .C1(n22275), .C2(n22226), .A(n22225), .B(n22224), .ZN(
        P1_U3112) );
  OAI22_X1 U23807 ( .A1(n22240), .A2(n22269), .B1(n22228), .B2(n22227), .ZN(
        n22229) );
  INV_X1 U23808 ( .A(n22229), .ZN(n22233) );
  AOI22_X1 U23809 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22231), .B1(
        n22230), .B2(n22258), .ZN(n22232) );
  OAI211_X1 U23810 ( .C1(n22234), .C2(n22247), .A(n22233), .B(n22232), .ZN(
        P1_U3120) );
  AOI22_X1 U23811 ( .A1(n22236), .A2(n22265), .B1(n22264), .B2(n22235), .ZN(
        n22239) );
  AOI22_X1 U23812 ( .A1(n22237), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n22242), .B2(n22243), .ZN(n22238) );
  OAI211_X1 U23813 ( .C1(n22275), .C2(n22240), .A(n22239), .B(n22238), .ZN(
        P1_U3128) );
  AOI22_X1 U23814 ( .A1(n22251), .A2(n22242), .B1(n22264), .B2(n22241), .ZN(
        n22246) );
  AOI22_X1 U23815 ( .A1(n22244), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n22258), .B2(n22243), .ZN(n22245) );
  OAI211_X1 U23816 ( .C1(n22248), .C2(n22247), .A(n22246), .B(n22245), .ZN(
        P1_U3136) );
  AOI22_X1 U23817 ( .A1(n22265), .A2(n22250), .B1(n22264), .B2(n22249), .ZN(
        n22254) );
  AOI22_X1 U23818 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22252), .B1(
        n22251), .B2(n22258), .ZN(n22253) );
  OAI211_X1 U23819 ( .C1(n22269), .C2(n22255), .A(n22254), .B(n22253), .ZN(
        P1_U3144) );
  AOI22_X1 U23820 ( .A1(n22264), .A2(n22257), .B1(n22265), .B2(n22256), .ZN(
        n22262) );
  AOI22_X1 U23821 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22260), .B1(
        n22259), .B2(n22258), .ZN(n22261) );
  OAI211_X1 U23822 ( .C1(n22269), .C2(n22274), .A(n22262), .B(n22261), .ZN(
        P1_U3152) );
  AOI22_X1 U23823 ( .A1(n22266), .A2(n22265), .B1(n22264), .B2(n22263), .ZN(
        n22273) );
  INV_X1 U23824 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n22267) );
  OAI22_X1 U23825 ( .A1(n22270), .A2(n22269), .B1(n22268), .B2(n22267), .ZN(
        n22271) );
  INV_X1 U23826 ( .A(n22271), .ZN(n22272) );
  OAI211_X1 U23827 ( .C1(n22275), .C2(n22274), .A(n22273), .B(n22272), .ZN(
        P1_U3160) );
  INV_X1 U23828 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22278) );
  AOI22_X1 U23829 ( .A1(n22279), .A2(n22278), .B1(n22277), .B2(n22276), .ZN(
        P1_U3486) );
  BUF_X1 U11094 ( .A(n12964), .Z(n13799) );
  BUF_X2 U11332 ( .A(n12474), .Z(n17659) );
  OR2_X1 U22581 ( .A1(n20555), .A2(n11194), .ZN(n20566) );
  BUF_X1 U11163 ( .A(n13305), .Z(n10957) );
  CLKBUF_X1 U11091 ( .A(n11871), .Z(n12320) );
  CLKBUF_X1 U11113 ( .A(n11573), .Z(n14056) );
  NAND2_X1 U11117 ( .A1(n21214), .A2(n20808), .ZN(n12430) );
  NAND2_X1 U11123 ( .A1(n14568), .A2(n12777), .ZN(n11695) );
  CLKBUF_X1 U11137 ( .A(n13748), .Z(n10955) );
  INV_X1 U11157 ( .A(n10954), .ZN(n11663) );
  CLKBUF_X1 U11182 ( .A(n15826), .Z(n20018) );
  CLKBUF_X1 U11187 ( .A(n14320), .Z(n15297) );
  NAND2_X2 U11254 ( .A1(n12978), .A2(n12977), .ZN(n13024) );
  CLKBUF_X1 U11371 ( .A(n13090), .Z(n14978) );
  CLKBUF_X1 U11440 ( .A(n15608), .Z(n10978) );
  OR2_X2 U12094 ( .A1(n11513), .A2(n11512), .ZN(n15576) );
  CLKBUF_X1 U12451 ( .A(n17254), .Z(n17264) );
  CLKBUF_X1 U12740 ( .A(n14994), .Z(n10973) );
  INV_X2 U12888 ( .A(n20097), .ZN(n21253) );
  INV_X2 U12952 ( .A(n14141), .ZN(n18559) );
endmodule

