

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6548, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867;

  OR2_X1 U7277 ( .A1(n14759), .A2(n14761), .ZN(n14760) );
  OAI21_X1 U7278 ( .B1(n14758), .B2(n7789), .A(n7173), .ZN(n6897) );
  AND4_X1 U7279 ( .A1(n8607), .A2(n8606), .A3(n8605), .A4(n8604), .ZN(n10364)
         );
  CLKBUF_X3 U7282 ( .A(n10133), .Z(n10310) );
  CLKBUF_X2 U7284 ( .A(n8784), .Z(n9317) );
  CLKBUF_X2 U7285 ( .A(n8089), .Z(n6534) );
  CLKBUF_X3 U7286 ( .A(n6548), .Z(n9973) );
  NOR2_X2 U7287 ( .A1(n11696), .A2(n10080), .ZN(n13643) );
  NAND2_X1 U7288 ( .A1(n9602), .A2(n6754), .ZN(n12388) );
  XNOR2_X1 U7289 ( .A(n8597), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8598) );
  CLKBUF_X1 U7290 ( .A(n13324), .Z(n6529) );
  NOR2_X1 U7291 ( .A1(n11769), .A2(n15512), .ZN(n13324) );
  OAI21_X1 U7292 ( .B1(n6753), .B2(n6751), .A(n7536), .ZN(n13772) );
  INV_X1 U7293 ( .A(n10115), .ZN(n10309) );
  NAND2_X1 U7294 ( .A1(n6787), .A2(n6786), .ZN(n13179) );
  BUF_X1 U7295 ( .A(n9668), .Z(n9732) );
  OR2_X1 U7296 ( .A1(n9932), .A2(n13587), .ZN(n9946) );
  NAND2_X1 U7297 ( .A1(n11793), .A2(n11792), .ZN(n11890) );
  INV_X1 U7298 ( .A(n10134), .ZN(n10190) );
  INV_X1 U7299 ( .A(n10310), .ZN(n10316) );
  INV_X1 U7300 ( .A(n14967), .ZN(n14961) );
  INV_X1 U7301 ( .A(n11421), .ZN(n12462) );
  CLKBUF_X3 U7302 ( .A(n8089), .Z(n6535) );
  NAND2_X1 U7303 ( .A1(n11153), .A2(n7998), .ZN(n11152) );
  OR2_X1 U7304 ( .A1(n9946), .A2(n13530), .ZN(n9959) );
  AND2_X1 U7306 ( .A1(n10039), .A2(n10038), .ZN(n13953) );
  NAND2_X1 U7307 ( .A1(n8841), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n8878) );
  NAND2_X1 U7308 ( .A1(n9485), .A2(n8800), .ZN(n15275) );
  INV_X1 U7309 ( .A(n13833), .ZN(n10080) );
  INV_X1 U7310 ( .A(n9653), .ZN(n12536) );
  INV_X1 U7311 ( .A(n9973), .ZN(n10089) );
  AND2_X1 U7312 ( .A1(n9648), .A2(n9679), .ZN(n10649) );
  XNOR2_X1 U7313 ( .A(n9285), .B(n9284), .ZN(n15156) );
  NAND2_X1 U7314 ( .A1(n10511), .A2(n10510), .ZN(n10556) );
  AND2_X1 U7315 ( .A1(n8877), .A2(n8876), .ZN(n15251) );
  XNOR2_X1 U7316 ( .A(n10557), .B(n10556), .ZN(n10555) );
  NAND2_X1 U7317 ( .A1(n10685), .A2(n9581), .ZN(n9645) );
  INV_X1 U7318 ( .A(n14568), .ZN(n10150) );
  NAND2_X2 U7319 ( .A1(n11850), .A2(n11849), .ZN(n11848) );
  NAND3_X2 U7320 ( .A1(n7351), .A2(n8148), .A3(n7349), .ZN(n11850) );
  NOR2_X2 U7321 ( .A1(n10686), .A2(n13640), .ZN(n13641) );
  AOI21_X2 U7322 ( .B1(n12368), .B2(n7296), .A(n6618), .ZN(n15194) );
  NAND3_X2 U7323 ( .A1(n6740), .A2(n6739), .A3(n9494), .ZN(n14959) );
  OR2_X1 U7324 ( .A1(n14569), .A2(n15315), .ZN(n9485) );
  BUF_X2 U7325 ( .A(n9184), .Z(n6530) );
  BUF_X1 U7326 ( .A(n9184), .Z(n6531) );
  NAND2_X1 U7327 ( .A1(n9404), .A2(n9403), .ZN(n9184) );
  NOR2_X2 U7328 ( .A1(n14139), .A2(n14262), .ZN(n14112) );
  NAND2_X1 U7329 ( .A1(n13638), .A2(n9912), .ZN(n6532) );
  NAND2_X1 U7330 ( .A1(n13638), .A2(n9912), .ZN(n6533) );
  INV_X2 U7331 ( .A(n13792), .ZN(n13810) );
  XNOR2_X2 U7332 ( .A(n10152), .B(n10270), .ZN(n14462) );
  OR2_X2 U7333 ( .A1(n15506), .A2(n15497), .ZN(n11644) );
  OAI21_X2 U7334 ( .B1(n11301), .B2(n9437), .A(n9436), .ZN(n11584) );
  INV_X1 U7335 ( .A(n11659), .ZN(n7381) );
  XNOR2_X1 U7336 ( .A(n13168), .B(n13339), .ZN(n13159) );
  NAND4_X2 U7337 ( .A1(n8448), .A2(n8447), .A3(n8446), .A4(n8445), .ZN(n13168)
         );
  NAND3_X2 U7339 ( .A1(n8617), .A2(n8616), .A3(n8768), .ZN(n8828) );
  NAND2_X1 U7340 ( .A1(n9655), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U7341 ( .A1(n13484), .A2(n8055), .ZN(n8089) );
  AND2_X2 U7342 ( .A1(n9667), .A2(n9716), .ZN(n10664) );
  BUF_X4 U7344 ( .A(n9645), .Z(n6537) );
  XNOR2_X2 U7345 ( .A(n9701), .B(P2_IR_REG_6__SCAN_IN), .ZN(n15377) );
  NOR2_X2 U7346 ( .A1(n7899), .A2(n7855), .ZN(n7874) );
  NAND2_X2 U7347 ( .A1(n6798), .A2(n7808), .ZN(n14525) );
  BUF_X4 U7348 ( .A(n8622), .Z(n6545) );
  CLKBUF_X3 U7349 ( .A(n9654), .Z(n6548) );
  NAND2_X4 U7350 ( .A1(n10108), .A2(n10107), .ZN(n10115) );
  NAND2_X2 U7351 ( .A1(n9401), .A2(n10533), .ZN(n10108) );
  OAI22_X2 U7352 ( .A1(n11632), .A2(n11631), .B1(n8010), .B2(n6938), .ZN(
        n11828) );
  AOI21_X2 U7353 ( .B1(n11379), .B2(n8009), .A(n11365), .ZN(n11632) );
  XNOR2_X2 U7354 ( .A(n7958), .B(n8046), .ZN(n7986) );
  NAND2_X2 U7355 ( .A1(n12748), .A2(n12747), .ZN(n12745) );
  CLKBUF_X1 U7356 ( .A(n14392), .Z(n7102) );
  OAI21_X1 U7357 ( .B1(n13595), .B2(n13592), .A(n13593), .ZN(n9968) );
  AOI21_X1 U7358 ( .B1(n7596), .B2(n7595), .A(n6643), .ZN(n7594) );
  NAND2_X1 U7359 ( .A1(n7752), .A2(n7753), .ZN(n7200) );
  XNOR2_X1 U7360 ( .A(n8032), .B(n8325), .ZN(n13094) );
  NAND2_X1 U7361 ( .A1(n6994), .A2(n9892), .ZN(n13560) );
  OR2_X1 U7362 ( .A1(n15416), .A2(n15415), .ZN(n15417) );
  OAI22_X1 U7363 ( .A1(n11860), .A2(n11855), .B1(n12205), .B2(n14563), .ZN(
        n11518) );
  OR2_X1 U7364 ( .A1(n10196), .A2(n10195), .ZN(n7848) );
  NAND2_X1 U7365 ( .A1(n9798), .A2(n9797), .ZN(n14297) );
  NAND2_X1 U7366 ( .A1(n9037), .A2(n9036), .ZN(n15055) );
  NAND2_X1 U7367 ( .A1(n6976), .A2(n8671), .ZN(n9167) );
  NAND2_X1 U7368 ( .A1(n9812), .A2(n9811), .ZN(n14292) );
  INV_X2 U7369 ( .A(n14987), .ZN(n6538) );
  NOR2_X1 U7370 ( .A1(n8443), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8457) );
  INV_X1 U7371 ( .A(n13903), .ZN(n13675) );
  OR2_X1 U7372 ( .A1(n9835), .A2(n9834), .ZN(n9851) );
  INV_X2 U7373 ( .A(n12752), .ZN(n12742) );
  INV_X1 U7374 ( .A(n14567), .ZN(n11396) );
  CLKBUF_X1 U7375 ( .A(n10108), .Z(n10409) );
  NAND4_X1 U7376 ( .A1(n8078), .A2(n8077), .A3(n8076), .A4(n8075), .ZN(n15506)
         );
  AND2_X1 U7377 ( .A1(n9639), .A2(n9640), .ZN(n7593) );
  CLKBUF_X3 U7378 ( .A(n9732), .Z(n6540) );
  INV_X2 U7379 ( .A(n9296), .ZN(n8870) );
  CLKBUF_X2 U7380 ( .A(n8775), .Z(n9324) );
  INV_X1 U7381 ( .A(n9878), .ZN(n9663) );
  CLKBUF_X2 U7382 ( .A(n8101), .Z(n12563) );
  OR2_X1 U7383 ( .A1(n9668), .A2(n9277), .ZN(n9629) );
  NAND2_X1 U7384 ( .A1(n9393), .A2(n9392), .ZN(n12106) );
  INV_X2 U7385 ( .A(n6535), .ZN(n6539) );
  INV_X2 U7386 ( .A(n12562), .ZN(n8473) );
  CLKBUF_X1 U7387 ( .A(n8969), .Z(n8655) );
  CLKBUF_X2 U7388 ( .A(n8736), .Z(n9314) );
  OAI21_X1 U7389 ( .B1(n7764), .B2(n9394), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8712) );
  OR2_X1 U7390 ( .A1(n9721), .A2(n15585), .ZN(n9737) );
  NOR2_X1 U7391 ( .A1(n9561), .A2(n9578), .ZN(n9568) );
  AOI21_X1 U7392 ( .B1(n9377), .B2(n9376), .A(n9352), .ZN(n9378) );
  NOR2_X1 U7393 ( .A1(n7322), .A2(n7321), .ZN(n7320) );
  OR2_X1 U7394 ( .A1(n15108), .A2(n9548), .ZN(n6888) );
  AOI21_X1 U7395 ( .B1(n13946), .B2(n12541), .A(n12540), .ZN(n12542) );
  OR2_X1 U7396 ( .A1(n13946), .A2(n6968), .ZN(n6966) );
  NAND2_X1 U7397 ( .A1(n7566), .A2(n6636), .ZN(n13946) );
  AOI21_X1 U7398 ( .B1(n13962), .B2(n14180), .A(n7134), .ZN(n14217) );
  MUX2_X1 U7399 ( .A(n13120), .B(P3_REG0_REG_28__SCAN_IN), .S(n15539), .Z(
        n8544) );
  AOI211_X1 U7400 ( .C1(n14194), .C2(n14206), .A(n13957), .B(n13956), .ZN(
        n13958) );
  AND2_X1 U7401 ( .A1(n14208), .A2(n7112), .ZN(n7111) );
  NOR2_X1 U7402 ( .A1(n13334), .A2(n6563), .ZN(n13398) );
  OR2_X1 U7403 ( .A1(n14210), .A2(n14319), .ZN(n7112) );
  MUX2_X1 U7404 ( .A(n13401), .B(n13400), .S(n15540), .Z(n13402) );
  OR3_X1 U7405 ( .A1(n14245), .A2(n14244), .A3(n14243), .ZN(n14329) );
  XNOR2_X1 U7406 ( .A(n6897), .B(n10367), .ZN(n12396) );
  NOR2_X1 U7407 ( .A1(n13337), .A2(n7078), .ZN(n13400) );
  OR2_X1 U7408 ( .A1(n7609), .A2(n7623), .ZN(n6984) );
  OR2_X1 U7409 ( .A1(n7102), .A2(n14393), .ZN(n7825) );
  NAND2_X1 U7410 ( .A1(n7079), .A2(n13125), .ZN(n8505) );
  AND2_X1 U7411 ( .A1(n14777), .A2(n14776), .ZN(n15015) );
  AND2_X1 U7412 ( .A1(n6844), .A2(n6843), .ZN(n10363) );
  OAI21_X1 U7413 ( .B1(n13981), .B2(n7597), .A(n7594), .ZN(n6834) );
  NAND2_X1 U7414 ( .A1(n14819), .A2(n6632), .ZN(n14803) );
  OAI21_X1 U7415 ( .B1(n7200), .B2(n6842), .A(n6840), .ZN(n6844) );
  NAND2_X1 U7416 ( .A1(n12366), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n12368) );
  NAND2_X1 U7417 ( .A1(n12518), .A2(n12517), .ZN(n14203) );
  NAND2_X1 U7418 ( .A1(n9326), .A2(n9325), .ZN(n12491) );
  NAND2_X1 U7419 ( .A1(n14010), .A2(n12511), .ZN(n13987) );
  NAND2_X1 U7420 ( .A1(n7387), .A2(n8420), .ZN(n13167) );
  NAND2_X1 U7421 ( .A1(n8488), .A2(n8487), .ZN(n8579) );
  AND2_X1 U7422 ( .A1(n14834), .A2(n6682), .ZN(n14746) );
  XNOR2_X1 U7423 ( .A(n9323), .B(n9322), .ZN(n14352) );
  NAND2_X1 U7424 ( .A1(n14026), .A2(n12509), .ZN(n14028) );
  XNOR2_X1 U7425 ( .A(n13333), .B(n13143), .ZN(n13125) );
  OAI21_X1 U7426 ( .B1(n7758), .B2(n9512), .A(n9511), .ZN(n7020) );
  NAND2_X1 U7427 ( .A1(n8472), .A2(n8471), .ZN(n13333) );
  OAI21_X1 U7428 ( .B1(n13560), .B2(n7634), .A(n7632), .ZN(n6997) );
  NAND2_X1 U7429 ( .A1(n9295), .A2(n9294), .ZN(n13800) );
  NAND2_X1 U7430 ( .A1(n6836), .A2(n6835), .ZN(n14026) );
  NAND2_X1 U7431 ( .A1(n14129), .A2(n7254), .ZN(n6836) );
  NOR2_X1 U7432 ( .A1(n8449), .A2(n7386), .ZN(n7385) );
  NAND2_X1 U7433 ( .A1(n14825), .A2(n9503), .ZN(n14812) );
  NAND2_X1 U7434 ( .A1(n10013), .A2(n10012), .ZN(n14220) );
  OR2_X1 U7435 ( .A1(n9293), .A2(n9292), .ZN(n9295) );
  NAND2_X1 U7436 ( .A1(n9248), .A2(n9247), .ZN(n14753) );
  NAND2_X1 U7437 ( .A1(n9227), .A2(n9226), .ZN(n14765) );
  NAND2_X1 U7438 ( .A1(n14131), .A2(n14130), .ZN(n14129) );
  NAND2_X1 U7439 ( .A1(n10008), .A2(n10007), .ZN(n14225) );
  NAND2_X1 U7440 ( .A1(n14411), .A2(n10210), .ZN(n14479) );
  NAND2_X1 U7441 ( .A1(n12319), .A2(n7626), .ZN(n13503) );
  XNOR2_X1 U7442 ( .A(n9263), .B(n9262), .ZN(n12378) );
  XNOR2_X1 U7443 ( .A(n9246), .B(n9245), .ZN(n12351) );
  NAND2_X1 U7444 ( .A1(n6953), .A2(n12522), .ZN(n14159) );
  NOR2_X1 U7445 ( .A1(n7257), .A2(n7602), .ZN(n7254) );
  AND2_X1 U7446 ( .A1(n6569), .A2(n6686), .ZN(n6890) );
  NAND2_X1 U7447 ( .A1(n6991), .A2(n6989), .ZN(n12319) );
  NAND2_X1 U7448 ( .A1(n9213), .A2(n9212), .ZN(n15117) );
  INV_X1 U7449 ( .A(n6735), .ZN(n6734) );
  INV_X1 U7450 ( .A(n7787), .ZN(n7786) );
  AOI21_X1 U7451 ( .B1(n6553), .B2(n8565), .A(n7403), .ZN(n7402) );
  NAND2_X1 U7452 ( .A1(n7347), .A2(n7345), .ZN(n13242) );
  NOR2_X1 U7453 ( .A1(n10222), .A2(n10221), .ZN(n14426) );
  OAI21_X1 U7454 ( .B1(n9464), .B2(n6556), .A(n9466), .ZN(n7787) );
  NAND2_X1 U7455 ( .A1(n9199), .A2(n9198), .ZN(n14800) );
  NAND2_X1 U7456 ( .A1(n6881), .A2(n6879), .ZN(n13268) );
  NAND2_X1 U7457 ( .A1(n8684), .A2(n8683), .ZN(n9211) );
  OAI21_X1 U7458 ( .B1(n7599), .B2(n6559), .A(n6654), .ZN(n7257) );
  OR2_X1 U7459 ( .A1(n7239), .A2(n7592), .ZN(n6839) );
  NAND2_X1 U7460 ( .A1(n6558), .A2(n14948), .ZN(n14931) );
  AND2_X1 U7461 ( .A1(n9368), .A2(n9499), .ZN(n9500) );
  NAND2_X1 U7462 ( .A1(n9173), .A2(n9172), .ZN(n9519) );
  NOR2_X1 U7463 ( .A1(n7848), .A2(n7804), .ZN(n7803) );
  NAND2_X1 U7464 ( .A1(n15164), .A2(n6531), .ZN(n14817) );
  NAND2_X2 U7465 ( .A1(n7065), .A2(n6697), .ZN(n14246) );
  AND2_X1 U7466 ( .A1(n14828), .A2(n9355), .ZN(n14855) );
  AND2_X1 U7467 ( .A1(n9849), .A2(n9848), .ZN(n14280) );
  OAI21_X1 U7468 ( .B1(n9956), .B2(n7284), .A(n8680), .ZN(n9197) );
  XNOR2_X1 U7469 ( .A(n14875), .B(n14557), .ZN(n9368) );
  NAND2_X1 U7470 ( .A1(n12722), .A2(n12723), .ZN(n13218) );
  OR2_X1 U7471 ( .A1(n14858), .A2(n14401), .ZN(n14828) );
  NAND2_X1 U7472 ( .A1(n9915), .A2(n9914), .ZN(n14257) );
  NAND2_X1 U7473 ( .A1(n6875), .A2(n7392), .ZN(n13313) );
  OAI21_X1 U7474 ( .B1(n13697), .B2(n6743), .A(n6744), .ZN(n13702) );
  NAND2_X1 U7475 ( .A1(n9931), .A2(n9930), .ZN(n14252) );
  NAND2_X2 U7476 ( .A1(n8986), .A2(n8985), .ZN(n14875) );
  NAND2_X1 U7477 ( .A1(n11511), .A2(n9286), .ZN(n8986) );
  NAND2_X1 U7478 ( .A1(n9063), .A2(n9062), .ZN(n11059) );
  NAND2_X1 U7479 ( .A1(n9867), .A2(n9866), .ZN(n14274) );
  NAND2_X1 U7480 ( .A1(n7178), .A2(n7177), .ZN(n11175) );
  OAI211_X1 U7481 ( .C1(n8676), .C2(n6597), .A(n6957), .B(n6956), .ZN(n9956)
         );
  INV_X1 U7482 ( .A(n14115), .ZN(n14262) );
  NAND2_X2 U7483 ( .A1(n9024), .A2(n9023), .ZN(n15060) );
  NAND2_X1 U7484 ( .A1(n8998), .A2(n8997), .ZN(n15048) );
  OR2_X1 U7485 ( .A1(n9317), .A2(n14735), .ZN(n8605) );
  XNOR2_X1 U7486 ( .A(n6849), .B(n8983), .ZN(n11511) );
  AOI21_X1 U7487 ( .B1(n7755), .B2(n7025), .A(n6598), .ZN(n7024) );
  AOI21_X1 U7488 ( .B1(n11418), .B2(n13785), .A(n7093), .ZN(n14115) );
  NAND2_X1 U7489 ( .A1(n11005), .A2(n8870), .ZN(n9024) );
  NAND2_X1 U7490 ( .A1(n8978), .A2(n8977), .ZN(n14974) );
  NAND2_X1 U7491 ( .A1(n9167), .A2(n8673), .ZN(n8676) );
  XNOR2_X1 U7492 ( .A(n9018), .B(n9017), .ZN(n11005) );
  OAI21_X1 U7493 ( .B1(n8994), .B2(n8979), .A(n8980), .ZN(n6849) );
  OAI21_X1 U7494 ( .B1(n9046), .B2(n7179), .A(n7175), .ZN(n7174) );
  AND2_X1 U7495 ( .A1(n10948), .A2(n10947), .ZN(n10951) );
  INV_X1 U7496 ( .A(n15096), .ZN(n12301) );
  NAND2_X1 U7497 ( .A1(n8959), .A2(n8958), .ZN(n14507) );
  NAND2_X1 U7498 ( .A1(n9780), .A2(n9779), .ZN(n13711) );
  INV_X1 U7499 ( .A(n9509), .ZN(n14747) );
  OR2_X1 U7500 ( .A1(n9044), .A2(n10860), .ZN(n9046) );
  XNOR2_X1 U7501 ( .A(n8973), .B(n8972), .ZN(n10715) );
  AND2_X1 U7502 ( .A1(n9223), .A2(n9222), .ZN(n9509) );
  OR2_X1 U7503 ( .A1(n10927), .A2(n10926), .ZN(n10948) );
  NAND2_X1 U7504 ( .A1(n9090), .A2(n9089), .ZN(n14984) );
  OAI21_X1 U7505 ( .B1(n9044), .B2(n9014), .A(n9013), .ZN(n9016) );
  INV_X2 U7506 ( .A(n14135), .ZN(n14186) );
  OR2_X1 U7507 ( .A1(n11592), .A2(n11576), .ZN(n11593) );
  XNOR2_X1 U7508 ( .A(n8971), .B(n8970), .ZN(n10697) );
  OAI21_X1 U7509 ( .B1(n8971), .B2(n8970), .A(n8969), .ZN(n8973) );
  OAI21_X2 U7510 ( .B1(n10570), .B2(n9629), .A(n9764), .ZN(n14302) );
  NAND2_X1 U7511 ( .A1(n6797), .A2(n8658), .ZN(n9044) );
  NAND2_X1 U7512 ( .A1(n10924), .A2(n10923), .ZN(n10927) );
  NAND2_X1 U7513 ( .A1(n9085), .A2(n9086), .ZN(n6797) );
  NAND2_X1 U7514 ( .A1(n9751), .A2(n9750), .ZN(n14307) );
  NAND2_X1 U7515 ( .A1(n9734), .A2(n9733), .ZN(n14314) );
  NAND2_X1 U7516 ( .A1(n8933), .A2(n8954), .ZN(n8971) );
  NOR2_X1 U7517 ( .A1(n14458), .A2(n14907), .ZN(n14538) );
  AND2_X1 U7518 ( .A1(n8434), .A2(n8433), .ZN(n13181) );
  INV_X1 U7519 ( .A(n8476), .ZN(n8474) );
  OAI21_X1 U7520 ( .B1(n13649), .B2(n13648), .A(n13647), .ZN(n13652) );
  AND2_X1 U7521 ( .A1(n9147), .A2(n9146), .ZN(n14401) );
  AND2_X1 U7522 ( .A1(n12689), .A2(n12688), .ZN(n13316) );
  NAND2_X1 U7523 ( .A1(n9868), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9883) );
  NAND2_X1 U7524 ( .A1(n8908), .A2(n8907), .ZN(n8906) );
  NOR2_X1 U7525 ( .A1(n10540), .A2(n10742), .ZN(n15244) );
  NAND2_X1 U7526 ( .A1(n15262), .A2(n14567), .ZN(n7831) );
  INV_X1 U7527 ( .A(n13692), .ZN(n6832) );
  XNOR2_X2 U7528 ( .A(n13906), .B(n10867), .ZN(n13650) );
  INV_X1 U7529 ( .A(n9870), .ZN(n9868) );
  AND2_X1 U7530 ( .A1(n8365), .A2(n8364), .ZN(n13233) );
  AND3_X2 U7531 ( .A1(n8778), .A2(n8777), .A3(n8776), .ZN(n15306) );
  NAND2_X1 U7532 ( .A1(n8351), .A2(n8350), .ZN(n13243) );
  AND3_X2 U7533 ( .A1(n8797), .A2(n8796), .A3(n8795), .ZN(n15315) );
  INV_X1 U7534 ( .A(n11788), .ZN(n13900) );
  NAND2_X1 U7535 ( .A1(n9635), .A2(n9636), .ZN(n10867) );
  AND2_X1 U7536 ( .A1(n9742), .A2(n9741), .ZN(n13692) );
  NAND2_X1 U7537 ( .A1(n9651), .A2(n9650), .ZN(n13662) );
  INV_X2 U7538 ( .A(n15294), .ZN(n10117) );
  NAND2_X1 U7539 ( .A1(n11261), .A2(n11260), .ZN(n11421) );
  INV_X2 U7540 ( .A(n15482), .ZN(n7378) );
  OAI211_X1 U7541 ( .C1(n9296), .C2(n12473), .A(n7763), .B(n7762), .ZN(n15294)
         );
  NOR2_X2 U7542 ( .A1(n9001), .A2(n8987), .ZN(n9141) );
  OR2_X1 U7543 ( .A1(n12971), .A2(n12216), .ZN(n12658) );
  AND3_X1 U7544 ( .A1(n8289), .A2(n8288), .A3(n8287), .ZN(n13272) );
  BUF_X1 U7545 ( .A(n10822), .Z(n6543) );
  INV_X1 U7546 ( .A(n14565), .ZN(n11491) );
  AOI21_X1 U7547 ( .B1(n7694), .B2(n7696), .A(n6665), .ZN(n7693) );
  OR2_X1 U7548 ( .A1(n6792), .A2(n6791), .ZN(n11770) );
  INV_X1 U7549 ( .A(n9629), .ZN(n6550) );
  AND2_X2 U7550 ( .A1(n11763), .A2(n12766), .ZN(n12752) );
  INV_X2 U7551 ( .A(n9629), .ZN(n13785) );
  NAND4_X1 U7552 ( .A1(n8139), .A2(n8138), .A3(n8137), .A4(n8136), .ZN(n12972)
         );
  AOI21_X1 U7553 ( .B1(n9913), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n9634), .ZN(
        n9635) );
  NAND4_X2 U7554 ( .A1(n8125), .A2(n8124), .A3(n8123), .A4(n8122), .ZN(n12971)
         );
  NAND4_X2 U7555 ( .A1(n8812), .A2(n8811), .A3(n8810), .A4(n8809), .ZN(n14568)
         );
  NAND4_X1 U7556 ( .A1(n8093), .A2(n8092), .A3(n8091), .A4(n8090), .ZN(n11659)
         );
  OAI21_X1 U7557 ( .B1(n13489), .B2(P3_REG2_REG_0__SCAN_IN), .A(n7996), .ZN(
        n11288) );
  AND2_X1 U7558 ( .A1(n9400), .A2(n9399), .ZN(n10533) );
  NAND4_X1 U7559 ( .A1(n8789), .A2(n8788), .A3(n8787), .A4(n8786), .ZN(n14569)
         );
  AND2_X1 U7560 ( .A1(n8064), .A2(n8063), .ZN(n15513) );
  NOR4_X1 U7561 ( .A1(n8285), .A2(n7026), .A3(P3_REG3_REG_16__SCAN_IN), .A4(
        P3_REG3_REG_18__SCAN_IN), .ZN(n7028) );
  NAND4_X1 U7562 ( .A1(n8106), .A2(n8105), .A3(n8104), .A4(n8103), .ZN(n12973)
         );
  AOI21_X1 U7563 ( .B1(n8891), .B2(n6964), .A(n6963), .ZN(n6962) );
  INV_X1 U7564 ( .A(n6848), .ZN(n9013) );
  INV_X2 U7565 ( .A(n6531), .ZN(n10537) );
  AND2_X1 U7566 ( .A1(n8934), .A2(n7699), .ZN(n7698) );
  OR2_X1 U7567 ( .A1(n8804), .A2(n10125), .ZN(n8737) );
  MUX2_X1 U7568 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9398), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9400) );
  NAND2_X4 U7569 ( .A1(n6530), .A2(n9277), .ZN(n9296) );
  AND2_X1 U7570 ( .A1(n7117), .A2(n8642), .ZN(n8866) );
  AND2_X1 U7571 ( .A1(n7185), .A2(n8954), .ZN(n8934) );
  XNOR2_X1 U7572 ( .A(n9574), .B(n15600), .ZN(n11924) );
  NAND2_X1 U7573 ( .A1(n9571), .A2(n9570), .ZN(n11696) );
  NAND2_X1 U7574 ( .A1(n6814), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8730) );
  NAND2_X2 U7575 ( .A1(n8054), .A2(n8055), .ZN(n8510) );
  INV_X1 U7576 ( .A(n12388), .ZN(n6974) );
  XNOR2_X1 U7577 ( .A(n9396), .B(P1_IR_REG_26__SCAN_IN), .ZN(n10532) );
  XNOR2_X1 U7578 ( .A(n8720), .B(n8719), .ZN(n9520) );
  INV_X2 U7579 ( .A(n8019), .ZN(n6541) );
  AND3_X2 U7580 ( .A1(n9612), .A2(n9611), .A3(n9613), .ZN(n14354) );
  NAND2_X1 U7581 ( .A1(n7099), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9767) );
  INV_X1 U7582 ( .A(n9737), .ZN(n7099) );
  AND2_X1 U7583 ( .A1(n9019), .A2(n8727), .ZN(n9021) );
  AND2_X1 U7584 ( .A1(n8611), .A2(SI_0_), .ZN(n8753) );
  CLKBUF_X1 U7585 ( .A(n9403), .Z(n15163) );
  OR2_X1 U7586 ( .A1(n9681), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9716) );
  OAI21_X1 U7587 ( .B1(n7830), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U7588 ( .A1(n8648), .A2(SI_10_), .ZN(n8954) );
  OAI21_X1 U7589 ( .B1(n9828), .B2(n9578), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9579) );
  INV_X8 U7590 ( .A(n6545), .ZN(n9277) );
  INV_X1 U7591 ( .A(n7946), .ZN(n6945) );
  AND3_X1 U7592 ( .A1(n9568), .A2(n9584), .A3(n9576), .ZN(n10059) );
  AND2_X1 U7593 ( .A1(n8724), .A2(n9380), .ZN(n9384) );
  NAND2_X2 U7594 ( .A1(n6546), .A2(P3_U3151), .ZN(n13487) );
  OR2_X1 U7595 ( .A1(n9794), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9828) );
  NAND2_X2 U7596 ( .A1(n6545), .A2(P2_U3088), .ZN(n14360) );
  INV_X1 U7597 ( .A(n8622), .ZN(n8609) );
  OR2_X1 U7598 ( .A1(n9647), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9679) );
  XNOR2_X1 U7599 ( .A(n7888), .B(P3_IR_REG_2__SCAN_IN), .ZN(n11161) );
  NAND2_X1 U7600 ( .A1(n9590), .A2(n9630), .ZN(n10597) );
  AND4_X1 U7601 ( .A1(n9565), .A2(n9564), .A3(n9563), .A4(n9562), .ZN(n9567)
         );
  AND2_X1 U7602 ( .A1(n9589), .A2(n9566), .ZN(n9632) );
  AND2_X1 U7603 ( .A1(n6999), .A2(n6998), .ZN(n9577) );
  AND3_X1 U7604 ( .A1(n9383), .A2(n9390), .A3(n8585), .ZN(n8710) );
  NOR2_X1 U7605 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n8584) );
  NOR2_X1 U7606 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n8583) );
  NOR2_X2 U7607 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7891) );
  INV_X1 U7608 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7902) );
  INV_X1 U7609 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8719) );
  NOR2_X1 U7610 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7422) );
  INV_X1 U7611 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9383) );
  INV_X1 U7612 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9064) );
  INV_X1 U7613 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7886) );
  NOR2_X1 U7614 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n8588) );
  NOR2_X1 U7615 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8587) );
  INV_X1 U7616 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8729) );
  NOR2_X1 U7617 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n8590) );
  NOR2_X1 U7618 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n8707) );
  NOR2_X1 U7619 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7303) );
  INV_X2 U7620 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7621 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n9565) );
  NOR2_X1 U7622 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n7301) );
  INV_X1 U7623 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10076) );
  NOR2_X1 U7624 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n7300) );
  NOR2_X1 U7625 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n8702) );
  NOR2_X1 U7626 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n9559) );
  NOR2_X2 U7627 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8749) );
  NOR2_X1 U7628 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n9560) );
  NOR2_X1 U7629 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6999) );
  NOR2_X1 U7630 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6998) );
  INV_X4 U7631 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7632 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9829) );
  NOR2_X2 U7633 ( .A1(n14095), .A2(n14252), .ZN(n12543) );
  NAND2_X1 U7634 ( .A1(n8508), .A2(n9277), .ZN(n6542) );
  NAND4_X1 U7635 ( .A1(n9617), .A2(n9616), .A3(n9615), .A4(n9614), .ZN(n10822)
         );
  OAI21_X2 U7636 ( .B1(n14876), .B2(n9317), .A(n8992), .ZN(n14557) );
  NAND2_X2 U7637 ( .A1(n7986), .A2(n8019), .ZN(n8508) );
  NOR2_X2 U7638 ( .A1(n9189), .A2(n14384), .ZN(n9202) );
  OAI21_X2 U7639 ( .B1(n14056), .B2(n6660), .A(n7558), .ZN(n7557) );
  NAND2_X2 U7640 ( .A1(n14079), .A2(n7843), .ZN(n14056) );
  NOR2_X1 U7641 ( .A1(n9668), .A2(n9277), .ZN(n6544) );
  NOR2_X2 U7642 ( .A1(n14929), .A2(n15055), .ZN(n14906) );
  INV_X4 U7643 ( .A(n9878), .ZN(n9913) );
  OAI21_X1 U7644 ( .B1(n8609), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n7272), .ZN(
        n8614) );
  CLKBUF_X1 U7645 ( .A(n10687), .Z(n13846) );
  NOR2_X2 U7646 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n15561) );
  NOR2_X2 U7647 ( .A1(n8878), .A2(n8600), .ZN(n8896) );
  XNOR2_X2 U7648 ( .A(n9579), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9912) );
  AND2_X4 U7649 ( .A1(n6974), .A2(n14354), .ZN(n9653) );
  OAI21_X2 U7650 ( .B1(n14479), .B2(n7796), .A(n7794), .ZN(n14442) );
  AOI211_X2 U7651 ( .C1(n14224), .C2(n14194), .A(n14002), .B(n14001), .ZN(
        n14003) );
  BUF_X4 U7652 ( .A(n8622), .Z(n6546) );
  AND2_X2 U7653 ( .A1(n6847), .A2(n6846), .ZN(n8622) );
  NOR2_X1 U7655 ( .A1(n12388), .A2(n14354), .ZN(n9654) );
  NAND4_X4 U7656 ( .A1(n9623), .A2(n9622), .A3(n9621), .A4(n9620), .ZN(n10686)
         );
  AOI21_X2 U7657 ( .B1(n14125), .B2(n12525), .A(n7106), .ZN(n14105) );
  OAI21_X2 U7658 ( .B1(n11059), .B2(n9296), .A(n9070), .ZN(n14957) );
  AND2_X2 U7659 ( .A1(n9141), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9157) );
  NAND2_X1 U7660 ( .A1(n7007), .A2(n7530), .ZN(n9668) );
  AND2_X1 U7661 ( .A1(n7476), .A2(n7475), .ZN(n7896) );
  INV_X1 U7662 ( .A(n8355), .ZN(n7655) );
  AND2_X1 U7663 ( .A1(n7721), .A2(n7723), .ZN(n7714) );
  INV_X1 U7664 ( .A(n12770), .ZN(n8055) );
  NAND2_X1 U7665 ( .A1(n11036), .A2(n6637), .ZN(n7224) );
  INV_X1 U7666 ( .A(n7385), .ZN(n7384) );
  NAND2_X1 U7667 ( .A1(n7095), .A2(n8428), .ZN(n8479) );
  NAND2_X1 U7668 ( .A1(n7959), .A2(n7451), .ZN(n6793) );
  AND2_X1 U7669 ( .A1(n8053), .A2(n7841), .ZN(n7961) );
  NOR2_X1 U7670 ( .A1(n7960), .A2(n15816), .ZN(n7451) );
  AND2_X1 U7671 ( .A1(n13844), .A2(n7604), .ZN(n7603) );
  NAND2_X1 U7672 ( .A1(n12506), .A2(n12507), .ZN(n7604) );
  NAND2_X1 U7673 ( .A1(n10108), .A2(n10106), .ZN(n10133) );
  AOI21_X1 U7674 ( .B1(n7749), .B2(n11878), .A(n7748), .ZN(n7747) );
  AND2_X1 U7675 ( .A1(n8586), .A2(n8710), .ZN(n8593) );
  AND2_X1 U7676 ( .A1(n7746), .A2(n7745), .ZN(n8586) );
  NOR2_X1 U7677 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7746) );
  NOR2_X1 U7678 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n7745) );
  NOR2_X1 U7679 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n8591) );
  NAND2_X1 U7680 ( .A1(n6942), .A2(n12445), .ZN(n12793) );
  NAND2_X1 U7681 ( .A1(n7144), .A2(n7142), .ZN(n6942) );
  AOI21_X1 U7682 ( .B1(n7145), .B2(n7148), .A(n7143), .ZN(n7142) );
  NAND2_X1 U7684 ( .A1(n8508), .A2(n9277), .ZN(n8177) );
  NOR2_X1 U7685 ( .A1(n10393), .A2(n10392), .ZN(n7372) );
  OAI21_X1 U7686 ( .B1(n10379), .B2(n7681), .A(n7679), .ZN(n12556) );
  INV_X1 U7687 ( .A(n7682), .ZN(n7681) );
  AOI21_X1 U7688 ( .B1(n7680), .B2(n7682), .A(n6731), .ZN(n7679) );
  INV_X1 U7689 ( .A(n7683), .ZN(n7680) );
  OR2_X1 U7690 ( .A1(n14075), .A2(n14057), .ZN(n7843) );
  NAND2_X1 U7691 ( .A1(n8599), .A2(n8598), .ZN(n8784) );
  INV_X1 U7692 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7182) );
  AOI21_X1 U7693 ( .B1(n7332), .B2(n7331), .A(n7329), .ZN(n7328) );
  NAND2_X1 U7694 ( .A1(n12691), .A2(n12690), .ZN(n7314) );
  NAND2_X1 U7695 ( .A1(n13752), .A2(n13754), .ZN(n7531) );
  OAI21_X1 U7696 ( .B1(n13751), .B2(n13750), .A(n6657), .ZN(n6746) );
  AOI21_X1 U7697 ( .B1(n13751), .B2(n13750), .A(n13749), .ZN(n6745) );
  NAND2_X1 U7698 ( .A1(n9155), .A2(n7703), .ZN(n7701) );
  NAND2_X1 U7699 ( .A1(n9175), .A2(n7704), .ZN(n7703) );
  INV_X1 U7700 ( .A(n13764), .ZN(n6752) );
  NAND2_X1 U7701 ( .A1(n13761), .A2(n13763), .ZN(n7535) );
  AND2_X1 U7702 ( .A1(n8653), .A2(n8972), .ZN(n8654) );
  NAND2_X1 U7703 ( .A1(n8655), .A2(n7698), .ZN(n7697) );
  INV_X1 U7704 ( .A(n8647), .ZN(n7699) );
  INV_X1 U7705 ( .A(n11094), .ZN(n7226) );
  INV_X1 U7706 ( .A(n13780), .ZN(n7524) );
  NOR2_X1 U7707 ( .A1(n7560), .A2(n6594), .ZN(n7559) );
  INV_X1 U7708 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U7709 ( .A1(n8705), .A2(n8706), .ZN(n8717) );
  AOI21_X1 U7710 ( .B1(n6848), .B2(n9015), .A(n8664), .ZN(n8665) );
  NAND2_X1 U7711 ( .A1(n10461), .A2(n10460), .ZN(n7055) );
  OAI21_X1 U7712 ( .B1(n12587), .B2(n13108), .A(n12572), .ZN(n12583) );
  NAND2_X1 U7713 ( .A1(n7969), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U7714 ( .A1(n7898), .A2(n7226), .ZN(n7225) );
  NAND2_X1 U7715 ( .A1(n11375), .A2(n7908), .ZN(n7221) );
  INV_X1 U7716 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7880) );
  NAND2_X1 U7717 ( .A1(n6935), .A2(n6934), .ZN(n7920) );
  NAND2_X1 U7718 ( .A1(n7480), .A2(n6587), .ZN(n6935) );
  AOI21_X1 U7719 ( .B1(n12097), .B2(n12096), .A(n6710), .ZN(n6934) );
  AND2_X1 U7720 ( .A1(n7917), .A2(n7481), .ZN(n7480) );
  NAND2_X1 U7721 ( .A1(n7219), .A2(n7214), .ZN(n7937) );
  OAI211_X1 U7722 ( .C1(n7217), .C2(n7213), .A(n7212), .B(n7211), .ZN(n7214)
         );
  NAND2_X1 U7723 ( .A1(n13020), .A2(n6701), .ZN(n7219) );
  NAND2_X1 U7724 ( .A1(n7215), .A2(n8280), .ZN(n7212) );
  NAND2_X1 U7725 ( .A1(n8474), .A2(n8475), .ZN(n8491) );
  NAND2_X1 U7726 ( .A1(n13154), .A2(n8574), .ZN(n12739) );
  INV_X1 U7727 ( .A(n8420), .ZN(n7386) );
  NAND2_X1 U7728 ( .A1(n7029), .A2(n8428), .ZN(n8459) );
  NAND2_X1 U7729 ( .A1(n13411), .A2(n13208), .ZN(n6786) );
  OR2_X1 U7730 ( .A1(n13197), .A2(n8398), .ZN(n6787) );
  NAND2_X1 U7731 ( .A1(n8319), .A2(n8318), .ZN(n7347) );
  OR2_X1 U7732 ( .A1(n12972), .A2(n11770), .ZN(n12647) );
  NAND2_X1 U7733 ( .A1(n11644), .A2(n8545), .ZN(n11643) );
  NOR2_X1 U7734 ( .A1(n8382), .A2(n7376), .ZN(n7375) );
  INV_X1 U7735 ( .A(n8366), .ZN(n7376) );
  OR2_X1 U7736 ( .A1(n13423), .A2(n13233), .ZN(n12722) );
  OR2_X1 U7737 ( .A1(n13469), .A2(n13306), .ZN(n12689) );
  NAND2_X1 U7738 ( .A1(n11528), .A2(n9414), .ZN(n9421) );
  INV_X1 U7739 ( .A(n13493), .ZN(n8520) );
  AND2_X1 U7740 ( .A1(n7864), .A2(n7736), .ZN(n7735) );
  INV_X1 U7741 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7861) );
  NOR2_X1 U7742 ( .A1(n7655), .A2(n7651), .ZN(n7650) );
  INV_X1 U7743 ( .A(n8339), .ZN(n7651) );
  INV_X1 U7744 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7857) );
  NOR2_X1 U7745 ( .A1(n14119), .A2(n7600), .ZN(n7599) );
  INV_X1 U7746 ( .A(n12503), .ZN(n7600) );
  NAND2_X1 U7747 ( .A1(n12500), .A2(n12499), .ZN(n7096) );
  NOR2_X1 U7748 ( .A1(n12040), .A2(n7243), .ZN(n7242) );
  INV_X1 U7749 ( .A(n11888), .ZN(n7243) );
  NAND2_X1 U7750 ( .A1(n11627), .A2(n13900), .ZN(n11784) );
  NAND2_X1 U7751 ( .A1(n11623), .A2(n15438), .ZN(n7556) );
  AND2_X1 U7752 ( .A1(n11900), .A2(n10173), .ZN(n7805) );
  XNOR2_X1 U7753 ( .A(n10116), .B(n10190), .ZN(n10129) );
  INV_X1 U7754 ( .A(n10190), .ZN(n10303) );
  AND3_X1 U7755 ( .A1(n10320), .A2(n11298), .A3(n11296), .ZN(n10331) );
  INV_X1 U7756 ( .A(n8703), .ZN(n8706) );
  NOR2_X1 U7757 ( .A1(n12491), .A2(n14738), .ZN(n7497) );
  AOI21_X1 U7758 ( .B1(n7786), .B2(n6556), .A(n7785), .ZN(n7784) );
  OR2_X1 U7759 ( .A1(n7201), .A2(n7019), .ZN(n6845) );
  AND2_X1 U7760 ( .A1(n9461), .A2(n7776), .ZN(n7775) );
  OR2_X1 U7761 ( .A1(n7778), .A2(n7777), .ZN(n7776) );
  OR2_X1 U7762 ( .A1(n14957), .A2(n14480), .ZN(n9495) );
  NAND2_X1 U7763 ( .A1(n15274), .A2(n8781), .ZN(n9357) );
  NOR2_X1 U7764 ( .A1(n14875), .A2(n15048), .ZN(n7506) );
  OAI21_X1 U7765 ( .B1(n9263), .B2(n8695), .A(n8694), .ZN(n8700) );
  NAND2_X1 U7766 ( .A1(n7262), .A2(n7259), .ZN(n9263) );
  AND2_X1 U7767 ( .A1(n7261), .A2(n7260), .ZN(n7259) );
  NAND2_X1 U7768 ( .A1(n8688), .A2(n7263), .ZN(n7262) );
  NAND2_X1 U7769 ( .A1(n7266), .A2(n7268), .ZN(n7261) );
  NAND2_X1 U7770 ( .A1(n9211), .A2(n8685), .ZN(n8688) );
  INV_X1 U7771 ( .A(n9210), .ZN(n8685) );
  NAND2_X1 U7772 ( .A1(n9384), .A2(n9383), .ZN(n9389) );
  NOR2_X1 U7773 ( .A1(n12940), .A2(n6634), .ZN(n7721) );
  NOR2_X1 U7774 ( .A1(n12451), .A2(n12913), .ZN(n7160) );
  INV_X1 U7775 ( .A(n7727), .ZN(n7726) );
  OAI21_X1 U7776 ( .B1(n12232), .B2(n6557), .A(n12256), .ZN(n7727) );
  OR2_X1 U7777 ( .A1(n8510), .A2(n13106), .ZN(n12567) );
  AND2_X1 U7778 ( .A1(n8381), .A2(n8380), .ZN(n12443) );
  OAI21_X1 U7779 ( .B1(n13489), .B2(P3_REG2_REG_2__SCAN_IN), .A(n7988), .ZN(
        n7989) );
  OR2_X1 U7780 ( .A1(n7968), .A2(n10451), .ZN(n7970) );
  NOR2_X1 U7781 ( .A1(n7898), .A2(n7897), .ZN(n11036) );
  NAND2_X1 U7782 ( .A1(n8015), .A2(n12094), .ZN(n7447) );
  NAND2_X1 U7783 ( .A1(n7235), .A2(n6912), .ZN(n7234) );
  NAND2_X1 U7784 ( .A1(n6932), .A2(n6931), .ZN(n7206) );
  INV_X1 U7785 ( .A(n6717), .ZN(n6931) );
  NAND2_X1 U7786 ( .A1(n13044), .A2(n13377), .ZN(n6932) );
  OAI21_X1 U7787 ( .B1(n7216), .B2(n8023), .A(n6933), .ZN(n13044) );
  AOI21_X1 U7788 ( .B1(n7218), .B2(n8021), .A(n8280), .ZN(n6933) );
  AND2_X1 U7789 ( .A1(n7428), .A2(n13068), .ZN(n7427) );
  OR2_X1 U7790 ( .A1(n13056), .A2(n7429), .ZN(n7428) );
  INV_X1 U7791 ( .A(n8028), .ZN(n7429) );
  INV_X1 U7792 ( .A(n6923), .ZN(n6922) );
  OAI22_X1 U7793 ( .A1(n13079), .A2(n6924), .B1(n7985), .B2(n6925), .ZN(n6923)
         );
  INV_X1 U7794 ( .A(n12739), .ZN(n7420) );
  OR2_X1 U7795 ( .A1(n8574), .A2(n13154), .ZN(n12738) );
  AOI21_X1 U7796 ( .B1(n7400), .B2(n7402), .A(n7399), .ZN(n7398) );
  INV_X1 U7797 ( .A(n12728), .ZN(n7399) );
  AND3_X1 U7798 ( .A1(n8317), .A2(n8316), .A3(n8315), .ZN(n13273) );
  NAND2_X1 U7799 ( .A1(n12627), .A2(n9408), .ZN(n15512) );
  AND4_X1 U7800 ( .A1(n8481), .A2(n8480), .A3(n8479), .A4(n8478), .ZN(n13143)
         );
  NAND2_X1 U7801 ( .A1(n7366), .A2(n6613), .ZN(n7367) );
  NAND2_X1 U7802 ( .A1(n13339), .A2(n8572), .ZN(n8573) );
  NAND2_X1 U7803 ( .A1(n8509), .A2(n12752), .ZN(n15492) );
  INV_X1 U7804 ( .A(n7361), .ZN(n7360) );
  OAI21_X1 U7805 ( .B1(n8275), .B2(n7362), .A(n8274), .ZN(n7361) );
  NAND2_X1 U7806 ( .A1(n8231), .A2(n8230), .ZN(n7362) );
  OR2_X1 U7807 ( .A1(n13301), .A2(n12593), .ZN(n8564) );
  INV_X1 U7808 ( .A(n12569), .ZN(n8342) );
  INV_X1 U7809 ( .A(n7080), .ZN(n8341) );
  AND2_X1 U7810 ( .A1(n11256), .A2(n12752), .ZN(n13320) );
  NOR3_X1 U7811 ( .A1(n7899), .A2(n7855), .A3(P3_IR_REG_27__SCAN_IN), .ZN(
        n6866) );
  NOR2_X1 U7812 ( .A1(n12552), .A2(n7684), .ZN(n7683) );
  INV_X1 U7813 ( .A(n10378), .ZN(n7684) );
  NAND2_X1 U7814 ( .A1(n6945), .A2(n7735), .ZN(n7959) );
  INV_X1 U7815 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n15810) );
  NAND2_X1 U7816 ( .A1(n8401), .A2(n8400), .ZN(n7645) );
  NAND2_X1 U7817 ( .A1(n6945), .A2(n7857), .ZN(n8499) );
  NAND2_X1 U7818 ( .A1(n7011), .A2(n6706), .ZN(n8338) );
  NAND2_X1 U7819 ( .A1(n8307), .A2(n7641), .ZN(n7011) );
  NAND2_X1 U7820 ( .A1(n8247), .A2(n8246), .ZN(n8235) );
  AND2_X1 U7821 ( .A1(n10550), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U7822 ( .A1(n10520), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8129) );
  NAND2_X1 U7823 ( .A1(n8140), .A2(n8141), .ZN(n8144) );
  NAND2_X1 U7824 ( .A1(n7646), .A2(n6631), .ZN(n8127) );
  NAND2_X1 U7825 ( .A1(n7904), .A2(n7905), .ZN(n8004) );
  NAND2_X1 U7826 ( .A1(n9967), .A2(n7610), .ZN(n7609) );
  NOR2_X1 U7827 ( .A1(n7614), .A2(n9996), .ZN(n7610) );
  NAND2_X1 U7828 ( .A1(n10995), .A2(n7081), .ZN(n11109) );
  NOR2_X1 U7829 ( .A1(n11111), .A2(n7625), .ZN(n7081) );
  INV_X1 U7830 ( .A(n9644), .ZN(n7625) );
  NAND2_X1 U7831 ( .A1(n13503), .A2(n6995), .ZN(n6994) );
  AND2_X1 U7832 ( .A1(n10022), .A2(n10021), .ZN(n13782) );
  INV_X1 U7833 ( .A(n14354), .ZN(n6975) );
  INV_X1 U7834 ( .A(n10597), .ZN(n9591) );
  NOR2_X1 U7835 ( .A1(n13953), .A2(n13793), .ZN(n12515) );
  NAND2_X1 U7836 ( .A1(n6834), .A2(n13955), .ZN(n13954) );
  AND2_X1 U7837 ( .A1(n13994), .A2(n6971), .ZN(n6970) );
  OR2_X1 U7838 ( .A1(n14005), .A2(n6972), .ZN(n6971) );
  NAND2_X1 U7839 ( .A1(n14028), .A2(n12510), .ZN(n14010) );
  NAND2_X1 U7840 ( .A1(n7064), .A2(n6647), .ZN(n7253) );
  NAND2_X1 U7841 ( .A1(n7603), .A2(n7601), .ZN(n7064) );
  XNOR2_X1 U7842 ( .A(n14049), .B(n14058), .ZN(n14044) );
  INV_X1 U7843 ( .A(n7571), .ZN(n7570) );
  OAI21_X1 U7844 ( .B1(n7572), .B2(n12528), .A(n14076), .ZN(n7571) );
  NAND2_X1 U7845 ( .A1(n14137), .A2(n13742), .ZN(n14139) );
  NOR2_X1 U7846 ( .A1(n6545), .A2(n7529), .ZN(n7526) );
  INV_X1 U7847 ( .A(n9586), .ZN(n7529) );
  NAND2_X1 U7848 ( .A1(n12520), .A2(n13866), .ZN(n6953) );
  OR2_X1 U7849 ( .A1(n12036), .A2(n13898), .ZN(n7835) );
  INV_X1 U7850 ( .A(n14094), .ZN(n14108) );
  NAND2_X1 U7851 ( .A1(n7008), .A2(n7528), .ZN(n7007) );
  NAND2_X1 U7852 ( .A1(n9586), .A2(n6658), .ZN(n7528) );
  AND2_X1 U7853 ( .A1(n10686), .A2(n11717), .ZN(n10865) );
  AND2_X1 U7854 ( .A1(n11924), .A2(n11696), .ZN(n10826) );
  NAND2_X1 U7855 ( .A1(n7818), .A2(n7817), .ZN(n7812) );
  NAND2_X1 U7856 ( .A1(n14803), .A2(n7770), .ZN(n14781) );
  AND2_X1 U7857 ( .A1(n14773), .A2(n9468), .ZN(n7770) );
  NAND2_X1 U7858 ( .A1(n7200), .A2(n7198), .ZN(n14775) );
  AOI21_X1 U7859 ( .B1(n14967), .B2(n7744), .A(n7743), .ZN(n7742) );
  INV_X1 U7860 ( .A(n14960), .ZN(n7744) );
  INV_X1 U7861 ( .A(n9495), .ZN(n7743) );
  OR2_X1 U7862 ( .A1(n7747), .A2(n7197), .ZN(n6739) );
  AND2_X1 U7863 ( .A1(n9450), .A2(n9448), .ZN(n7781) );
  INV_X1 U7864 ( .A(n14907), .ZN(n14939) );
  INV_X1 U7865 ( .A(n14909), .ZN(n14940) );
  NAND2_X1 U7866 ( .A1(n7077), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8597) );
  AND2_X1 U7867 ( .A1(n8718), .A2(n15718), .ZN(n7189) );
  INV_X1 U7868 ( .A(n9955), .ZN(n7284) );
  NAND2_X1 U7869 ( .A1(n10506), .A2(n10465), .ZN(n10509) );
  NAND2_X1 U7870 ( .A1(n10783), .A2(n10782), .ZN(n10999) );
  NAND2_X1 U7871 ( .A1(n8470), .A2(n7380), .ZN(n7379) );
  INV_X1 U7872 ( .A(n10452), .ZN(n7380) );
  NAND2_X1 U7873 ( .A1(n10034), .A2(n10033), .ZN(n13891) );
  INV_X1 U7874 ( .A(n15420), .ZN(n15398) );
  INV_X1 U7875 ( .A(n9507), .ZN(n14552) );
  NAND2_X1 U7876 ( .A1(n10755), .A2(n10756), .ZN(n14640) );
  NAND2_X1 U7877 ( .A1(n10369), .A2(n10370), .ZN(n12397) );
  INV_X1 U7878 ( .A(n12363), .ZN(n7290) );
  NAND2_X1 U7879 ( .A1(n12364), .A2(n12363), .ZN(n12367) );
  NAND2_X1 U7880 ( .A1(n15181), .A2(n15180), .ZN(n15195) );
  OAI21_X1 U7881 ( .B1(n8822), .B2(n7105), .A(n7104), .ZN(n8779) );
  INV_X1 U7882 ( .A(n9479), .ZN(n7105) );
  NAND2_X1 U7883 ( .A1(n8822), .A2(n9481), .ZN(n7104) );
  OR2_X1 U7884 ( .A1(n8864), .A2(n7340), .ZN(n7339) );
  INV_X1 U7885 ( .A(n8863), .ZN(n7340) );
  NAND2_X1 U7886 ( .A1(n6743), .A2(n6744), .ZN(n6741) );
  INV_X1 U7887 ( .A(n13723), .ZN(n7541) );
  AND2_X1 U7888 ( .A1(n7543), .A2(n13715), .ZN(n7538) );
  OR2_X1 U7889 ( .A1(n15060), .A2(n9330), .ZN(n9110) );
  NAND2_X1 U7890 ( .A1(n14941), .A2(n9151), .ZN(n7131) );
  NAND2_X1 U7891 ( .A1(n15060), .A2(n9091), .ZN(n7132) );
  OAI21_X1 U7892 ( .B1(n8903), .B2(n7332), .A(n6809), .ZN(n8923) );
  AND2_X1 U7893 ( .A1(n7331), .A2(n7329), .ZN(n6809) );
  NOR2_X1 U7894 ( .A1(n8946), .A2(n8943), .ZN(n7342) );
  INV_X1 U7895 ( .A(n8943), .ZN(n7341) );
  INV_X1 U7896 ( .A(n8960), .ZN(n6807) );
  NAND2_X1 U7897 ( .A1(n9008), .A2(n9368), .ZN(n9137) );
  NAND2_X1 U7898 ( .A1(n7092), .A2(n7089), .ZN(n9059) );
  AOI21_X1 U7899 ( .B1(n7306), .B2(n7305), .A(n6862), .ZN(n6861) );
  NAND2_X1 U7900 ( .A1(n13281), .A2(n6863), .ZN(n6862) );
  INV_X1 U7901 ( .A(n12700), .ZN(n6863) );
  NAND2_X1 U7902 ( .A1(n7313), .A2(n7312), .ZN(n7311) );
  NOR2_X1 U7903 ( .A1(n12731), .A2(n7317), .ZN(n7316) );
  NAND2_X1 U7904 ( .A1(n6816), .A2(n7333), .ZN(n9230) );
  NAND2_X1 U7905 ( .A1(n9216), .A2(n9214), .ZN(n7333) );
  OAI21_X1 U7906 ( .B1(n9186), .B2(n6819), .A(n6817), .ZN(n6816) );
  INV_X1 U7907 ( .A(n9032), .ZN(n8667) );
  INV_X1 U7908 ( .A(n12583), .ZN(n12755) );
  NAND2_X1 U7909 ( .A1(n8023), .A2(n13035), .ZN(n7215) );
  NAND2_X1 U7910 ( .A1(n13457), .A2(n12346), .ZN(n12693) );
  NAND2_X1 U7911 ( .A1(n7128), .A2(n6615), .ZN(n7127) );
  INV_X1 U7912 ( .A(n14895), .ZN(n7128) );
  INV_X1 U7913 ( .A(n9249), .ZN(n7691) );
  INV_X1 U7914 ( .A(n9496), .ZN(n7202) );
  NAND2_X1 U7915 ( .A1(n8655), .A2(n8934), .ZN(n7700) );
  OAI21_X1 U7916 ( .B1(n9277), .B2(n10526), .A(n7119), .ZN(n8639) );
  NAND2_X1 U7917 ( .A1(n9277), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7119) );
  NAND2_X1 U7918 ( .A1(n6885), .A2(n6884), .ZN(n8612) );
  NAND2_X1 U7919 ( .A1(n7288), .A2(n7289), .ZN(n10504) );
  NOR2_X1 U7920 ( .A1(n7718), .A2(n7717), .ZN(n7712) );
  INV_X1 U7921 ( .A(n7721), .ZN(n7718) );
  INV_X1 U7922 ( .A(n12918), .ZN(n7147) );
  INV_X1 U7923 ( .A(n12822), .ZN(n7731) );
  NOR2_X1 U7924 ( .A1(n7732), .A2(n7150), .ZN(n7149) );
  INV_X1 U7925 ( .A(n12439), .ZN(n7150) );
  INV_X1 U7926 ( .A(n7733), .ZN(n7732) );
  AND2_X1 U7927 ( .A1(n8521), .A2(n11259), .ZN(n6948) );
  AND2_X1 U7928 ( .A1(n10396), .A2(n12576), .ZN(n12550) );
  INV_X1 U7929 ( .A(n6666), .ZN(n6909) );
  NAND2_X1 U7930 ( .A1(n6909), .A2(n6911), .ZN(n6906) );
  NOR2_X1 U7931 ( .A1(n11101), .A2(n6578), .ZN(n6908) );
  NOR2_X1 U7932 ( .A1(n11379), .A2(n6903), .ZN(n6902) );
  NAND2_X1 U7933 ( .A1(n7489), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7488) );
  NAND2_X1 U7934 ( .A1(n11835), .A2(n7076), .ZN(n7973) );
  OR2_X1 U7935 ( .A1(n11838), .A2(n12071), .ZN(n7076) );
  NAND2_X1 U7936 ( .A1(n12091), .A2(n6703), .ZN(n7975) );
  NOR2_X1 U7937 ( .A1(n12977), .A2(n7449), .ZN(n7448) );
  INV_X1 U7938 ( .A(n12083), .ZN(n7449) );
  INV_X1 U7939 ( .A(n7448), .ZN(n7440) );
  OR2_X1 U7940 ( .A1(n8462), .A2(n13152), .ZN(n13139) );
  NAND2_X1 U7941 ( .A1(n13179), .A2(n13185), .ZN(n7387) );
  INV_X1 U7942 ( .A(n8101), .ZN(n8392) );
  NAND2_X1 U7943 ( .A1(n11929), .A2(n8196), .ZN(n8198) );
  AND2_X1 U7944 ( .A1(n8146), .A2(n11817), .ZN(n7353) );
  NAND2_X1 U7945 ( .A1(n15561), .A2(n8133), .ZN(n8135) );
  NAND2_X1 U7946 ( .A1(n8548), .A2(n12634), .ZN(n11645) );
  NAND2_X1 U7947 ( .A1(n11659), .A2(n15482), .ZN(n12634) );
  OR2_X1 U7948 ( .A1(n10396), .A2(n12576), .ZN(n12751) );
  AND2_X1 U7949 ( .A1(n12738), .A2(n12739), .ZN(n12735) );
  AOI21_X1 U7950 ( .B1(n13281), .B2(n12699), .A(n7408), .ZN(n7407) );
  INV_X1 U7951 ( .A(n12705), .ZN(n7408) );
  NOR2_X1 U7952 ( .A1(n7409), .A2(n7406), .ZN(n7405) );
  INV_X1 U7953 ( .A(n7411), .ZN(n7406) );
  INV_X1 U7954 ( .A(n12693), .ZN(n12593) );
  NAND2_X1 U7955 ( .A1(n12680), .A2(n12674), .ZN(n7394) );
  INV_X1 U7956 ( .A(n12679), .ZN(n7396) );
  NAND2_X1 U7957 ( .A1(n8180), .A2(n6783), .ZN(n6782) );
  INV_X1 U7958 ( .A(n8163), .ZN(n6783) );
  OAI21_X1 U7959 ( .B1(n11762), .B2(n12652), .A(n8556), .ZN(n11846) );
  NAND2_X1 U7960 ( .A1(n8087), .A2(n8086), .ZN(n11647) );
  INV_X1 U7961 ( .A(n12766), .ZN(n9408) );
  OAI21_X1 U7962 ( .B1(n8353), .B2(n7655), .A(n8368), .ZN(n7654) );
  NAND2_X1 U7963 ( .A1(n8338), .A2(n8337), .ZN(n8340) );
  NOR2_X1 U7964 ( .A1(n6867), .A2(n7875), .ZN(n6790) );
  NOR2_X1 U7965 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7302) );
  NOR2_X1 U7966 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n7299) );
  NOR2_X1 U7967 ( .A1(n8237), .A2(n7665), .ZN(n7664) );
  INV_X1 U7968 ( .A(n8234), .ZN(n7665) );
  INV_X1 U7969 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8652) );
  OAI21_X1 U7970 ( .B1(n7671), .B2(n7670), .A(n8183), .ZN(n7669) );
  NOR2_X1 U7971 ( .A1(n8157), .A2(n7675), .ZN(n7674) );
  INV_X1 U7972 ( .A(n8129), .ZN(n7675) );
  INV_X1 U7973 ( .A(n8156), .ZN(n8157) );
  NAND2_X1 U7974 ( .A1(n10515), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8126) );
  INV_X1 U7975 ( .A(n9995), .ZN(n7621) );
  NAND2_X1 U7976 ( .A1(n14235), .A2(n7586), .ZN(n7585) );
  INV_X1 U7977 ( .A(n7587), .ZN(n7586) );
  OR2_X1 U7978 ( .A1(n14049), .A2(n14246), .ZN(n7587) );
  NOR2_X1 U7979 ( .A1(n14089), .A2(n7573), .ZN(n7572) );
  INV_X1 U7980 ( .A(n12526), .ZN(n7573) );
  NAND2_X1 U7981 ( .A1(n7100), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9835) );
  AND2_X1 U7982 ( .A1(n12039), .A2(n6829), .ZN(n6828) );
  OR2_X1 U7983 ( .A1(n13856), .A2(n6831), .ZN(n6829) );
  NAND2_X1 U7984 ( .A1(n12177), .A2(n6630), .ZN(n7592) );
  AND2_X1 U7985 ( .A1(n11738), .A2(n6673), .ZN(n11617) );
  NAND2_X1 U7986 ( .A1(n11051), .A2(n13853), .ZN(n6973) );
  NAND3_X1 U7987 ( .A1(n9605), .A2(n9606), .A3(n9604), .ZN(n7530) );
  NAND2_X1 U7988 ( .A1(n11924), .A2(n13643), .ZN(n13836) );
  INV_X1 U7989 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9564) );
  INV_X1 U7990 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9563) );
  INV_X1 U7991 ( .A(n7824), .ZN(n7822) );
  NAND2_X1 U7992 ( .A1(n10234), .A2(n6801), .ZN(n7796) );
  OR2_X1 U7993 ( .A1(n14426), .A2(n7797), .ZN(n6801) );
  INV_X1 U7994 ( .A(n10217), .ZN(n7797) );
  INV_X1 U7995 ( .A(n14478), .ZN(n7798) );
  INV_X1 U7996 ( .A(n7805), .ZN(n7804) );
  INV_X1 U7997 ( .A(n7848), .ZN(n7801) );
  OR2_X1 U7998 ( .A1(n14462), .A2(n11566), .ZN(n10156) );
  NAND2_X1 U7999 ( .A1(n9305), .A2(n9304), .ZN(n9335) );
  NAND2_X1 U8000 ( .A1(n15107), .A2(n9330), .ZN(n9305) );
  INV_X1 U8001 ( .A(n6671), .ZN(n7276) );
  OR2_X1 U8002 ( .A1(n14717), .A2(n14719), .ZN(n7275) );
  NAND2_X1 U8003 ( .A1(n14717), .A2(n9307), .ZN(n7274) );
  NOR2_X1 U8004 ( .A1(n14773), .A2(n7199), .ZN(n7198) );
  INV_X1 U8005 ( .A(n9506), .ZN(n7199) );
  NOR2_X1 U8006 ( .A1(n14800), .A2(n7511), .ZN(n7510) );
  INV_X1 U8007 ( .A(n14844), .ZN(n7017) );
  NAND2_X1 U8008 ( .A1(n14855), .A2(n14846), .ZN(n7016) );
  INV_X1 U8009 ( .A(n9459), .ZN(n7777) );
  NAND2_X1 U8010 ( .A1(n11387), .A2(n9442), .ZN(n9449) );
  AND2_X1 U8011 ( .A1(n9447), .A2(n9441), .ZN(n9442) );
  NAND2_X1 U8012 ( .A1(n7023), .A2(n6737), .ZN(n11395) );
  NAND2_X1 U8013 ( .A1(n6669), .A2(n7831), .ZN(n7023) );
  NAND2_X1 U8014 ( .A1(n11302), .A2(n6625), .ZN(n6737) );
  NAND2_X1 U8015 ( .A1(n9308), .A2(n11544), .ZN(n10107) );
  NAND2_X1 U8016 ( .A1(n8757), .A2(n10117), .ZN(n9481) );
  AND2_X1 U8017 ( .A1(n14906), .A2(n6683), .ZN(n14856) );
  OR2_X1 U8018 ( .A1(n10863), .A2(n9521), .ZN(n10109) );
  AOI21_X1 U8019 ( .B1(n8699), .B2(n9275), .A(n7281), .ZN(n7280) );
  INV_X1 U8020 ( .A(n9322), .ZN(n7281) );
  INV_X1 U8021 ( .A(n9275), .ZN(n7278) );
  NAND2_X1 U8022 ( .A1(n7283), .A2(n7282), .ZN(n9276) );
  INV_X1 U8023 ( .A(n8699), .ZN(n7282) );
  AND2_X1 U8024 ( .A1(n8687), .A2(n7271), .ZN(n7270) );
  INV_X1 U8025 ( .A(n9224), .ZN(n7271) );
  NAND2_X1 U8026 ( .A1(n9197), .A2(n8682), .ZN(n8684) );
  OR2_X1 U8027 ( .A1(n8678), .A2(n6960), .ZN(n6959) );
  AND2_X1 U8028 ( .A1(n8670), .A2(n8981), .ZN(n8671) );
  NOR2_X1 U8029 ( .A1(n8717), .A2(n7829), .ZN(n7828) );
  NAND2_X1 U8030 ( .A1(n8718), .A2(n8715), .ZN(n7829) );
  NOR2_X1 U8031 ( .A1(n7827), .A2(n8717), .ZN(n7826) );
  AOI21_X1 U8032 ( .B1(n6670), .B2(n8665), .A(n6577), .ZN(n7695) );
  NAND2_X1 U8033 ( .A1(n6795), .A2(SI_8_), .ZN(n8643) );
  NAND2_X1 U8034 ( .A1(n8636), .A2(n8638), .ZN(n8855) );
  NAND2_X1 U8035 ( .A1(n10560), .A2(n10508), .ZN(n10561) );
  OR2_X1 U8036 ( .A1(n10507), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U8037 ( .A1(n11004), .A2(n11003), .ZN(n11319) );
  OR2_X1 U8038 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n11002), .ZN(n11003) );
  OR2_X1 U8039 ( .A1(n15187), .A2(n15186), .ZN(n15189) );
  INV_X1 U8040 ( .A(n13314), .ZN(n12336) );
  NAND2_X1 U8041 ( .A1(n8426), .A2(n8425), .ZN(n8443) );
  OR2_X1 U8042 ( .A1(n12856), .A2(n12431), .ZN(n6941) );
  NAND2_X1 U8043 ( .A1(n6943), .A2(n12227), .ZN(n12892) );
  NAND2_X1 U8044 ( .A1(n12863), .A2(n12221), .ZN(n6943) );
  AOI21_X1 U8045 ( .B1(n7726), .B2(n6570), .A(n7725), .ZN(n7724) );
  INV_X1 U8046 ( .A(n12341), .ZN(n7725) );
  NOR2_X1 U8047 ( .A1(n12762), .A2(n6853), .ZN(n7391) );
  AND4_X1 U8048 ( .A1(n8244), .A2(n8243), .A3(n8242), .A4(n8241), .ZN(n8273)
         );
  NAND2_X1 U8049 ( .A1(n7205), .A2(n7204), .ZN(n7476) );
  NAND2_X1 U8050 ( .A1(n7203), .A2(n7893), .ZN(n7205) );
  INV_X1 U8051 ( .A(n11190), .ZN(n7203) );
  NOR2_X1 U8052 ( .A1(n8003), .A2(n7437), .ZN(n7436) );
  INV_X1 U8053 ( .A(n11043), .ZN(n7437) );
  AOI21_X1 U8054 ( .B1(n7474), .B2(n7970), .A(n11098), .ZN(n11101) );
  INV_X1 U8055 ( .A(n11091), .ZN(n7433) );
  AND2_X1 U8056 ( .A1(n7908), .A2(n7907), .ZN(n11216) );
  OAI21_X1 U8057 ( .B1(n7221), .B2(n6590), .A(n6936), .ZN(n7912) );
  INV_X1 U8058 ( .A(n6937), .ZN(n6936) );
  OAI21_X1 U8059 ( .B1(n7220), .B2(n6590), .A(n6938), .ZN(n6937) );
  NAND2_X1 U8060 ( .A1(n6601), .A2(n10454), .ZN(n7487) );
  OAI21_X1 U8061 ( .B1(n6901), .B2(n6900), .A(n7452), .ZN(n11835) );
  INV_X1 U8062 ( .A(n7454), .ZN(n6900) );
  AOI21_X1 U8063 ( .B1(n7455), .B2(n7454), .A(n7453), .ZN(n7452) );
  NAND2_X1 U8064 ( .A1(n6938), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7454) );
  AND3_X1 U8065 ( .A1(n7487), .A2(n7912), .A3(P3_REG1_REG_7__SCAN_IN), .ZN(
        n11840) );
  AND2_X1 U8066 ( .A1(n7482), .A2(n6587), .ZN(n12098) );
  AND2_X1 U8067 ( .A1(n7917), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7482) );
  INV_X1 U8068 ( .A(n7921), .ZN(n10417) );
  AND2_X1 U8069 ( .A1(n10416), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7233) );
  NAND2_X1 U8070 ( .A1(n10417), .A2(n10416), .ZN(n7232) );
  NAND2_X1 U8071 ( .A1(n6913), .A2(n6912), .ZN(n6914) );
  INV_X1 U8072 ( .A(n7975), .ZN(n6913) );
  NAND2_X1 U8073 ( .A1(n6699), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n12978) );
  OAI21_X1 U8074 ( .B1(n12977), .B2(n7447), .A(n6698), .ZN(n7446) );
  NOR2_X1 U8075 ( .A1(n7446), .A2(n10415), .ZN(n7443) );
  NAND2_X1 U8076 ( .A1(n12084), .A2(n7448), .ZN(n7444) );
  NAND2_X1 U8077 ( .A1(n6918), .A2(n8280), .ZN(n6917) );
  NAND2_X1 U8078 ( .A1(n7980), .A2(n13035), .ZN(n13050) );
  OAI21_X1 U8079 ( .B1(n7478), .B2(n7209), .A(n7208), .ZN(n13098) );
  AOI21_X1 U8080 ( .B1(n7206), .B2(n7939), .A(n8309), .ZN(n7208) );
  NAND2_X1 U8081 ( .A1(n6551), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n13099) );
  NAND2_X1 U8082 ( .A1(n7466), .A2(n13081), .ZN(n13082) );
  INV_X1 U8083 ( .A(n7467), .ZN(n7466) );
  NAND2_X1 U8084 ( .A1(n7985), .A2(n6925), .ZN(n6924) );
  INV_X1 U8085 ( .A(n8491), .ZN(n8490) );
  AND4_X1 U8086 ( .A1(n8461), .A2(n8460), .A3(n8459), .A4(n8458), .ZN(n13154)
         );
  OR2_X2 U8087 ( .A1(n8390), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8412) );
  NAND2_X1 U8088 ( .A1(n7355), .A2(n7357), .ZN(n6789) );
  INV_X1 U8089 ( .A(n7358), .ZN(n7357) );
  OAI21_X1 U8090 ( .B1(n7360), .B2(n13281), .A(n8290), .ZN(n7358) );
  NAND2_X1 U8091 ( .A1(n8560), .A2(n12672), .ZN(n12113) );
  AND3_X1 U8092 ( .A1(n8132), .A2(n8131), .A3(n8130), .ZN(n12216) );
  OR2_X1 U8093 ( .A1(n12569), .A2(n10446), .ZN(n8131) );
  INV_X1 U8094 ( .A(n12627), .ZN(n11763) );
  OR2_X1 U8095 ( .A1(n11537), .A2(n12761), .ZN(n11769) );
  NAND2_X1 U8096 ( .A1(n7414), .A2(n7413), .ZN(n12591) );
  NAND2_X1 U8097 ( .A1(n7031), .A2(n12748), .ZN(n7413) );
  NAND2_X1 U8098 ( .A1(n7416), .A2(n12747), .ZN(n7031) );
  NAND2_X1 U8099 ( .A1(n12751), .A2(n12754), .ZN(n12611) );
  INV_X1 U8100 ( .A(n12726), .ZN(n7403) );
  AND2_X1 U8101 ( .A1(n12728), .A2(n12729), .ZN(n13196) );
  NAND2_X1 U8102 ( .A1(n13258), .A2(n13259), .ZN(n6882) );
  OR2_X1 U8103 ( .A1(n13247), .A2(n13232), .ZN(n13228) );
  NAND2_X1 U8104 ( .A1(n13242), .A2(n8335), .ZN(n13231) );
  NOR2_X1 U8105 ( .A1(n8275), .A2(n7365), .ZN(n7364) );
  INV_X1 U8106 ( .A(n8230), .ZN(n7365) );
  NOR2_X1 U8107 ( .A1(n12698), .A2(n7412), .ZN(n7411) );
  INV_X1 U8108 ( .A(n12694), .ZN(n7412) );
  NAND2_X1 U8109 ( .A1(n13313), .A2(n13316), .ZN(n8563) );
  NAND2_X1 U8110 ( .A1(n8562), .A2(n8561), .ZN(n12115) );
  INV_X1 U8111 ( .A(n12113), .ZN(n8562) );
  AND2_X1 U8112 ( .A1(n12684), .A2(n12685), .ZN(n12679) );
  CLKBUF_X1 U8113 ( .A(n12275), .Z(n12276) );
  AND2_X1 U8114 ( .A1(n12752), .A2(n12760), .ZN(n11179) );
  NOR2_X1 U8115 ( .A1(n9421), .A2(n8538), .ZN(n11249) );
  NOR2_X1 U8116 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  INV_X1 U8117 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7736) );
  AOI21_X1 U8118 ( .B1(n6585), .B2(n7683), .A(n6724), .ZN(n7682) );
  NAND2_X1 U8119 ( .A1(n13478), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U8120 ( .A1(n7009), .A2(n8485), .ZN(n10379) );
  INV_X1 U8121 ( .A(n7864), .ZN(n6944) );
  AND2_X1 U8122 ( .A1(n7738), .A2(n7858), .ZN(n7737) );
  AND2_X1 U8123 ( .A1(n7861), .A2(n7739), .ZN(n7738) );
  NAND2_X1 U8124 ( .A1(n7952), .A2(n7737), .ZN(n7872) );
  NAND2_X1 U8125 ( .A1(n8387), .A2(n8386), .ZN(n8401) );
  AND2_X1 U8126 ( .A1(n7952), .A2(n7858), .ZN(n7954) );
  NOR2_X1 U8127 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7166) );
  INV_X1 U8128 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7858) );
  INV_X1 U8129 ( .A(n8308), .ZN(n7642) );
  NAND2_X1 U8130 ( .A1(n8295), .A2(n8294), .ZN(n8307) );
  INV_X1 U8131 ( .A(n7659), .ZN(n7658) );
  NOR2_X1 U8132 ( .A1(n8278), .A2(n7662), .ZN(n7661) );
  INV_X1 U8133 ( .A(n8236), .ZN(n7662) );
  OAI21_X1 U8134 ( .B1(n8202), .B2(n6667), .A(n7014), .ZN(n8247) );
  NOR2_X1 U8135 ( .A1(n7637), .A2(n6596), .ZN(n7014) );
  XNOR2_X1 U8136 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .ZN(n8246) );
  OR2_X1 U8137 ( .A1(n7878), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U8138 ( .A1(n8204), .A2(n8205), .ZN(n8220) );
  NOR2_X1 U8139 ( .A1(n8174), .A2(n7672), .ZN(n7671) );
  INV_X1 U8140 ( .A(n7676), .ZN(n7672) );
  NAND2_X1 U8141 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n7677), .ZN(n7676) );
  INV_X1 U8142 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7677) );
  XNOR2_X1 U8143 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .ZN(n8156) );
  NAND2_X1 U8144 ( .A1(n8127), .A2(n8126), .ZN(n8140) );
  AND2_X1 U8145 ( .A1(n8129), .A2(n8128), .ZN(n8141) );
  NAND2_X1 U8146 ( .A1(n8097), .A2(n7647), .ZN(n7646) );
  NOR2_X1 U8147 ( .A1(n8108), .A2(n7648), .ZN(n7647) );
  INV_X1 U8148 ( .A(n8096), .ZN(n7648) );
  NOR2_X1 U8149 ( .A1(n13506), .A2(n7627), .ZN(n7626) );
  INV_X1 U8150 ( .A(n9827), .ZN(n7627) );
  NAND2_X1 U8151 ( .A1(n9997), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n10015) );
  INV_X1 U8152 ( .A(n9999), .ZN(n9997) );
  NAND2_X1 U8153 ( .A1(n9793), .A2(n6992), .ZN(n6991) );
  NOR2_X1 U8154 ( .A1(n12159), .A2(n6993), .ZN(n6992) );
  INV_X1 U8155 ( .A(n9792), .ZN(n6993) );
  INV_X1 U8156 ( .A(n9945), .ZN(n7608) );
  NAND2_X1 U8157 ( .A1(n9781), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9800) );
  NOR2_X1 U8158 ( .A1(n11774), .A2(n7631), .ZN(n7630) );
  INV_X1 U8159 ( .A(n9761), .ZN(n7631) );
  NAND2_X1 U8160 ( .A1(n11109), .A2(n9696), .ZN(n6987) );
  NAND2_X1 U8161 ( .A1(n9967), .A2(n7624), .ZN(n7622) );
  NOR2_X1 U8162 ( .A1(n10011), .A2(n10010), .ZN(n7615) );
  NAND2_X1 U8163 ( .A1(n13795), .A2(n13794), .ZN(n7525) );
  AOI22_X1 U8164 ( .A1(n7520), .A2(n7523), .B1(n7517), .B2(n7519), .ZN(n7516)
         );
  INV_X1 U8165 ( .A(n6576), .ZN(n7519) );
  AND2_X1 U8166 ( .A1(n6561), .A2(n6684), .ZN(n7515) );
  OR2_X1 U8167 ( .A1(n13828), .A2(n7837), .ZN(n7836) );
  AND2_X1 U8168 ( .A1(n10094), .A2(n10093), .ZN(n13799) );
  OR2_X1 U8169 ( .A1(n10597), .A2(n11508), .ZN(n7075) );
  OAI22_X1 U8170 ( .A1(n15397), .A2(n15396), .B1(n11472), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n15421) );
  NAND2_X1 U8171 ( .A1(n13981), .A2(n12514), .ZN(n7598) );
  NAND2_X1 U8172 ( .A1(n13973), .A2(n13968), .ZN(n13963) );
  AOI21_X1 U8173 ( .B1(n7563), .B2(n7561), .A(n6641), .ZN(n7560) );
  INV_X1 U8174 ( .A(n12529), .ZN(n7561) );
  NAND2_X1 U8175 ( .A1(n14056), .A2(n12529), .ZN(n7564) );
  AND2_X1 U8176 ( .A1(n7565), .A2(n14044), .ZN(n7563) );
  AND2_X1 U8177 ( .A1(n7564), .A2(n7565), .ZN(n14040) );
  NOR2_X1 U8178 ( .A1(n14071), .A2(n14246), .ZN(n14060) );
  NAND2_X1 U8179 ( .A1(n7101), .A2(n9919), .ZN(n9932) );
  OR2_X1 U8180 ( .A1(n14262), .A2(n14091), .ZN(n12526) );
  AND2_X1 U8181 ( .A1(n7574), .A2(n7572), .ZN(n14087) );
  AND2_X1 U8182 ( .A1(n14268), .A2(n13743), .ZN(n7106) );
  NAND2_X1 U8183 ( .A1(n7097), .A2(n7096), .ZN(n7248) );
  INV_X1 U8184 ( .A(n7577), .ZN(n7005) );
  INV_X1 U8185 ( .A(n14280), .ZN(n14170) );
  INV_X1 U8186 ( .A(n7096), .ZN(n14166) );
  NOR3_X1 U8187 ( .A1(n14183), .A2(n13724), .A3(n14292), .ZN(n14167) );
  OAI21_X1 U8188 ( .B1(n6952), .B2(n13861), .A(n6949), .ZN(n12520) );
  AOI21_X1 U8189 ( .B1(n12174), .B2(n6955), .A(n6614), .ZN(n6952) );
  AND2_X1 U8190 ( .A1(n6955), .A2(n6954), .ZN(n6950) );
  NAND2_X1 U8191 ( .A1(n13716), .A2(n13897), .ZN(n6955) );
  OR2_X1 U8192 ( .A1(n12175), .A2(n12174), .ZN(n6951) );
  NAND2_X1 U8193 ( .A1(n13858), .A2(n7242), .ZN(n7237) );
  INV_X1 U8194 ( .A(n7242), .ZN(n7238) );
  NAND2_X1 U8195 ( .A1(n6827), .A2(n11783), .ZN(n7589) );
  NAND2_X1 U8196 ( .A1(n11782), .A2(n13856), .ZN(n6827) );
  AND2_X1 U8197 ( .A1(n11791), .A2(n11790), .ZN(n11792) );
  INV_X1 U8198 ( .A(n13901), .ZN(n11736) );
  NAND2_X1 U8199 ( .A1(n7553), .A2(n7556), .ZN(n7551) );
  INV_X1 U8200 ( .A(n14106), .ZN(n14092) );
  NAND2_X1 U8201 ( .A1(n10574), .A2(n10580), .ZN(n14094) );
  NAND2_X1 U8202 ( .A1(n13872), .A2(n14180), .ZN(n6968) );
  NAND2_X1 U8203 ( .A1(n9732), .A2(n9591), .ZN(n9592) );
  INV_X1 U8204 ( .A(n9597), .ZN(n10058) );
  INV_X1 U8205 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n14343) );
  INV_X1 U8206 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n15600) );
  INV_X1 U8207 ( .A(n10059), .ZN(n9601) );
  NAND2_X1 U8208 ( .A1(n6545), .A2(SI_0_), .ZN(n9618) );
  NAND2_X1 U8209 ( .A1(n14512), .A2(n10255), .ZN(n14392) );
  NAND2_X1 U8210 ( .A1(n11545), .A2(n7805), .ZN(n11898) );
  OR2_X1 U8211 ( .A1(n10286), .A2(n10285), .ZN(n10287) );
  AOI21_X1 U8212 ( .B1(n14393), .B2(n7824), .A(n14473), .ZN(n7823) );
  NAND2_X1 U8213 ( .A1(n6530), .A2(n6546), .ZN(n8775) );
  INV_X1 U8214 ( .A(n10432), .ZN(n10145) );
  NAND2_X1 U8215 ( .A1(n14420), .A2(n7814), .ZN(n7813) );
  INV_X1 U8216 ( .A(n10287), .ZN(n7814) );
  NOR2_X1 U8217 ( .A1(n6607), .A2(n7807), .ZN(n7806) );
  INV_X1 U8218 ( .A(n14383), .ZN(n7807) );
  NOR2_X1 U8219 ( .A1(n7815), .A2(n7810), .ZN(n7809) );
  OR2_X1 U8220 ( .A1(n14454), .A2(n7817), .ZN(n7810) );
  NAND2_X1 U8221 ( .A1(n9344), .A2(n9341), .ZN(n9347) );
  NAND2_X1 U8222 ( .A1(n6803), .A2(n7129), .ZN(n9271) );
  NAND2_X1 U8223 ( .A1(n9266), .A2(n9268), .ZN(n7129) );
  AND2_X1 U8224 ( .A1(n9209), .A2(n9208), .ZN(n9507) );
  AND4_X1 U8225 ( .A1(n8919), .A2(n8918), .A3(n8917), .A4(n8916), .ZN(n11522)
         );
  INV_X1 U8226 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n15554) );
  AND2_X1 U8227 ( .A1(n14624), .A2(n10729), .ZN(n14643) );
  NAND2_X1 U8228 ( .A1(n11022), .A2(n6766), .ZN(n11135) );
  NOR2_X1 U8229 ( .A1(n11025), .A2(n6767), .ZN(n6766) );
  INV_X1 U8230 ( .A(n11021), .ZN(n6767) );
  INV_X1 U8231 ( .A(n11951), .ZN(n6758) );
  NAND2_X1 U8232 ( .A1(n14682), .A2(n14681), .ZN(n14698) );
  NAND2_X1 U8233 ( .A1(n10372), .A2(n7492), .ZN(n7491) );
  AND2_X1 U8234 ( .A1(n7495), .A2(n7494), .ZN(n7492) );
  NAND2_X1 U8235 ( .A1(n7194), .A2(n9513), .ZN(n7193) );
  INV_X1 U8236 ( .A(n9515), .ZN(n7194) );
  OR2_X1 U8237 ( .A1(n10362), .A2(n7789), .ZN(n7170) );
  OAI21_X1 U8238 ( .B1(n7173), .B2(n10362), .A(n9472), .ZN(n7172) );
  NAND2_X1 U8239 ( .A1(n10363), .A2(n10362), .ZN(n10361) );
  NAND2_X1 U8240 ( .A1(n14758), .A2(n14761), .ZN(n14757) );
  AND2_X1 U8241 ( .A1(n7754), .A2(n14806), .ZN(n7753) );
  NAND2_X1 U8242 ( .A1(n14820), .A2(n9504), .ZN(n7754) );
  NAND2_X1 U8243 ( .A1(n14834), .A2(n7510), .ZN(n14797) );
  NAND2_X1 U8244 ( .A1(n6895), .A2(n6893), .ZN(n14819) );
  AND2_X1 U8245 ( .A1(n7784), .A2(n6894), .ZN(n6893) );
  NAND2_X1 U8246 ( .A1(n7786), .A2(n9368), .ZN(n6894) );
  OR2_X1 U8247 ( .A1(n14812), .A2(n14820), .ZN(n14810) );
  NAND2_X1 U8248 ( .A1(n14850), .A2(n9464), .ZN(n14852) );
  OR2_X1 U8249 ( .A1(n15048), .A2(n14910), .ZN(n14870) );
  NOR2_X1 U8250 ( .A1(n7779), .A2(n9460), .ZN(n7778) );
  INV_X1 U8251 ( .A(n9458), .ZN(n7779) );
  AND3_X1 U8252 ( .A1(n9030), .A2(n9029), .A3(n9028), .ZN(n14884) );
  NAND2_X1 U8253 ( .A1(n7499), .A2(n7498), .ZN(n14929) );
  INV_X1 U8254 ( .A(n14931), .ZN(n7499) );
  NAND2_X1 U8255 ( .A1(n6892), .A2(n7183), .ZN(n14919) );
  OAI21_X1 U8256 ( .B1(n14983), .B2(n6891), .A(n6890), .ZN(n6892) );
  AOI21_X1 U8257 ( .B1(n9457), .B2(n7184), .A(n6664), .ZN(n7183) );
  NAND2_X1 U8258 ( .A1(n14959), .A2(n7742), .ZN(n6738) );
  AOI21_X1 U8259 ( .B1(n7742), .B2(n14961), .A(n9457), .ZN(n7740) );
  AND4_X1 U8260 ( .A1(n9077), .A2(n9076), .A3(n9075), .A4(n9074), .ZN(n14480)
         );
  INV_X1 U8261 ( .A(n9492), .ZN(n7751) );
  AND4_X1 U8262 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(n11861)
         );
  NAND2_X1 U8263 ( .A1(n9449), .A2(n9448), .ZN(n11856) );
  NAND2_X1 U8264 ( .A1(n11856), .A2(n11855), .ZN(n11854) );
  NAND2_X1 U8265 ( .A1(n15275), .A2(n7767), .ZN(n7766) );
  NAND2_X1 U8266 ( .A1(n10537), .A2(n14625), .ZN(n7514) );
  NAND2_X1 U8267 ( .A1(n15287), .A2(n15315), .ZN(n15286) );
  OR2_X1 U8268 ( .A1(n9525), .A2(n15163), .ZN(n14907) );
  INV_X1 U8269 ( .A(n15295), .ZN(n15335) );
  NAND2_X1 U8270 ( .A1(n9531), .A2(n9530), .ZN(n10531) );
  NAND2_X1 U8271 ( .A1(n7022), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7761) );
  INV_X1 U8272 ( .A(n9389), .ZN(n9391) );
  NAND2_X1 U8273 ( .A1(n6600), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6773) );
  AND2_X1 U8274 ( .A1(n8794), .A2(n8814), .ZN(n10486) );
  INV_X1 U8275 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8773) );
  XNOR2_X1 U8276 ( .A(n10561), .B(n14635), .ZN(n10557) );
  NOR2_X1 U8277 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10663), .ZN(n7049) );
  NAND2_X1 U8278 ( .A1(n7036), .A2(n11000), .ZN(n11315) );
  NAND2_X1 U8279 ( .A1(n7716), .A2(n7720), .ZN(n12784) );
  NAND2_X1 U8280 ( .A1(n8411), .A2(n8410), .ZN(n13189) );
  NAND2_X1 U8281 ( .A1(n12461), .A2(n13143), .ZN(n7722) );
  NAND2_X1 U8282 ( .A1(n7156), .A2(n12890), .ZN(n7153) );
  NAND2_X1 U8283 ( .A1(n7159), .A2(n7162), .ZN(n7158) );
  NAND2_X1 U8284 ( .A1(n6555), .A2(n7160), .ZN(n7157) );
  AOI21_X1 U8285 ( .B1(n12910), .B2(n13180), .A(n6659), .ZN(n12883) );
  AND3_X1 U8286 ( .A1(n8117), .A2(n8116), .A3(n8115), .ZN(n11436) );
  INV_X1 U8287 ( .A(n13243), .ZN(n12906) );
  XNOR2_X1 U8288 ( .A(n12793), .B(n12791), .ZN(n12910) );
  AND2_X1 U8289 ( .A1(n11243), .A2(n11536), .ZN(n12958) );
  INV_X1 U8290 ( .A(n12443), .ZN(n13222) );
  INV_X1 U8291 ( .A(n13233), .ZN(n13207) );
  OAI211_X1 U8292 ( .C1(n12563), .C2(n13441), .A(n8303), .B(n8302), .ZN(n13283) );
  INV_X1 U8293 ( .A(n8273), .ZN(n13305) );
  OR2_X1 U8294 ( .A1(n11183), .A2(n11154), .ZN(n7998) );
  NAND2_X1 U8295 ( .A1(n11042), .A2(n8002), .ZN(n7435) );
  NAND2_X1 U8296 ( .A1(n11152), .A2(n7436), .ZN(n7434) );
  INV_X1 U8297 ( .A(n7447), .ZN(n7445) );
  NAND2_X1 U8298 ( .A1(n7234), .A2(n7921), .ZN(n12984) );
  INV_X1 U8299 ( .A(n13090), .ZN(n13077) );
  OAI21_X1 U8300 ( .B1(n13057), .B2(n7429), .A(n7427), .ZN(n13067) );
  AND2_X1 U8301 ( .A1(P3_U3897), .A2(n7986), .ZN(n13095) );
  XNOR2_X1 U8302 ( .A(n7949), .B(n8033), .ZN(n7223) );
  NAND2_X1 U8303 ( .A1(n6929), .A2(n6572), .ZN(n7949) );
  AND2_X1 U8304 ( .A1(n8037), .A2(n13489), .ZN(n13100) );
  NAND2_X1 U8305 ( .A1(n7984), .A2(n6920), .ZN(n6919) );
  AND2_X1 U8306 ( .A1(n6714), .A2(n6922), .ZN(n6920) );
  NAND2_X1 U8307 ( .A1(n6922), .A2(n6924), .ZN(n6921) );
  NAND2_X1 U8308 ( .A1(n6878), .A2(n6876), .ZN(n13334) );
  INV_X1 U8309 ( .A(n6877), .ZN(n6876) );
  NAND2_X1 U8310 ( .A1(n13335), .A2(n15511), .ZN(n6878) );
  OAI21_X1 U8311 ( .B1(n13131), .B2(n15508), .A(n13130), .ZN(n6877) );
  NAND2_X1 U8312 ( .A1(n6779), .A2(n6777), .ZN(n13337) );
  INV_X1 U8313 ( .A(n6778), .ZN(n6777) );
  NAND2_X1 U8314 ( .A1(n6780), .A2(n13308), .ZN(n6779) );
  OAI22_X1 U8315 ( .A1(n8572), .A2(n15492), .B1(n13143), .B2(n15491), .ZN(
        n6778) );
  AND2_X1 U8316 ( .A1(n13187), .A2(n13186), .ZN(n13348) );
  INV_X1 U8317 ( .A(n15500), .ZN(n15519) );
  INV_X1 U8318 ( .A(n15486), .ZN(n15516) );
  NOR2_X1 U8319 ( .A1(n7834), .A2(n9424), .ZN(n9425) );
  NAND2_X1 U8320 ( .A1(n12571), .A2(n12570), .ZN(n13395) );
  NOR2_X1 U8321 ( .A1(n7369), .A2(n13115), .ZN(n7368) );
  INV_X1 U8322 ( .A(n7372), .ZN(n7369) );
  NAND2_X1 U8323 ( .A1(n7415), .A2(n7416), .ZN(n10397) );
  NAND2_X1 U8324 ( .A1(n13138), .A2(n7418), .ZN(n7415) );
  NAND2_X1 U8325 ( .A1(n8373), .A2(n8372), .ZN(n13417) );
  NAND2_X1 U8326 ( .A1(n8357), .A2(n8356), .ZN(n13423) );
  NAND2_X1 U8327 ( .A1(n8344), .A2(n8343), .ZN(n13432) );
  NAND2_X1 U8328 ( .A1(n8311), .A2(n8310), .ZN(n13436) );
  NAND2_X1 U8329 ( .A1(n8282), .A2(n8281), .ZN(n13446) );
  NAND2_X1 U8330 ( .A1(n8239), .A2(n8238), .ZN(n13452) );
  OR2_X1 U8331 ( .A1(n10879), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8524) );
  INV_X1 U8332 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13475) );
  XNOR2_X1 U8333 ( .A(n7895), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10451) );
  INV_X1 U8334 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7853) );
  NAND2_X1 U8335 ( .A1(n6898), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7888) );
  INV_X1 U8336 ( .A(n7891), .ZN(n6898) );
  AND2_X1 U8337 ( .A1(n10048), .A2(n10047), .ZN(n13793) );
  OR2_X1 U8338 ( .A1(n13950), .A2(n10089), .ZN(n10048) );
  NAND2_X1 U8339 ( .A1(n12319), .A2(n9827), .ZN(n13505) );
  NAND2_X1 U8340 ( .A1(n9983), .A2(n9982), .ZN(n14034) );
  NAND2_X1 U8341 ( .A1(n7609), .A2(n6982), .ZN(n6981) );
  NAND2_X1 U8342 ( .A1(n6982), .A2(n7623), .ZN(n6980) );
  AND2_X1 U8343 ( .A1(n9991), .A2(n9990), .ZN(n13597) );
  NAND2_X1 U8344 ( .A1(n6997), .A2(n13519), .ZN(n13585) );
  INV_X1 U8345 ( .A(n7633), .ZN(n7632) );
  OAI21_X1 U8346 ( .B1(n7635), .B2(n7634), .A(n13520), .ZN(n7633) );
  NAND2_X1 U8347 ( .A1(n10082), .A2(n14146), .ZN(n13623) );
  OR2_X1 U8348 ( .A1(n10096), .A2(n10079), .ZN(n13625) );
  INV_X1 U8349 ( .A(n13880), .ZN(n13840) );
  NAND2_X1 U8350 ( .A1(n9980), .A2(n9979), .ZN(n13998) );
  INV_X1 U8351 ( .A(n13597), .ZN(n14041) );
  NAND2_X1 U8352 ( .A1(n9966), .A2(n9965), .ZN(n14058) );
  OAI21_X1 U8353 ( .B1(n14061), .B2(n10089), .A(n9952), .ZN(n14081) );
  NAND2_X1 U8354 ( .A1(n9939), .A2(n9938), .ZN(n14057) );
  NAND2_X1 U8355 ( .A1(n9906), .A2(n9905), .ZN(n13892) );
  NAND2_X1 U8356 ( .A1(n9653), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9620) );
  INV_X1 U8357 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n12424) );
  AOI22_X1 U8358 ( .A1(n12418), .A2(n15394), .B1(n15398), .B2(n12419), .ZN(
        n12422) );
  AOI21_X1 U8359 ( .B1(n12421), .B2(n15394), .A(n14152), .ZN(n7071) );
  INV_X1 U8360 ( .A(n12420), .ZN(n7072) );
  NAND2_X1 U8361 ( .A1(n7258), .A2(n13959), .ZN(n14214) );
  NAND2_X1 U8362 ( .A1(n7598), .A2(n6592), .ZN(n7258) );
  NAND2_X1 U8363 ( .A1(n7598), .A2(n7596), .ZN(n14213) );
  NAND2_X1 U8364 ( .A1(n7136), .A2(n7135), .ZN(n7134) );
  NAND2_X1 U8365 ( .A1(n13999), .A2(n14106), .ZN(n7135) );
  OR2_X1 U8366 ( .A1(n15434), .A2(n10682), .ZN(n14146) );
  NAND2_X1 U8367 ( .A1(n10063), .A2(n10062), .ZN(n15431) );
  AOI21_X1 U8368 ( .B1(n14525), .B2(n14526), .A(n10300), .ZN(n14365) );
  OR2_X1 U8369 ( .A1(n10273), .A2(n10272), .ZN(n10274) );
  NAND2_X1 U8370 ( .A1(n7816), .A2(n10287), .ZN(n7118) );
  NAND2_X1 U8371 ( .A1(n7812), .A2(n7811), .ZN(n7816) );
  INV_X1 U8372 ( .A(n7812), .ZN(n14453) );
  AND4_X1 U8373 ( .A1(n8932), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(n12206)
         );
  AND2_X1 U8374 ( .A1(n10330), .A2(n15280), .ZN(n14524) );
  NAND2_X1 U8375 ( .A1(n10334), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14528) );
  INV_X1 U8376 ( .A(n14524), .ZN(n14544) );
  NOR2_X1 U8377 ( .A1(n7688), .A2(n11926), .ZN(n7338) );
  NAND2_X1 U8378 ( .A1(n6671), .A2(n7689), .ZN(n7688) );
  INV_X1 U8379 ( .A(n9350), .ZN(n7689) );
  INV_X1 U8380 ( .A(n14884), .ZN(n14925) );
  NAND2_X1 U8381 ( .A1(n10759), .A2(n10758), .ZN(n14659) );
  NAND2_X1 U8382 ( .A1(n10769), .A2(n10768), .ZN(n10798) );
  AND2_X1 U8383 ( .A1(n11950), .A2(n6588), .ZN(n11952) );
  OAI21_X1 U8384 ( .B1(n14713), .B2(n14712), .A(n6762), .ZN(n6761) );
  OR2_X1 U8385 ( .A1(n14715), .A2(n14714), .ZN(n6762) );
  OAI211_X1 U8386 ( .C1(n14711), .C2(n14712), .A(n14710), .B(n14709), .ZN(
        n6765) );
  AND2_X1 U8387 ( .A1(n7082), .A2(n14760), .ZN(n14763) );
  NOR2_X1 U8388 ( .A1(n12397), .A2(n6889), .ZN(n15108) );
  NAND2_X1 U8389 ( .A1(n10375), .A2(n10374), .ZN(n6889) );
  INV_X1 U8390 ( .A(n12401), .ZN(n10374) );
  NOR2_X1 U8391 ( .A1(n15008), .A2(n7085), .ZN(n15112) );
  NAND2_X1 U8392 ( .A1(n7087), .A2(n7086), .ZN(n7085) );
  INV_X1 U8393 ( .A(n15009), .ZN(n7086) );
  NAND2_X1 U8394 ( .A1(n15010), .A2(n15339), .ZN(n7087) );
  NAND2_X1 U8395 ( .A1(n10564), .A2(n10563), .ZN(n10783) );
  NAND2_X1 U8396 ( .A1(n7039), .A2(n7038), .ZN(n12149) );
  OR2_X1 U8397 ( .A1(n7045), .A2(n7042), .ZN(n7038) );
  INV_X1 U8398 ( .A(n7040), .ZN(n7039) );
  OAI211_X1 U8399 ( .C1(n11556), .C2(n7041), .A(n7044), .B(n7294), .ZN(n7040)
         );
  NAND2_X1 U8400 ( .A1(n11920), .A2(n11919), .ZN(n12150) );
  NAND2_X1 U8401 ( .A1(n11910), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7295) );
  AND2_X1 U8402 ( .A1(n12367), .A2(n6674), .ZN(n7296) );
  NAND2_X1 U8403 ( .A1(n7297), .A2(n7107), .ZN(n15181) );
  NOR2_X1 U8404 ( .A1(n15179), .A2(n6649), .ZN(n7107) );
  INV_X1 U8405 ( .A(n8846), .ZN(n6826) );
  INV_X1 U8406 ( .A(n8848), .ZN(n6823) );
  NAND2_X1 U8407 ( .A1(n13696), .A2(n13699), .ZN(n6744) );
  NOR2_X1 U8408 ( .A1(n13699), .A2(n13696), .ZN(n6743) );
  NAND2_X1 U8409 ( .A1(n13697), .A2(n6744), .ZN(n6742) );
  OAI21_X1 U8410 ( .B1(n13719), .B2(n13718), .A(n13715), .ZN(n7542) );
  NAND2_X1 U8411 ( .A1(n8902), .A2(n8905), .ZN(n7331) );
  NAND2_X1 U8412 ( .A1(n8890), .A2(n8889), .ZN(n6810) );
  NAND2_X1 U8413 ( .A1(n8886), .A2(n8885), .ZN(n6811) );
  NOR2_X1 U8414 ( .A1(n8905), .A2(n8902), .ZN(n7332) );
  NAND2_X1 U8415 ( .A1(n9039), .A2(n9110), .ZN(n7091) );
  NAND2_X1 U8416 ( .A1(n7313), .A2(n12692), .ZN(n7307) );
  INV_X1 U8417 ( .A(n7314), .ZN(n7313) );
  INV_X1 U8418 ( .A(n9137), .ZN(n7686) );
  INV_X1 U8419 ( .A(n9097), .ZN(n7685) );
  NAND2_X1 U8420 ( .A1(n6806), .A2(n8960), .ZN(n6805) );
  OAI22_X1 U8421 ( .A1(n8944), .A2(n7342), .B1(n7341), .B2(n8945), .ZN(n8961)
         );
  AOI21_X1 U8422 ( .B1(n6604), .B2(n9123), .A(n9122), .ZN(n9136) );
  AOI21_X1 U8423 ( .B1(n6860), .B2(n12704), .A(n12703), .ZN(n12709) );
  NAND2_X1 U8424 ( .A1(n7309), .A2(n6861), .ZN(n6860) );
  NAND2_X1 U8425 ( .A1(n13745), .A2(n13748), .ZN(n7532) );
  NOR2_X1 U8426 ( .A1(n13748), .A2(n13745), .ZN(n7533) );
  NAND2_X1 U8427 ( .A1(n13178), .A2(n12730), .ZN(n7317) );
  INV_X1 U8428 ( .A(n13171), .ZN(n12731) );
  NAND2_X1 U8429 ( .A1(n7706), .A2(n9201), .ZN(n7705) );
  NOR2_X1 U8430 ( .A1(n7334), .A2(n6818), .ZN(n6817) );
  NOR2_X1 U8431 ( .A1(n9201), .A2(n7706), .ZN(n6818) );
  AND2_X1 U8432 ( .A1(n9215), .A2(n7335), .ZN(n7334) );
  INV_X1 U8433 ( .A(n9214), .ZN(n7335) );
  AOI21_X1 U8434 ( .B1(n12741), .B2(n12740), .A(n13125), .ZN(n6858) );
  INV_X1 U8435 ( .A(n7265), .ZN(n7264) );
  OAI21_X1 U8436 ( .B1(n7270), .B2(n6584), .A(n9244), .ZN(n7265) );
  AND2_X1 U8437 ( .A1(n7695), .A2(n6677), .ZN(n7694) );
  AND2_X1 U8438 ( .A1(n12096), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7481) );
  AND2_X1 U8439 ( .A1(n12992), .A2(n7215), .ZN(n7210) );
  INV_X1 U8440 ( .A(n7215), .ZN(n7213) );
  NAND2_X1 U8441 ( .A1(n13139), .A2(n8463), .ZN(n7383) );
  NOR2_X1 U8442 ( .A1(n8211), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7033) );
  NAND2_X1 U8443 ( .A1(n12651), .A2(n8553), .ZN(n12652) );
  INV_X1 U8444 ( .A(n13473), .ZN(n11528) );
  NAND2_X1 U8445 ( .A1(n13767), .A2(n13769), .ZN(n7536) );
  INV_X1 U8446 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9562) );
  NAND2_X1 U8447 ( .A1(n14957), .A2(n10309), .ZN(n6802) );
  INV_X1 U8448 ( .A(n7267), .ZN(n7266) );
  OAI21_X1 U8449 ( .B1(n7270), .B2(n7268), .A(n13492), .ZN(n7267) );
  INV_X1 U8450 ( .A(n8692), .ZN(n7268) );
  OR2_X1 U8451 ( .A1(n7264), .A2(n7266), .ZN(n7263) );
  NAND2_X1 U8452 ( .A1(n7264), .A2(n6584), .ZN(n7260) );
  INV_X1 U8453 ( .A(n8672), .ZN(n6977) );
  NAND2_X1 U8454 ( .A1(n6797), .A2(n7694), .ZN(n7692) );
  XNOR2_X1 U8455 ( .A(n12462), .B(n7141), .ZN(n12224) );
  OAI21_X1 U8456 ( .B1(n12774), .B2(n12831), .A(n12223), .ZN(n12225) );
  INV_X1 U8457 ( .A(n12841), .ZN(n7143) );
  INV_X1 U8458 ( .A(n12758), .ZN(n12759) );
  OAI21_X1 U8459 ( .B1(n8019), .B2(P3_REG2_REG_1__SCAN_IN), .A(n7993), .ZN(
        n7995) );
  NAND2_X1 U8460 ( .A1(n8019), .A2(n15541), .ZN(n7993) );
  NAND2_X1 U8461 ( .A1(n7995), .A2(n7994), .ZN(n7997) );
  NOR2_X1 U8462 ( .A1(n6595), .A2(n11144), .ZN(n7968) );
  NAND2_X1 U8463 ( .A1(n7990), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7475) );
  NAND2_X1 U8464 ( .A1(n7473), .A2(n7970), .ZN(n11099) );
  INV_X1 U8465 ( .A(n7474), .ZN(n7473) );
  NAND2_X1 U8466 ( .A1(n8006), .A2(n11106), .ZN(n7438) );
  INV_X1 U8467 ( .A(n11374), .ZN(n7220) );
  INV_X1 U8468 ( .A(n11831), .ZN(n7453) );
  NOR2_X1 U8469 ( .A1(n6938), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7455) );
  NOR2_X1 U8470 ( .A1(n7233), .A2(n6583), .ZN(n7228) );
  INV_X1 U8471 ( .A(n7218), .ZN(n7217) );
  OAI21_X1 U8472 ( .B1(n13021), .B2(P3_REG1_REG_13__SCAN_IN), .A(n13022), .ZN(
        n7218) );
  NAND2_X1 U8473 ( .A1(n7925), .A2(n12992), .ZN(n7216) );
  INV_X1 U8474 ( .A(n8034), .ZN(n6925) );
  NAND2_X1 U8475 ( .A1(n10381), .A2(n10380), .ZN(n10396) );
  OR2_X1 U8476 ( .A1(n13189), .A2(n12913), .ZN(n12617) );
  NOR2_X1 U8477 ( .A1(n8412), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8426) );
  NOR2_X1 U8478 ( .A1(n6553), .A2(n12608), .ZN(n7400) );
  NAND2_X1 U8479 ( .A1(n8312), .A2(n7027), .ZN(n7026) );
  INV_X1 U8480 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7027) );
  AND2_X1 U8481 ( .A1(n7409), .A2(n7364), .ZN(n7356) );
  NAND2_X1 U8482 ( .A1(n7033), .A2(n7032), .ZN(n8250) );
  INV_X1 U8483 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n7032) );
  INV_X1 U8484 ( .A(n7033), .ZN(n8224) );
  NAND2_X1 U8485 ( .A1(n8190), .A2(n12026), .ZN(n8211) );
  INV_X1 U8486 ( .A(n13127), .ZN(n7079) );
  NAND2_X1 U8487 ( .A1(n7422), .A2(n7891), .ZN(n7899) );
  INV_X1 U8488 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7854) );
  OAI21_X1 U8489 ( .B1(n8401), .B2(n7644), .A(n7012), .ZN(n8437) );
  AOI21_X1 U8490 ( .B1(n7643), .B2(n8399), .A(n7013), .ZN(n7012) );
  INV_X1 U8491 ( .A(n8421), .ZN(n7013) );
  NAND2_X1 U8492 ( .A1(n7954), .A2(n7861), .ZN(n7870) );
  AOI21_X1 U8493 ( .B1(n8305), .B2(n8308), .A(n8321), .ZN(n7641) );
  NAND2_X1 U8494 ( .A1(n7641), .A2(n7642), .ZN(n7639) );
  OR2_X1 U8495 ( .A1(n7940), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n7942) );
  OAI21_X1 U8496 ( .B1(n7661), .B2(n7660), .A(n8292), .ZN(n7659) );
  NOR2_X1 U8497 ( .A1(n7638), .A2(n8219), .ZN(n7637) );
  INV_X1 U8498 ( .A(n8232), .ZN(n7638) );
  INV_X1 U8499 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7856) );
  CLKBUF_X1 U8500 ( .A(n7899), .Z(n7900) );
  NOR2_X1 U8501 ( .A1(n9893), .A2(n6996), .ZN(n6995) );
  INV_X1 U8502 ( .A(n9845), .ZN(n6996) );
  INV_X1 U8503 ( .A(n6537), .ZN(n10014) );
  NAND2_X1 U8504 ( .A1(n7518), .A2(n6576), .ZN(n7523) );
  NOR2_X1 U8505 ( .A1(n7522), .A2(n7518), .ZN(n7517) );
  AOI21_X1 U8506 ( .B1(n7518), .B2(n7522), .A(n7521), .ZN(n7520) );
  INV_X1 U8507 ( .A(n13783), .ZN(n7521) );
  AOI22_X1 U8508 ( .A1(n12406), .A2(n12405), .B1(P2_REG1_REG_17__SCAN_IN), 
        .B2(n12410), .ZN(n12407) );
  NOR2_X1 U8509 ( .A1(n7559), .A2(n12530), .ZN(n7558) );
  INV_X1 U8510 ( .A(n12507), .ZN(n7601) );
  NOR2_X1 U8511 ( .A1(n12528), .A2(n7569), .ZN(n7568) );
  INV_X1 U8512 ( .A(n7850), .ZN(n7569) );
  NAND2_X1 U8513 ( .A1(n9605), .A2(n9604), .ZN(n10083) );
  NAND2_X1 U8514 ( .A1(n14280), .A2(n7578), .ZN(n7577) );
  INV_X1 U8515 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9834) );
  INV_X1 U8516 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9799) );
  INV_X1 U8517 ( .A(n7100), .ZN(n9814) );
  NAND2_X1 U8518 ( .A1(n6833), .A2(n6832), .ZN(n11785) );
  AND2_X1 U8519 ( .A1(n10869), .A2(n13659), .ZN(n7576) );
  NOR2_X1 U8520 ( .A1(n14280), .A2(n13894), .ZN(n12523) );
  NAND2_X1 U8521 ( .A1(n7001), .A2(n13674), .ZN(n11706) );
  INV_X1 U8522 ( .A(n11056), .ZN(n7001) );
  INV_X1 U8523 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9558) );
  OR2_X1 U8524 ( .A1(n9846), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n9859) );
  OR2_X1 U8525 ( .A1(n9762), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n9777) );
  INV_X1 U8526 ( .A(n10133), .ZN(n10307) );
  NAND2_X1 U8527 ( .A1(n9334), .A2(n7066), .ZN(n9338) );
  INV_X1 U8528 ( .A(n9333), .ZN(n7066) );
  AND2_X1 U8529 ( .A1(n9367), .A2(n7126), .ZN(n9369) );
  NOR2_X1 U8530 ( .A1(n14918), .A2(n7127), .ZN(n7126) );
  NAND2_X1 U8531 ( .A1(n9250), .A2(n7691), .ZN(n7690) );
  NOR2_X1 U8532 ( .A1(n6552), .A2(n6575), .ZN(n7130) );
  NAND2_X1 U8533 ( .A1(n7068), .A2(n7067), .ZN(n9333) );
  NAND2_X1 U8534 ( .A1(n14549), .A2(n9307), .ZN(n7067) );
  NAND2_X1 U8535 ( .A1(n12491), .A2(n9091), .ZN(n7068) );
  NAND2_X1 U8536 ( .A1(n14761), .A2(n9510), .ZN(n7758) );
  INV_X1 U8537 ( .A(n6841), .ZN(n6840) );
  OAI21_X1 U8538 ( .B1(n7198), .B2(n6842), .A(n7759), .ZN(n6841) );
  NOR2_X1 U8539 ( .A1(n9512), .A2(n7760), .ZN(n7759) );
  INV_X1 U8540 ( .A(n9510), .ZN(n7760) );
  INV_X1 U8541 ( .A(n9508), .ZN(n6842) );
  NOR2_X1 U8542 ( .A1(n15117), .A2(n7509), .ZN(n7508) );
  INV_X1 U8543 ( .A(n7510), .ZN(n7509) );
  NAND2_X1 U8544 ( .A1(n9157), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9176) );
  INV_X1 U8545 ( .A(n9454), .ZN(n6891) );
  NOR2_X1 U8546 ( .A1(n14975), .A2(n7502), .ZN(n7501) );
  OR2_X1 U8547 ( .A1(n14974), .A2(n14984), .ZN(n7502) );
  OR2_X1 U8548 ( .A1(n8927), .A2(n8601), .ZN(n8948) );
  AND2_X1 U8549 ( .A1(n11457), .A2(n15251), .ZN(n7505) );
  INV_X1 U8550 ( .A(n11593), .ZN(n7504) );
  INV_X1 U8551 ( .A(n9434), .ZN(n7767) );
  OR2_X1 U8552 ( .A1(n8598), .A2(n8735), .ZN(n7326) );
  NAND2_X1 U8553 ( .A1(n7325), .A2(n8603), .ZN(n7324) );
  AND2_X1 U8554 ( .A1(n15160), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7325) );
  INV_X1 U8555 ( .A(n10539), .ZN(n9525) );
  OR2_X1 U8556 ( .A1(n10531), .A2(n9544), .ZN(n11296) );
  INV_X1 U8557 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n15815) );
  NAND2_X1 U8558 ( .A1(n8676), .A2(n8675), .ZN(n6961) );
  AND2_X1 U8559 ( .A1(n8718), .A2(n8709), .ZN(n9380) );
  INV_X1 U8560 ( .A(n9148), .ZN(n9165) );
  XNOR2_X1 U8561 ( .A(n9167), .B(SI_20_), .ZN(n9166) );
  INV_X1 U8562 ( .A(n8993), .ZN(n8979) );
  NAND2_X1 U8563 ( .A1(n7692), .A2(n7693), .ZN(n6978) );
  NAND2_X1 U8564 ( .A1(n8659), .A2(n10974), .ZN(n9015) );
  NAND2_X1 U8565 ( .A1(n7179), .A2(n8663), .ZN(n6848) );
  AND2_X1 U8566 ( .A1(n9060), .A2(n10860), .ZN(n9014) );
  NAND2_X1 U8567 ( .A1(n8724), .A2(n8725), .ZN(n8726) );
  NAND2_X1 U8568 ( .A1(n9045), .A2(n6611), .ZN(n7175) );
  INV_X1 U8569 ( .A(n9047), .ZN(n7179) );
  NAND2_X1 U8570 ( .A1(n9045), .A2(n8662), .ZN(n7180) );
  XNOR2_X1 U8571 ( .A(n8657), .B(SI_13_), .ZN(n9086) );
  NAND2_X1 U8572 ( .A1(n8650), .A2(n10546), .ZN(n8969) );
  NAND2_X1 U8573 ( .A1(n6883), .A2(n10440), .ZN(n8751) );
  INV_X1 U8574 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6799) );
  INV_X1 U8575 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n6800) );
  INV_X1 U8576 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7181) );
  XNOR2_X1 U8577 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n10470) );
  XNOR2_X1 U8578 ( .A(n7055), .B(n7287), .ZN(n10467) );
  INV_X1 U8579 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7287) );
  INV_X1 U8580 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n10463) );
  OAI21_X1 U8581 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n10780), .A(n10779), .ZN(
        n11002) );
  NAND2_X1 U8582 ( .A1(n11321), .A2(n11320), .ZN(n11558) );
  NAND2_X1 U8583 ( .A1(n11560), .A2(n11559), .ZN(n11563) );
  OR2_X1 U8584 ( .A1(n11558), .A2(n11557), .ZN(n11560) );
  OR2_X1 U8585 ( .A1(n11563), .A2(n11562), .ZN(n11913) );
  OR2_X1 U8586 ( .A1(n15174), .A2(n15173), .ZN(n15177) );
  NAND2_X1 U8587 ( .A1(n8491), .A2(n8477), .ZN(n7095) );
  NOR2_X1 U8588 ( .A1(n7714), .A2(n6562), .ZN(n7720) );
  NAND2_X1 U8589 ( .A1(n12799), .A2(n12232), .ZN(n12801) );
  XNOR2_X1 U8590 ( .A(n11423), .B(n11659), .ZN(n12814) );
  NAND2_X1 U8591 ( .A1(n7711), .A2(n7713), .ZN(n7710) );
  NAND2_X1 U8592 ( .A1(n7714), .A2(n12785), .ZN(n7713) );
  NOR2_X1 U8593 ( .A1(n7712), .A2(n6650), .ZN(n7711) );
  INV_X1 U8594 ( .A(n7720), .ZN(n7719) );
  XNOR2_X1 U8595 ( .A(n12224), .B(n12969), .ZN(n12831) );
  AND2_X1 U8596 ( .A1(n7146), .A2(n7730), .ZN(n7145) );
  AOI21_X1 U8597 ( .B1(n7733), .B2(n7731), .A(n6621), .ZN(n7730) );
  NAND2_X1 U8598 ( .A1(n7149), .A2(n7147), .ZN(n7146) );
  INV_X1 U8599 ( .A(n7149), .ZN(n7148) );
  NAND2_X1 U8600 ( .A1(n12215), .A2(n12214), .ZN(n12864) );
  INV_X1 U8601 ( .A(n7160), .ZN(n7159) );
  XNOR2_X1 U8602 ( .A(n11421), .B(n7378), .ZN(n11423) );
  NOR2_X1 U8603 ( .A1(n12903), .A2(n7734), .ZN(n7733) );
  INV_X1 U8604 ( .A(n12441), .ZN(n7734) );
  INV_X1 U8605 ( .A(n12234), .ZN(n7728) );
  NAND2_X1 U8606 ( .A1(n12801), .A2(n12234), .ZN(n12327) );
  AND4_X1 U8607 ( .A1(n12567), .A2(n12566), .A3(n12565), .A4(n12564), .ZN(
        n13108) );
  AND4_X1 U8608 ( .A1(n8497), .A2(n8496), .A3(n8495), .A4(n8494), .ZN(n10391)
         );
  OR2_X1 U8609 ( .A1(n12563), .A2(n15737), .ZN(n6859) );
  NAND2_X1 U8610 ( .A1(n6868), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n6874) );
  INV_X1 U8611 ( .A(n12562), .ZN(n6868) );
  OAI21_X1 U8612 ( .B1(n11197), .B2(n7892), .A(n7893), .ZN(n11191) );
  NOR2_X1 U8613 ( .A1(n11191), .A2(n15541), .ZN(n11190) );
  NOR2_X1 U8614 ( .A1(n11188), .A2(n11189), .ZN(n11187) );
  XNOR2_X1 U8615 ( .A(n11161), .B(n6899), .ZN(n11146) );
  NOR2_X1 U8616 ( .A1(n11145), .A2(n11146), .ZN(n11144) );
  NAND2_X1 U8617 ( .A1(n7968), .A2(n10451), .ZN(n7969) );
  NAND2_X1 U8618 ( .A1(n11036), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U8619 ( .A1(n7224), .A2(n7225), .ZN(n11097) );
  NAND2_X1 U8620 ( .A1(n7483), .A2(n6911), .ZN(n7908) );
  NAND2_X1 U8621 ( .A1(n11216), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n11375) );
  AND2_X1 U8622 ( .A1(n7221), .A2(n7220), .ZN(n11373) );
  AOI21_X1 U8623 ( .B1(n11101), .B2(n6911), .A(n6905), .ZN(n6904) );
  INV_X1 U8624 ( .A(n6908), .ZN(n6907) );
  NAND2_X1 U8625 ( .A1(n6906), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U8626 ( .A1(n7972), .A2(n10454), .ZN(n7456) );
  NAND2_X1 U8627 ( .A1(n6901), .A2(n6938), .ZN(n7457) );
  NOR2_X1 U8628 ( .A1(n7458), .A2(n11832), .ZN(n11833) );
  NAND2_X1 U8629 ( .A1(n7456), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7458) );
  INV_X1 U8630 ( .A(n7912), .ZN(n11841) );
  AND2_X1 U8631 ( .A1(n11839), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7486) );
  NAND2_X1 U8632 ( .A1(n7470), .A2(n7472), .ZN(n7471) );
  AND3_X1 U8633 ( .A1(n7234), .A2(n7921), .A3(P3_REG1_REG_11__SCAN_IN), .ZN(
        n12983) );
  NAND2_X1 U8634 ( .A1(n7232), .A2(n7230), .ZN(n7923) );
  OAI21_X1 U8635 ( .B1(n7921), .B2(n6583), .A(n7227), .ZN(n7230) );
  AOI21_X1 U8636 ( .B1(n7235), .B2(n7229), .A(n7228), .ZN(n7227) );
  NOR2_X1 U8637 ( .A1(n6583), .A2(n12982), .ZN(n7229) );
  AOI21_X1 U8638 ( .B1(n7443), .B2(n7440), .A(n6705), .ZN(n7439) );
  INV_X1 U8639 ( .A(n7443), .ZN(n7441) );
  AND2_X1 U8640 ( .A1(n13015), .A2(n6599), .ZN(n13001) );
  OR2_X1 U8641 ( .A1(n7926), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7929) );
  NOR2_X1 U8642 ( .A1(n13009), .A2(n13010), .ZN(n13008) );
  NAND2_X1 U8643 ( .A1(n13001), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n13017) );
  NAND2_X1 U8644 ( .A1(n7462), .A2(n7461), .ZN(n7460) );
  INV_X1 U8645 ( .A(n13016), .ZN(n7461) );
  NAND2_X1 U8646 ( .A1(n13001), .A2(n7463), .ZN(n7459) );
  NOR2_X1 U8647 ( .A1(n13016), .A2(n13309), .ZN(n7463) );
  INV_X1 U8648 ( .A(n7937), .ZN(n13039) );
  NAND2_X1 U8649 ( .A1(n13057), .A2(n13056), .ZN(n13055) );
  NAND2_X1 U8650 ( .A1(n13039), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n13045) );
  NAND2_X1 U8651 ( .A1(n6580), .A2(n6917), .ZN(n13052) );
  NAND2_X1 U8652 ( .A1(n13055), .A2(n8028), .ZN(n13069) );
  AOI21_X1 U8653 ( .B1(n7427), .B2(n7429), .A(n6707), .ZN(n7425) );
  NAND2_X1 U8654 ( .A1(n6928), .A2(n6927), .ZN(n6926) );
  INV_X1 U8655 ( .A(n13098), .ZN(n6928) );
  NAND2_X1 U8656 ( .A1(n6551), .A2(n6586), .ZN(n6929) );
  OR2_X1 U8657 ( .A1(n8474), .A2(n7030), .ZN(n7029) );
  INV_X1 U8658 ( .A(n13142), .ZN(n6780) );
  AOI21_X1 U8659 ( .B1(n7387), .B2(n7385), .A(n6785), .ZN(n13141) );
  INV_X1 U8660 ( .A(n13139), .ZN(n6785) );
  NOR2_X1 U8661 ( .A1(n13159), .A2(n7122), .ZN(n13152) );
  INV_X1 U8662 ( .A(n13150), .ZN(n7122) );
  AND2_X1 U8663 ( .A1(n12618), .A2(n12620), .ZN(n13171) );
  AND2_X1 U8664 ( .A1(n8358), .A2(n8374), .ZN(n7034) );
  NOR2_X2 U8665 ( .A1(n8345), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8359) );
  NOR2_X1 U8666 ( .A1(n7348), .A2(n7346), .ZN(n7345) );
  INV_X1 U8667 ( .A(n8320), .ZN(n7346) );
  NAND2_X1 U8668 ( .A1(n7347), .A2(n8320), .ZN(n13240) );
  NOR3_X1 U8669 ( .A1(n8285), .A2(P3_REG3_REG_16__SCAN_IN), .A3(
        P3_REG3_REG_15__SCAN_IN), .ZN(n8313) );
  INV_X1 U8670 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8312) );
  NOR2_X1 U8671 ( .A1(n8285), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8300) );
  OR2_X1 U8672 ( .A1(n8263), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8285) );
  NOR2_X1 U8673 ( .A1(n8250), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8261) );
  INV_X1 U8674 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U8675 ( .A1(n8261), .A2(n8260), .ZN(n8263) );
  NAND2_X1 U8676 ( .A1(n11848), .A2(n8163), .ZN(n11970) );
  INV_X1 U8677 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8164) );
  AND2_X1 U8678 ( .A1(n8165), .A2(n8164), .ZN(n8190) );
  INV_X1 U8679 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7035) );
  NOR2_X1 U8680 ( .A1(n8149), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8165) );
  XNOR2_X1 U8681 ( .A(n12970), .B(n12777), .ZN(n12656) );
  NAND2_X1 U8682 ( .A1(n7352), .A2(n8099), .ZN(n7354) );
  AND2_X1 U8683 ( .A1(n11645), .A2(n8118), .ZN(n7352) );
  OAI22_X1 U8684 ( .A1(n8177), .A2(n10447), .B1(n8508), .B2(n11215), .ZN(n6792) );
  NOR2_X1 U8685 ( .A1(n12569), .A2(SI_5_), .ZN(n6791) );
  AOI21_X1 U8686 ( .B1(n12634), .B2(n8550), .A(n8549), .ZN(n8551) );
  AND2_X1 U8687 ( .A1(n11245), .A2(n13374), .ZN(n11536) );
  INV_X1 U8688 ( .A(n11643), .ZN(n15489) );
  NAND2_X1 U8689 ( .A1(n8578), .A2(n8577), .ZN(n15511) );
  INV_X1 U8690 ( .A(n13471), .ZN(n9414) );
  NOR2_X1 U8691 ( .A1(n7419), .A2(n13125), .ZN(n7418) );
  NOR2_X1 U8692 ( .A1(n7420), .A2(n12738), .ZN(n7419) );
  AOI21_X1 U8693 ( .B1(n7418), .B2(n7420), .A(n7417), .ZN(n7416) );
  INV_X1 U8694 ( .A(n12746), .ZN(n7417) );
  INV_X1 U8695 ( .A(n12735), .ZN(n13140) );
  OAI21_X1 U8696 ( .B1(n13221), .B2(n7374), .A(n7373), .ZN(n13197) );
  AOI21_X1 U8697 ( .B1(n7375), .B2(n13220), .A(n6642), .ZN(n7373) );
  INV_X1 U8698 ( .A(n7375), .ZN(n7374) );
  OR2_X1 U8699 ( .A1(n8567), .A2(n8566), .ZN(n13216) );
  AND2_X1 U8700 ( .A1(n12711), .A2(n12715), .ZN(n13259) );
  AOI21_X1 U8701 ( .B1(n7405), .B2(n12593), .A(n6880), .ZN(n6879) );
  NAND2_X1 U8702 ( .A1(n13301), .A2(n7405), .ZN(n6881) );
  INV_X1 U8703 ( .A(n7407), .ZN(n6880) );
  OR2_X1 U8704 ( .A1(n12275), .A2(n8231), .ZN(n7359) );
  INV_X1 U8705 ( .A(n7393), .ZN(n7392) );
  NAND2_X1 U8706 ( .A1(n7395), .A2(n12113), .ZN(n6875) );
  OAI21_X1 U8707 ( .B1(n7396), .B2(n7394), .A(n12684), .ZN(n7393) );
  INV_X1 U8708 ( .A(n8180), .ZN(n6784) );
  AND2_X1 U8709 ( .A1(n6782), .A2(n8182), .ZN(n6781) );
  AND2_X1 U8710 ( .A1(n12672), .A2(n12671), .ZN(n12594) );
  NAND2_X1 U8711 ( .A1(n8535), .A2(n9419), .ZN(n11247) );
  NAND2_X1 U8712 ( .A1(n8519), .A2(n8520), .ZN(n10879) );
  AND2_X1 U8713 ( .A1(n7957), .A2(P3_STATE_REG_SCAN_IN), .ZN(n7950) );
  NAND2_X1 U8714 ( .A1(n7010), .A2(n8469), .ZN(n8484) );
  XNOR2_X1 U8715 ( .A(n8437), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n8435) );
  INV_X1 U8716 ( .A(n7654), .ZN(n7653) );
  INV_X1 U8717 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n15823) );
  OR2_X1 U8718 ( .A1(n7883), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7913) );
  INV_X1 U8719 ( .A(n7669), .ZN(n7668) );
  CLKBUF_X1 U8720 ( .A(n7891), .Z(n7964) );
  OR2_X1 U8721 ( .A1(n9959), .A2(n13596), .ZN(n9984) );
  NAND2_X1 U8722 ( .A1(n9971), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9986) );
  INV_X1 U8723 ( .A(n9984), .ZN(n9971) );
  AND2_X1 U8724 ( .A1(n6581), .A2(n13496), .ZN(n6982) );
  XNOR2_X1 U8725 ( .A(n9645), .B(n10871), .ZN(n9626) );
  NAND2_X1 U8726 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9686) );
  OR2_X1 U8727 ( .A1(n11753), .A2(n11754), .ZN(n11751) );
  NOR2_X1 U8728 ( .A1(n13611), .A2(n7636), .ZN(n7635) );
  INV_X1 U8729 ( .A(n9897), .ZN(n7636) );
  INV_X1 U8730 ( .A(n9911), .ZN(n7634) );
  OR2_X1 U8731 ( .A1(n13585), .A2(n13586), .ZN(n13583) );
  NAND2_X1 U8732 ( .A1(n7098), .A2(n9765), .ZN(n9783) );
  AND2_X1 U8733 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n9765) );
  INV_X1 U8734 ( .A(n9767), .ZN(n7098) );
  NAND2_X1 U8735 ( .A1(n13560), .A2(n7635), .ZN(n13608) );
  NAND2_X1 U8736 ( .A1(n7620), .A2(n7613), .ZN(n7611) );
  NAND2_X1 U8737 ( .A1(n13503), .A2(n9845), .ZN(n13546) );
  INV_X1 U8738 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9850) );
  AND2_X1 U8739 ( .A1(n9755), .A2(n9754), .ZN(n11788) );
  NAND2_X1 U8740 ( .A1(n15354), .A2(n15353), .ZN(n15352) );
  NAND2_X1 U8741 ( .A1(n15365), .A2(n15366), .ZN(n15364) );
  NAND2_X1 U8742 ( .A1(n15379), .A2(n15380), .ZN(n15378) );
  OR2_X1 U8743 ( .A1(n10934), .A2(n10933), .ZN(n10944) );
  NAND2_X1 U8744 ( .A1(n15393), .A2(n11465), .ZN(n15416) );
  AOI21_X1 U8745 ( .B1(n11473), .B2(P2_REG1_REG_13__SCAN_IN), .A(n15419), .ZN(
        n11983) );
  OR2_X1 U8746 ( .A1(n12414), .A2(n12413), .ZN(n12416) );
  NOR2_X1 U8747 ( .A1(n7581), .A2(n14203), .ZN(n7580) );
  NAND2_X1 U8748 ( .A1(n13953), .A2(n13968), .ZN(n7581) );
  NAND2_X1 U8749 ( .A1(n13961), .A2(n14108), .ZN(n7136) );
  AND2_X1 U8750 ( .A1(n10040), .A2(n10016), .ZN(n13979) );
  NAND2_X1 U8751 ( .A1(n12543), .A2(n6573), .ZN(n14013) );
  INV_X1 U8752 ( .A(n7585), .ZN(n7584) );
  NAND2_X1 U8753 ( .A1(n14006), .A2(n14005), .ZN(n14004) );
  NOR2_X1 U8754 ( .A1(n14071), .A2(n7587), .ZN(n14047) );
  NAND2_X1 U8755 ( .A1(n7255), .A2(n7256), .ZN(n14070) );
  INV_X1 U8756 ( .A(n7257), .ZN(n7256) );
  OR2_X1 U8757 ( .A1(n14129), .A2(n6559), .ZN(n7255) );
  INV_X1 U8758 ( .A(n7101), .ZN(n9918) );
  INV_X1 U8759 ( .A(n12039), .ZN(n7241) );
  NAND2_X1 U8760 ( .A1(n6830), .A2(n6828), .ZN(n7240) );
  AOI21_X1 U8761 ( .B1(n7591), .B2(n12178), .A(n6655), .ZN(n7590) );
  INV_X1 U8762 ( .A(n7592), .ZN(n7591) );
  NOR2_X1 U8763 ( .A1(n14183), .A2(n14292), .ZN(n14182) );
  AND2_X1 U8764 ( .A1(n9788), .A2(n9787), .ZN(n13709) );
  AOI22_X1 U8765 ( .A1(n11890), .A2(n13858), .B1(n11891), .B2(n14302), .ZN(
        n12037) );
  NAND2_X1 U8766 ( .A1(n11889), .A2(n12036), .ZN(n12045) );
  AND2_X1 U8767 ( .A1(n11795), .A2(n11799), .ZN(n11889) );
  NAND2_X1 U8768 ( .A1(n11730), .A2(n7002), .ZN(n11743) );
  NOR2_X1 U8769 ( .A1(n14314), .A2(n13687), .ZN(n7002) );
  NOR2_X1 U8770 ( .A1(n11743), .A2(n14307), .ZN(n11795) );
  NAND2_X1 U8771 ( .A1(n11785), .A2(n11789), .ZN(n11738) );
  INV_X1 U8772 ( .A(n11725), .ZN(n7549) );
  NAND2_X1 U8773 ( .A1(n9704), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9721) );
  INV_X1 U8774 ( .A(n9705), .ZN(n9704) );
  INV_X1 U8775 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n15585) );
  NOR2_X2 U8776 ( .A1(n11706), .A2(n15438), .ZN(n11730) );
  NAND2_X1 U8777 ( .A1(n11730), .A2(n15452), .ZN(n11745) );
  INV_X1 U8778 ( .A(n13662), .ZN(n13659) );
  NAND2_X1 U8779 ( .A1(n11340), .A2(n7576), .ZN(n10985) );
  OAI21_X1 U8780 ( .B1(n13846), .B2(n10865), .A(n10866), .ZN(n10868) );
  OR2_X1 U8781 ( .A1(n6543), .A2(n11068), .ZN(n10872) );
  INV_X1 U8782 ( .A(n13650), .ZN(n13848) );
  NOR2_X1 U8783 ( .A1(n10871), .A2(n11717), .ZN(n10869) );
  INV_X1 U8784 ( .A(n14315), .ZN(n15451) );
  OAI21_X1 U8785 ( .B1(n10410), .B2(n12354), .A(n11907), .ZN(n10098) );
  INV_X1 U8786 ( .A(n9599), .ZN(n9600) );
  XNOR2_X1 U8787 ( .A(n10060), .B(P2_IR_REG_26__SCAN_IN), .ZN(n10411) );
  OR2_X1 U8788 ( .A1(n9863), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n9898) );
  AND2_X1 U8789 ( .A1(n9796), .A2(n9828), .ZN(n11472) );
  NOR2_X1 U8790 ( .A1(n9236), .A2(n14527), .ZN(n9252) );
  AOI21_X1 U8791 ( .B1(n14479), .B2(n14478), .A(n10217), .ZN(n14375) );
  OR2_X1 U8792 ( .A1(n9176), .A2(n14494), .ZN(n9189) );
  AND2_X1 U8793 ( .A1(n11898), .A2(n10183), .ZN(n12289) );
  NAND2_X1 U8794 ( .A1(n7820), .A2(n6622), .ZN(n14398) );
  NOR2_X1 U8795 ( .A1(n6593), .A2(n7822), .ZN(n7821) );
  NOR2_X1 U8796 ( .A1(n9054), .A2(n9009), .ZN(n9025) );
  NOR2_X1 U8797 ( .A1(n7796), .A2(n6633), .ZN(n7795) );
  NAND2_X1 U8798 ( .A1(n14442), .A2(n14444), .ZN(n14441) );
  OR2_X1 U8799 ( .A1(n10310), .A2(n10150), .ZN(n10151) );
  NAND2_X1 U8800 ( .A1(n8896), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8927) );
  AND2_X1 U8801 ( .A1(n8963), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9078) );
  NAND2_X1 U8802 ( .A1(n7802), .A2(n7799), .ZN(n14501) );
  NAND2_X1 U8803 ( .A1(n7801), .A2(n7800), .ZN(n7799) );
  NAND2_X1 U8804 ( .A1(n10197), .A2(n10183), .ZN(n7800) );
  INV_X1 U8805 ( .A(n10314), .ZN(n10305) );
  AND2_X1 U8806 ( .A1(n15165), .A2(n9308), .ZN(n10539) );
  NAND2_X1 U8807 ( .A1(n7276), .A2(n7273), .ZN(n9348) );
  AND2_X1 U8808 ( .A1(n9007), .A2(n9006), .ZN(n14910) );
  OR2_X1 U8809 ( .A1(n9257), .A2(n10749), .ZN(n8763) );
  OR2_X1 U8810 ( .A1(n10838), .A2(n10837), .ZN(n11029) );
  NAND2_X1 U8811 ( .A1(n11029), .A2(n11028), .ZN(n11030) );
  NAND2_X1 U8812 ( .A1(n11135), .A2(n11134), .ZN(n11137) );
  OR2_X1 U8813 ( .A1(n11201), .A2(n11202), .ZN(n11804) );
  OR2_X1 U8814 ( .A1(n11137), .A2(n11136), .ZN(n11210) );
  OR2_X1 U8815 ( .A1(n11960), .A2(n11959), .ZN(n12198) );
  NAND2_X1 U8816 ( .A1(n10372), .A2(n12472), .ZN(n10350) );
  NAND2_X1 U8817 ( .A1(n7792), .A2(n9470), .ZN(n7789) );
  INV_X1 U8818 ( .A(n14529), .ZN(n14749) );
  NAND2_X1 U8819 ( .A1(n9202), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U8820 ( .A1(n14834), .A2(n7508), .ZN(n14783) );
  INV_X1 U8821 ( .A(n9465), .ZN(n7788) );
  OAI21_X1 U8822 ( .B1(n7015), .B2(n6736), .A(n14827), .ZN(n6735) );
  INV_X1 U8823 ( .A(n14828), .ZN(n6736) );
  AOI21_X1 U8824 ( .B1(n7775), .B2(n7777), .A(n7773), .ZN(n7772) );
  INV_X1 U8825 ( .A(n9462), .ZN(n7773) );
  NAND2_X1 U8826 ( .A1(n14906), .A2(n14894), .ZN(n14889) );
  NAND2_X1 U8827 ( .A1(n9078), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9080) );
  INV_X1 U8828 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9071) );
  OR2_X1 U8829 ( .A1(n9080), .A2(n9071), .ZN(n9073) );
  NAND2_X1 U8830 ( .A1(n14959), .A2(n14960), .ZN(n7741) );
  INV_X1 U8831 ( .A(n7501), .ZN(n14977) );
  NAND2_X1 U8832 ( .A1(n14983), .A2(n14982), .ZN(n14981) );
  NAND2_X1 U8833 ( .A1(n12057), .A2(n7748), .ZN(n12056) );
  NAND2_X1 U8834 ( .A1(n11516), .A2(n9492), .ZN(n11874) );
  AND2_X1 U8835 ( .A1(n11858), .A2(n12301), .ZN(n11880) );
  OR2_X1 U8836 ( .A1(n10549), .A2(n9296), .ZN(n8913) );
  INV_X1 U8837 ( .A(n9488), .ZN(n7025) );
  NAND2_X1 U8838 ( .A1(n7504), .A2(n6603), .ZN(n11857) );
  NAND2_X1 U8839 ( .A1(n11938), .A2(n9488), .ZN(n7757) );
  NOR2_X1 U8840 ( .A1(n11593), .A2(n11605), .ZN(n11944) );
  NAND2_X1 U8841 ( .A1(n9439), .A2(n9438), .ZN(n11582) );
  NAND2_X1 U8842 ( .A1(n11302), .A2(n9486), .ZN(n11586) );
  AND2_X1 U8843 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8841) );
  NOR2_X2 U8844 ( .A1(n11443), .A2(n11362), .ZN(n15287) );
  INV_X1 U8845 ( .A(n9357), .ZN(n11360) );
  OR2_X1 U8846 ( .A1(n15323), .A2(n8984), .ZN(n10332) );
  OR2_X1 U8847 ( .A1(n9525), .A2(n14587), .ZN(n14909) );
  NAND2_X1 U8848 ( .A1(n9297), .A2(n9286), .ZN(n9299) );
  INV_X1 U8849 ( .A(n14753), .ZN(n15002) );
  NAND2_X1 U8850 ( .A1(n14906), .A2(n7506), .ZN(n14857) );
  AND2_X1 U8851 ( .A1(n14936), .A2(n9496), .ZN(n14923) );
  INV_X1 U8852 ( .A(n14507), .ZN(n15087) );
  AND2_X1 U8853 ( .A1(n9524), .A2(n9523), .ZN(n15295) );
  AND3_X1 U8854 ( .A1(n10319), .A2(n10332), .A3(n11296), .ZN(n9551) );
  INV_X1 U8855 ( .A(n9394), .ZN(n9395) );
  AND2_X1 U8856 ( .A1(n10409), .A2(n10408), .ZN(n10536) );
  AOI21_X1 U8857 ( .B1(n7280), .B2(n7278), .A(n6708), .ZN(n7277) );
  INV_X1 U8858 ( .A(n7280), .ZN(n7279) );
  AND2_X1 U8859 ( .A1(n8718), .A2(n7187), .ZN(n7186) );
  AND2_X1 U8860 ( .A1(n15718), .A2(n8595), .ZN(n7187) );
  NAND2_X1 U8861 ( .A1(n9276), .A2(n9275), .ZN(n9323) );
  NAND2_X1 U8862 ( .A1(n9276), .A2(n8701), .ZN(n14355) );
  NAND2_X1 U8863 ( .A1(n7269), .A2(n8692), .ZN(n9246) );
  NAND2_X1 U8864 ( .A1(n8688), .A2(n7270), .ZN(n7269) );
  NAND2_X1 U8865 ( .A1(n8688), .A2(n8687), .ZN(n9225) );
  INV_X1 U8866 ( .A(n6958), .ZN(n6957) );
  OAI21_X1 U8867 ( .B1(n8675), .B2(n6597), .A(n6959), .ZN(n6958) );
  XNOR2_X1 U8868 ( .A(n8733), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9308) );
  NAND2_X1 U8869 ( .A1(n7830), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8733) );
  AND2_X1 U8870 ( .A1(n8723), .A2(n7830), .ZN(n9521) );
  NAND2_X1 U8871 ( .A1(n8716), .A2(n7828), .ZN(n8721) );
  AND2_X1 U8872 ( .A1(n8728), .A2(n6813), .ZN(n6812) );
  NAND2_X1 U8873 ( .A1(n9021), .A2(n8728), .ZN(n6815) );
  XNOR2_X1 U8874 ( .A(n9069), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11805) );
  OR2_X1 U8875 ( .A1(n8956), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n8957) );
  NAND2_X1 U8876 ( .A1(n8649), .A2(n10528), .ZN(n7185) );
  INV_X1 U8877 ( .A(n8643), .ZN(n6963) );
  INV_X1 U8878 ( .A(n8642), .ZN(n6964) );
  AND2_X1 U8879 ( .A1(n8647), .A2(n8646), .ZN(n8907) );
  OR2_X1 U8880 ( .A1(n8910), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U8881 ( .A1(n8892), .A2(n8891), .ZN(n8893) );
  OR2_X1 U8882 ( .A1(n8859), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8872) );
  NAND2_X1 U8883 ( .A1(n8874), .A2(n8873), .ZN(n8910) );
  INV_X1 U8884 ( .A(n8872), .ZN(n8874) );
  NAND2_X1 U8885 ( .A1(n8716), .A2(n8715), .ZN(n8859) );
  INV_X1 U8886 ( .A(n8854), .ZN(n8856) );
  INV_X1 U8887 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10473) );
  AND2_X1 U8888 ( .A1(n10473), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10471) );
  AND2_X1 U8889 ( .A1(n10460), .A2(n10459), .ZN(n10468) );
  NAND2_X1 U8890 ( .A1(n11317), .A2(n11316), .ZN(n11552) );
  INV_X1 U8891 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7042) );
  AND2_X1 U8892 ( .A1(n11555), .A2(n6656), .ZN(n7045) );
  OR2_X1 U8893 ( .A1(n11555), .A2(n6656), .ZN(n7044) );
  INV_X1 U8894 ( .A(n11919), .ZN(n7294) );
  AND2_X1 U8895 ( .A1(n6656), .A2(n7042), .ZN(n7041) );
  INV_X1 U8896 ( .A(n7095), .ZN(n13132) );
  NAND2_X1 U8897 ( .A1(n7140), .A2(n7724), .ZN(n12344) );
  NAND2_X1 U8898 ( .A1(n12799), .A2(n6560), .ZN(n7140) );
  NAND2_X1 U8899 ( .A1(n12344), .A2(n12343), .ZN(n12428) );
  AND2_X1 U8900 ( .A1(n8334), .A2(n8333), .ZN(n13232) );
  NAND2_X1 U8901 ( .A1(n12823), .A2(n12822), .ZN(n12821) );
  NAND2_X1 U8902 ( .A1(n12917), .A2(n12439), .ZN(n12823) );
  AND4_X1 U8903 ( .A1(n12567), .A2(n8513), .A3(n8512), .A4(n8511), .ZN(n12576)
         );
  OAI21_X1 U8904 ( .B1(n12793), .B2(n12446), .A(n12450), .ZN(n12457) );
  OAI21_X1 U8905 ( .B1(n12454), .B2(n12453), .A(n12452), .ZN(n12455) );
  INV_X1 U8906 ( .A(n11770), .ZN(n12868) );
  NAND2_X1 U8907 ( .A1(n6941), .A2(n12433), .ZN(n12875) );
  NAND2_X1 U8908 ( .A1(n6941), .A2(n6554), .ZN(n12876) );
  NAND2_X1 U8909 ( .A1(n12821), .A2(n12441), .ZN(n12902) );
  OR2_X1 U8910 ( .A1(n12569), .A2(SI_2_), .ZN(n8084) );
  OR2_X1 U8911 ( .A1(n11257), .A2(n11256), .ZN(n12922) );
  NAND2_X1 U8912 ( .A1(n6940), .A2(n6939), .ZN(n12919) );
  AOI21_X1 U8913 ( .B1(n6554), .B2(n12431), .A(n6709), .ZN(n6939) );
  NAND2_X1 U8914 ( .A1(n12856), .A2(n6554), .ZN(n6940) );
  NAND2_X1 U8915 ( .A1(n12919), .A2(n12918), .ZN(n12917) );
  NAND2_X1 U8916 ( .A1(n8327), .A2(n8326), .ZN(n13247) );
  AND2_X1 U8917 ( .A1(n11255), .A2(n11256), .ZN(n12933) );
  INV_X1 U8918 ( .A(n12922), .ZN(n12951) );
  NAND2_X1 U8919 ( .A1(n11242), .A2(n11241), .ZN(n12952) );
  OR2_X1 U8920 ( .A1(n7724), .A2(n7139), .ZN(n7137) );
  NAND2_X1 U8921 ( .A1(n7388), .A2(n6646), .ZN(n7321) );
  INV_X1 U8922 ( .A(n7389), .ZN(n7322) );
  AND4_X1 U8923 ( .A1(n12567), .A2(n10388), .A3(n10387), .A4(n10386), .ZN(
        n12584) );
  INV_X1 U8924 ( .A(n13154), .ZN(n13129) );
  OR2_X1 U8925 ( .A1(n12562), .A2(n8442), .ZN(n8447) );
  INV_X1 U8926 ( .A(n13181), .ZN(n12965) );
  INV_X1 U8927 ( .A(n13232), .ZN(n13261) );
  INV_X1 U8928 ( .A(n13272), .ZN(n13295) );
  OR2_X1 U8929 ( .A1(n12562), .A2(n15544), .ZN(n8137) );
  INV_X1 U8930 ( .A(n7205), .ZN(n11150) );
  NAND2_X1 U8931 ( .A1(n7487), .A2(n7912), .ZN(n11634) );
  OAI21_X1 U8932 ( .B1(n12098), .B2(n12097), .A(n12096), .ZN(n12095) );
  AND2_X1 U8933 ( .A1(n7232), .A2(n7231), .ZN(n10419) );
  AOI21_X1 U8934 ( .B1(n10420), .B2(n7465), .A(n6718), .ZN(n7464) );
  NAND2_X1 U8935 ( .A1(n7444), .A2(n7442), .ZN(n10414) );
  INV_X1 U8936 ( .A(n7446), .ZN(n7442) );
  NAND2_X1 U8937 ( .A1(n7924), .A2(n7925), .ZN(n12992) );
  OR2_X1 U8938 ( .A1(n7923), .A2(n12998), .ZN(n7924) );
  NAND2_X1 U8939 ( .A1(n7459), .A2(n7460), .ZN(n13019) );
  NAND2_X1 U8940 ( .A1(n6917), .A2(n13050), .ZN(n13029) );
  INV_X1 U8941 ( .A(n7206), .ZN(n7479) );
  NAND2_X1 U8942 ( .A1(n6915), .A2(n13049), .ZN(n13054) );
  NAND2_X1 U8943 ( .A1(n6916), .A2(n13050), .ZN(n6915) );
  NAND2_X1 U8944 ( .A1(n6917), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U8945 ( .A1(n6929), .A2(n6926), .ZN(n13102) );
  NAND2_X1 U8946 ( .A1(n7984), .A2(n13079), .ZN(n13084) );
  INV_X1 U8947 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n7121) );
  XNOR2_X1 U8948 ( .A(n13126), .B(n13125), .ZN(n13335) );
  XNOR2_X1 U8949 ( .A(n6789), .B(n6788), .ZN(n13271) );
  INV_X1 U8950 ( .A(n13270), .ZN(n6788) );
  NAND2_X1 U8951 ( .A1(n8298), .A2(n8297), .ZN(n13373) );
  INV_X1 U8952 ( .A(n6529), .ZN(n15483) );
  NAND2_X2 U8953 ( .A1(n11537), .A2(n15486), .ZN(n15500) );
  AND2_X1 U8954 ( .A1(n8574), .A2(n13374), .ZN(n7078) );
  AND2_X1 U8955 ( .A1(n13348), .A2(n13347), .ZN(n13406) );
  NAND2_X1 U8956 ( .A1(n7397), .A2(n7402), .ZN(n13195) );
  NAND2_X1 U8957 ( .A1(n13214), .A2(n6553), .ZN(n7397) );
  NAND2_X1 U8958 ( .A1(n7377), .A2(n8366), .ZN(n13206) );
  NAND2_X1 U8959 ( .A1(n13221), .A2(n13218), .ZN(n7377) );
  NAND2_X1 U8960 ( .A1(n7404), .A2(n8569), .ZN(n13204) );
  OR2_X1 U8961 ( .A1(n13214), .A2(n8565), .ZN(n7404) );
  NAND2_X1 U8962 ( .A1(n7363), .A2(n7360), .ZN(n13282) );
  NAND2_X1 U8963 ( .A1(n12276), .A2(n7364), .ZN(n7363) );
  NAND2_X1 U8964 ( .A1(n7410), .A2(n12697), .ZN(n13280) );
  NAND2_X1 U8965 ( .A1(n8564), .A2(n7411), .ZN(n7410) );
  NAND2_X1 U8966 ( .A1(n8564), .A2(n12694), .ZN(n13289) );
  NAND2_X1 U8967 ( .A1(n8249), .A2(n8248), .ZN(n13469) );
  NAND2_X1 U8968 ( .A1(n12115), .A2(n7395), .ZN(n12278) );
  INV_X1 U8969 ( .A(n11436), .ZN(n15472) );
  INV_X1 U8970 ( .A(n7950), .ZN(n13472) );
  XNOR2_X1 U8971 ( .A(n12559), .B(n12558), .ZN(n13481) );
  NAND2_X1 U8972 ( .A1(n12556), .A2(n12555), .ZN(n12559) );
  AND2_X1 U8973 ( .A1(n7864), .A2(n6865), .ZN(n6864) );
  AND2_X1 U8974 ( .A1(n8046), .A2(n7736), .ZN(n6865) );
  NAND2_X1 U8975 ( .A1(n7678), .A2(n7682), .ZN(n12568) );
  OAI21_X1 U8976 ( .B1(n8049), .B2(n13475), .A(n8048), .ZN(n8050) );
  NAND2_X1 U8977 ( .A1(n7867), .A2(n7959), .ZN(n13493) );
  INV_X1 U8978 ( .A(SI_25_), .ZN(n12285) );
  XNOR2_X1 U8979 ( .A(n7868), .B(n15810), .ZN(n12286) );
  NAND2_X1 U8980 ( .A1(n6947), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7868) );
  AND2_X1 U8981 ( .A1(n7737), .A2(n7860), .ZN(n6946) );
  NAND2_X1 U8982 ( .A1(n7872), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U8983 ( .A1(n7645), .A2(n7643), .ZN(n8422) );
  NAND2_X1 U8984 ( .A1(n7645), .A2(n8403), .ZN(n8408) );
  XNOR2_X1 U8985 ( .A(n7956), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12766) );
  NAND2_X1 U8986 ( .A1(n7167), .A2(n7165), .ZN(n12627) );
  OR2_X1 U8987 ( .A1(n7953), .A2(n7858), .ZN(n7167) );
  NOR2_X1 U8988 ( .A1(n7954), .A2(n7166), .ZN(n7165) );
  NAND2_X1 U8989 ( .A1(n8502), .A2(n8501), .ZN(n11385) );
  NAND2_X1 U8990 ( .A1(n7652), .A2(n8355), .ZN(n8369) );
  NAND2_X1 U8991 ( .A1(n8354), .A2(n8353), .ZN(n7652) );
  INV_X1 U8992 ( .A(SI_19_), .ZN(n11163) );
  NAND2_X1 U8993 ( .A1(n7948), .A2(n8499), .ZN(n12613) );
  INV_X1 U8994 ( .A(SI_18_), .ZN(n15667) );
  INV_X1 U8995 ( .A(n7640), .ZN(n8322) );
  AOI21_X1 U8996 ( .B1(n8307), .B2(n8306), .A(n7642), .ZN(n7640) );
  INV_X1 U8997 ( .A(SI_15_), .ZN(n10974) );
  INV_X1 U8998 ( .A(n7657), .ZN(n8293) );
  AOI21_X1 U8999 ( .B1(n7663), .B2(n7661), .A(n7660), .ZN(n7657) );
  INV_X1 U9000 ( .A(SI_14_), .ZN(n10860) );
  NAND2_X1 U9001 ( .A1(n7663), .A2(n8236), .ZN(n8279) );
  NAND2_X1 U9002 ( .A1(n8235), .A2(n8234), .ZN(n8257) );
  INV_X1 U9003 ( .A(SI_12_), .ZN(n10568) );
  INV_X1 U9004 ( .A(SI_11_), .ZN(n10546) );
  NAND2_X1 U9005 ( .A1(n8220), .A2(n8219), .ZN(n8233) );
  INV_X1 U9006 ( .A(SI_10_), .ZN(n10528) );
  INV_X1 U9007 ( .A(SI_9_), .ZN(n10496) );
  INV_X1 U9008 ( .A(n7667), .ZN(n8184) );
  AOI21_X1 U9009 ( .B1(n7673), .B2(n7671), .A(n7670), .ZN(n7667) );
  NAND2_X1 U9010 ( .A1(n7673), .A2(n7676), .ZN(n8175) );
  NAND2_X1 U9011 ( .A1(n8144), .A2(n8129), .ZN(n8158) );
  NAND2_X1 U9012 ( .A1(n7646), .A2(n8107), .ZN(n8113) );
  NAND2_X1 U9013 ( .A1(n8097), .A2(n8096), .ZN(n8109) );
  NAND2_X1 U9014 ( .A1(n11119), .A2(n9715), .ZN(n11167) );
  OR2_X1 U9015 ( .A1(n11059), .A2(n9629), .ZN(n9833) );
  NAND2_X1 U9016 ( .A1(n11751), .A2(n9761), .ZN(n11775) );
  NAND2_X1 U9017 ( .A1(n10995), .A2(n9644), .ZN(n11112) );
  NAND2_X1 U9018 ( .A1(n13608), .A2(n9911), .ZN(n13521) );
  NAND2_X1 U9019 ( .A1(n13583), .A2(n9945), .ZN(n13529) );
  NAND2_X1 U9020 ( .A1(n11694), .A2(n13785), .ZN(n7065) );
  AND2_X1 U9021 ( .A1(n9821), .A2(n9820), .ZN(n13720) );
  NAND2_X1 U9022 ( .A1(n7618), .A2(n9995), .ZN(n13536) );
  AND2_X1 U9023 ( .A1(n9881), .A2(n9880), .ZN(n13742) );
  NAND2_X1 U9024 ( .A1(n9619), .A2(n7245), .ZN(n13640) );
  NAND2_X1 U9025 ( .A1(n7247), .A2(n7246), .ZN(n7245) );
  INV_X1 U9026 ( .A(n7845), .ZN(n7246) );
  INV_X1 U9027 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13587) );
  NOR2_X1 U9028 ( .A1(n12317), .A2(n6990), .ZN(n6989) );
  INV_X1 U9029 ( .A(n12160), .ZN(n6990) );
  NAND2_X1 U9030 ( .A1(n6991), .A2(n12160), .ZN(n12318) );
  NAND2_X1 U9031 ( .A1(n7607), .A2(n7605), .ZN(n13595) );
  AOI21_X1 U9032 ( .B1(n13586), .B2(n6602), .A(n7606), .ZN(n7605) );
  NOR2_X1 U9033 ( .A1(n9954), .A2(n9953), .ZN(n7606) );
  AOI21_X1 U9034 ( .B1(n7630), .B2(n11754), .A(n6579), .ZN(n7628) );
  NAND2_X1 U9035 ( .A1(n13560), .A2(n9897), .ZN(n13610) );
  AND2_X1 U9036 ( .A1(n9925), .A2(n9924), .ZN(n13607) );
  AND2_X1 U9037 ( .A1(n6985), .A2(n6987), .ZN(n11121) );
  NOR2_X1 U9038 ( .A1(n9695), .A2(n6986), .ZN(n6985) );
  INV_X1 U9039 ( .A(n13891), .ZN(n13978) );
  NAND2_X1 U9040 ( .A1(n13550), .A2(n14108), .ZN(n13621) );
  NAND2_X1 U9041 ( .A1(n6984), .A2(n7611), .ZN(n13615) );
  INV_X1 U9042 ( .A(n7615), .ZN(n7612) );
  NAND2_X1 U9043 ( .A1(n7622), .A2(n7619), .ZN(n7617) );
  INV_X1 U9044 ( .A(n13625), .ZN(n13627) );
  NAND2_X1 U9045 ( .A1(n6748), .A2(n6747), .ZN(n13880) );
  NOR2_X1 U9046 ( .A1(n7836), .A2(n6651), .ZN(n6747) );
  NAND2_X1 U9047 ( .A1(n13778), .A2(n7515), .ZN(n6748) );
  INV_X1 U9048 ( .A(n13793), .ZN(n13961) );
  NAND2_X1 U9049 ( .A1(n10006), .A2(n10005), .ZN(n14007) );
  INV_X1 U9050 ( .A(n13607), .ZN(n14109) );
  INV_X1 U9051 ( .A(n13720), .ZN(n13896) );
  INV_X1 U9052 ( .A(n13709), .ZN(n13898) );
  INV_X1 U9053 ( .A(n6750), .ZN(n6749) );
  OAI21_X1 U9054 ( .B1(n12536), .B2(n11729), .A(n9720), .ZN(n6750) );
  NAND2_X1 U9055 ( .A1(n15357), .A2(n15356), .ZN(n15355) );
  NAND2_X1 U9056 ( .A1(n15368), .A2(n15369), .ZN(n15367) );
  NAND2_X1 U9057 ( .A1(n15382), .A2(n15383), .ZN(n15381) );
  OR2_X1 U9058 ( .A1(n10634), .A2(n10633), .ZN(n10924) );
  XNOR2_X1 U9059 ( .A(n11978), .B(n11981), .ZN(n11976) );
  AND2_X1 U9060 ( .A1(n10578), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15408) );
  AND2_X1 U9061 ( .A1(n10589), .A2(n10582), .ZN(n15394) );
  NAND2_X1 U9062 ( .A1(n13802), .A2(n13801), .ZN(n13942) );
  OR2_X1 U9063 ( .A1(n13800), .A2(n9629), .ZN(n13802) );
  XNOR2_X1 U9064 ( .A(n12519), .B(n13872), .ZN(n14205) );
  AND2_X1 U9065 ( .A1(n7583), .A2(n7582), .ZN(n14202) );
  OAI22_X1 U9066 ( .A1(n13963), .A2(n7579), .B1(n15453), .B2(n14203), .ZN(
        n7583) );
  NAND2_X1 U9067 ( .A1(n13953), .A2(n14308), .ZN(n7579) );
  AND2_X1 U9068 ( .A1(n13948), .A2(n7004), .ZN(n14206) );
  AOI21_X1 U9069 ( .B1(n13973), .B2(n7003), .A(n15453), .ZN(n7004) );
  NOR2_X1 U9070 ( .A1(n14207), .A2(n14211), .ZN(n7003) );
  OAI21_X1 U9071 ( .B1(n6834), .B2(n13955), .A(n13954), .ZN(n14210) );
  OAI21_X1 U9072 ( .B1(n7562), .B2(n14056), .A(n7560), .ZN(n14022) );
  AND2_X1 U9073 ( .A1(n7252), .A2(n12508), .ZN(n6835) );
  NAND2_X1 U9074 ( .A1(n7563), .A2(n7564), .ZN(n14039) );
  INV_X1 U9075 ( .A(n14246), .ZN(n14064) );
  NAND2_X1 U9076 ( .A1(n7574), .A2(n12526), .ZN(n14088) );
  NAND2_X1 U9077 ( .A1(n14116), .A2(n12505), .ZN(n14086) );
  NAND2_X1 U9078 ( .A1(n14129), .A2(n12503), .ZN(n14118) );
  INV_X1 U9079 ( .A(n9900), .ZN(n7093) );
  INV_X1 U9080 ( .A(n13742), .ZN(n14268) );
  AND2_X1 U9081 ( .A1(n14164), .A2(n12501), .ZN(n14154) );
  OAI21_X1 U9082 ( .B1(n12179), .B2(n12178), .A(n12177), .ZN(n14190) );
  NAND2_X1 U9083 ( .A1(n6951), .A2(n6955), .ZN(n14177) );
  NAND2_X1 U9084 ( .A1(n7244), .A2(n11888), .ZN(n12041) );
  NAND2_X1 U9085 ( .A1(n7589), .A2(n11887), .ZN(n7244) );
  NAND2_X1 U9086 ( .A1(n7550), .A2(n7551), .ZN(n11727) );
  INV_X1 U9087 ( .A(n10867), .ZN(n11340) );
  NAND2_X1 U9088 ( .A1(n14135), .A2(n11329), .ZN(n14188) );
  INV_X1 U9089 ( .A(n13640), .ZN(n11717) );
  INV_X1 U9090 ( .A(n14188), .ZN(n14169) );
  NAND2_X1 U9091 ( .A1(n14217), .A2(n7133), .ZN(n14324) );
  AND2_X1 U9092 ( .A1(n14215), .A2(n14216), .ZN(n7133) );
  INV_X1 U9093 ( .A(n15434), .ZN(n15432) );
  OR2_X1 U9094 ( .A1(n10098), .A2(P2_U3088), .ZN(n15434) );
  OR2_X1 U9095 ( .A1(n9610), .A2(n9609), .ZN(n9611) );
  INV_X1 U9096 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12124) );
  XNOR2_X1 U9097 ( .A(n10056), .B(n10055), .ZN(n12125) );
  OAI21_X1 U9098 ( .B1(n10054), .B2(P2_IR_REG_24__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10056) );
  XNOR2_X1 U9099 ( .A(n10053), .B(n10052), .ZN(n12109) );
  INV_X1 U9100 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n10052) );
  OR2_X1 U9101 ( .A1(n10051), .A2(n9573), .ZN(n9574) );
  XNOR2_X1 U9102 ( .A(n9956), .B(n9955), .ZN(n11922) );
  INV_X1 U9103 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12380) );
  INV_X1 U9104 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11419) );
  INV_X1 U9105 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n15707) );
  INV_X1 U9106 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n15748) );
  INV_X1 U9107 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n11080) );
  INV_X1 U9108 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10832) );
  INV_X1 U9109 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10700) );
  INV_X1 U9110 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10571) );
  INV_X1 U9111 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10548) );
  INV_X1 U9112 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10543) );
  INV_X1 U9113 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10493) );
  INV_X1 U9114 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10495) );
  INV_X1 U9115 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10487) );
  INV_X1 U9116 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10503) );
  NAND2_X1 U9117 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n9588) );
  XNOR2_X1 U9118 ( .A(n9618), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n7845) );
  OR2_X1 U9119 ( .A1(n9324), .A2(n10489), .ZN(n8796) );
  AND2_X1 U9120 ( .A1(n11545), .A2(n10173), .ZN(n11899) );
  OR2_X1 U9121 ( .A1(n6531), .A2(n12477), .ZN(n7762) );
  OR2_X1 U9122 ( .A1(n8775), .A2(n12475), .ZN(n7763) );
  AND3_X1 U9124 ( .A1(n9057), .A2(n9056), .A3(n9055), .ZN(n14435) );
  INV_X1 U9125 ( .A(n15262), .ZN(n11576) );
  NAND2_X1 U9126 ( .A1(n7102), .A2(n7824), .ZN(n7819) );
  CLKBUF_X1 U9127 ( .A(n12478), .Z(n12479) );
  INV_X1 U9128 ( .A(n14458), .ZN(n14497) );
  INV_X1 U9129 ( .A(n14546), .ZN(n14515) );
  NOR2_X1 U9130 ( .A1(n14458), .A2(n14909), .ZN(n14521) );
  NAND2_X1 U9131 ( .A1(n10430), .A2(n6617), .ZN(n7793) );
  NOR2_X1 U9132 ( .A1(n6640), .A2(n7809), .ZN(n7808) );
  NAND2_X1 U9133 ( .A1(n14382), .A2(n7806), .ZN(n6798) );
  NAND2_X1 U9134 ( .A1(n9260), .A2(n9259), .ZN(n14748) );
  INV_X1 U9135 ( .A(n14910), .ZN(n14558) );
  NAND2_X1 U9136 ( .A1(n10725), .A2(n10724), .ZN(n14622) );
  NAND2_X1 U9137 ( .A1(n14655), .A2(n14654), .ZN(n14668) );
  NAND2_X1 U9138 ( .A1(n6756), .A2(n10760), .ZN(n14674) );
  NAND2_X1 U9139 ( .A1(n14659), .A2(n14658), .ZN(n6756) );
  NAND2_X1 U9140 ( .A1(n10767), .A2(n10766), .ZN(n10813) );
  OR2_X1 U9141 ( .A1(n10806), .A2(n10807), .ZN(n10804) );
  NAND2_X1 U9142 ( .A1(n6755), .A2(n10795), .ZN(n10845) );
  NAND2_X1 U9143 ( .A1(n10798), .A2(n10797), .ZN(n6755) );
  NAND2_X1 U9144 ( .A1(n11022), .A2(n11021), .ZN(n11024) );
  NAND2_X1 U9145 ( .A1(n6588), .A2(n6771), .ZN(n11808) );
  NAND2_X1 U9146 ( .A1(n11952), .A2(n11951), .ZN(n12193) );
  OAI21_X1 U9147 ( .B1(n11952), .B2(n6759), .A(n6725), .ZN(n14682) );
  INV_X1 U9148 ( .A(n12192), .ZN(n6759) );
  NAND2_X1 U9149 ( .A1(n6758), .A2(n12192), .ZN(n6757) );
  NAND2_X1 U9150 ( .A1(n7496), .A2(n14717), .ZN(n7490) );
  OR2_X1 U9151 ( .A1(n10372), .A2(n7494), .ZN(n7493) );
  NAND2_X1 U9152 ( .A1(n9515), .A2(n9514), .ZN(n7192) );
  NAND2_X1 U9153 ( .A1(n14760), .A2(n9510), .ZN(n14743) );
  NAND2_X1 U9154 ( .A1(n14757), .A2(n9470), .ZN(n14742) );
  NAND2_X1 U9155 ( .A1(n14803), .A2(n9468), .ZN(n14779) );
  NAND2_X1 U9156 ( .A1(n7200), .A2(n9506), .ZN(n14772) );
  NAND2_X1 U9157 ( .A1(n14810), .A2(n9504), .ZN(n14792) );
  NAND2_X1 U9158 ( .A1(n14819), .A2(n9467), .ZN(n14805) );
  NAND2_X1 U9159 ( .A1(n14834), .A2(n14817), .ZN(n14799) );
  AND2_X1 U9160 ( .A1(n14813), .A2(n10110), .ZN(n15024) );
  NAND2_X1 U9161 ( .A1(n14852), .A2(n9465), .ZN(n14824) );
  NAND2_X1 U9162 ( .A1(n7774), .A2(n9459), .ZN(n14896) );
  NAND2_X1 U9163 ( .A1(n14917), .A2(n7778), .ZN(n7774) );
  NAND2_X1 U9164 ( .A1(n14917), .A2(n9458), .ZN(n14902) );
  INV_X1 U9165 ( .A(n9456), .ZN(n14948) );
  OAI21_X1 U9166 ( .B1(n14959), .B2(n14961), .A(n7742), .ZN(n14937) );
  OAI21_X1 U9167 ( .B1(n11516), .B2(n11878), .A(n7749), .ZN(n12052) );
  NAND2_X1 U9168 ( .A1(n11854), .A2(n9450), .ZN(n11514) );
  INV_X1 U9169 ( .A(n7513), .ZN(n7512) );
  OAI21_X1 U9170 ( .B1(n9324), .B2(n10515), .A(n7514), .ZN(n7513) );
  NAND2_X1 U9171 ( .A1(n7769), .A2(n9434), .ZN(n15271) );
  NAND2_X1 U9172 ( .A1(n11351), .A2(n9432), .ZN(n7769) );
  OR2_X1 U9173 ( .A1(n12487), .A2(n14731), .ZN(n15265) );
  INV_X1 U9174 ( .A(n15283), .ZN(n14752) );
  NAND2_X1 U9175 ( .A1(n8741), .A2(n11445), .ZN(n11347) );
  NAND2_X1 U9176 ( .A1(n10329), .A2(n10536), .ZN(n15280) );
  INV_X1 U9177 ( .A(n10332), .ZN(n10329) );
  NOR2_X1 U9178 ( .A1(n6538), .A2(n15276), .ZN(n14905) );
  INV_X1 U9179 ( .A(n9519), .ZN(n15127) );
  INV_X1 U9180 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n15152) );
  INV_X1 U9181 ( .A(n8598), .ZN(n15160) );
  INV_X1 U9182 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n12379) );
  CLKBUF_X1 U9183 ( .A(n9404), .Z(n14586) );
  INV_X1 U9184 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15628) );
  INV_X1 U9185 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12126) );
  INV_X1 U9186 ( .A(n10533), .ZN(n12128) );
  AND2_X1 U9187 ( .A1(n9397), .A2(n7842), .ZN(n9392) );
  OR2_X1 U9188 ( .A1(n9388), .A2(n9390), .ZN(n9393) );
  INV_X1 U9189 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12382) );
  INV_X1 U9190 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11543) );
  INV_X1 U9191 ( .A(n9521), .ZN(n11544) );
  INV_X1 U9192 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n15666) );
  INV_X1 U9193 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n15783) );
  INV_X1 U9194 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n15681) );
  INV_X1 U9195 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11178) );
  INV_X1 U9196 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n11060) );
  INV_X1 U9197 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10818) );
  INV_X1 U9198 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10698) );
  INV_X1 U9199 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10569) );
  INV_X1 U9200 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10550) );
  INV_X1 U9201 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10524) );
  INV_X1 U9202 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10520) );
  XNOR2_X1 U9203 ( .A(n8820), .B(P1_IR_REG_4__SCAN_IN), .ZN(n14625) );
  NAND2_X1 U9204 ( .A1(n6773), .A2(n15551), .ZN(n8819) );
  XNOR2_X1 U9205 ( .A(n6773), .B(n15551), .ZN(n14612) );
  XNOR2_X1 U9206 ( .A(n8774), .B(n8773), .ZN(n14596) );
  XNOR2_X1 U9207 ( .A(n10509), .B(n10466), .ZN(n10484) );
  NAND2_X1 U9208 ( .A1(n7052), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7051) );
  XNOR2_X1 U9209 ( .A(n10999), .B(n10784), .ZN(n10785) );
  NAND2_X1 U9210 ( .A1(n10785), .A2(n10786), .ZN(n7036) );
  XNOR2_X1 U9211 ( .A(n11315), .B(n11313), .ZN(n11312) );
  NAND2_X1 U9212 ( .A1(n7045), .A2(n11556), .ZN(n11910) );
  INV_X1 U9213 ( .A(n7043), .ZN(n11911) );
  AOI21_X1 U9214 ( .B1(n11556), .B2(n11555), .A(n6656), .ZN(n7043) );
  INV_X1 U9215 ( .A(n12155), .ZN(n7293) );
  NAND2_X1 U9216 ( .A1(n12151), .A2(n12150), .ZN(n12156) );
  AND2_X1 U9217 ( .A1(n15194), .A2(n15193), .ZN(n15196) );
  NOR2_X1 U9218 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n15219), .ZN(n7088) );
  NOR2_X1 U9219 ( .A1(n12883), .A2(n7155), .ZN(n7154) );
  NAND2_X1 U9220 ( .A1(n6672), .A2(n12890), .ZN(n7155) );
  AOI21_X1 U9221 ( .B1(n11152), .B2(n11043), .A(n11042), .ZN(n11045) );
  NAND2_X1 U9222 ( .A1(n7434), .A2(n7435), .ZN(n11092) );
  AOI21_X1 U9223 ( .B1(n12084), .B2(n12083), .A(n7445), .ZN(n12976) );
  NAND2_X1 U9224 ( .A1(n7468), .A2(n13081), .ZN(n13066) );
  OAI211_X1 U9225 ( .C1(n7984), .C2(n6921), .A(n6919), .B(n13090), .ZN(n8044)
         );
  NAND2_X1 U9226 ( .A1(n7223), .A2(n13100), .ZN(n7222) );
  OAI21_X1 U9227 ( .B1(n13120), .B2(n15519), .A(n7120), .ZN(n13123) );
  NAND2_X1 U9228 ( .A1(n15519), .A2(n7121), .ZN(n7120) );
  INV_X1 U9229 ( .A(n9426), .ZN(n9427) );
  OAI21_X1 U9230 ( .B1(n13124), .B2(n13386), .A(n9425), .ZN(n9426) );
  AOI21_X1 U9231 ( .B1(n13333), .B2(n13383), .A(n7114), .ZN(n7113) );
  NOR2_X1 U9232 ( .A1(n15549), .A2(n13336), .ZN(n7114) );
  NAND2_X1 U9233 ( .A1(n6776), .A2(n6774), .ZN(P3_U3485) );
  INV_X1 U9234 ( .A(n6775), .ZN(n6774) );
  OR2_X1 U9235 ( .A1(n13400), .A2(n15546), .ZN(n6776) );
  OAI22_X1 U9236 ( .A1(n13403), .A2(n13386), .B1(n15549), .B2(n13338), .ZN(
        n6775) );
  NAND2_X1 U9237 ( .A1(n7370), .A2(n15540), .ZN(n10407) );
  AOI21_X1 U9238 ( .B1(n13333), .B2(n13458), .A(n7116), .ZN(n7115) );
  NOR2_X1 U9239 ( .A1(n15540), .A2(n13399), .ZN(n7116) );
  XNOR2_X1 U9240 ( .A(n6983), .B(n6606), .ZN(n10105) );
  NAND2_X1 U9241 ( .A1(n7073), .A2(n7070), .ZN(n12423) );
  NAND2_X1 U9242 ( .A1(n7072), .A2(n7071), .ZN(n7070) );
  NAND2_X1 U9243 ( .A1(n12422), .A2(n14152), .ZN(n7073) );
  INV_X1 U9244 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7059) );
  NAND2_X1 U9245 ( .A1(n15460), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7124) );
  XNOR2_X1 U9246 ( .A(n7118), .B(n7815), .ZN(n14425) );
  OAI21_X1 U9247 ( .B1(n7103), .B2(n14546), .A(n14460), .ZN(P1_U3229) );
  XNOR2_X1 U9248 ( .A(n14453), .B(n7811), .ZN(n7103) );
  AOI21_X1 U9249 ( .B1(n9379), .B2(n7338), .A(n7337), .ZN(n7336) );
  INV_X1 U9250 ( .A(n9407), .ZN(n7337) );
  AOI21_X1 U9251 ( .B1(n15244), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n14716), .ZN(
        n6763) );
  NAND2_X1 U9252 ( .A1(n6765), .A2(n14731), .ZN(n6764) );
  NAND2_X1 U9253 ( .A1(n6761), .A2(n8984), .ZN(n6760) );
  NAND2_X1 U9254 ( .A1(n6888), .A2(n6886), .ZN(P1_U3555) );
  NOR2_X1 U9255 ( .A1(n6887), .A2(n6704), .ZN(n6886) );
  NOR2_X1 U9256 ( .A1(n15348), .A2(n10376), .ZN(n6887) );
  NAND2_X1 U9257 ( .A1(n7084), .A2(n7083), .ZN(n15011) );
  OR2_X1 U9258 ( .A1(n15348), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U9259 ( .A1(n15112), .A2(n15348), .ZN(n7084) );
  AOI21_X1 U9260 ( .B1(n10373), .B2(n7110), .A(n7109), .ZN(n7108) );
  NOR2_X1 U9261 ( .A1(n15342), .A2(n15109), .ZN(n7109) );
  NAND2_X1 U9262 ( .A1(n12368), .A2(n12367), .ZN(n15169) );
  INV_X1 U9263 ( .A(n13792), .ZN(n13808) );
  OR2_X1 U9264 ( .A1(n14868), .A2(n9368), .ZN(n14850) );
  AND2_X1 U9265 ( .A1(n13098), .A2(n7207), .ZN(n6551) );
  AND2_X1 U9266 ( .A1(n9267), .A2(n7323), .ZN(n6552) );
  NAND2_X2 U9267 ( .A1(n8734), .A2(n10107), .ZN(n8760) );
  NAND2_X2 U9268 ( .A1(n14308), .A2(n14152), .ZN(n9652) );
  INV_X1 U9269 ( .A(n10454), .ZN(n6938) );
  XNOR2_X2 U9270 ( .A(n8730), .B(n8729), .ZN(n8984) );
  AND2_X1 U9271 ( .A1(n8569), .A2(n6610), .ZN(n6553) );
  AND2_X1 U9272 ( .A1(n12434), .A2(n12433), .ZN(n6554) );
  XOR2_X1 U9273 ( .A(n12886), .B(n13181), .Z(n6555) );
  OR2_X1 U9274 ( .A1(n14827), .A2(n7788), .ZN(n6556) );
  OR2_X1 U9275 ( .A1(n12257), .A2(n7728), .ZN(n6557) );
  AND2_X1 U9276 ( .A1(n7501), .A2(n7500), .ZN(n6558) );
  NAND2_X1 U9277 ( .A1(n6662), .A2(n12505), .ZN(n6559) );
  INV_X1 U9278 ( .A(n10177), .ZN(n15336) );
  INV_X1 U9279 ( .A(n13872), .ZN(n12539) );
  XNOR2_X1 U9280 ( .A(n14203), .B(n13799), .ZN(n13872) );
  AND4_X1 U9281 ( .A1(n8716), .A2(n8705), .A3(n8706), .A4(n8715), .ZN(n8724)
         );
  AND2_X1 U9282 ( .A1(n7726), .A2(n6722), .ZN(n6560) );
  AND4_X1 U9283 ( .A1(n13841), .A2(n13809), .A3(n13822), .A4(n13824), .ZN(
        n6561) );
  NOR2_X1 U9284 ( .A1(n12459), .A2(n13129), .ZN(n6562) );
  INV_X1 U9285 ( .A(n11483), .ZN(n6872) );
  AND2_X1 U9286 ( .A1(n13335), .A2(n6716), .ZN(n6563) );
  AND3_X1 U9287 ( .A1(n9373), .A2(n10362), .A3(n9515), .ZN(n6564) );
  NAND2_X1 U9288 ( .A1(n8264), .A2(n6619), .ZN(n13319) );
  OR3_X1 U9289 ( .A1(n14183), .A2(n7577), .A3(n13724), .ZN(n6565) );
  OR3_X1 U9290 ( .A1(n8285), .A2(n7026), .A3(P3_REG3_REG_16__SCAN_IN), .ZN(
        n6566) );
  INV_X1 U9291 ( .A(n13784), .ZN(n7518) );
  AND2_X1 U9292 ( .A1(n6681), .A2(n11215), .ZN(n6567) );
  AND3_X1 U9293 ( .A1(n12591), .A2(n12613), .A3(n12751), .ZN(n6568) );
  AND2_X1 U9294 ( .A1(n9457), .A2(n9455), .ZN(n6569) );
  AND2_X1 U9295 ( .A1(n6557), .A2(n6722), .ZN(n6570) );
  INV_X1 U9296 ( .A(n9996), .ZN(n7624) );
  AND2_X1 U9297 ( .A1(n7168), .A2(n6695), .ZN(n6571) );
  AND2_X1 U9298 ( .A1(n6926), .A2(n7945), .ZN(n6572) );
  AND2_X1 U9299 ( .A1(n7584), .A2(n7588), .ZN(n6573) );
  NAND2_X1 U9300 ( .A1(n14129), .A2(n7599), .ZN(n14116) );
  AND2_X1 U9301 ( .A1(n8675), .A2(SI_22_), .ZN(n6574) );
  AND2_X1 U9302 ( .A1(n9251), .A2(n9249), .ZN(n6575) );
  NAND2_X1 U9303 ( .A1(n8913), .A2(n8912), .ZN(n11991) );
  INV_X1 U9304 ( .A(n11991), .ZN(n12205) );
  NAND2_X1 U9305 ( .A1(n13779), .A2(n7524), .ZN(n6576) );
  AND2_X1 U9306 ( .A1(n8666), .A2(n11077), .ZN(n6577) );
  NAND2_X1 U9307 ( .A1(n6666), .A2(n11215), .ZN(n6578) );
  AND2_X1 U9308 ( .A1(n9496), .A2(n9356), .ZN(n14952) );
  AND2_X1 U9309 ( .A1(n9776), .A2(n9775), .ZN(n6579) );
  AND2_X1 U9310 ( .A1(n13050), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6580) );
  AND2_X1 U9311 ( .A1(n7611), .A2(n10025), .ZN(n6581) );
  OAI211_X1 U9312 ( .C1(n6555), .C2(n7158), .A(n7163), .B(n7157), .ZN(n7156)
         );
  AND2_X1 U9313 ( .A1(n11120), .A2(n9700), .ZN(n6582) );
  INV_X1 U9314 ( .A(n15147), .ZN(n7110) );
  NOR2_X1 U9315 ( .A1(n7976), .A2(n13387), .ZN(n6583) );
  NAND2_X1 U9316 ( .A1(n15549), .A2(n13374), .ZN(n13391) );
  NAND2_X1 U9317 ( .A1(n8692), .A2(SI_26_), .ZN(n6584) );
  INV_X1 U9318 ( .A(n7939), .ZN(n7209) );
  NAND2_X1 U9319 ( .A1(n8389), .A2(n8388), .ZN(n13411) );
  AND2_X1 U9320 ( .A1(n15840), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6585) );
  INV_X1 U9321 ( .A(n9668), .ZN(n7247) );
  INV_X1 U9322 ( .A(n13097), .ZN(n6927) );
  AND2_X1 U9323 ( .A1(n6927), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n6586) );
  OAI21_X1 U9324 ( .B1(n11101), .B2(n6909), .A(n6911), .ZN(n6910) );
  INV_X1 U9325 ( .A(n12543), .ZN(n14071) );
  OR2_X1 U9326 ( .A1(n7916), .A2(n12028), .ZN(n6587) );
  NAND2_X1 U9327 ( .A1(n11807), .A2(n6768), .ZN(n6588) );
  NAND2_X1 U9328 ( .A1(n8235), .A2(n7664), .ZN(n7663) );
  NAND2_X1 U9329 ( .A1(n8144), .A2(n7674), .ZN(n7673) );
  NAND2_X1 U9330 ( .A1(n9958), .A2(n9957), .ZN(n14049) );
  NAND2_X1 U9331 ( .A1(n7359), .A2(n8230), .ZN(n13290) );
  AND2_X1 U9332 ( .A1(n9638), .A2(n9637), .ZN(n6589) );
  AND2_X1 U9333 ( .A1(n10445), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n6590) );
  INV_X1 U9334 ( .A(n14454), .ZN(n7811) );
  NAND2_X1 U9335 ( .A1(n7923), .A2(n12998), .ZN(n7925) );
  INV_X1 U9336 ( .A(n14420), .ZN(n7815) );
  INV_X1 U9337 ( .A(n14820), .ZN(n7785) );
  NAND2_X1 U9338 ( .A1(n6882), .A2(n12715), .ZN(n13214) );
  NAND2_X1 U9339 ( .A1(n14919), .A2(n14918), .ZN(n14917) );
  NAND2_X1 U9340 ( .A1(n8456), .A2(n8455), .ZN(n8574) );
  NAND2_X1 U9341 ( .A1(n13432), .A2(n13243), .ZN(n6591) );
  NAND2_X1 U9342 ( .A1(n14981), .A2(n9454), .ZN(n14949) );
  NOR2_X1 U9343 ( .A1(n12992), .A2(n15767), .ZN(n12991) );
  INV_X1 U9344 ( .A(n12053), .ZN(n7748) );
  OR2_X1 U9345 ( .A1(n8579), .A2(n10391), .ZN(n12748) );
  OR2_X1 U9346 ( .A1(n14220), .A2(n13999), .ZN(n6592) );
  AND2_X1 U9347 ( .A1(n9495), .A2(n9102), .ZN(n14967) );
  XNOR2_X1 U9348 ( .A(n14302), .B(n13899), .ZN(n13858) );
  AND2_X1 U9349 ( .A1(n10263), .A2(n10262), .ZN(n6593) );
  AND2_X1 U9350 ( .A1(n14034), .A2(n13597), .ZN(n6594) );
  AND2_X1 U9351 ( .A1(n7990), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6595) );
  INV_X1 U9352 ( .A(n15055), .ZN(n7090) );
  NAND4_X1 U9353 ( .A1(n8765), .A2(n8764), .A3(n8763), .A4(n8762), .ZN(n9433)
         );
  INV_X1 U9354 ( .A(n12785), .ZN(n7717) );
  AND2_X1 U9355 ( .A1(n10698), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U9356 ( .A1(n8678), .A2(n6960), .ZN(n6597) );
  XNOR2_X1 U9357 ( .A(n11991), .B(n11522), .ZN(n11855) );
  NAND2_X1 U9358 ( .A1(n8441), .A2(n8440), .ZN(n13339) );
  AND2_X1 U9359 ( .A1(n15336), .A2(n14564), .ZN(n6598) );
  INV_X1 U9360 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10513) );
  OR2_X1 U9361 ( .A1(n7977), .A2(n12998), .ZN(n6599) );
  NAND2_X1 U9362 ( .A1(n8749), .A2(n8773), .ZN(n6600) );
  NOR2_X1 U9363 ( .A1(n11373), .A2(n6590), .ZN(n6601) );
  AND2_X1 U9364 ( .A1(n6975), .A2(n12388), .ZN(n9674) );
  INV_X1 U9365 ( .A(n9674), .ZN(n9707) );
  NAND2_X1 U9366 ( .A1(n12561), .A2(n12560), .ZN(n12587) );
  NOR2_X1 U9367 ( .A1(n13528), .A2(n7608), .ZN(n6602) );
  BUF_X1 U9368 ( .A(n8870), .Z(n9286) );
  INV_X1 U9369 ( .A(n10362), .ZN(n10367) );
  XNOR2_X1 U9370 ( .A(n10373), .B(n14748), .ZN(n10362) );
  OAI21_X1 U9371 ( .B1(n13214), .B2(n7401), .A(n7398), .ZN(n13184) );
  AND2_X1 U9372 ( .A1(n7505), .A2(n15336), .ZN(n6603) );
  INV_X1 U9373 ( .A(n14817), .ZN(n7511) );
  NAND2_X1 U9374 ( .A1(n10027), .A2(n10026), .ZN(n14211) );
  AND2_X1 U9375 ( .A1(n9059), .A2(n9058), .ZN(n6604) );
  AND2_X1 U9376 ( .A1(n7435), .A2(n7433), .ZN(n6605) );
  XOR2_X1 U9377 ( .A(n13953), .B(n10050), .Z(n6606) );
  OR2_X1 U9378 ( .A1(n7815), .A2(n14454), .ZN(n6607) );
  NAND2_X1 U9379 ( .A1(n8714), .A2(n8713), .ZN(n14738) );
  NAND2_X1 U9380 ( .A1(n14921), .A2(n9497), .ZN(n14842) );
  NAND2_X1 U9381 ( .A1(n15170), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6608) );
  AND2_X1 U9382 ( .A1(n9567), .A2(n9632), .ZN(n9576) );
  NAND2_X1 U9383 ( .A1(n8821), .A2(n7512), .ZN(n14464) );
  INV_X1 U9384 ( .A(n14464), .ZN(n15322) );
  OR2_X1 U9385 ( .A1(n8508), .A2(n10451), .ZN(n6609) );
  NAND2_X1 U9386 ( .A1(n9288), .A2(n9287), .ZN(n14717) );
  INV_X1 U9387 ( .A(n14717), .ZN(n7494) );
  OR2_X1 U9388 ( .A1(n13417), .A2(n12443), .ZN(n6610) );
  XNOR2_X1 U9389 ( .A(n7859), .B(P3_IR_REG_24__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U9390 ( .A1(n9150), .A2(n9149), .ZN(n14858) );
  AOI21_X1 U9391 ( .B1(n13793), .B2(n13953), .A(n12515), .ZN(n13955) );
  AND2_X1 U9392 ( .A1(n9047), .A2(n8662), .ZN(n6611) );
  NAND2_X1 U9393 ( .A1(n6738), .A2(n7740), .ZN(n14936) );
  AND4_X1 U9394 ( .A1(n13178), .A2(n12609), .A3(n13196), .A4(n13205), .ZN(
        n6612) );
  NAND2_X1 U9395 ( .A1(n7018), .A2(n7015), .ZN(n14826) );
  AND2_X1 U9396 ( .A1(n10382), .A2(n13308), .ZN(n6613) );
  NAND2_X1 U9397 ( .A1(n14936), .A2(n7201), .ZN(n14921) );
  AND2_X1 U9398 ( .A1(n14292), .A2(n13720), .ZN(n6614) );
  NOR2_X1 U9399 ( .A1(n14918), .A2(n7202), .ZN(n7201) );
  INV_X1 U9400 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n15718) );
  NAND2_X1 U9401 ( .A1(n13228), .A2(n12714), .ZN(n13254) );
  INV_X1 U9402 ( .A(n13254), .ZN(n7348) );
  XNOR2_X1 U9403 ( .A(n14211), .B(n13891), .ZN(n13959) );
  AND2_X1 U9404 ( .A1(n14952), .A2(n14901), .ZN(n6615) );
  OR2_X1 U9405 ( .A1(n14071), .A2(n7585), .ZN(n6616) );
  AND2_X1 U9406 ( .A1(n10155), .A2(n10149), .ZN(n6617) );
  AND2_X1 U9407 ( .A1(n6649), .A2(n15179), .ZN(n6618) );
  AND3_X1 U9408 ( .A1(n8266), .A2(n8265), .A3(n6859), .ZN(n6619) );
  NAND2_X1 U9409 ( .A1(n14775), .A2(n9508), .ZN(n14759) );
  AND2_X1 U9410 ( .A1(n10559), .A2(n7053), .ZN(n6620) );
  NAND2_X1 U9411 ( .A1(n7964), .A2(n7853), .ZN(n7894) );
  INV_X1 U9412 ( .A(n8202), .ZN(n8204) );
  AND2_X1 U9413 ( .A1(n12442), .A2(n13233), .ZN(n6621) );
  INV_X1 U9414 ( .A(n15048), .ZN(n14894) );
  OR2_X1 U9415 ( .A1(n7823), .A2(n6593), .ZN(n6622) );
  AND2_X1 U9416 ( .A1(n7819), .A2(n7823), .ZN(n6623) );
  NAND2_X1 U9417 ( .A1(n7741), .A2(n14967), .ZN(n14958) );
  OR2_X1 U9418 ( .A1(n10930), .A2(n10929), .ZN(n6624) );
  AND2_X1 U9419 ( .A1(n7831), .A2(n9486), .ZN(n6625) );
  INV_X1 U9420 ( .A(n11783), .ZN(n6831) );
  AND2_X1 U9421 ( .A1(n14738), .A2(n14550), .ZN(n6626) );
  INV_X1 U9422 ( .A(n8173), .ZN(n7670) );
  INV_X1 U9423 ( .A(n8962), .ZN(n6806) );
  INV_X1 U9424 ( .A(n9470), .ZN(n7791) );
  AND2_X1 U9425 ( .A1(n12821), .A2(n7733), .ZN(n6627) );
  NOR2_X1 U9426 ( .A1(n7524), .A2(n13779), .ZN(n7522) );
  AND2_X1 U9427 ( .A1(n9458), .A2(n9366), .ZN(n14918) );
  AND2_X1 U9428 ( .A1(n7697), .A2(n8654), .ZN(n6628) );
  AND2_X1 U9429 ( .A1(n7460), .A2(n7979), .ZN(n6629) );
  NAND2_X1 U9430 ( .A1(n14292), .A2(n13896), .ZN(n6630) );
  AND2_X1 U9431 ( .A1(n8111), .A2(n8107), .ZN(n6631) );
  AND2_X1 U9432 ( .A1(n14793), .A2(n9467), .ZN(n6632) );
  NOR2_X1 U9433 ( .A1(n14426), .A2(n7798), .ZN(n6633) );
  NOR2_X1 U9434 ( .A1(n12848), .A2(n7723), .ZN(n6634) );
  OR2_X1 U9435 ( .A1(n8865), .A2(n8863), .ZN(n6635) );
  AND2_X1 U9436 ( .A1(n13871), .A2(n12533), .ZN(n6636) );
  INV_X1 U9437 ( .A(n14297), .ZN(n13716) );
  AND2_X1 U9438 ( .A1(n7226), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n6637) );
  INV_X1 U9439 ( .A(n9700), .ZN(n6986) );
  NAND2_X1 U9440 ( .A1(n7525), .A2(n7516), .ZN(n6638) );
  INV_X1 U9441 ( .A(n13861), .ZN(n6954) );
  NAND2_X1 U9442 ( .A1(n8579), .A2(n10391), .ZN(n12747) );
  AND2_X1 U9443 ( .A1(n12524), .A2(n13893), .ZN(n6639) );
  NAND2_X1 U9444 ( .A1(n7813), .A2(n10294), .ZN(n6640) );
  NOR2_X1 U9445 ( .A1(n14024), .A2(n14049), .ZN(n6641) );
  NOR2_X1 U9446 ( .A1(n13417), .A2(n13222), .ZN(n6642) );
  NOR2_X1 U9447 ( .A1(n13978), .A2(n13968), .ZN(n6643) );
  INV_X1 U9448 ( .A(n6794), .ZN(n8891) );
  OAI21_X1 U9449 ( .B1(n6795), .B2(SI_8_), .A(n8643), .ZN(n6794) );
  XOR2_X1 U9450 ( .A(n12745), .B(n12462), .Z(n6644) );
  NAND2_X1 U9451 ( .A1(n9299), .A2(n9298), .ZN(n14725) );
  INV_X1 U9452 ( .A(n14725), .ZN(n15107) );
  AND2_X1 U9453 ( .A1(n7054), .A2(n10559), .ZN(n6645) );
  AND2_X1 U9454 ( .A1(n12590), .A2(n7833), .ZN(n6646) );
  OR2_X1 U9455 ( .A1(n14246), .A2(n14081), .ZN(n6647) );
  AND4_X1 U9456 ( .A1(n8749), .A2(n8702), .A3(n8773), .A4(n8707), .ZN(n6648)
         );
  INV_X1 U9457 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10545) );
  INV_X1 U9458 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n15651) );
  INV_X1 U9459 ( .A(n7614), .ZN(n7613) );
  OR2_X1 U9460 ( .A1(n13616), .A2(n7615), .ZN(n7614) );
  AND2_X1 U9461 ( .A1(n15172), .A2(n15171), .ZN(n6649) );
  AND2_X1 U9462 ( .A1(n12785), .A2(n6562), .ZN(n6650) );
  AND2_X1 U9463 ( .A1(n6561), .A2(n6638), .ZN(n6651) );
  NAND2_X1 U9464 ( .A1(n10347), .A2(n10346), .ZN(n6652) );
  NAND2_X1 U9465 ( .A1(n12542), .A2(n6966), .ZN(n6653) );
  INV_X1 U9466 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7960) );
  OR2_X1 U9467 ( .A1(n14098), .A2(n13607), .ZN(n6654) );
  NOR2_X1 U9468 ( .A1(n14292), .A2(n13896), .ZN(n6655) );
  NAND2_X1 U9469 ( .A1(n11913), .A2(n11564), .ZN(n6656) );
  OR2_X1 U9470 ( .A1(n13754), .A2(n13752), .ZN(n6657) );
  INV_X1 U9471 ( .A(n7756), .ZN(n7755) );
  NAND2_X1 U9472 ( .A1(n9491), .A2(n9490), .ZN(n7756) );
  NAND3_X1 U9473 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .A3(P2_IR_REG_31__SCAN_IN), .ZN(n6658) );
  AND2_X1 U9474 ( .A1(n12793), .A2(n12792), .ZN(n6659) );
  INV_X1 U9475 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10526) );
  OR2_X1 U9476 ( .A1(n7562), .A2(n6594), .ZN(n6660) );
  AND2_X1 U9477 ( .A1(n7423), .A2(n8043), .ZN(n6661) );
  INV_X1 U9478 ( .A(n13953), .ZN(n14207) );
  OR2_X1 U9479 ( .A1(n14257), .A2(n14109), .ZN(n6662) );
  INV_X1 U9480 ( .A(n7597), .ZN(n7596) );
  NAND2_X1 U9481 ( .A1(n13970), .A2(n6592), .ZN(n7597) );
  AND2_X1 U9482 ( .A1(n8962), .A2(n6807), .ZN(n6663) );
  AND2_X1 U9483 ( .A1(n14948), .A2(n14435), .ZN(n6664) );
  AND2_X1 U9484 ( .A1(n8667), .A2(SI_17_), .ZN(n6665) );
  NOR2_X1 U9485 ( .A1(n7896), .A2(n10451), .ZN(n7898) );
  NAND2_X1 U9486 ( .A1(n8004), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6666) );
  AND2_X1 U9487 ( .A1(n12701), .A2(n12705), .ZN(n13281) );
  INV_X1 U9488 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10491) );
  NAND2_X1 U9489 ( .A1(n8205), .A2(n8232), .ZN(n6667) );
  NOR2_X1 U9490 ( .A1(n7396), .A2(n12675), .ZN(n7395) );
  AND2_X1 U9491 ( .A1(n8660), .A2(n9015), .ZN(n6668) );
  NAND2_X1 U9492 ( .A1(n11585), .A2(n7832), .ZN(n6669) );
  NAND2_X1 U9493 ( .A1(n6668), .A2(n8658), .ZN(n6670) );
  AND2_X1 U9494 ( .A1(n9329), .A2(n9328), .ZN(n6671) );
  INV_X1 U9495 ( .A(n7620), .ZN(n7619) );
  NOR2_X1 U9496 ( .A1(n6555), .A2(n7160), .ZN(n6672) );
  INV_X1 U9497 ( .A(n13864), .ZN(n14153) );
  INV_X1 U9498 ( .A(n7496), .ZN(n7495) );
  NAND2_X1 U9499 ( .A1(n15107), .A2(n7497), .ZN(n7496) );
  OR2_X1 U9500 ( .A1(n13901), .A2(n13687), .ZN(n6673) );
  INV_X1 U9501 ( .A(n12343), .ZN(n7139) );
  INV_X1 U9502 ( .A(n8922), .ZN(n7329) );
  AND2_X1 U9503 ( .A1(n6608), .A2(n15179), .ZN(n6674) );
  AND2_X1 U9504 ( .A1(n11619), .A2(n11783), .ZN(n6675) );
  OR2_X1 U9505 ( .A1(n12663), .A2(n12662), .ZN(n6676) );
  INV_X1 U9506 ( .A(n12745), .ZN(n7315) );
  OR2_X1 U9507 ( .A1(n8667), .A2(SI_17_), .ZN(n6677) );
  OR2_X1 U9508 ( .A1(n7326), .A2(n8603), .ZN(n6678) );
  AND2_X1 U9509 ( .A1(n7418), .A2(n12748), .ZN(n6679) );
  AND2_X1 U9510 ( .A1(n6984), .A2(n6581), .ZN(n6680) );
  NAND2_X1 U9511 ( .A1(n8004), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6681) );
  AND2_X1 U9512 ( .A1(n7508), .A2(n7507), .ZN(n6682) );
  AND2_X1 U9513 ( .A1(n7506), .A2(n15036), .ZN(n6683) );
  OR2_X1 U9514 ( .A1(n7520), .A2(n7517), .ZN(n6684) );
  AND2_X1 U9515 ( .A1(n7674), .A2(n8173), .ZN(n6685) );
  OR2_X1 U9516 ( .A1(n14982), .A2(n6891), .ZN(n6686) );
  NOR2_X1 U9517 ( .A1(n13724), .A2(n14274), .ZN(n6687) );
  AND2_X1 U9518 ( .A1(n11622), .A2(n7556), .ZN(n6688) );
  INV_X1 U9519 ( .A(n13178), .ZN(n13185) );
  AND2_X1 U9520 ( .A1(n12617), .A2(n12621), .ZN(n13178) );
  AND2_X1 U9521 ( .A1(n13411), .A2(n13180), .ZN(n12608) );
  OR2_X1 U9522 ( .A1(n13769), .A2(n13767), .ZN(n6689) );
  AND2_X1 U9523 ( .A1(n8520), .A2(n7729), .ZN(n6690) );
  AND2_X1 U9524 ( .A1(n7353), .A2(n8118), .ZN(n6691) );
  OR2_X1 U9525 ( .A1(n13761), .A2(n13763), .ZN(n6692) );
  INV_X1 U9526 ( .A(n13995), .ZN(n6972) );
  INV_X1 U9527 ( .A(n13281), .ZN(n7409) );
  AND2_X1 U9528 ( .A1(n7857), .A2(n7164), .ZN(n6693) );
  AND2_X1 U9529 ( .A1(n7750), .A2(n9493), .ZN(n7749) );
  NAND2_X1 U9530 ( .A1(n10037), .A2(n10036), .ZN(n6694) );
  INV_X1 U9531 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8046) );
  NAND2_X1 U9532 ( .A1(n8656), .A2(n10568), .ZN(n6695) );
  INV_X1 U9533 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6813) );
  INV_X1 U9534 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9390) );
  INV_X1 U9535 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10518) );
  INV_X1 U9536 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7739) );
  INV_X1 U9537 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9584) );
  INV_X1 U9538 ( .A(n8665), .ZN(n7696) );
  INV_X1 U9539 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10541) );
  INV_X1 U9540 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10489) );
  INV_X1 U9541 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7164) );
  INV_X1 U9542 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n7477) );
  INV_X1 U9543 ( .A(n14957), .ZN(n7500) );
  INV_X1 U9544 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8299) );
  OAI21_X1 U9545 ( .B1(n11616), .B2(n11615), .A(n11614), .ZN(n11723) );
  INV_X1 U9546 ( .A(n12960), .ZN(n7163) );
  INV_X1 U9547 ( .A(n14765), .ZN(n7507) );
  AND2_X1 U9548 ( .A1(n8522), .A2(n8521), .ZN(n13473) );
  NAND2_X1 U9549 ( .A1(n6973), .A2(n11052), .ZN(n11621) );
  NAND2_X1 U9550 ( .A1(n15540), .A2(n13374), .ZN(n13470) );
  INV_X1 U9551 ( .A(n13470), .ZN(n13458) );
  NAND2_X1 U9552 ( .A1(n7504), .A2(n7505), .ZN(n11489) );
  NAND2_X1 U9553 ( .A1(n14164), .A2(n7097), .ZN(n14155) );
  AND2_X1 U9554 ( .A1(n8099), .A2(n11645), .ZN(n6696) );
  OR2_X1 U9555 ( .A1(n12892), .A2(n12893), .ZN(n12799) );
  NAND2_X1 U9556 ( .A1(n9663), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6697) );
  INV_X1 U9557 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n6899) );
  OR2_X1 U9558 ( .A1(n8016), .A2(n12982), .ZN(n6698) );
  NAND2_X1 U9559 ( .A1(n7757), .A2(n7755), .ZN(n11495) );
  NAND2_X1 U9560 ( .A1(n11393), .A2(n9487), .ZN(n11938) );
  NAND2_X1 U9561 ( .A1(n15273), .A2(n9485), .ZN(n11302) );
  OAI21_X1 U9562 ( .B1(n12799), .B2(n6557), .A(n7726), .ZN(n12342) );
  NAND2_X1 U9563 ( .A1(n9793), .A2(n9792), .ZN(n12158) );
  AND2_X1 U9564 ( .A1(n6914), .A2(n10420), .ZN(n6699) );
  NAND2_X1 U9565 ( .A1(n9970), .A2(n9969), .ZN(n14230) );
  INV_X1 U9566 ( .A(n14230), .ZN(n7588) );
  AND2_X1 U9567 ( .A1(n10430), .A2(n10149), .ZN(n6700) );
  NAND2_X1 U9568 ( .A1(n11874), .A2(n11873), .ZN(n11872) );
  NAND2_X1 U9569 ( .A1(n9483), .A2(n9484), .ZN(n15273) );
  AND2_X1 U9570 ( .A1(n8397), .A2(n8396), .ZN(n13180) );
  INV_X1 U9571 ( .A(n13180), .ZN(n13208) );
  INV_X1 U9572 ( .A(n7006), .ZN(n14183) );
  NOR2_X1 U9573 ( .A1(n12045), .A2(n14297), .ZN(n7006) );
  NAND2_X1 U9574 ( .A1(n7757), .A2(n9490), .ZN(n11496) );
  AND2_X1 U9575 ( .A1(n8280), .A2(n8021), .ZN(n6701) );
  AND2_X1 U9576 ( .A1(n7444), .A2(n7443), .ZN(n6702) );
  OR2_X1 U9577 ( .A1(n12094), .A2(n12270), .ZN(n6703) );
  NAND2_X1 U9578 ( .A1(n14153), .A2(n12501), .ZN(n7251) );
  INV_X1 U9579 ( .A(n7251), .ZN(n7097) );
  NOR2_X1 U9580 ( .A1(n15110), .A2(n15086), .ZN(n6704) );
  INV_X1 U9581 ( .A(n12913), .ZN(n13198) );
  AND2_X1 U9582 ( .A1(n8419), .A2(n8418), .ZN(n12913) );
  INV_X1 U9583 ( .A(n7503), .ZN(n11858) );
  INV_X1 U9584 ( .A(n7162), .ZN(n7161) );
  NOR2_X1 U9585 ( .A1(n13198), .A2(n12884), .ZN(n7162) );
  INV_X1 U9586 ( .A(n8277), .ZN(n7660) );
  AND3_X1 U9587 ( .A1(n6687), .A2(n7006), .A3(n7005), .ZN(n14137) );
  AND2_X1 U9588 ( .A1(n8017), .A2(n10567), .ZN(n6705) );
  AND2_X1 U9589 ( .A1(n7639), .A2(n8323), .ZN(n6706) );
  INV_X1 U9590 ( .A(n10373), .ZN(n15110) );
  NAND2_X1 U9591 ( .A1(n9265), .A2(n9264), .ZN(n10373) );
  NOR2_X1 U9592 ( .A1(n8309), .A2(n8030), .ZN(n6707) );
  AND2_X1 U9593 ( .A1(n9278), .A2(n15777), .ZN(n6708) );
  AND2_X1 U9594 ( .A1(n12436), .A2(n12857), .ZN(n6709) );
  INV_X1 U9595 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10515) );
  INV_X1 U9596 ( .A(n7644), .ZN(n7643) );
  NAND2_X1 U9597 ( .A1(n8406), .A2(n8403), .ZN(n7644) );
  NOR2_X1 U9598 ( .A1(n12094), .A2(n12306), .ZN(n6710) );
  INV_X1 U9599 ( .A(n8510), .ZN(n8428) );
  AND2_X1 U9600 ( .A1(n7664), .A2(n8277), .ZN(n6711) );
  AND2_X1 U9601 ( .A1(n12115), .A2(n12674), .ZN(n6712) );
  INV_X1 U9602 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7053) );
  AND2_X1 U9603 ( .A1(n6555), .A2(n7161), .ZN(n6713) );
  NAND2_X1 U9604 ( .A1(n14246), .A2(n13600), .ZN(n7565) );
  INV_X1 U9605 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U9606 ( .A1(n13079), .A2(n8034), .ZN(n6714) );
  AND2_X1 U9607 ( .A1(n11556), .A2(n7285), .ZN(SUB_1596_U54) );
  NOR2_X1 U9608 ( .A1(n15514), .A2(n12766), .ZN(n6716) );
  AND2_X1 U9609 ( .A1(n8179), .A2(n8178), .ZN(n12219) );
  INV_X1 U9610 ( .A(n12219), .ZN(n7141) );
  INV_X1 U9611 ( .A(n14292), .ZN(n7578) );
  NAND2_X1 U9612 ( .A1(n9684), .A2(n9683), .ZN(n13670) );
  INV_X1 U9613 ( .A(n13670), .ZN(n7575) );
  NAND2_X1 U9614 ( .A1(n6907), .A2(n6904), .ZN(n11217) );
  INV_X2 U9615 ( .A(n15546), .ZN(n15549) );
  CLKBUF_X1 U9616 ( .A(n10118), .Z(n12392) );
  INV_X1 U9617 ( .A(n10118), .ZN(n8742) );
  XOR2_X1 U9618 ( .A(n8296), .B(P3_REG1_REG_16__SCAN_IN), .Z(n6717) );
  INV_X1 U9619 ( .A(n14314), .ZN(n6833) );
  XOR2_X1 U9620 ( .A(n10567), .B(n13321), .Z(n6718) );
  AND2_X1 U9621 ( .A1(n6732), .A2(n8536), .ZN(n15508) );
  INV_X1 U9622 ( .A(n15508), .ZN(n13308) );
  NAND2_X1 U9623 ( .A1(n9481), .A2(n9479), .ZN(n11444) );
  INV_X1 U9624 ( .A(n15060), .ZN(n7498) );
  INV_X1 U9625 ( .A(n14319), .ZN(n15458) );
  AND2_X1 U9626 ( .A1(n13803), .A2(n10688), .ZN(n14162) );
  INV_X1 U9627 ( .A(n14162), .ZN(n14180) );
  INV_X1 U9628 ( .A(n8280), .ZN(n13035) );
  AND2_X1 U9629 ( .A1(n7936), .A2(n7940), .ZN(n8280) );
  AND2_X1 U9630 ( .A1(n11940), .A2(n15310), .ZN(n15100) );
  OR2_X1 U9631 ( .A1(n7971), .A2(n6908), .ZN(n6719) );
  AND2_X1 U9632 ( .A1(n12088), .A2(n7471), .ZN(n6720) );
  NAND2_X1 U9633 ( .A1(n7484), .A2(n7485), .ZN(n6721) );
  NAND2_X1 U9634 ( .A1(n12258), .A2(n12346), .ZN(n6722) );
  AND2_X1 U9635 ( .A1(n6605), .A2(n7434), .ZN(n6723) );
  AND2_X1 U9636 ( .A1(n15158), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6724) );
  AND2_X1 U9637 ( .A1(n12190), .A2(n6757), .ZN(n6725) );
  AND2_X1 U9638 ( .A1(n7457), .A2(n7456), .ZN(n6726) );
  NAND2_X1 U9639 ( .A1(n6987), .A2(n6988), .ZN(n6727) );
  AND2_X1 U9640 ( .A1(n11340), .A2(n10869), .ZN(n6728) );
  INV_X1 U9641 ( .A(n6901), .ZN(n7972) );
  OR2_X1 U9642 ( .A1(n11368), .A2(n6902), .ZN(n6901) );
  AND2_X1 U9643 ( .A1(n7939), .A2(n8309), .ZN(n6729) );
  INV_X1 U9644 ( .A(SI_22_), .ZN(n6960) );
  AND2_X1 U9645 ( .A1(n7037), .A2(n7036), .ZN(SUB_1596_U56) );
  XNOR2_X1 U9646 ( .A(n7906), .B(P3_IR_REG_5__SCAN_IN), .ZN(n11215) );
  XNOR2_X1 U9647 ( .A(n7884), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11838) );
  INV_X1 U9648 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U9649 ( .A1(n6837), .A2(n8893), .ZN(n6896) );
  XOR2_X1 U9650 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .Z(n6731) );
  OR2_X1 U9651 ( .A1(n12627), .A2(n11385), .ZN(n6732) );
  NAND2_X1 U9652 ( .A1(n6870), .A2(n6871), .ZN(n15505) );
  INV_X1 U9653 ( .A(n15505), .ZN(n6869) );
  NAND2_X1 U9654 ( .A1(n7970), .A2(n7969), .ZN(n6733) );
  INV_X1 U9655 ( .A(n12768), .ZN(n7390) );
  INV_X1 U9656 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n6903) );
  INV_X1 U9657 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n7465) );
  INV_X1 U9658 ( .A(n12028), .ZN(n7472) );
  NAND2_X1 U9659 ( .A1(n7973), .A2(n12028), .ZN(n12088) );
  INV_X1 U9660 ( .A(n12982), .ZN(n6912) );
  NAND2_X1 U9661 ( .A1(n7920), .A2(n12982), .ZN(n7921) );
  NAND2_X1 U9662 ( .A1(n7975), .A2(n12982), .ZN(n10420) );
  OAI21_X2 U9663 ( .B1(n7018), .B2(n6736), .A(n6734), .ZN(n14825) );
  XNOR2_X1 U9664 ( .A(n7761), .B(n15718), .ZN(n9403) );
  XNOR2_X1 U9665 ( .A(n8712), .B(n8711), .ZN(n9404) );
  NAND3_X1 U9666 ( .A1(n11516), .A2(n7749), .A3(n14978), .ZN(n6740) );
  NAND3_X1 U9667 ( .A1(n6742), .A2(n13703), .A3(n6741), .ZN(n13701) );
  OAI21_X1 U9668 ( .B1(n6746), .B2(n6745), .A(n7531), .ZN(n13757) );
  NAND2_X2 U9669 ( .A1(n9725), .A2(n6749), .ZN(n13901) );
  AOI21_X1 U9670 ( .B1(n13765), .B2(n13766), .A(n6752), .ZN(n6751) );
  OAI21_X1 U9671 ( .B1(n13765), .B2(n13766), .A(n6689), .ZN(n6753) );
  AOI21_X1 U9672 ( .B1(n7840), .B2(n10059), .A(n9600), .ZN(n6754) );
  NAND2_X1 U9673 ( .A1(n10845), .A2(n10844), .ZN(n10842) );
  NAND2_X1 U9674 ( .A1(n14674), .A2(n14673), .ZN(n10763) );
  NAND3_X1 U9675 ( .A1(n6764), .A2(n6763), .A3(n6760), .ZN(P1_U3262) );
  NAND3_X1 U9676 ( .A1(n6588), .A2(n6771), .A3(n6770), .ZN(n11950) );
  NAND2_X1 U9677 ( .A1(n11807), .A2(n11806), .ZN(n6772) );
  NOR2_X1 U9678 ( .A1(n6769), .A2(n11812), .ZN(n6768) );
  INV_X1 U9679 ( .A(n11806), .ZN(n6769) );
  INV_X1 U9680 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n6770) );
  NAND2_X1 U9681 ( .A1(n6772), .A2(n11812), .ZN(n6771) );
  OAI21_X2 U9682 ( .B1(n11848), .B2(n6784), .A(n6781), .ZN(n11929) );
  OAI22_X2 U9683 ( .A1(n6789), .A2(n8304), .B1(n13283), .B2(n13373), .ZN(
        n13260) );
  OAI22_X2 U9684 ( .A1(n13231), .A2(n8352), .B1(n12906), .B2(n13432), .ZN(
        n13221) );
  NAND2_X1 U9685 ( .A1(n7874), .A2(n6790), .ZN(n7946) );
  AND2_X1 U9686 ( .A1(n6866), .A2(n6790), .ZN(n7421) );
  NAND2_X2 U9687 ( .A1(n8508), .A2(n6546), .ZN(n12569) );
  NAND2_X2 U9688 ( .A1(n7961), .A2(n6793), .ZN(n8019) );
  OAI21_X1 U9689 ( .B1(n6545), .B2(n10541), .A(n6796), .ZN(n6795) );
  NAND2_X1 U9690 ( .A1(n6545), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6796) );
  OAI21_X1 U9691 ( .B1(n6797), .B2(n7696), .A(n7695), .ZN(n9031) );
  NAND2_X2 U9692 ( .A1(n14488), .A2(n10274), .ZN(n14382) );
  NAND4_X1 U9693 ( .A1(n12424), .A2(P3_ADDR_REG_19__SCAN_IN), .A3(n6800), .A4(
        n6799), .ZN(n6847) );
  NAND2_X1 U9694 ( .A1(n6802), .A2(n10218), .ZN(n10219) );
  AOI21_X1 U9695 ( .B1(n9271), .B2(n9270), .A(n9269), .ZN(n9272) );
  NAND2_X1 U9696 ( .A1(n6804), .A2(n7130), .ZN(n6803) );
  NAND3_X1 U9697 ( .A1(n9235), .A2(n9234), .A3(n7690), .ZN(n6804) );
  OAI21_X1 U9698 ( .B1(n8961), .B2(n6663), .A(n6805), .ZN(n6808) );
  AOI21_X1 U9699 ( .B1(n6808), .B2(n9099), .A(n9098), .ZN(n9100) );
  NAND2_X1 U9700 ( .A1(n6811), .A2(n6810), .ZN(n8903) );
  NAND2_X1 U9701 ( .A1(n9021), .A2(n6812), .ZN(n6814) );
  NAND2_X1 U9702 ( .A1(n6815), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8995) );
  OAI21_X1 U9703 ( .B1(n9188), .B2(n9187), .A(n7705), .ZN(n6819) );
  INV_X1 U9704 ( .A(n8847), .ZN(n6824) );
  NAND2_X1 U9705 ( .A1(n6826), .A2(n8848), .ZN(n6825) );
  NAND2_X1 U9706 ( .A1(n6820), .A2(n7339), .ZN(n8887) );
  NAND3_X1 U9707 ( .A1(n6822), .A2(n6821), .A3(n6635), .ZN(n6820) );
  NAND2_X1 U9708 ( .A1(n6823), .A2(n8846), .ZN(n6821) );
  NAND2_X1 U9709 ( .A1(n6824), .A2(n6825), .ZN(n6822) );
  NAND2_X1 U9710 ( .A1(n11620), .A2(n11619), .ZN(n11782) );
  NAND2_X1 U9711 ( .A1(n11620), .A2(n6675), .ZN(n6830) );
  NAND2_X1 U9712 ( .A1(n14314), .A2(n13692), .ZN(n11789) );
  NAND2_X1 U9713 ( .A1(n6836), .A2(n7252), .ZN(n14045) );
  NAND3_X1 U9714 ( .A1(n6837), .A2(n8893), .A3(n13785), .ZN(n9734) );
  INV_X1 U9715 ( .A(n8892), .ZN(n6838) );
  NAND2_X1 U9716 ( .A1(n6838), .A2(n6794), .ZN(n6837) );
  NAND3_X1 U9717 ( .A1(n6839), .A2(n7590), .A3(n12180), .ZN(n12500) );
  NAND2_X1 U9718 ( .A1(n6839), .A2(n7590), .ZN(n12181) );
  INV_X1 U9719 ( .A(n7020), .ZN(n6843) );
  OAI211_X2 U9720 ( .C1(n14936), .C2(n7019), .A(n6845), .B(n9500), .ZN(n7018)
         );
  MUX2_X1 U9721 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n6546), .Z(n8661) );
  NAND4_X1 U9722 ( .A1(n7182), .A2(n7181), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n6846) );
  NAND2_X1 U9723 ( .A1(n6850), .A2(n13159), .ZN(n12736) );
  NAND2_X1 U9724 ( .A1(n6851), .A2(n7316), .ZN(n6850) );
  NAND3_X1 U9725 ( .A1(n6852), .A2(n12727), .A3(n13196), .ZN(n6851) );
  NAND3_X1 U9726 ( .A1(n12725), .A2(n13205), .A3(n12724), .ZN(n6852) );
  OAI21_X1 U9727 ( .B1(n6855), .B2(n9412), .A(n6854), .ZN(n6853) );
  NAND2_X1 U9728 ( .A1(n6855), .A2(n12761), .ZN(n6854) );
  NAND2_X1 U9729 ( .A1(n7304), .A2(n12759), .ZN(n6855) );
  OAI211_X1 U9730 ( .C1(n6857), .C2(n12752), .A(n12751), .B(n6856), .ZN(n12753) );
  NAND2_X1 U9731 ( .A1(n6857), .A2(n12750), .ZN(n6856) );
  OAI21_X1 U9732 ( .B1(n6858), .B2(n12744), .A(n7315), .ZN(n6857) );
  NAND2_X1 U9733 ( .A1(n7421), .A2(n6864), .ZN(n13478) );
  NAND2_X1 U9734 ( .A1(n7735), .A2(n7421), .ZN(n8053) );
  NAND4_X1 U9735 ( .A1(n7302), .A2(n7299), .A3(n7301), .A4(n7300), .ZN(n6867)
         );
  NAND4_X1 U9736 ( .A1(n7303), .A2(n7880), .A3(n7856), .A4(n7886), .ZN(n7875)
         );
  NAND2_X1 U9737 ( .A1(n6869), .A2(n6872), .ZN(n15502) );
  AND2_X1 U9738 ( .A1(n8066), .A2(n8067), .ZN(n6870) );
  INV_X1 U9739 ( .A(n6873), .ZN(n6871) );
  OAI21_X1 U9740 ( .B1(n8510), .B2(n11254), .A(n6874), .ZN(n6873) );
  NAND2_X1 U9741 ( .A1(n13268), .A2(n13270), .ZN(n13267) );
  INV_X1 U9742 ( .A(n8612), .ZN(n6883) );
  NAND2_X1 U9743 ( .A1(n6546), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U9744 ( .A1(n8609), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U9745 ( .A1(n14868), .A2(n7786), .ZN(n6895) );
  OAI21_X2 U9746 ( .B1(n6896), .B2(n9296), .A(n8895), .ZN(n10177) );
  INV_X1 U9747 ( .A(n6910), .ZN(n7971) );
  INV_X1 U9748 ( .A(n11215), .ZN(n6911) );
  NAND2_X1 U9749 ( .A1(n7464), .A2(n6914), .ZN(n10422) );
  INV_X1 U9750 ( .A(n7980), .ZN(n6918) );
  INV_X1 U9751 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n6930) );
  NAND3_X1 U9752 ( .A1(n7225), .A2(n7224), .A3(n6681), .ZN(n7483) );
  NAND3_X1 U9753 ( .A1(n7224), .A2(n7225), .A3(n6567), .ZN(n7907) );
  INV_X1 U9754 ( .A(n7204), .ZN(n11151) );
  XNOR2_X1 U9755 ( .A(n11161), .B(P3_REG1_REG_2__SCAN_IN), .ZN(n7204) );
  NAND3_X1 U9756 ( .A1(n12812), .A2(n12814), .A3(n12811), .ZN(n12813) );
  OR2_X1 U9757 ( .A1(n7946), .A2(n6944), .ZN(n7866) );
  NAND2_X1 U9758 ( .A1(n7952), .A2(n6946), .ZN(n6947) );
  NAND2_X1 U9759 ( .A1(n8522), .A2(n6948), .ZN(n11261) );
  NAND2_X1 U9760 ( .A1(n12175), .A2(n6950), .ZN(n6949) );
  NAND2_X1 U9761 ( .A1(n8676), .A2(n6574), .ZN(n6956) );
  NAND2_X1 U9762 ( .A1(n6961), .A2(n8678), .ZN(n8679) );
  NAND2_X1 U9763 ( .A1(n8869), .A2(n8642), .ZN(n8892) );
  OAI21_X2 U9764 ( .B1(n8869), .B2(n6794), .A(n6962), .ZN(n8908) );
  NAND2_X1 U9765 ( .A1(n6965), .A2(n15458), .ZN(n6967) );
  INV_X1 U9766 ( .A(n14205), .ZN(n6965) );
  NAND4_X1 U9767 ( .A1(n6967), .A2(n12542), .A3(n14204), .A4(n6966), .ZN(
        n14323) );
  INV_X1 U9768 ( .A(n7557), .ZN(n14006) );
  NAND2_X1 U9769 ( .A1(n6969), .A2(n6970), .ZN(n13993) );
  NAND2_X1 U9770 ( .A1(n7557), .A2(n13995), .ZN(n6969) );
  NAND3_X1 U9771 ( .A1(n6973), .A2(n6688), .A3(n11052), .ZN(n7550) );
  NAND3_X1 U9772 ( .A1(n7692), .A2(n6977), .A3(n7693), .ZN(n6976) );
  NAND2_X1 U9773 ( .A1(n6978), .A2(SI_18_), .ZN(n8980) );
  XNOR2_X1 U9774 ( .A(n6978), .B(SI_18_), .ZN(n8994) );
  NAND2_X1 U9775 ( .A1(n6979), .A2(n10991), .ZN(n10995) );
  NAND2_X1 U9776 ( .A1(n11065), .A2(n10992), .ZN(n6979) );
  NAND2_X1 U9777 ( .A1(n11067), .A2(n11066), .ZN(n11065) );
  XNOR2_X1 U9778 ( .A(n9626), .B(n9627), .ZN(n11066) );
  AND2_X1 U9779 ( .A1(n9624), .A2(n9625), .ZN(n11067) );
  NAND3_X1 U9780 ( .A1(n6981), .A2(n6980), .A3(n6694), .ZN(n6983) );
  NAND3_X1 U9781 ( .A1(n6988), .A2(n6987), .A3(n6582), .ZN(n11119) );
  INV_X1 U9782 ( .A(n9695), .ZN(n6988) );
  NAND2_X1 U9783 ( .A1(n9568), .A2(n9576), .ZN(n9603) );
  NOR2_X2 U9784 ( .A1(n9601), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n10051) );
  MUX2_X1 U9785 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n7000), .S(n15466), .Z(
        P2_U3527) );
  MUX2_X1 U9786 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n7000), .S(n15462), .Z(
        P2_U3495) );
  NAND2_X1 U9787 ( .A1(n7111), .A2(n14209), .ZN(n7000) );
  NAND3_X1 U9788 ( .A1(n11340), .A2(n7575), .A3(n7576), .ZN(n11056) );
  NOR2_X2 U9789 ( .A1(n14013), .A2(n14225), .ZN(n13988) );
  NAND3_X1 U9790 ( .A1(n9605), .A2(n9586), .A3(n9604), .ZN(n7008) );
  NAND2_X1 U9791 ( .A1(n8484), .A2(n8483), .ZN(n7009) );
  NAND2_X1 U9792 ( .A1(n8468), .A2(n8467), .ZN(n7010) );
  INV_X1 U9793 ( .A(n9500), .ZN(n14843) );
  AOI21_X1 U9794 ( .B1(n9500), .B2(n7017), .A(n7016), .ZN(n7015) );
  INV_X1 U9795 ( .A(n9497), .ZN(n7019) );
  NAND3_X1 U9796 ( .A1(n8584), .A2(n8583), .A3(n9064), .ZN(n8704) );
  NAND2_X1 U9797 ( .A1(n8749), .A2(n8707), .ZN(n7021) );
  NOR2_X2 U9798 ( .A1(n7021), .A2(n8704), .ZN(n8594) );
  NAND4_X1 U9799 ( .A1(n8594), .A2(n8718), .A3(n8593), .A4(n8592), .ZN(n7022)
         );
  NAND2_X1 U9800 ( .A1(n11395), .A2(n11394), .ZN(n11393) );
  OAI21_X2 U9801 ( .B1(n11938), .B2(n7756), .A(n7024), .ZN(n11860) );
  INV_X1 U9802 ( .A(n7028), .ZN(n8345) );
  INV_X1 U9803 ( .A(n7029), .ZN(n13144) );
  NOR2_X1 U9804 ( .A1(n8457), .A2(n12941), .ZN(n7030) );
  AND2_X1 U9805 ( .A1(n8359), .A2(n8358), .ZN(n8375) );
  NAND2_X1 U9806 ( .A1(n8359), .A2(n7034), .ZN(n8390) );
  NAND3_X1 U9807 ( .A1(n15561), .A2(n8133), .A3(n7035), .ZN(n8149) );
  OR2_X1 U9808 ( .A1(n10785), .A2(n10786), .ZN(n7037) );
  NAND2_X1 U9809 ( .A1(n10555), .A2(n10663), .ZN(n7054) );
  NAND3_X1 U9810 ( .A1(n7048), .A2(n7046), .A3(n7051), .ZN(n10564) );
  NAND2_X1 U9811 ( .A1(n7047), .A2(n6620), .ZN(n7046) );
  INV_X1 U9812 ( .A(n10555), .ZN(n7047) );
  AOI22_X1 U9813 ( .A1(n10555), .A2(n7050), .B1(n10559), .B2(n7049), .ZN(n7048) );
  AND2_X1 U9814 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10663), .ZN(n7050) );
  INV_X1 U9815 ( .A(n10559), .ZN(n7052) );
  NAND2_X1 U9816 ( .A1(n7055), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n7289) );
  AND3_X1 U9817 ( .A1(n15201), .A2(n7056), .A3(n15200), .ZN(n15209) );
  NAND2_X1 U9818 ( .A1(n15201), .A2(n15200), .ZN(n7057) );
  INV_X1 U9819 ( .A(n15206), .ZN(n7056) );
  NAND2_X1 U9820 ( .A1(n7057), .A2(n15206), .ZN(n15210) );
  NAND3_X1 U9821 ( .A1(n12151), .A2(n12150), .A3(n7293), .ZN(n12355) );
  NAND2_X1 U9822 ( .A1(n12355), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U9823 ( .A1(n7060), .A2(n7058), .ZN(P2_U3528) );
  OR2_X1 U9824 ( .A1(n15466), .A2(n7059), .ZN(n7058) );
  NAND2_X1 U9825 ( .A1(n14323), .A2(n15466), .ZN(n7060) );
  AOI21_X1 U9826 ( .B1(n7254), .B2(n6559), .A(n7253), .ZN(n7252) );
  NAND2_X1 U9827 ( .A1(n8633), .A2(n8632), .ZN(n8854) );
  OAI21_X2 U9828 ( .B1(n7542), .B2(n13714), .A(n7540), .ZN(n13727) );
  NAND2_X1 U9829 ( .A1(n8935), .A2(n8934), .ZN(n8933) );
  MUX2_X1 U9830 ( .A(n13717), .B(n13716), .S(n13810), .Z(n13718) );
  OAI21_X2 U9831 ( .B1(n13746), .B2(n7533), .A(n7532), .ZN(n13751) );
  NAND3_X1 U9832 ( .A1(n8828), .A2(n8833), .A3(n8827), .ZN(n8633) );
  NAND3_X1 U9833 ( .A1(n7062), .A2(n7061), .A3(n6692), .ZN(n7534) );
  NAND2_X1 U9834 ( .A1(n13760), .A2(n13759), .ZN(n7061) );
  NAND2_X1 U9835 ( .A1(n13756), .A2(n13755), .ZN(n7062) );
  NAND2_X1 U9836 ( .A1(n7063), .A2(n10457), .ZN(n10469) );
  NAND2_X1 U9837 ( .A1(n10471), .A2(n10470), .ZN(n7063) );
  NAND2_X1 U9838 ( .A1(n8614), .A2(n8608), .ZN(n8769) );
  NAND3_X1 U9839 ( .A1(n7550), .A2(n7551), .A3(n7549), .ZN(n7123) );
  NAND2_X1 U9840 ( .A1(n7629), .A2(n7628), .ZN(n12007) );
  MUX2_X2 U9841 ( .A(n12470), .B(n12469), .S(n15348), .Z(n12471) );
  INV_X1 U9842 ( .A(n8700), .ZN(n7283) );
  INV_X1 U9843 ( .A(n7172), .ZN(n7171) );
  NOR2_X1 U9844 ( .A1(n9346), .A2(n9347), .ZN(n7273) );
  INV_X1 U9845 ( .A(n7069), .ZN(n7790) );
  OAI21_X1 U9846 ( .B1(n7791), .B2(n14761), .A(n14744), .ZN(n7069) );
  NAND2_X1 U9847 ( .A1(n13960), .A2(n13959), .ZN(n7566) );
  NAND3_X1 U9848 ( .A1(n7075), .A2(n7074), .A3(n10584), .ZN(n10619) );
  NAND2_X1 U9849 ( .A1(n10597), .A2(n11508), .ZN(n7074) );
  INV_X1 U9850 ( .A(n7563), .ZN(n7562) );
  OAI22_X1 U9851 ( .A1(n7702), .A2(n7701), .B1(n7704), .B2(n9175), .ZN(n9188)
         );
  AOI21_X1 U9852 ( .B1(n9274), .B2(n9273), .A(n9272), .ZN(n9379) );
  INV_X1 U9853 ( .A(n9043), .ZN(n7092) );
  NAND2_X1 U9854 ( .A1(n7424), .A2(n13095), .ZN(n7423) );
  AOI22_X2 U9855 ( .A1(n11828), .A2(n11827), .B1(n11838), .B2(n8012), .ZN(
        n12024) );
  NOR2_X1 U9856 ( .A1(n11185), .A2(n11184), .ZN(n11183) );
  NOR2_X1 U9857 ( .A1(n11367), .A2(n11366), .ZN(n11365) );
  NAND3_X1 U9858 ( .A1(n6661), .A2(n8044), .A3(n7222), .ZN(P3_U3201) );
  NAND2_X1 U9859 ( .A1(n7468), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7467) );
  NAND3_X1 U9860 ( .A1(n7471), .A2(P3_REG2_REG_9__SCAN_IN), .A3(n12088), .ZN(
        n12025) );
  AOI21_X1 U9861 ( .B1(n11217), .B2(n6910), .A(n11369), .ZN(n11368) );
  NAND3_X1 U9862 ( .A1(n7188), .A2(n7189), .A3(n8594), .ZN(n7077) );
  OR2_X2 U9863 ( .A1(n8510), .A2(n12463), .ZN(n8495) );
  NAND2_X1 U9864 ( .A1(n7391), .A2(n7320), .ZN(n7319) );
  OAI21_X2 U9865 ( .B1(n12037), .B2(n13862), .A(n7835), .ZN(n12175) );
  INV_X1 U9866 ( .A(n7370), .ZN(n10403) );
  NAND2_X1 U9867 ( .A1(n13585), .A2(n6602), .ZN(n7607) );
  INV_X2 U9868 ( .A(n13836), .ZN(n13638) );
  NAND2_X1 U9869 ( .A1(n11873), .A2(n7751), .ZN(n7750) );
  NAND2_X1 U9870 ( .A1(n14759), .A2(n14761), .ZN(n7082) );
  AOI21_X1 U9871 ( .B1(n15222), .B2(n15221), .A(n7088), .ZN(n15230) );
  AND2_X1 U9872 ( .A1(n12367), .A2(n6608), .ZN(n7298) );
  AOI21_X1 U9873 ( .B1(n7091), .B2(n7090), .A(n9117), .ZN(n7089) );
  OAI211_X1 U9874 ( .C1(n13718), .C2(n7543), .A(n13719), .B(n13715), .ZN(n7539) );
  NAND2_X1 U9875 ( .A1(n7094), .A2(n12767), .ZN(P3_U3296) );
  NAND3_X1 U9876 ( .A1(n7318), .A2(n7319), .A3(n7390), .ZN(n7094) );
  OAI22_X2 U9877 ( .A1(n12024), .A2(n12023), .B1(n8013), .B2(n12028), .ZN(
        n12084) );
  NAND2_X1 U9878 ( .A1(n7236), .A2(n10910), .ZN(n10912) );
  XNOR2_X1 U9879 ( .A(n8036), .B(n8035), .ZN(n7424) );
  OAI21_X1 U9880 ( .B1(n6605), .B2(n7432), .A(n7430), .ZN(n11224) );
  NAND2_X1 U9881 ( .A1(n9671), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9705) );
  NOR2_X2 U9882 ( .A1(n9800), .A2(n9799), .ZN(n7100) );
  NOR2_X2 U9883 ( .A1(n9883), .A2(n9882), .ZN(n7101) );
  NOR2_X1 U9884 ( .A1(n7795), .A2(n10240), .ZN(n7794) );
  MUX2_X1 U9885 ( .A(n10515), .B(n10495), .S(n6546), .Z(n8626) );
  NAND2_X1 U9886 ( .A1(n8626), .A2(n8618), .ZN(n8816) );
  NAND2_X1 U9887 ( .A1(n7292), .A2(n12356), .ZN(n12364) );
  XNOR2_X1 U9888 ( .A(n8984), .B(n8731), .ZN(n8734) );
  AOI21_X2 U9889 ( .B1(n14148), .B2(n13864), .A(n6639), .ZN(n14125) );
  NAND2_X1 U9890 ( .A1(n13993), .A2(n12531), .ZN(n13975) );
  NAND2_X1 U9891 ( .A1(n8624), .A2(SI_3_), .ZN(n8813) );
  INV_X1 U9892 ( .A(n7603), .ZN(n7602) );
  INV_X1 U9893 ( .A(n13015), .ZN(n7462) );
  NAND2_X1 U9894 ( .A1(n7469), .A2(n8309), .ZN(n7468) );
  XNOR2_X1 U9895 ( .A(n7889), .B(n7890), .ZN(n11197) );
  NAND2_X1 U9896 ( .A1(n12025), .A2(n12088), .ZN(n7974) );
  INV_X1 U9897 ( .A(n9230), .ZN(n9233) );
  NAND3_X1 U9898 ( .A1(n7780), .A2(n11517), .A3(n7783), .ZN(n11513) );
  NAND2_X1 U9899 ( .A1(n7291), .A2(n7290), .ZN(n12366) );
  OR2_X1 U9900 ( .A1(n8908), .A2(n8907), .ZN(n8909) );
  OAI21_X1 U9901 ( .B1(n15108), .B2(n9554), .A(n7108), .ZN(P1_U3523) );
  OAI22_X2 U9902 ( .A1(n14159), .A2(n12523), .B1(n13733), .B2(n14170), .ZN(
        n14148) );
  AOI21_X2 U9903 ( .B1(n13947), .B2(n13946), .A(n13945), .ZN(n14209) );
  NAND2_X1 U9904 ( .A1(n7666), .A2(n7668), .ZN(n8186) );
  NAND2_X1 U9905 ( .A1(n8340), .A2(n8339), .ZN(n8354) );
  OAI21_X1 U9906 ( .B1(n13398), .B2(n15546), .A(n7113), .ZN(P3_U3486) );
  OAI21_X1 U9907 ( .B1(n13398), .B2(n15539), .A(n7115), .ZN(P3_U3454) );
  NAND2_X1 U9908 ( .A1(n7402), .A2(n12729), .ZN(n7401) );
  AOI21_X1 U9909 ( .B1(n8081), .B2(n8080), .A(n7839), .ZN(n8095) );
  NAND2_X1 U9910 ( .A1(n8641), .A2(n8640), .ZN(n7117) );
  INV_X1 U9911 ( .A(n9968), .ZN(n7623) );
  NOR2_X1 U9912 ( .A1(n13687), .A2(n11736), .ZN(n11725) );
  AOI21_X1 U9913 ( .B1(n7385), .B2(n13178), .A(n7383), .ZN(n7382) );
  NAND2_X1 U9914 ( .A1(n7123), .A2(n11724), .ZN(n11786) );
  NAND2_X1 U9915 ( .A1(n12532), .A2(n13842), .ZN(n13960) );
  NAND2_X1 U9916 ( .A1(n7125), .A2(n7124), .ZN(P2_U3496) );
  NAND2_X1 U9917 ( .A1(n14323), .A2(n15462), .ZN(n7125) );
  NAND4_X2 U9918 ( .A1(n9678), .A2(n9677), .A3(n9676), .A4(n9675), .ZN(n13903)
         );
  NAND3_X1 U9919 ( .A1(n8654), .A2(n7697), .A3(n7700), .ZN(n7168) );
  INV_X1 U9920 ( .A(n7180), .ZN(n7176) );
  OR4_X1 U9921 ( .A1(n14773), .A2(n14793), .A3(n14820), .A4(n9370), .ZN(n9371)
         );
  NAND3_X1 U9922 ( .A1(n9372), .A2(n6564), .A3(n9353), .ZN(n9374) );
  OAI22_X1 U9923 ( .A1(n8824), .A2(n7344), .B1(n8825), .B2(n7343), .ZN(n8847)
         );
  OR2_X4 U9924 ( .A1(n8603), .A2(n8598), .ZN(n9257) );
  AND2_X1 U9925 ( .A1(n8592), .A2(n8593), .ZN(n7188) );
  NAND2_X1 U9926 ( .A1(n8887), .A2(n8888), .ZN(n8886) );
  INV_X1 U9927 ( .A(n7982), .ZN(n7469) );
  NAND2_X1 U9928 ( .A1(n7391), .A2(n6732), .ZN(n7318) );
  NAND4_X1 U9929 ( .A1(n12735), .A2(n13159), .A3(n13171), .A4(n6612), .ZN(
        n12610) );
  NAND2_X1 U9931 ( .A1(n7132), .A2(n7131), .ZN(n9118) );
  INV_X1 U9932 ( .A(n12364), .ZN(n7291) );
  NAND2_X1 U9933 ( .A1(n7286), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n11556) );
  NAND2_X1 U9934 ( .A1(n12149), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U9935 ( .A1(n7687), .A2(n7336), .ZN(P1_U3242) );
  INV_X1 U9936 ( .A(n9156), .ZN(n7702) );
  NAND2_X1 U9937 ( .A1(n8767), .A2(n8756), .ZN(n12473) );
  NAND2_X1 U9938 ( .A1(n12430), .A2(n12429), .ZN(n12856) );
  NAND3_X1 U9939 ( .A1(n7138), .A2(n12427), .A3(n7137), .ZN(n12950) );
  NAND3_X1 U9940 ( .A1(n12799), .A2(n6560), .A3(n12343), .ZN(n7138) );
  OAI21_X1 U9941 ( .B1(n12919), .B2(n7148), .A(n7145), .ZN(n12840) );
  NAND2_X1 U9942 ( .A1(n12919), .A2(n7145), .ZN(n7144) );
  NAND2_X1 U9943 ( .A1(n7151), .A2(n7153), .ZN(n7152) );
  NAND3_X1 U9944 ( .A1(n12883), .A2(n6713), .A3(n12890), .ZN(n7151) );
  NOR2_X1 U9945 ( .A1(n7154), .A2(n7152), .ZN(P3_U3169) );
  XNOR2_X1 U9946 ( .A(n12883), .B(n12884), .ZN(n12885) );
  NAND2_X1 U9947 ( .A1(n6945), .A2(n6693), .ZN(n8501) );
  INV_X1 U9948 ( .A(n8501), .ZN(n7952) );
  NAND2_X1 U9949 ( .A1(n7169), .A2(n6571), .ZN(n9085) );
  NAND2_X1 U9950 ( .A1(n8906), .A2(n6628), .ZN(n7169) );
  NOR2_X2 U9951 ( .A1(n10347), .A2(n10346), .ZN(n10348) );
  OAI21_X1 U9952 ( .B1(n14758), .B2(n7170), .A(n7171), .ZN(n10347) );
  OR2_X2 U9953 ( .A1(n7790), .A2(n9471), .ZN(n7173) );
  INV_X1 U9954 ( .A(n7174), .ZN(n7178) );
  NAND2_X1 U9955 ( .A1(n7176), .A2(n9046), .ZN(n9063) );
  NAND2_X1 U9956 ( .A1(n9046), .A2(n9045), .ZN(n9061) );
  NAND3_X1 U9957 ( .A1(n9046), .A2(n7179), .A3(n7180), .ZN(n7177) );
  NOR2_X1 U9958 ( .A1(n14961), .A2(n14950), .ZN(n7184) );
  NAND2_X1 U9959 ( .A1(n15151), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8596) );
  NAND4_X1 U9960 ( .A1(n8594), .A2(n8592), .A3(n8593), .A4(n7186), .ZN(n15151)
         );
  NAND3_X1 U9961 ( .A1(n7191), .A2(n7190), .A3(n7192), .ZN(n12496) );
  NAND2_X1 U9962 ( .A1(n10355), .A2(n9515), .ZN(n7190) );
  OR2_X1 U9963 ( .A1(n10355), .A2(n7193), .ZN(n7191) );
  NAND3_X1 U9964 ( .A1(n9528), .A2(n7851), .A3(n7195), .ZN(n9553) );
  NAND2_X1 U9965 ( .A1(n12496), .A2(n15331), .ZN(n7195) );
  NAND2_X1 U9966 ( .A1(n7196), .A2(n7747), .ZN(n12051) );
  NAND2_X1 U9967 ( .A1(n11516), .A2(n7749), .ZN(n7196) );
  INV_X1 U9968 ( .A(n14978), .ZN(n7197) );
  AND3_X1 U9969 ( .A1(n7476), .A2(n7475), .A3(n10451), .ZN(n7897) );
  NAND2_X1 U9970 ( .A1(n13048), .A2(n6729), .ZN(n7207) );
  NAND2_X1 U9971 ( .A1(n7478), .A2(n7479), .ZN(n13048) );
  NAND2_X1 U9972 ( .A1(n7925), .A2(n7210), .ZN(n7211) );
  NAND2_X1 U9973 ( .A1(n7217), .A2(n7216), .ZN(n13020) );
  NAND3_X1 U9974 ( .A1(n7234), .A2(n7233), .A3(n7921), .ZN(n7231) );
  INV_X1 U9975 ( .A(n7920), .ZN(n7235) );
  OAI21_X1 U9976 ( .B1(n10868), .B2(n13848), .A(n7236), .ZN(n11336) );
  NAND2_X1 U9977 ( .A1(n10868), .A2(n13848), .ZN(n7236) );
  OAI211_X1 U9978 ( .C1(n7589), .C2(n7238), .A(n7237), .B(n12039), .ZN(n12179)
         );
  OAI22_X1 U9979 ( .A1(n7240), .A2(n13858), .B1(n7242), .B2(n7241), .ZN(n7239)
         );
  NAND2_X1 U9980 ( .A1(n7249), .A2(n7248), .ZN(n14131) );
  INV_X1 U9981 ( .A(n7250), .ZN(n7249) );
  OAI21_X1 U9982 ( .B1(n7251), .B2(n14165), .A(n12502), .ZN(n7250) );
  NAND2_X1 U9983 ( .A1(n14166), .A2(n14165), .ZN(n14164) );
  AOI21_X2 U9984 ( .B1(n13987), .B2(n12513), .A(n12512), .ZN(n13981) );
  NAND2_X1 U9985 ( .A1(n8609), .A2(n10518), .ZN(n7272) );
  NAND3_X1 U9986 ( .A1(n7275), .A2(n9331), .A3(n7274), .ZN(n9344) );
  OAI21_X1 U9987 ( .B1(n8700), .B2(n7279), .A(n7277), .ZN(n9293) );
  OR2_X1 U9988 ( .A1(n7286), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7285) );
  XNOR2_X1 U9989 ( .A(n11552), .B(n11553), .ZN(n7286) );
  NAND2_X1 U9990 ( .A1(n10467), .A2(n10462), .ZN(n7288) );
  NAND2_X1 U9991 ( .A1(n7295), .A2(n11911), .ZN(n11920) );
  NAND2_X1 U9992 ( .A1(n7298), .A2(n12368), .ZN(n7297) );
  NAND3_X1 U9993 ( .A1(n12753), .A2(n12755), .A3(n12754), .ZN(n7304) );
  INV_X1 U9994 ( .A(n12695), .ZN(n7305) );
  OAI211_X1 U9995 ( .C1(n7314), .C2(n7308), .A(n7307), .B(n12696), .ZN(n7306)
         );
  OR2_X1 U9996 ( .A1(n12682), .A2(n12683), .ZN(n7308) );
  NAND2_X1 U9997 ( .A1(n12664), .A2(n7310), .ZN(n7309) );
  NOR2_X1 U9998 ( .A1(n12682), .A2(n7311), .ZN(n7310) );
  NOR2_X1 U9999 ( .A1(n12695), .A2(n6676), .ZN(n7312) );
  INV_X1 U10000 ( .A(n9266), .ZN(n7323) );
  AND3_X1 U10001 ( .A1(n8738), .A2(n6678), .A3(n7324), .ZN(n7327) );
  NAND2_X2 U10002 ( .A1(n8603), .A2(n15160), .ZN(n9316) );
  INV_X1 U10003 ( .A(n8603), .ZN(n8599) );
  NAND2_X1 U10004 ( .A1(n8737), .A2(n7327), .ZN(n10118) );
  NAND2_X1 U10005 ( .A1(n7330), .A2(n7328), .ZN(n8921) );
  NAND2_X1 U10006 ( .A1(n8903), .A2(n7331), .ZN(n7330) );
  INV_X1 U10007 ( .A(n8823), .ZN(n7343) );
  NOR2_X1 U10008 ( .A1(n8826), .A2(n8823), .ZN(n7344) );
  NAND2_X1 U10009 ( .A1(n7350), .A2(n7353), .ZN(n7349) );
  INV_X1 U10010 ( .A(n8119), .ZN(n7350) );
  NAND3_X1 U10011 ( .A1(n8099), .A2(n6691), .A3(n11645), .ZN(n7351) );
  NAND2_X1 U10012 ( .A1(n7354), .A2(n8119), .ZN(n11764) );
  NAND2_X1 U10013 ( .A1(n12275), .A2(n7356), .ZN(n7355) );
  NAND2_X1 U10014 ( .A1(n10395), .A2(n10394), .ZN(n7371) );
  NAND3_X1 U10015 ( .A1(n7367), .A2(n7368), .A3(n7371), .ZN(n7370) );
  INV_X1 U10016 ( .A(n10395), .ZN(n7366) );
  NAND3_X1 U10017 ( .A1(n7371), .A2(n7372), .A3(n7367), .ZN(n13116) );
  NAND2_X1 U10018 ( .A1(n7381), .A2(n7378), .ZN(n8548) );
  OAI211_X2 U10019 ( .C1(SI_3_), .C2(n12569), .A(n7379), .B(n6609), .ZN(n15482) );
  OAI21_X1 U10020 ( .B1(n13179), .B2(n7384), .A(n7382), .ZN(n8465) );
  NAND2_X1 U10021 ( .A1(n6568), .A2(n12756), .ZN(n7388) );
  OAI21_X1 U10022 ( .B1(n12575), .B2(n12574), .A(n12573), .ZN(n7389) );
  NAND2_X1 U10023 ( .A1(n13138), .A2(n6679), .ZN(n7414) );
  AOI21_X1 U10024 ( .B1(n13138), .B2(n12738), .A(n7420), .ZN(n13126) );
  NAND2_X1 U10025 ( .A1(n13057), .A2(n7427), .ZN(n7426) );
  NAND2_X2 U10026 ( .A1(n7426), .A2(n7425), .ZN(n8032) );
  NAND2_X1 U10027 ( .A1(n11152), .A2(n7431), .ZN(n7430) );
  AND2_X1 U10028 ( .A1(n7436), .A2(n7438), .ZN(n7431) );
  INV_X1 U10029 ( .A(n7438), .ZN(n7432) );
  OAI21_X1 U10030 ( .B1(n12084), .B2(n7441), .A(n7439), .ZN(n7450) );
  INV_X1 U10031 ( .A(n7450), .ZN(n12995) );
  INV_X1 U10032 ( .A(n7457), .ZN(n11832) );
  NAND2_X1 U10033 ( .A1(n7459), .A2(n6629), .ZN(n7980) );
  NAND2_X1 U10034 ( .A1(n7467), .A2(n13081), .ZN(n7984) );
  INV_X1 U10035 ( .A(n7973), .ZN(n7470) );
  INV_X1 U10036 ( .A(n7476), .ZN(n11149) );
  NAND2_X1 U10037 ( .A1(n7937), .A2(n13044), .ZN(n7478) );
  NAND2_X1 U10038 ( .A1(n6587), .A2(n7917), .ZN(n12029) );
  NAND2_X1 U10039 ( .A1(n11841), .A2(n11839), .ZN(n7484) );
  NAND3_X1 U10040 ( .A1(n7484), .A2(n7485), .A3(n7488), .ZN(n7916) );
  NAND3_X1 U10041 ( .A1(n7912), .A2(n7487), .A3(n7486), .ZN(n7485) );
  INV_X1 U10042 ( .A(n11838), .ZN(n7489) );
  NAND2_X1 U10043 ( .A1(n10372), .A2(n7497), .ZN(n14724) );
  NAND3_X1 U10044 ( .A1(n7493), .A2(n7491), .A3(n7490), .ZN(n14718) );
  NAND3_X1 U10045 ( .A1(n7504), .A2(n6603), .A3(n12205), .ZN(n7503) );
  MUX2_X1 U10047 ( .A(n6543), .B(n10871), .S(n6532), .Z(n13648) );
  NAND2_X4 U10048 ( .A1(n13638), .A2(n9912), .ZN(n13792) );
  INV_X1 U10049 ( .A(n10083), .ZN(n7527) );
  OAI211_X2 U10050 ( .C1(n6658), .C2(n7527), .A(n7530), .B(n7526), .ZN(n9878)
         );
  NAND2_X1 U10051 ( .A1(n7534), .A2(n7535), .ZN(n13765) );
  INV_X1 U10052 ( .A(n13713), .ZN(n7543) );
  AND2_X1 U10053 ( .A1(n7539), .A2(n7537), .ZN(n7540) );
  AOI21_X1 U10054 ( .B1(n7538), .B2(n13718), .A(n7541), .ZN(n7537) );
  NAND3_X1 U10055 ( .A1(n7546), .A2(n13695), .A3(n7544), .ZN(n13697) );
  NAND3_X1 U10056 ( .A1(n7545), .A2(n13690), .A3(n13691), .ZN(n7544) );
  INV_X1 U10057 ( .A(n13688), .ZN(n7545) );
  NAND3_X1 U10058 ( .A1(n13689), .A2(n13691), .A3(n7547), .ZN(n7546) );
  NAND2_X1 U10059 ( .A1(n7548), .A2(n13688), .ZN(n7547) );
  INV_X1 U10060 ( .A(n13690), .ZN(n7548) );
  NAND2_X1 U10061 ( .A1(n7552), .A2(n11622), .ZN(n11700) );
  NAND2_X1 U10062 ( .A1(n11621), .A2(n13852), .ZN(n7552) );
  NAND2_X1 U10063 ( .A1(n7554), .A2(n13680), .ZN(n7553) );
  NAND2_X1 U10064 ( .A1(n7555), .A2(n11622), .ZN(n7554) );
  INV_X1 U10065 ( .A(n13852), .ZN(n7555) );
  NAND2_X1 U10066 ( .A1(n7566), .A2(n12533), .ZN(n13944) );
  NAND2_X1 U10067 ( .A1(n14105), .A2(n7850), .ZN(n7574) );
  NAND2_X1 U10068 ( .A1(n7567), .A2(n7570), .ZN(n14079) );
  NAND2_X1 U10069 ( .A1(n14105), .A2(n7568), .ZN(n7567) );
  NAND2_X1 U10070 ( .A1(n13973), .A2(n7580), .ZN(n7582) );
  INV_X1 U10071 ( .A(n7582), .ZN(n13938) );
  XNOR2_X1 U10072 ( .A(n7589), .B(n11887), .ZN(n14306) );
  INV_X1 U10073 ( .A(n12514), .ZN(n7595) );
  OAI21_X1 U10074 ( .B1(n14070), .B2(n12506), .A(n12507), .ZN(n14066) );
  NAND2_X1 U10075 ( .A1(n7623), .A2(n7619), .ZN(n7616) );
  NAND3_X1 U10076 ( .A1(n7617), .A2(n7616), .A3(n7612), .ZN(n13617) );
  OR2_X1 U10077 ( .A1(n7623), .A2(n7622), .ZN(n7618) );
  OR2_X1 U10078 ( .A1(n13535), .A2(n7621), .ZN(n7620) );
  NAND2_X1 U10079 ( .A1(n9968), .A2(n9967), .ZN(n13568) );
  NAND2_X1 U10080 ( .A1(n11753), .A2(n7630), .ZN(n7629) );
  NAND2_X1 U10081 ( .A1(n7649), .A2(n7653), .ZN(n8371) );
  NAND2_X1 U10082 ( .A1(n8340), .A2(n7650), .ZN(n7649) );
  NAND2_X1 U10083 ( .A1(n7656), .A2(n7658), .ZN(n8295) );
  NAND2_X1 U10084 ( .A1(n8235), .A2(n6711), .ZN(n7656) );
  NAND2_X1 U10085 ( .A1(n8144), .A2(n6685), .ZN(n7666) );
  NAND2_X1 U10086 ( .A1(n10379), .A2(n7683), .ZN(n7678) );
  OAI21_X1 U10087 ( .B1(n10379), .B2(n6585), .A(n10378), .ZN(n12553) );
  NAND3_X1 U10088 ( .A1(n7686), .A2(n7685), .A3(n6604), .ZN(n9098) );
  NAND2_X1 U10089 ( .A1(n9387), .A2(n9386), .ZN(n7687) );
  NAND2_X1 U10090 ( .A1(n8906), .A2(n8647), .ZN(n8935) );
  INV_X1 U10091 ( .A(n9174), .ZN(n7704) );
  INV_X1 U10092 ( .A(n9200), .ZN(n7706) );
  OAI21_X1 U10093 ( .B1(n11270), .B2(n7707), .A(n12812), .ZN(n11271) );
  NAND2_X1 U10094 ( .A1(n11270), .A2(n7707), .ZN(n12812) );
  XNOR2_X1 U10095 ( .A(n11422), .B(n15506), .ZN(n7707) );
  NAND3_X1 U10096 ( .A1(n7709), .A2(n7722), .A3(n7708), .ZN(n7715) );
  NAND2_X1 U10097 ( .A1(n7719), .A2(n7710), .ZN(n7708) );
  NAND2_X1 U10098 ( .A1(n12847), .A2(n7710), .ZN(n7709) );
  NAND2_X1 U10099 ( .A1(n12847), .A2(n7721), .ZN(n7716) );
  AOI21_X1 U10100 ( .B1(n12847), .B2(n12848), .A(n7723), .ZN(n12939) );
  XNOR2_X1 U10101 ( .A(n7715), .B(n6644), .ZN(n12468) );
  AND2_X1 U10102 ( .A1(n12458), .A2(n8572), .ZN(n7723) );
  NAND2_X1 U10103 ( .A1(n8519), .A2(n6690), .ZN(n8522) );
  INV_X1 U10104 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7729) );
  NAND2_X1 U10105 ( .A1(n14812), .A2(n9504), .ZN(n7752) );
  INV_X1 U10106 ( .A(n8717), .ZN(n7765) );
  NAND3_X1 U10107 ( .A1(n8718), .A2(n8709), .A3(n8710), .ZN(n9394) );
  AND3_X2 U10108 ( .A1(n8749), .A2(n8702), .A3(n8773), .ZN(n8716) );
  NAND2_X1 U10109 ( .A1(n7765), .A2(n6648), .ZN(n7764) );
  NAND3_X1 U10110 ( .A1(n7768), .A2(n9435), .A3(n7766), .ZN(n11301) );
  NAND3_X1 U10111 ( .A1(n11351), .A2(n15275), .A3(n9432), .ZN(n7768) );
  NAND2_X1 U10112 ( .A1(n14917), .A2(n7775), .ZN(n7771) );
  NAND2_X1 U10113 ( .A1(n7771), .A2(n7772), .ZN(n14868) );
  NAND2_X1 U10114 ( .A1(n9449), .A2(n7781), .ZN(n7780) );
  NAND2_X1 U10115 ( .A1(n9450), .A2(n7782), .ZN(n7783) );
  INV_X1 U10116 ( .A(n11855), .ZN(n7782) );
  OAI21_X1 U10117 ( .B1(n14850), .B2(n6556), .A(n7786), .ZN(n14821) );
  INV_X1 U10118 ( .A(n9471), .ZN(n7792) );
  NAND2_X1 U10119 ( .A1(n10161), .A2(n7793), .ZN(n11603) );
  NAND2_X1 U10120 ( .A1(n10146), .A2(n10145), .ZN(n10430) );
  NAND2_X1 U10121 ( .A1(n11545), .A2(n7803), .ZN(n7802) );
  NAND2_X1 U10122 ( .A1(n14382), .A2(n14383), .ZN(n7818) );
  NAND2_X1 U10123 ( .A1(n10280), .A2(n10279), .ZN(n7817) );
  NAND2_X1 U10124 ( .A1(n14392), .A2(n7821), .ZN(n7820) );
  AND2_X1 U10125 ( .A1(n7825), .A2(n7824), .ZN(n14474) );
  INV_X1 U10126 ( .A(n7825), .ZN(n14391) );
  NAND2_X1 U10127 ( .A1(n10257), .A2(n10258), .ZN(n7824) );
  NAND2_X1 U10128 ( .A1(n8716), .A2(n7826), .ZN(n7830) );
  NAND3_X1 U10129 ( .A1(n8718), .A2(n8715), .A3(n8589), .ZN(n7827) );
  CLKBUF_X1 U10130 ( .A(n11929), .Z(n11930) );
  NAND2_X1 U10131 ( .A1(n8505), .A2(n8504), .ZN(n10395) );
  NAND2_X2 U10132 ( .A1(n9703), .A2(n9702), .ZN(n15438) );
  INV_X1 U10133 ( .A(n13942), .ZN(n14201) );
  NAND2_X1 U10134 ( .A1(n9747), .A2(n11408), .ZN(n11753) );
  OR2_X1 U10135 ( .A1(n13167), .A2(n13149), .ZN(n13153) );
  AND2_X1 U10136 ( .A1(n10826), .A2(n13835), .ZN(n14315) );
  NAND2_X1 U10137 ( .A1(n12396), .A2(n15320), .ZN(n10375) );
  NAND2_X1 U10138 ( .A1(n12396), .A2(n10368), .ZN(n10369) );
  OAI21_X1 U10139 ( .B1(n13119), .B2(n13386), .A(n10399), .ZN(n10400) );
  NAND2_X1 U10140 ( .A1(n9652), .A2(n13906), .ZN(n9642) );
  NAND2_X1 U10141 ( .A1(n9605), .A2(n7846), .ZN(n9612) );
  OR2_X1 U10142 ( .A1(n8437), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8438) );
  INV_X1 U10143 ( .A(n11924), .ZN(n13884) );
  INV_X1 U10144 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U10145 ( .A1(n9518), .A2(n15322), .ZN(n11592) );
  INV_X1 U10146 ( .A(n15286), .ZN(n9518) );
  INV_X1 U10147 ( .A(n14738), .ZN(n12472) );
  INV_X1 U10148 ( .A(n8708), .ZN(n8709) );
  NAND2_X1 U10149 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), 
        .ZN(n7889) );
  CLKBUF_X1 U10150 ( .A(n11846), .Z(n11847) );
  NAND2_X2 U10151 ( .A1(n13037), .A2(n7847), .ZN(n13057) );
  NAND2_X1 U10152 ( .A1(n8053), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7958) );
  OAI21_X1 U10153 ( .B1(n13840), .B2(n7849), .A(n13839), .ZN(n13888) );
  NAND2_X1 U10154 ( .A1(n13840), .A2(n13838), .ZN(n13839) );
  INV_X1 U10155 ( .A(n8054), .ZN(n13484) );
  NAND2_X1 U10156 ( .A1(n9140), .A2(n9139), .ZN(n9154) );
  AND2_X1 U10157 ( .A1(n10122), .A2(n10121), .ZN(n10852) );
  CLKBUF_X1 U10158 ( .A(n14409), .Z(n14500) );
  INV_X1 U10159 ( .A(n9308), .ZN(n12384) );
  OAI21_X1 U10160 ( .B1(n6546), .B2(n10489), .A(n8619), .ZN(n8624) );
  OAI21_X1 U10161 ( .B1(n9379), .B2(n7844), .A(n9378), .ZN(n9387) );
  INV_X1 U10162 ( .A(n8704), .ZN(n8705) );
  NOR2_X1 U10163 ( .A1(n12220), .A2(n12831), .ZN(n12221) );
  INV_X1 U10164 ( .A(n14137), .ZN(n14144) );
  INV_X1 U10165 ( .A(n9520), .ZN(n15165) );
  NAND2_X1 U10166 ( .A1(n9732), .A2(n10676), .ZN(n9619) );
  NAND2_X1 U10167 ( .A1(n9480), .A2(n9479), .ZN(n9482) );
  NAND3_X1 U10168 ( .A1(n8053), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_IR_REG_30__SCAN_IN), .ZN(n8051) );
  NOR2_X2 U10169 ( .A1(n10348), .A2(n6626), .ZN(n9473) );
  INV_X1 U10170 ( .A(n11926), .ZN(n9386) );
  NAND2_X2 U10171 ( .A1(n12487), .A2(n15280), .ZN(n14987) );
  INV_X1 U10172 ( .A(n15342), .ZN(n9554) );
  AND2_X2 U10173 ( .A1(n9551), .A2(n9547), .ZN(n15348) );
  OR2_X1 U10174 ( .A1(n15262), .A2(n14567), .ZN(n7832) );
  OR2_X1 U10175 ( .A1(n12756), .A2(n12613), .ZN(n7833) );
  INV_X1 U10176 ( .A(n11789), .ZN(n11787) );
  AND2_X1 U10177 ( .A1(n8579), .A2(n13383), .ZN(n7834) );
  NOR2_X1 U10178 ( .A1(n13832), .A2(n13831), .ZN(n7837) );
  OR2_X1 U10179 ( .A1(n12472), .A2(n15147), .ZN(n7838) );
  AND2_X1 U10180 ( .A1(n10503), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7839) );
  AND4_X1 U10181 ( .A1(n10058), .A2(n9606), .A3(n9595), .A4(n14344), .ZN(n7840) );
  OR2_X1 U10182 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7841) );
  OR2_X1 U10183 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7842) );
  INV_X1 U10184 ( .A(n10532), .ZN(n9532) );
  INV_X2 U10185 ( .A(n12966), .ZN(P3_U3897) );
  INV_X1 U10186 ( .A(n11940), .ZN(n10368) );
  INV_X1 U10187 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n15816) );
  OR2_X1 U10188 ( .A1(n9347), .A2(n9346), .ZN(n7844) );
  INV_X1 U10189 ( .A(n14119), .ZN(n12504) );
  INV_X1 U10190 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8732) );
  INV_X1 U10191 ( .A(n8726), .ZN(n9019) );
  AND3_X1 U10192 ( .A1(n9604), .A2(P2_IR_REG_29__SCAN_IN), .A3(n9606), .ZN(
        n7846) );
  OR2_X1 U10193 ( .A1(n8025), .A2(n8280), .ZN(n7847) );
  AND2_X1 U10194 ( .A1(n11385), .A2(n12613), .ZN(n12760) );
  INV_X1 U10195 ( .A(n13320), .ZN(n15491) );
  AND2_X1 U10196 ( .A1(n13834), .A2(n9912), .ZN(n7849) );
  NAND2_X1 U10197 ( .A1(n10958), .A2(n15431), .ZN(n15460) );
  NAND2_X2 U10198 ( .A1(n11667), .A2(n14146), .ZN(n14135) );
  INV_X1 U10199 ( .A(n11276), .ZN(n11265) );
  OR2_X1 U10200 ( .A1(n14115), .A2(n13892), .ZN(n7850) );
  AND4_X1 U10201 ( .A1(n12494), .A2(n9527), .A3(n12488), .A4(n12486), .ZN(
        n7851) );
  INV_X1 U10202 ( .A(n13168), .ZN(n8572) );
  NOR2_X1 U10203 ( .A1(n13218), .A2(n13216), .ZN(n7852) );
  OR2_X1 U10204 ( .A1(n9422), .A2(n11531), .ZN(n15546) );
  INV_X2 U10205 ( .A(n15539), .ZN(n15540) );
  NAND2_X1 U10206 ( .A1(n13665), .A2(n13664), .ZN(n13666) );
  AND2_X1 U10207 ( .A1(n13853), .A2(n13666), .ZN(n13667) );
  OAI21_X1 U10208 ( .B1(n13741), .B2(n13740), .A(n13739), .ZN(n13746) );
  OAI21_X1 U10209 ( .B1(n9154), .B2(n9153), .A(n9152), .ZN(n9156) );
  MUX2_X1 U10210 ( .A(n12623), .B(n12622), .S(n12752), .Z(n12737) );
  INV_X1 U10211 ( .A(n9250), .ZN(n9251) );
  INV_X1 U10212 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U10213 ( .A1(n11787), .A2(n11788), .ZN(n11790) );
  NAND2_X1 U10214 ( .A1(n9303), .A2(n8760), .ZN(n9304) );
  NAND2_X1 U10215 ( .A1(n8588), .A2(n8587), .ZN(n8703) );
  NOR2_X1 U10216 ( .A1(n12791), .A2(n13208), .ZN(n12446) );
  INV_X1 U10217 ( .A(n13293), .ZN(n8268) );
  INV_X1 U10218 ( .A(n11647), .ZN(n8099) );
  NAND2_X1 U10219 ( .A1(n7902), .A2(n7854), .ZN(n7855) );
  INV_X1 U10220 ( .A(n11587), .ZN(n9438) );
  NOR2_X1 U10221 ( .A1(n8703), .A2(n8708), .ZN(n8592) );
  INV_X1 U10222 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8715) );
  OR2_X1 U10223 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14649), .ZN(n10777) );
  OAI21_X1 U10224 ( .B1(n12757), .B2(n12962), .A(n12756), .ZN(n12758) );
  NAND2_X1 U10225 ( .A1(n13489), .A2(n7477), .ZN(n7988) );
  OR2_X1 U10226 ( .A1(n8027), .A2(n8296), .ZN(n8028) );
  INV_X1 U10227 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U10228 ( .A1(n12695), .A2(n8268), .ZN(n8275) );
  AND2_X1 U10229 ( .A1(n10489), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8108) );
  OAI21_X1 U10230 ( .B1(n10239), .B2(n14428), .A(n14430), .ZN(n10240) );
  INV_X1 U10231 ( .A(n9335), .ZN(n9313) );
  INV_X1 U10232 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U10233 ( .A1(n8742), .A2(n11441), .ZN(n9480) );
  INV_X1 U10234 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U10235 ( .A1(n6546), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U10236 ( .A1(n11319), .A2(n11318), .ZN(n11321) );
  OR2_X1 U10237 ( .A1(n12358), .A2(n12357), .ZN(n12361) );
  INV_X1 U10238 ( .A(n11432), .ZN(n11429) );
  NAND2_X1 U10239 ( .A1(n7916), .A2(n12028), .ZN(n7917) );
  NOR2_X1 U10240 ( .A1(n13008), .A2(n8024), .ZN(n8025) );
  AND2_X1 U10241 ( .A1(n12752), .A2(n9412), .ZN(n11532) );
  OR2_X1 U10242 ( .A1(n10879), .A2(n8534), .ZN(n9419) );
  INV_X1 U10243 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10244 ( .A1(n10524), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8173) );
  INV_X1 U10245 ( .A(n8112), .ZN(n8111) );
  INV_X1 U10246 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9882) );
  INV_X1 U10247 ( .A(n14159), .ZN(n14160) );
  INV_X1 U10248 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n14345) );
  AND2_X1 U10249 ( .A1(n10216), .A2(n10215), .ZN(n10217) );
  NAND2_X1 U10250 ( .A1(n10307), .A2(n12392), .ZN(n10124) );
  INV_X1 U10251 ( .A(n11604), .ZN(n10164) );
  NAND2_X1 U10252 ( .A1(n9313), .A2(n9337), .ZN(n9329) );
  INV_X1 U10253 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9009) );
  OR2_X1 U10254 ( .A1(n10531), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9546) );
  OR2_X1 U10255 ( .A1(n10531), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9534) );
  OAI21_X1 U10256 ( .B1(n6545), .B2(n8068), .A(n8610), .ZN(n8611) );
  NAND2_X1 U10257 ( .A1(n12361), .A2(n12360), .ZN(n12371) );
  OAI21_X1 U10258 ( .B1(n11421), .B2(n11265), .A(n11264), .ZN(n11280) );
  INV_X1 U10259 ( .A(n12455), .ZN(n12456) );
  INV_X1 U10260 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n12026) );
  AND2_X1 U10261 ( .A1(n11245), .A2(n11179), .ZN(n12764) );
  INV_X1 U10262 ( .A(n12680), .ZN(n8561) );
  NAND2_X1 U10263 ( .A1(n12658), .A2(n12651), .ZN(n11817) );
  INV_X1 U10264 ( .A(n12613), .ZN(n12579) );
  OR2_X1 U10265 ( .A1(n13411), .A2(n13180), .ZN(n12728) );
  NOR2_X1 U10266 ( .A1(n8568), .A2(n7852), .ZN(n8569) );
  INV_X1 U10267 ( .A(n11645), .ZN(n12595) );
  AND2_X1 U10268 ( .A1(n11235), .A2(n7950), .ZN(n11245) );
  AND2_X1 U10269 ( .A1(n8219), .A2(n8203), .ZN(n8205) );
  INV_X1 U10270 ( .A(n13894), .ZN(n13733) );
  OR2_X1 U10271 ( .A1(n10096), .A2(n10095), .ZN(n13632) );
  INV_X1 U10272 ( .A(n11696), .ZN(n13877) );
  OR2_X1 U10273 ( .A1(n14031), .A2(n10089), .ZN(n9991) );
  INV_X1 U10274 ( .A(n14211), .ZN(n13968) );
  INV_X1 U10275 ( .A(n14257), .ZN(n14098) );
  AND2_X1 U10276 ( .A1(n13884), .A2(n13877), .ZN(n10574) );
  NAND2_X1 U10277 ( .A1(n10977), .A2(n10976), .ZN(n10979) );
  OR2_X1 U10278 ( .A1(n13861), .A2(n6614), .ZN(n14189) );
  OR2_X1 U10279 ( .A1(n12125), .A2(n12109), .ZN(n10410) );
  OR2_X1 U10280 ( .A1(n10075), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n10054) );
  AND2_X1 U10281 ( .A1(n10338), .A2(n14515), .ZN(n10326) );
  NAND2_X1 U10282 ( .A1(n10126), .A2(n10134), .ZN(n10127) );
  NAND2_X1 U10283 ( .A1(n9025), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9026) );
  NAND2_X1 U10284 ( .A1(n10208), .A2(n10209), .ZN(n10210) );
  NAND2_X1 U10285 ( .A1(n10165), .A2(n10164), .ZN(n11601) );
  INV_X1 U10286 ( .A(n9317), .ZN(n9238) );
  INV_X1 U10287 ( .A(n9257), .ZN(n9315) );
  INV_X1 U10288 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14572) );
  INV_X1 U10289 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15556) );
  INV_X1 U10290 ( .A(n15244), .ZN(n14650) );
  INV_X1 U10291 ( .A(n8984), .ZN(n14731) );
  NAND2_X1 U10292 ( .A1(n9546), .A2(n10553), .ZN(n11297) );
  AND2_X1 U10294 ( .A1(n10538), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10408) );
  NAND2_X1 U10295 ( .A1(n9295), .A2(n9282), .ZN(n9285) );
  INV_X1 U10296 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8711) );
  OR2_X1 U10297 ( .A1(n11247), .A2(n11246), .ZN(n11251) );
  OR2_X1 U10298 ( .A1(n7869), .A2(n12286), .ZN(n11235) );
  NAND2_X1 U10299 ( .A1(n8473), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8058) );
  INV_X1 U10300 ( .A(n15467), .ZN(n13007) );
  AND2_X1 U10301 ( .A1(n8037), .A2(n7987), .ZN(n13090) );
  OR2_X1 U10302 ( .A1(n13214), .A2(n13254), .ZN(n13365) );
  INV_X1 U10303 ( .A(n11817), .ZN(n12597) );
  AND2_X1 U10304 ( .A1(n11385), .A2(n12579), .ZN(n12761) );
  INV_X1 U10305 ( .A(n12761), .ZN(n15514) );
  INV_X1 U10306 ( .A(n13391), .ZN(n13383) );
  INV_X1 U10307 ( .A(n12691), .ZN(n13303) );
  INV_X1 U10308 ( .A(n15492), .ZN(n15504) );
  OR2_X1 U10309 ( .A1(n15511), .A2(n6716), .ZN(n15537) );
  OR2_X1 U10310 ( .A1(n11247), .A2(n8537), .ZN(n8543) );
  INV_X1 U10311 ( .A(n15512), .ZN(n13374) );
  NOR2_X1 U10312 ( .A1(n10880), .A2(n13472), .ZN(n10887) );
  INV_X1 U10313 ( .A(n13632), .ZN(n13550) );
  INV_X1 U10314 ( .A(n13599), .ZN(n13634) );
  OR2_X1 U10315 ( .A1(n13989), .A2(n10089), .ZN(n10006) );
  INV_X1 U10316 ( .A(n10578), .ZN(n10589) );
  AND2_X1 U10317 ( .A1(n10574), .A2(n10088), .ZN(n14106) );
  AND2_X1 U10318 ( .A1(n11668), .A2(n14152), .ZN(n14194) );
  INV_X1 U10319 ( .A(n15431), .ZN(n10684) );
  INV_X1 U10320 ( .A(n14308), .ZN(n15453) );
  OR2_X1 U10321 ( .A1(n13642), .A2(n10080), .ZN(n14301) );
  AND2_X1 U10322 ( .A1(n10685), .A2(n14301), .ZN(n14319) );
  AND2_X1 U10323 ( .A1(n15433), .A2(n10683), .ZN(n10958) );
  AND2_X1 U10324 ( .A1(n10061), .A2(n10411), .ZN(n15427) );
  AND2_X1 U10325 ( .A1(n9864), .A2(n9898), .ZN(n12141) );
  OR2_X1 U10326 ( .A1(n10335), .A2(n10853), .ZN(n14458) );
  INV_X1 U10327 ( .A(n14528), .ZN(n14539) );
  INV_X1 U10328 ( .A(n14714), .ZN(n14708) );
  INV_X1 U10329 ( .A(n14709), .ZN(n14653) );
  INV_X1 U10330 ( .A(n14712), .ZN(n14677) );
  XNOR2_X1 U10331 ( .A(n14765), .B(n9509), .ZN(n14761) );
  AND3_X1 U10332 ( .A1(n14959), .A2(n15331), .A3(n14979), .ZN(n15076) );
  NAND2_X1 U10333 ( .A1(n9517), .A2(n9516), .ZN(n15331) );
  INV_X1 U10334 ( .A(n15265), .ZN(n15289) );
  INV_X1 U10335 ( .A(n14953), .ZN(n14990) );
  INV_X1 U10336 ( .A(n15348), .ZN(n9548) );
  INV_X1 U10337 ( .A(n15331), .ZN(n15276) );
  INV_X1 U10338 ( .A(n15100), .ZN(n15339) );
  AND2_X1 U10339 ( .A1(n9022), .A2(n9034), .ZN(n12196) );
  AND2_X1 U10340 ( .A1(n8040), .A2(n8039), .ZN(n15467) );
  INV_X1 U10341 ( .A(n12958), .ZN(n12926) );
  AND2_X1 U10342 ( .A1(n11251), .A2(n11250), .ZN(n12960) );
  OR2_X1 U10343 ( .A1(n11235), .A2(n13472), .ZN(n12966) );
  MUX2_X1 U10344 ( .A(n8038), .B(n12966), .S(n12763), .Z(n13088) );
  INV_X1 U10345 ( .A(n13095), .ZN(n13030) );
  INV_X1 U10346 ( .A(n13100), .ZN(n13046) );
  NAND2_X1 U10347 ( .A1(n15500), .A2(n15477), .ZN(n13327) );
  NAND2_X1 U10348 ( .A1(n11536), .A2(n12761), .ZN(n15486) );
  INV_X1 U10349 ( .A(n10400), .ZN(n10401) );
  NAND2_X1 U10350 ( .A1(n15549), .A2(n15537), .ZN(n13386) );
  NAND2_X1 U10351 ( .A1(n15540), .A2(n15537), .ZN(n13461) );
  AND2_X1 U10352 ( .A1(n8543), .A2(n8542), .ZN(n15539) );
  AND2_X1 U10353 ( .A1(n8524), .A2(n8523), .ZN(n13471) );
  INV_X1 U10354 ( .A(SI_16_), .ZN(n11077) );
  INV_X1 U10355 ( .A(SI_13_), .ZN(n10573) );
  INV_X1 U10356 ( .A(n13480), .ZN(n13495) );
  AND2_X1 U10357 ( .A1(n10103), .A2(n10102), .ZN(n10104) );
  NAND2_X1 U10358 ( .A1(n10962), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13599) );
  INV_X1 U10359 ( .A(n13623), .ZN(n13637) );
  INV_X1 U10360 ( .A(n13782), .ZN(n13999) );
  OR2_X1 U10361 ( .A1(n15349), .A2(P2_U3088), .ZN(n15412) );
  INV_X1 U10362 ( .A(n15394), .ZN(n15414) );
  NAND2_X1 U10363 ( .A1(n14135), .A2(n11502), .ZN(n14191) );
  AND2_X2 U10364 ( .A1(n10958), .A2(n10684), .ZN(n15466) );
  AND3_X1 U10365 ( .A1(n15448), .A2(n15447), .A3(n15446), .ZN(n15463) );
  NOR2_X1 U10366 ( .A1(n15434), .A2(n15427), .ZN(n15428) );
  INV_X1 U10367 ( .A(n15428), .ZN(n15429) );
  INV_X1 U10368 ( .A(n10411), .ZN(n12354) );
  INV_X1 U10369 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10820) );
  OR2_X1 U10370 ( .A1(n10328), .A2(n10321), .ZN(n14546) );
  INV_X1 U10371 ( .A(n10365), .ZN(n14551) );
  INV_X1 U10372 ( .A(n11861), .ZN(n14564) );
  AND2_X1 U10373 ( .A1(n14943), .A2(n14942), .ZN(n15066) );
  OR2_X1 U10374 ( .A1(n6538), .A2(n11300), .ZN(n14953) );
  NAND2_X1 U10375 ( .A1(n15348), .A2(n15295), .ZN(n15086) );
  NAND2_X1 U10376 ( .A1(n15342), .A2(n15295), .ZN(n15147) );
  AND2_X2 U10377 ( .A1(n9552), .A2(n9551), .ZN(n15342) );
  NAND2_X1 U10378 ( .A1(n10536), .A2(n10531), .ZN(n15859) );
  OR4_X1 U10379 ( .A1(n10428), .A2(n10427), .A3(n10426), .A4(n10425), .ZN(
        P3_U3194) );
  OAI21_X1 U10380 ( .B1(n9428), .B2(n15546), .A(n9427), .ZN(P3_U3487) );
  NAND2_X1 U10381 ( .A1(n8582), .A2(n8581), .ZN(P3_U3455) );
  NOR2_X1 U10382 ( .A1(P2_U3088), .A2(n10577), .ZN(P2_U3947) );
  INV_X1 U10383 ( .A(n14570), .ZN(P1_U4016) );
  NAND4_X1 U10384 ( .A1(n7164), .A2(n15810), .A3(n7857), .A4(n7739), .ZN(n7863) );
  NAND3_X1 U10385 ( .A1(n7861), .A2(n7860), .A3(n7858), .ZN(n7862) );
  NAND2_X1 U10386 ( .A1(n7866), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7865) );
  MUX2_X1 U10387 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7865), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n7867) );
  NAND2_X1 U10388 ( .A1(n8517), .A2(n8520), .ZN(n7869) );
  NAND2_X1 U10389 ( .A1(n7870), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7871) );
  MUX2_X1 U10390 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7871), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n7873) );
  NAND2_X1 U10391 ( .A1(n7873), .A2(n7872), .ZN(n7957) );
  INV_X1 U10392 ( .A(n7874), .ZN(n7885) );
  OR2_X1 U10393 ( .A1(n7885), .A2(n7875), .ZN(n7918) );
  INV_X1 U10394 ( .A(n7918), .ZN(n7876) );
  NAND2_X1 U10395 ( .A1(n7876), .A2(n15823), .ZN(n7878) );
  NAND2_X1 U10396 ( .A1(n7878), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7877) );
  MUX2_X1 U10397 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7877), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n7879) );
  NAND2_X1 U10398 ( .A1(n7879), .A2(n7926), .ZN(n10567) );
  INV_X1 U10399 ( .A(n10567), .ZN(n7976) );
  INV_X1 U10400 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n13387) );
  AND2_X1 U10401 ( .A1(n7874), .A2(n7886), .ZN(n7909) );
  NAND2_X1 U10402 ( .A1(n7909), .A2(n7880), .ZN(n7883) );
  OAI21_X1 U10403 ( .B1(n7913), .B2(P3_IR_REG_9__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7882) );
  INV_X1 U10404 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7881) );
  XNOR2_X1 U10405 ( .A(n7882), .B(n7881), .ZN(n10529) );
  INV_X1 U10406 ( .A(n10529), .ZN(n12094) );
  INV_X1 U10407 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12306) );
  NAND2_X1 U10408 ( .A1(n7883), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7884) );
  INV_X1 U10409 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n12111) );
  NAND2_X1 U10410 ( .A1(n7885), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7887) );
  XNOR2_X1 U10411 ( .A(n7887), .B(n7886), .ZN(n10445) );
  INV_X1 U10412 ( .A(n11161), .ZN(n7990) );
  INV_X1 U10413 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7890) );
  INV_X1 U10414 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11181) );
  NOR2_X1 U10415 ( .A1(n11181), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U10416 ( .A1(n7964), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7893) );
  INV_X1 U10417 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15541) );
  NAND2_X1 U10418 ( .A1(n7894), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7895) );
  INV_X1 U10419 ( .A(n7898), .ZN(n11093) );
  NAND2_X1 U10420 ( .A1(n7900), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7901) );
  MUX2_X1 U10421 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7901), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7904) );
  INV_X1 U10422 ( .A(n7900), .ZN(n7903) );
  NAND2_X1 U10423 ( .A1(n7903), .A2(n7902), .ZN(n7905) );
  XNOR2_X1 U10424 ( .A(n8004), .B(P3_REG1_REG_4__SCAN_IN), .ZN(n11094) );
  NAND2_X1 U10425 ( .A1(n7905), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7906) );
  XNOR2_X1 U10426 ( .A(n10445), .B(P3_REG1_REG_6__SCAN_IN), .ZN(n11374) );
  INV_X1 U10427 ( .A(n7909), .ZN(n7910) );
  NAND2_X1 U10428 ( .A1(n7910), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7911) );
  XNOR2_X1 U10429 ( .A(n7911), .B(P3_IR_REG_7__SCAN_IN), .ZN(n10454) );
  INV_X1 U10430 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15571) );
  XNOR2_X1 U10431 ( .A(n11838), .B(P3_REG1_REG_8__SCAN_IN), .ZN(n11839) );
  NAND2_X1 U10432 ( .A1(n7913), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7915) );
  INV_X1 U10433 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7914) );
  XNOR2_X1 U10434 ( .A(n7915), .B(n7914), .ZN(n12028) );
  INV_X1 U10435 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n12066) );
  INV_X1 U10436 ( .A(n7917), .ZN(n12097) );
  XNOR2_X1 U10437 ( .A(n10529), .B(n12306), .ZN(n12096) );
  NAND2_X1 U10438 ( .A1(n7918), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7919) );
  XNOR2_X1 U10439 ( .A(n7919), .B(n15823), .ZN(n12982) );
  INV_X1 U10440 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n15739) );
  XNOR2_X1 U10441 ( .A(n10567), .B(n13387), .ZN(n10416) );
  NAND2_X1 U10442 ( .A1(n7926), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7922) );
  INV_X1 U10443 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n15595) );
  XNOR2_X1 U10444 ( .A(n7922), .B(n15595), .ZN(n12998) );
  INV_X1 U10445 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15767) );
  INV_X1 U10446 ( .A(n7925), .ZN(n13021) );
  NAND2_X1 U10447 ( .A1(n7929), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7927) );
  XNOR2_X1 U10448 ( .A(n7927), .B(P3_IR_REG_14__SCAN_IN), .ZN(n13013) );
  INV_X1 U10449 ( .A(n13013), .ZN(n10858) );
  NAND2_X1 U10450 ( .A1(n10858), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8021) );
  INV_X1 U10451 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13380) );
  NAND2_X1 U10452 ( .A1(n13013), .A2(n13380), .ZN(n7928) );
  AND2_X1 U10453 ( .A1(n8021), .A2(n7928), .ZN(n13022) );
  INV_X1 U10454 ( .A(n7929), .ZN(n7931) );
  INV_X1 U10455 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10456 ( .A1(n7931), .A2(n7930), .ZN(n7933) );
  NAND2_X1 U10457 ( .A1(n7933), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7932) );
  MUX2_X1 U10458 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7932), .S(
        P3_IR_REG_15__SCAN_IN), .Z(n7936) );
  INV_X1 U10459 ( .A(n7933), .ZN(n7935) );
  INV_X1 U10460 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U10461 ( .A1(n7935), .A2(n7934), .ZN(n7940) );
  NAND2_X1 U10462 ( .A1(n7940), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7938) );
  XNOR2_X1 U10463 ( .A(n7938), .B(P3_IR_REG_16__SCAN_IN), .ZN(n8296) );
  INV_X1 U10464 ( .A(n8296), .ZN(n13061) );
  NAND2_X1 U10465 ( .A1(n13061), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U10466 ( .A1(n7942), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7941) );
  XNOR2_X1 U10467 ( .A(n7941), .B(P3_IR_REG_17__SCAN_IN), .ZN(n8309) );
  INV_X1 U10468 ( .A(n8309), .ZN(n13073) );
  OAI21_X1 U10469 ( .B1(n7942), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7943) );
  XNOR2_X1 U10470 ( .A(n7943), .B(P3_IR_REG_18__SCAN_IN), .ZN(n8325) );
  INV_X1 U10471 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n8031) );
  OR2_X1 U10472 ( .A1(n8325), .A2(n8031), .ZN(n7945) );
  NAND2_X1 U10473 ( .A1(n8325), .A2(n8031), .ZN(n7944) );
  NAND2_X1 U10474 ( .A1(n7945), .A2(n7944), .ZN(n13097) );
  NAND2_X1 U10475 ( .A1(n7946), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7947) );
  MUX2_X1 U10476 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7947), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n7948) );
  XNOR2_X1 U10477 ( .A(n12579), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n8033) );
  INV_X1 U10478 ( .A(n11245), .ZN(n7951) );
  INV_X1 U10479 ( .A(n7957), .ZN(n11232) );
  NAND2_X1 U10480 ( .A1(n11232), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12768) );
  NAND2_X1 U10481 ( .A1(n7951), .A2(n12768), .ZN(n8040) );
  NAND2_X1 U10482 ( .A1(n8501), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7953) );
  INV_X1 U10483 ( .A(n7954), .ZN(n7955) );
  NAND2_X1 U10484 ( .A1(n7955), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7956) );
  NAND2_X1 U10485 ( .A1(n12752), .A2(n7957), .ZN(n7962) );
  NAND2_X1 U10486 ( .A1(n7962), .A2(n7080), .ZN(n8039) );
  INV_X1 U10487 ( .A(n8039), .ZN(n7963) );
  AND2_X1 U10488 ( .A1(n8040), .A2(n7963), .ZN(n8037) );
  INV_X1 U10489 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n13321) );
  INV_X1 U10490 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12270) );
  INV_X1 U10491 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n12071) );
  INV_X1 U10492 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11539) );
  NOR2_X1 U10493 ( .A1(n11539), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n7965) );
  NAND2_X1 U10494 ( .A1(n7964), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7966) );
  OAI21_X1 U10495 ( .B1(n11197), .B2(n7965), .A(n7966), .ZN(n11188) );
  INV_X1 U10496 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11189) );
  INV_X1 U10497 ( .A(n7966), .ZN(n7967) );
  NOR2_X1 U10498 ( .A1(n11187), .A2(n7967), .ZN(n11145) );
  XNOR2_X1 U10499 ( .A(n8004), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n11098) );
  XNOR2_X1 U10500 ( .A(n10445), .B(P3_REG2_REG_6__SCAN_IN), .ZN(n11369) );
  XNOR2_X1 U10501 ( .A(n11838), .B(P3_REG2_REG_8__SCAN_IN), .ZN(n11831) );
  INV_X1 U10502 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12078) );
  XNOR2_X1 U10503 ( .A(n10529), .B(n12270), .ZN(n12087) );
  NAND2_X1 U10504 ( .A1(n7974), .A2(n12087), .ZN(n12091) );
  OAI21_X1 U10505 ( .B1(n7976), .B2(n13321), .A(n10422), .ZN(n7977) );
  NAND2_X1 U10506 ( .A1(n7977), .A2(n12998), .ZN(n13015) );
  NAND2_X1 U10507 ( .A1(n10858), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7979) );
  INV_X1 U10508 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13297) );
  NAND2_X1 U10509 ( .A1(n13013), .A2(n13297), .ZN(n7978) );
  NAND2_X1 U10510 ( .A1(n7979), .A2(n7978), .ZN(n13016) );
  INV_X1 U10511 ( .A(n7979), .ZN(n8022) );
  INV_X1 U10512 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13285) );
  XNOR2_X1 U10513 ( .A(n8296), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n13049) );
  INV_X1 U10514 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13276) );
  OR2_X1 U10515 ( .A1(n8296), .A2(n13276), .ZN(n7981) );
  NAND2_X1 U10516 ( .A1(n13054), .A2(n7981), .ZN(n7982) );
  NAND2_X1 U10517 ( .A1(n7982), .A2(n13073), .ZN(n13081) );
  INV_X1 U10518 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13250) );
  OR2_X1 U10519 ( .A1(n8325), .A2(n13250), .ZN(n7985) );
  NAND2_X1 U10520 ( .A1(n8325), .A2(n13250), .ZN(n7983) );
  AND2_X1 U10521 ( .A1(n7985), .A2(n7983), .ZN(n13079) );
  INV_X1 U10522 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13236) );
  XNOR2_X1 U10523 ( .A(n12613), .B(n13236), .ZN(n8034) );
  OR2_X1 U10524 ( .A1(n7986), .A2(n8019), .ZN(n8507) );
  INV_X1 U10525 ( .A(n8507), .ZN(n7987) );
  MUX2_X1 U10526 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n8019), .Z(n8018) );
  INV_X4 U10527 ( .A(n6541), .ZN(n13489) );
  MUX2_X1 U10528 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13489), .Z(n8017) );
  INV_X1 U10529 ( .A(n10445), .ZN(n11379) );
  MUX2_X1 U10530 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13489), .Z(n8008) );
  INV_X1 U10531 ( .A(n8008), .ZN(n8009) );
  INV_X1 U10532 ( .A(n8004), .ZN(n11106) );
  MUX2_X1 U10533 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n8019), .Z(n8005) );
  INV_X1 U10534 ( .A(n8005), .ZN(n8006) );
  NAND2_X1 U10535 ( .A1(n7989), .A2(n11161), .ZN(n11043) );
  INV_X1 U10536 ( .A(n7989), .ZN(n7991) );
  NAND2_X1 U10537 ( .A1(n7991), .A2(n7990), .ZN(n7992) );
  AND2_X1 U10538 ( .A1(n11043), .A2(n7992), .ZN(n11153) );
  INV_X1 U10539 ( .A(n11197), .ZN(n7994) );
  OAI21_X1 U10540 ( .B1(n7995), .B2(n7994), .A(n7997), .ZN(n11185) );
  NAND2_X1 U10541 ( .A1(n8019), .A2(n11181), .ZN(n7996) );
  NAND2_X1 U10542 ( .A1(n11288), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11184) );
  INV_X1 U10543 ( .A(n7997), .ZN(n11154) );
  INV_X1 U10544 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n15480) );
  INV_X1 U10545 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11652) );
  MUX2_X1 U10546 ( .A(n15480), .B(n11652), .S(n8019), .Z(n7999) );
  NAND2_X1 U10547 ( .A1(n7999), .A2(n10451), .ZN(n8002) );
  INV_X1 U10548 ( .A(n7999), .ZN(n8000) );
  INV_X1 U10549 ( .A(n10451), .ZN(n11048) );
  NAND2_X1 U10550 ( .A1(n8000), .A2(n11048), .ZN(n8001) );
  NAND2_X1 U10551 ( .A1(n8002), .A2(n8001), .ZN(n11042) );
  INV_X1 U10552 ( .A(n8002), .ZN(n8003) );
  XNOR2_X1 U10553 ( .A(n8005), .B(n8004), .ZN(n11091) );
  INV_X1 U10554 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15795) );
  INV_X1 U10555 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15544) );
  MUX2_X1 U10556 ( .A(n15795), .B(n15544), .S(n13489), .Z(n8007) );
  NOR2_X1 U10557 ( .A1(n8007), .A2(n11215), .ZN(n11225) );
  NOR2_X1 U10558 ( .A1(n11224), .A2(n11225), .ZN(n11223) );
  AND2_X1 U10559 ( .A1(n8007), .A2(n11215), .ZN(n11227) );
  NOR2_X1 U10560 ( .A1(n11223), .A2(n11227), .ZN(n11367) );
  XNOR2_X1 U10561 ( .A(n8008), .B(n10445), .ZN(n11366) );
  MUX2_X1 U10562 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13489), .Z(n8010) );
  XOR2_X1 U10563 ( .A(n10454), .B(n8010), .Z(n11631) );
  MUX2_X1 U10564 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13489), .Z(n8011) );
  XNOR2_X1 U10565 ( .A(n8011), .B(n11838), .ZN(n11827) );
  INV_X1 U10566 ( .A(n8011), .ZN(n8012) );
  MUX2_X1 U10567 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13489), .Z(n8013) );
  XNOR2_X1 U10568 ( .A(n8013), .B(n12028), .ZN(n12023) );
  MUX2_X1 U10569 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n8019), .Z(n8014) );
  XOR2_X1 U10570 ( .A(n10529), .B(n8014), .Z(n12083) );
  INV_X1 U10571 ( .A(n8014), .ZN(n8015) );
  MUX2_X1 U10572 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13489), .Z(n8016) );
  XNOR2_X1 U10573 ( .A(n8016), .B(n12982), .ZN(n12977) );
  XNOR2_X1 U10574 ( .A(n8017), .B(n10567), .ZN(n10415) );
  XOR2_X1 U10575 ( .A(n12998), .B(n8018), .Z(n12994) );
  NAND2_X1 U10576 ( .A1(n12995), .A2(n12994), .ZN(n12993) );
  OAI21_X1 U10577 ( .B1(n8018), .B2(n12998), .A(n12993), .ZN(n13009) );
  INV_X1 U10578 ( .A(n13022), .ZN(n8020) );
  MUX2_X1 U10579 ( .A(n8020), .B(n13016), .S(n6541), .Z(n13010) );
  INV_X1 U10580 ( .A(n8021), .ZN(n8023) );
  MUX2_X1 U10581 ( .A(n8023), .B(n8022), .S(n6541), .Z(n8024) );
  XNOR2_X1 U10582 ( .A(n8025), .B(n8280), .ZN(n13032) );
  INV_X1 U10583 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13377) );
  MUX2_X1 U10584 ( .A(n13285), .B(n13377), .S(n13489), .Z(n13031) );
  OR2_X2 U10585 ( .A1(n13032), .A2(n13031), .ZN(n13037) );
  MUX2_X1 U10586 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n13489), .Z(n8026) );
  XNOR2_X1 U10587 ( .A(n8296), .B(n8026), .ZN(n13056) );
  INV_X1 U10588 ( .A(n8026), .ZN(n8027) );
  MUX2_X1 U10589 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13489), .Z(n8029) );
  XNOR2_X1 U10590 ( .A(n8309), .B(n8029), .ZN(n13068) );
  INV_X1 U10591 ( .A(n8029), .ZN(n8030) );
  INV_X1 U10592 ( .A(n8325), .ZN(n13087) );
  MUX2_X1 U10593 ( .A(n13250), .B(n8031), .S(n13489), .Z(n13093) );
  NAND2_X1 U10594 ( .A1(n13094), .A2(n13093), .ZN(n13092) );
  OAI21_X1 U10595 ( .B1(n8032), .B2(n13087), .A(n13092), .ZN(n8036) );
  MUX2_X1 U10596 ( .A(n8034), .B(n8033), .S(n13489), .Z(n8035) );
  INV_X1 U10597 ( .A(n8037), .ZN(n8038) );
  INV_X1 U10598 ( .A(n7986), .ZN(n12763) );
  AND2_X1 U10599 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12824) );
  AOI21_X1 U10600 ( .B1(n15467), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n12824), 
        .ZN(n8041) );
  OAI21_X1 U10601 ( .B1(n13088), .B2(n12613), .A(n8041), .ZN(n8042) );
  INV_X1 U10602 ( .A(n8042), .ZN(n8043) );
  XNOR2_X2 U10603 ( .A(n8045), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8054) );
  INV_X1 U10604 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n13474) );
  NAND2_X1 U10605 ( .A1(n8046), .A2(n13474), .ZN(n8049) );
  INV_X1 U10606 ( .A(n8049), .ZN(n8047) );
  NAND2_X1 U10607 ( .A1(n8047), .A2(n13475), .ZN(n8052) );
  XNOR2_X1 U10608 ( .A(P3_IR_REG_31__SCAN_IN), .B(P3_IR_REG_30__SCAN_IN), .ZN(
        n8048) );
  OAI211_X2 U10609 ( .C1(n8053), .C2(n8052), .A(n8051), .B(n8050), .ZN(n12770)
         );
  NAND2_X1 U10610 ( .A1(n6539), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8059) );
  NAND2_X2 U10611 ( .A1(n8054), .A2(n12770), .ZN(n12562) );
  INV_X1 U10612 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11284) );
  OR2_X1 U10613 ( .A1(n8510), .A2(n11284), .ZN(n8057) );
  NAND2_X1 U10614 ( .A1(n13484), .A2(n12770), .ZN(n8101) );
  INV_X1 U10615 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15598) );
  OR2_X1 U10616 ( .A1(n8101), .A2(n15598), .ZN(n8056) );
  NAND4_X4 U10617 ( .A1(n8059), .A2(n8058), .A3(n8057), .A4(n8056), .ZN(n12974) );
  OR2_X1 U10618 ( .A1(n8508), .A2(n11197), .ZN(n8064) );
  XNOR2_X1 U10619 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n8080) );
  NAND2_X1 U10620 ( .A1(n10545), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8079) );
  XNOR2_X1 U10621 ( .A(n8080), .B(n8079), .ZN(n10441) );
  NAND2_X1 U10622 ( .A1(n10441), .A2(n9277), .ZN(n8061) );
  INV_X1 U10623 ( .A(SI_1_), .ZN(n10440) );
  NAND2_X1 U10624 ( .A1(n6545), .A2(n10440), .ZN(n8060) );
  AND2_X1 U10625 ( .A1(n8061), .A2(n8060), .ZN(n8062) );
  OAI21_X1 U10626 ( .B1(n12763), .B2(n6541), .A(n8062), .ZN(n8063) );
  XNOR2_X2 U10627 ( .A(n12974), .B(n15513), .ZN(n11276) );
  INV_X1 U10628 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n11254) );
  INV_X1 U10629 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8065) );
  OR2_X1 U10630 ( .A1(n8101), .A2(n8065), .ZN(n8067) );
  OR2_X1 U10631 ( .A1(n6535), .A2(n11539), .ZN(n8066) );
  INV_X1 U10632 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n8072) );
  INV_X1 U10633 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8068) );
  NAND2_X1 U10634 ( .A1(n8068), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U10635 ( .A1(n8079), .A2(n8069), .ZN(n8070) );
  NAND2_X1 U10636 ( .A1(n9277), .A2(n8070), .ZN(n8071) );
  AND2_X1 U10637 ( .A1(n8071), .A2(n9618), .ZN(n10439) );
  MUX2_X1 U10638 ( .A(n8072), .B(n10439), .S(n8508), .Z(n11483) );
  NAND2_X1 U10639 ( .A1(n15505), .A2(n6872), .ZN(n11279) );
  NAND2_X1 U10640 ( .A1(n11276), .A2(n11279), .ZN(n8074) );
  INV_X1 U10641 ( .A(n15513), .ZN(n11267) );
  OR2_X1 U10642 ( .A1(n12974), .A2(n11267), .ZN(n8073) );
  NAND2_X1 U10643 ( .A1(n8074), .A2(n8073), .ZN(n15487) );
  NAND2_X1 U10644 ( .A1(n8392), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8078) );
  OR2_X1 U10645 ( .A1(n12562), .A2(n7477), .ZN(n8077) );
  INV_X1 U10646 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11274) );
  OR2_X1 U10647 ( .A1(n8510), .A2(n11274), .ZN(n8076) );
  OR2_X1 U10648 ( .A1(n6534), .A2(n6899), .ZN(n8075) );
  INV_X1 U10649 ( .A(n8079), .ZN(n8081) );
  INV_X1 U10650 ( .A(n8095), .ZN(n8083) );
  XNOR2_X1 U10651 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8082) );
  XNOR2_X1 U10652 ( .A(n8083), .B(n8082), .ZN(n10442) );
  OR2_X1 U10653 ( .A1(n8177), .A2(n10442), .ZN(n8085) );
  OAI211_X1 U10654 ( .C1(n11161), .C2(n8508), .A(n8085), .B(n8084), .ZN(n15497) );
  NAND2_X1 U10655 ( .A1(n15506), .A2(n15497), .ZN(n8545) );
  NAND2_X1 U10656 ( .A1(n15487), .A2(n11643), .ZN(n8087) );
  INV_X1 U10657 ( .A(n15497), .ZN(n11262) );
  OR2_X1 U10658 ( .A1(n15506), .A2(n11262), .ZN(n8086) );
  NAND2_X1 U10659 ( .A1(n8473), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8093) );
  OR2_X1 U10660 ( .A1(n8510), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8092) );
  INV_X1 U10661 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8088) );
  OR2_X1 U10662 ( .A1(n8101), .A2(n8088), .ZN(n8091) );
  OR2_X1 U10663 ( .A1(n6534), .A2(n15480), .ZN(n8090) );
  NAND2_X1 U10664 ( .A1(n10491), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10665 ( .A1(n8095), .A2(n8094), .ZN(n8097) );
  NAND2_X1 U10666 ( .A1(n10518), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8096) );
  XNOR2_X1 U10667 ( .A(n10489), .B(P1_DATAO_REG_3__SCAN_IN), .ZN(n8098) );
  XNOR2_X1 U10668 ( .A(n8109), .B(n8098), .ZN(n10452) );
  NAND2_X1 U10669 ( .A1(n8473), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8106) );
  INV_X1 U10670 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n15475) );
  OR2_X1 U10671 ( .A1(n6535), .A2(n15475), .ZN(n8105) );
  AND2_X1 U10672 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8100) );
  NOR2_X1 U10673 ( .A1(n15561), .A2(n8100), .ZN(n15470) );
  OR2_X1 U10674 ( .A1(n8510), .A2(n15470), .ZN(n8104) );
  INV_X1 U10675 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8102) );
  OR2_X1 U10676 ( .A1(n8101), .A2(n8102), .ZN(n8103) );
  OR2_X1 U10677 ( .A1(n12569), .A2(SI_4_), .ZN(n8117) );
  NAND2_X1 U10678 ( .A1(n10487), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8107) );
  NAND2_X1 U10679 ( .A1(n10495), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U10680 ( .A1(n8126), .A2(n8110), .ZN(n8112) );
  NAND2_X1 U10681 ( .A1(n8113), .A2(n8112), .ZN(n8114) );
  AND2_X1 U10682 ( .A1(n8127), .A2(n8114), .ZN(n10449) );
  OR2_X1 U10683 ( .A1(n6542), .A2(n10449), .ZN(n8116) );
  OR2_X1 U10684 ( .A1(n8508), .A2(n11106), .ZN(n8115) );
  OR2_X1 U10685 ( .A1(n12973), .A2(n11436), .ZN(n8118) );
  AND2_X1 U10686 ( .A1(n7378), .A2(n11659), .ZN(n11657) );
  AOI22_X1 U10687 ( .A1(n11657), .A2(n8118), .B1(n11436), .B2(n12973), .ZN(
        n8119) );
  NAND2_X1 U10688 ( .A1(n6539), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8125) );
  INV_X1 U10689 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15547) );
  OR2_X1 U10690 ( .A1(n12562), .A2(n15547), .ZN(n8124) );
  NAND2_X1 U10691 ( .A1(n8135), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8120) );
  AND2_X1 U10692 ( .A1(n8149), .A2(n8120), .ZN(n11824) );
  OR2_X1 U10693 ( .A1(n8510), .A2(n11824), .ZN(n8123) );
  INV_X1 U10694 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8121) );
  OR2_X1 U10695 ( .A1(n8101), .A2(n8121), .ZN(n8122) );
  NAND2_X1 U10696 ( .A1(n10493), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8128) );
  XNOR2_X1 U10697 ( .A(n8158), .B(n8156), .ZN(n10444) );
  OR2_X1 U10698 ( .A1(n6542), .A2(n10444), .ZN(n8132) );
  INV_X1 U10699 ( .A(SI_6_), .ZN(n10446) );
  OR2_X1 U10700 ( .A1(n8508), .A2(n10445), .ZN(n8130) );
  NAND2_X1 U10701 ( .A1(n12971), .A2(n12216), .ZN(n12651) );
  NAND2_X1 U10702 ( .A1(n8392), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8139) );
  OR2_X1 U10703 ( .A1(n6534), .A2(n15795), .ZN(n8138) );
  OR2_X1 U10704 ( .A1(n15561), .A2(n8133), .ZN(n8134) );
  AND2_X1 U10705 ( .A1(n8135), .A2(n8134), .ZN(n11771) );
  OR2_X1 U10706 ( .A1(n8510), .A2(n11771), .ZN(n8136) );
  INV_X1 U10707 ( .A(n8140), .ZN(n8143) );
  INV_X1 U10708 ( .A(n8141), .ZN(n8142) );
  NAND2_X1 U10709 ( .A1(n8143), .A2(n8142), .ZN(n8145) );
  AND2_X1 U10710 ( .A1(n8145), .A2(n8144), .ZN(n10447) );
  OR2_X1 U10711 ( .A1(n12972), .A2(n12868), .ZN(n8146) );
  INV_X1 U10712 ( .A(n8146), .ZN(n11819) );
  NAND2_X1 U10713 ( .A1(n12972), .A2(n11770), .ZN(n8553) );
  NAND2_X1 U10714 ( .A1(n12647), .A2(n8553), .ZN(n12645) );
  NOR2_X1 U10715 ( .A1(n11819), .A2(n12645), .ZN(n8147) );
  INV_X1 U10716 ( .A(n12216), .ZN(n12932) );
  AOI22_X1 U10717 ( .A1(n8147), .A2(n11817), .B1(n12971), .B2(n12932), .ZN(
        n8148) );
  NAND2_X1 U10718 ( .A1(n6539), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8155) );
  OR2_X1 U10719 ( .A1(n12562), .A2(n15571), .ZN(n8154) );
  AND2_X1 U10720 ( .A1(n8149), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8150) );
  NOR2_X1 U10721 ( .A1(n8165), .A2(n8150), .ZN(n12778) );
  OR2_X1 U10722 ( .A1(n8510), .A2(n12778), .ZN(n8153) );
  INV_X1 U10723 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8151) );
  OR2_X1 U10724 ( .A1(n8101), .A2(n8151), .ZN(n8152) );
  NAND4_X1 U10725 ( .A1(n8155), .A2(n8154), .A3(n8153), .A4(n8152), .ZN(n12970) );
  NAND2_X1 U10726 ( .A1(n10526), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U10727 ( .A1(n8173), .A2(n8159), .ZN(n8174) );
  INV_X1 U10728 ( .A(n8174), .ZN(n8160) );
  XNOR2_X1 U10729 ( .A(n8175), .B(n8160), .ZN(n10455) );
  OR2_X1 U10730 ( .A1(n10455), .A2(n6542), .ZN(n8162) );
  OR2_X1 U10731 ( .A1(n12569), .A2(SI_7_), .ZN(n8161) );
  OAI211_X1 U10732 ( .C1(n10454), .C2(n7080), .A(n8162), .B(n8161), .ZN(n12000) );
  INV_X1 U10733 ( .A(n12000), .ZN(n12777) );
  INV_X1 U10734 ( .A(n12656), .ZN(n11849) );
  NAND2_X1 U10735 ( .A1(n12777), .A2(n12970), .ZN(n8163) );
  NAND2_X1 U10736 ( .A1(n6539), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8172) );
  OR2_X1 U10737 ( .A1(n12562), .A2(n12111), .ZN(n8171) );
  NOR2_X1 U10738 ( .A1(n8165), .A2(n8164), .ZN(n8166) );
  OR2_X1 U10739 ( .A1(n8190), .A2(n8166), .ZN(n12835) );
  INV_X1 U10740 ( .A(n12835), .ZN(n8167) );
  OR2_X1 U10741 ( .A1(n8510), .A2(n8167), .ZN(n8170) );
  INV_X1 U10742 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8168) );
  OR2_X1 U10743 ( .A1(n12563), .A2(n8168), .ZN(n8169) );
  NAND4_X1 U10744 ( .A1(n8172), .A2(n8171), .A3(n8170), .A4(n8169), .ZN(n12969) );
  INV_X1 U10745 ( .A(n12969), .ZN(n8181) );
  XNOR2_X1 U10746 ( .A(n10543), .B(P2_DATAO_REG_8__SCAN_IN), .ZN(n8176) );
  XNOR2_X1 U10747 ( .A(n8184), .B(n8176), .ZN(n10500) );
  INV_X4 U10748 ( .A(n8177), .ZN(n8470) );
  NAND2_X1 U10749 ( .A1(n10500), .A2(n8470), .ZN(n8179) );
  AOI22_X1 U10750 ( .A1(n8342), .A2(SI_8_), .B1(n8341), .B2(n11838), .ZN(n8178) );
  NAND2_X1 U10751 ( .A1(n8181), .A2(n12219), .ZN(n8180) );
  OR2_X1 U10752 ( .A1(n8181), .A2(n12219), .ZN(n8182) );
  NAND2_X1 U10753 ( .A1(n10543), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U10754 ( .A1(n10541), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8185) );
  NAND2_X1 U10755 ( .A1(n8186), .A2(n8185), .ZN(n8201) );
  XNOR2_X1 U10756 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .ZN(n8187) );
  XNOR2_X1 U10757 ( .A(n8201), .B(n8187), .ZN(n10497) );
  NAND2_X1 U10758 ( .A1(n10497), .A2(n8470), .ZN(n8189) );
  AOI22_X1 U10759 ( .A1(n8342), .A2(n10496), .B1(n8341), .B2(n12028), .ZN(
        n8188) );
  NAND2_X1 U10760 ( .A1(n8189), .A2(n8188), .ZN(n12228) );
  NAND2_X1 U10761 ( .A1(n6539), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8195) );
  OR2_X1 U10762 ( .A1(n12562), .A2(n12066), .ZN(n8194) );
  OR2_X1 U10763 ( .A1(n8190), .A2(n12026), .ZN(n8191) );
  AND2_X1 U10764 ( .A1(n8211), .A2(n8191), .ZN(n12079) );
  OR2_X1 U10765 ( .A1(n8510), .A2(n12079), .ZN(n8193) );
  INV_X1 U10766 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n11933) );
  OR2_X1 U10767 ( .A1(n12563), .A2(n11933), .ZN(n8192) );
  NAND4_X1 U10768 ( .A1(n8195), .A2(n8194), .A3(n8193), .A4(n8192), .ZN(n12968) );
  OR2_X1 U10769 ( .A1(n12228), .A2(n12968), .ZN(n12672) );
  NAND2_X1 U10770 ( .A1(n12228), .A2(n12968), .ZN(n12671) );
  INV_X1 U10771 ( .A(n12594), .ZN(n8196) );
  INV_X1 U10772 ( .A(n12968), .ZN(n12230) );
  OR2_X1 U10773 ( .A1(n12228), .A2(n12230), .ZN(n8197) );
  NAND2_X1 U10774 ( .A1(n8198), .A2(n8197), .ZN(n12116) );
  NAND2_X1 U10775 ( .A1(n10548), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8199) );
  OAI21_X1 U10776 ( .B1(n8201), .B2(n8200), .A(n8199), .ZN(n8202) );
  NAND2_X1 U10777 ( .A1(n10569), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8219) );
  NAND2_X1 U10778 ( .A1(n10571), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8203) );
  INV_X1 U10779 ( .A(n8205), .ZN(n8206) );
  NAND2_X1 U10780 ( .A1(n8202), .A2(n8206), .ZN(n8207) );
  NAND2_X1 U10781 ( .A1(n8220), .A2(n8207), .ZN(n10530) );
  NAND2_X1 U10782 ( .A1(n10530), .A2(n8470), .ZN(n8209) );
  AOI22_X1 U10783 ( .A1(n8342), .A2(n10528), .B1(n8341), .B2(n10529), .ZN(
        n8208) );
  NAND2_X1 U10784 ( .A1(n8209), .A2(n8208), .ZN(n12308) );
  NAND2_X1 U10785 ( .A1(n8473), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8216) );
  INV_X1 U10786 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8210) );
  OR2_X1 U10787 ( .A1(n8101), .A2(n8210), .ZN(n8215) );
  NAND2_X1 U10788 ( .A1(n8211), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8212) );
  AND2_X1 U10789 ( .A1(n8224), .A2(n8212), .ZN(n12271) );
  OR2_X1 U10790 ( .A1(n8510), .A2(n12271), .ZN(n8214) );
  OR2_X1 U10791 ( .A1(n6534), .A2(n12270), .ZN(n8213) );
  NAND4_X1 U10792 ( .A1(n8216), .A2(n8215), .A3(n8214), .A4(n8213), .ZN(n12967) );
  OR2_X1 U10793 ( .A1(n12308), .A2(n12967), .ZN(n12673) );
  NAND2_X1 U10794 ( .A1(n12308), .A2(n12967), .ZN(n12674) );
  NAND2_X1 U10795 ( .A1(n12673), .A2(n12674), .ZN(n12680) );
  NAND2_X1 U10796 ( .A1(n12116), .A2(n12680), .ZN(n8218) );
  INV_X1 U10797 ( .A(n12967), .ZN(n12237) );
  OR2_X1 U10798 ( .A1(n12308), .A2(n12237), .ZN(n8217) );
  NAND2_X1 U10799 ( .A1(n8218), .A2(n8217), .ZN(n12275) );
  XNOR2_X1 U10800 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8221) );
  XNOR2_X1 U10801 ( .A(n8233), .B(n8221), .ZN(n10547) );
  NAND2_X1 U10802 ( .A1(n10547), .A2(n8470), .ZN(n8223) );
  AOI22_X1 U10803 ( .A1(n8342), .A2(n10546), .B1(n8341), .B2(n12982), .ZN(
        n8222) );
  NAND2_X1 U10804 ( .A1(n8223), .A2(n8222), .ZN(n12235) );
  NAND2_X1 U10805 ( .A1(n6539), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8229) );
  OR2_X1 U10806 ( .A1(n12562), .A2(n15739), .ZN(n8228) );
  NAND2_X1 U10807 ( .A1(n8224), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8225) );
  AND2_X1 U10808 ( .A1(n8250), .A2(n8225), .ZN(n12311) );
  OR2_X1 U10809 ( .A1(n8510), .A2(n12311), .ZN(n8227) );
  INV_X1 U10810 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n12281) );
  OR2_X1 U10811 ( .A1(n12563), .A2(n12281), .ZN(n8226) );
  NAND4_X1 U10812 ( .A1(n8229), .A2(n8228), .A3(n8227), .A4(n8226), .ZN(n13314) );
  NOR2_X1 U10813 ( .A1(n12235), .A2(n12336), .ZN(n8231) );
  NAND2_X1 U10814 ( .A1(n12235), .A2(n12336), .ZN(n8230) );
  NAND2_X1 U10815 ( .A1(n10700), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8232) );
  NAND2_X1 U10816 ( .A1(n8652), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8234) );
  AND2_X1 U10817 ( .A1(n10818), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8237) );
  NAND2_X1 U10818 ( .A1(n10820), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8236) );
  XNOR2_X1 U10819 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .ZN(n8276) );
  XNOR2_X1 U10820 ( .A(n8279), .B(n8276), .ZN(n10857) );
  NAND2_X1 U10821 ( .A1(n10857), .A2(n8470), .ZN(n8239) );
  AOI22_X1 U10822 ( .A1(n8342), .A2(SI_14_), .B1(n8341), .B2(n13013), .ZN(
        n8238) );
  NAND2_X1 U10823 ( .A1(n8263), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U10824 ( .A1(n8285), .A2(n8240), .ZN(n13298) );
  NAND2_X1 U10825 ( .A1(n8428), .A2(n13298), .ZN(n8244) );
  OR2_X1 U10826 ( .A1(n12562), .A2(n13380), .ZN(n8243) );
  INV_X1 U10827 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13451) );
  OR2_X1 U10828 ( .A1(n8101), .A2(n13451), .ZN(n8242) );
  OR2_X1 U10829 ( .A1(n6535), .A2(n13297), .ZN(n8241) );
  NOR2_X1 U10830 ( .A1(n13452), .A2(n8273), .ZN(n12698) );
  INV_X1 U10831 ( .A(n12698), .ZN(n8245) );
  NAND2_X1 U10832 ( .A1(n13452), .A2(n8273), .ZN(n12697) );
  NAND2_X1 U10833 ( .A1(n8245), .A2(n12697), .ZN(n12695) );
  XNOR2_X1 U10834 ( .A(n8247), .B(n8246), .ZN(n10566) );
  NAND2_X1 U10835 ( .A1(n10566), .A2(n8470), .ZN(n8249) );
  AOI22_X1 U10836 ( .A1(n8342), .A2(n10568), .B1(n8341), .B2(n10567), .ZN(
        n8248) );
  NAND2_X1 U10837 ( .A1(n8473), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8255) );
  OR2_X1 U10838 ( .A1(n6535), .A2(n13321), .ZN(n8254) );
  AND2_X1 U10839 ( .A1(n8250), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8251) );
  NOR2_X1 U10840 ( .A1(n8261), .A2(n8251), .ZN(n12333) );
  OR2_X1 U10841 ( .A1(n8510), .A2(n12333), .ZN(n8253) );
  INV_X1 U10842 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n13464) );
  OR2_X1 U10843 ( .A1(n12563), .A2(n13464), .ZN(n8252) );
  NAND4_X1 U10844 ( .A1(n8255), .A2(n8254), .A3(n8253), .A4(n8252), .ZN(n13306) );
  NAND2_X1 U10845 ( .A1(n13469), .A2(n13306), .ZN(n12688) );
  INV_X1 U10846 ( .A(n13316), .ZN(n12605) );
  XNOR2_X1 U10847 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .ZN(n8256) );
  XNOR2_X1 U10848 ( .A(n8257), .B(n8256), .ZN(n10572) );
  NAND2_X1 U10849 ( .A1(n10572), .A2(n8470), .ZN(n8259) );
  AOI22_X1 U10850 ( .A1(n8342), .A2(n10573), .B1(n8341), .B2(n12998), .ZN(
        n8258) );
  NAND2_X1 U10851 ( .A1(n8259), .A2(n8258), .ZN(n12263) );
  OR2_X1 U10852 ( .A1(n8261), .A2(n8260), .ZN(n8262) );
  NAND2_X1 U10853 ( .A1(n8263), .A2(n8262), .ZN(n13310) );
  NAND2_X1 U10854 ( .A1(n8428), .A2(n13310), .ZN(n8266) );
  INV_X1 U10855 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13309) );
  OR2_X1 U10856 ( .A1(n6535), .A2(n13309), .ZN(n8265) );
  OR2_X1 U10857 ( .A1(n12562), .A2(n15767), .ZN(n8264) );
  INV_X1 U10858 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n15737) );
  INV_X1 U10859 ( .A(n13319), .ZN(n12346) );
  NAND2_X1 U10860 ( .A1(n12263), .A2(n12346), .ZN(n8267) );
  NAND2_X1 U10861 ( .A1(n12605), .A2(n8267), .ZN(n13293) );
  INV_X1 U10862 ( .A(n12263), .ZN(n13457) );
  INV_X1 U10863 ( .A(n13306), .ZN(n12262) );
  OR2_X1 U10864 ( .A1(n13469), .A2(n12262), .ZN(n8270) );
  NAND2_X1 U10865 ( .A1(n8270), .A2(n12346), .ZN(n8269) );
  NAND2_X1 U10866 ( .A1(n13457), .A2(n8269), .ZN(n8272) );
  INV_X1 U10867 ( .A(n8270), .ZN(n13302) );
  NAND2_X1 U10868 ( .A1(n13302), .A2(n13319), .ZN(n8271) );
  NAND2_X1 U10869 ( .A1(n8272), .A2(n8271), .ZN(n13291) );
  AOI22_X1 U10870 ( .A1(n12695), .A2(n13291), .B1(n13305), .B2(n13452), .ZN(
        n8274) );
  INV_X1 U10871 ( .A(n8276), .ZN(n8278) );
  NAND2_X1 U10872 ( .A1(n11060), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8277) );
  XNOR2_X1 U10873 ( .A(n11178), .B(P1_DATAO_REG_15__SCAN_IN), .ZN(n8291) );
  XNOR2_X1 U10874 ( .A(n8293), .B(n8291), .ZN(n10972) );
  NAND2_X1 U10875 ( .A1(n10972), .A2(n8470), .ZN(n8282) );
  AOI22_X1 U10876 ( .A1(n8342), .A2(SI_15_), .B1(n8280), .B2(n8341), .ZN(n8281) );
  NAND2_X1 U10877 ( .A1(n8473), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U10878 ( .A1(n8392), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8283) );
  AND2_X1 U10879 ( .A1(n8284), .A2(n8283), .ZN(n8289) );
  AND2_X1 U10880 ( .A1(n8285), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8286) );
  OR2_X1 U10881 ( .A1(n8286), .A2(n8300), .ZN(n13286) );
  NAND2_X1 U10882 ( .A1(n13286), .A2(n8428), .ZN(n8288) );
  NAND2_X1 U10883 ( .A1(n6539), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8287) );
  OR2_X1 U10884 ( .A1(n13446), .A2(n13272), .ZN(n12701) );
  NAND2_X1 U10885 ( .A1(n13446), .A2(n13272), .ZN(n12705) );
  NAND2_X1 U10886 ( .A1(n13446), .A2(n13295), .ZN(n8290) );
  INV_X1 U10887 ( .A(n8291), .ZN(n8292) );
  NAND2_X1 U10888 ( .A1(n11178), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8294) );
  XNOR2_X1 U10889 ( .A(n15748), .B(P2_DATAO_REG_16__SCAN_IN), .ZN(n8305) );
  XNOR2_X1 U10890 ( .A(n8307), .B(n8305), .ZN(n11075) );
  NAND2_X1 U10891 ( .A1(n11075), .A2(n8470), .ZN(n8298) );
  AOI22_X1 U10892 ( .A1(n8341), .A2(n8296), .B1(n8342), .B2(SI_16_), .ZN(n8297) );
  INV_X1 U10893 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13441) );
  NOR2_X1 U10894 ( .A1(n8300), .A2(n8299), .ZN(n8301) );
  OR2_X1 U10895 ( .A1(n8313), .A2(n8301), .ZN(n13274) );
  NAND2_X1 U10896 ( .A1(n13274), .A2(n8428), .ZN(n8303) );
  AOI22_X1 U10897 ( .A1(n6539), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n8473), .B2(
        P3_REG1_REG_16__SCAN_IN), .ZN(n8302) );
  AND2_X1 U10898 ( .A1(n13373), .A2(n13283), .ZN(n8304) );
  INV_X1 U10899 ( .A(n13260), .ZN(n8319) );
  INV_X1 U10900 ( .A(n8305), .ZN(n8306) );
  NAND2_X1 U10901 ( .A1(n15681), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8308) );
  XNOR2_X1 U10902 ( .A(n15783), .B(P1_DATAO_REG_17__SCAN_IN), .ZN(n8321) );
  XNOR2_X1 U10903 ( .A(n8322), .B(n8321), .ZN(n11125) );
  NAND2_X1 U10904 ( .A1(n11125), .A2(n8470), .ZN(n8311) );
  AOI22_X1 U10905 ( .A1(n8309), .A2(n8341), .B1(n8342), .B2(SI_17_), .ZN(n8310) );
  OR2_X1 U10906 ( .A1(n8313), .A2(n8312), .ZN(n8314) );
  NAND2_X1 U10907 ( .A1(n6566), .A2(n8314), .ZN(n13264) );
  NAND2_X1 U10908 ( .A1(n13264), .A2(n8428), .ZN(n8317) );
  AOI22_X1 U10909 ( .A1(n8392), .A2(P3_REG0_REG_17__SCAN_IN), .B1(n8473), .B2(
        P3_REG1_REG_17__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10910 ( .A1(n6539), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8315) );
  OR2_X1 U10911 ( .A1(n13436), .A2(n13273), .ZN(n12711) );
  NAND2_X1 U10912 ( .A1(n13436), .A2(n13273), .ZN(n12715) );
  INV_X1 U10913 ( .A(n13259), .ZN(n8318) );
  INV_X1 U10914 ( .A(n13273), .ZN(n12857) );
  NAND2_X1 U10915 ( .A1(n13436), .A2(n12857), .ZN(n8320) );
  NAND2_X1 U10916 ( .A1(n15783), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8323) );
  XNOR2_X1 U10917 ( .A(n11419), .B(P2_DATAO_REG_18__SCAN_IN), .ZN(n8336) );
  XNOR2_X1 U10918 ( .A(n8338), .B(n8336), .ZN(n11173) );
  NAND2_X1 U10919 ( .A1(n11173), .A2(n8470), .ZN(n8327) );
  NOR2_X1 U10920 ( .A1(n12569), .A2(n15667), .ZN(n8324) );
  AOI21_X1 U10921 ( .B1(n8325), .B2(n8341), .A(n8324), .ZN(n8326) );
  NAND2_X1 U10922 ( .A1(n6566), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U10923 ( .A1(n8345), .A2(n8328), .ZN(n13248) );
  NAND2_X1 U10924 ( .A1(n13248), .A2(n8428), .ZN(n8334) );
  INV_X1 U10925 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10926 ( .A1(n8473), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U10927 ( .A1(n6539), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8329) );
  OAI211_X1 U10928 ( .C1(n8331), .C2(n12563), .A(n8330), .B(n8329), .ZN(n8332)
         );
  INV_X1 U10929 ( .A(n8332), .ZN(n8333) );
  NAND2_X1 U10930 ( .A1(n13247), .A2(n13232), .ZN(n12714) );
  OR2_X1 U10931 ( .A1(n13247), .A2(n13261), .ZN(n8335) );
  INV_X1 U10932 ( .A(n8336), .ZN(n8337) );
  NAND2_X1 U10933 ( .A1(n15666), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8339) );
  XNOR2_X1 U10934 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .ZN(n8353) );
  XNOR2_X1 U10935 ( .A(n8354), .B(n8353), .ZN(n11164) );
  NAND2_X1 U10936 ( .A1(n11164), .A2(n8470), .ZN(n8344) );
  AOI22_X1 U10937 ( .A1(n8342), .A2(n11163), .B1(n8341), .B2(n12613), .ZN(
        n8343) );
  AND2_X1 U10938 ( .A1(n8345), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8346) );
  OR2_X1 U10939 ( .A1(n8346), .A2(n8359), .ZN(n13237) );
  NAND2_X1 U10940 ( .A1(n13237), .A2(n8428), .ZN(n8351) );
  NAND2_X1 U10941 ( .A1(n8392), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10942 ( .A1(n8473), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8347) );
  OAI211_X1 U10943 ( .C1(n6534), .C2(n13236), .A(n8348), .B(n8347), .ZN(n8349)
         );
  INV_X1 U10944 ( .A(n8349), .ZN(n8350) );
  AND2_X1 U10945 ( .A1(n13432), .A2(n12906), .ZN(n8352) );
  INV_X1 U10946 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11654) );
  NAND2_X1 U10947 ( .A1(n11654), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8355) );
  XNOR2_X1 U10948 ( .A(n11543), .B(P1_DATAO_REG_20__SCAN_IN), .ZN(n8367) );
  XNOR2_X1 U10949 ( .A(n8369), .B(n8367), .ZN(n11383) );
  NAND2_X1 U10950 ( .A1(n11383), .A2(n8470), .ZN(n8357) );
  INV_X1 U10951 ( .A(SI_20_), .ZN(n11384) );
  OR2_X1 U10952 ( .A1(n12569), .A2(n11384), .ZN(n8356) );
  INV_X1 U10953 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n8358) );
  NOR2_X1 U10954 ( .A1(n8359), .A2(n8358), .ZN(n8360) );
  OR2_X1 U10955 ( .A1(n8375), .A2(n8360), .ZN(n13225) );
  NAND2_X1 U10956 ( .A1(n13225), .A2(n8428), .ZN(n8365) );
  INV_X1 U10957 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13422) );
  NAND2_X1 U10958 ( .A1(n6539), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10959 ( .A1(n8473), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8361) );
  OAI211_X1 U10960 ( .C1(n13422), .C2(n12563), .A(n8362), .B(n8361), .ZN(n8363) );
  INV_X1 U10961 ( .A(n8363), .ZN(n8364) );
  NAND2_X1 U10962 ( .A1(n13423), .A2(n13233), .ZN(n12723) );
  NAND2_X1 U10963 ( .A1(n13423), .A2(n13207), .ZN(n8366) );
  INV_X1 U10964 ( .A(n8367), .ZN(n8368) );
  NAND2_X1 U10965 ( .A1(n11543), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U10966 ( .A1(n8371), .A2(n8370), .ZN(n8385) );
  XNOR2_X1 U10967 ( .A(n12382), .B(P1_DATAO_REG_21__SCAN_IN), .ZN(n8383) );
  XNOR2_X1 U10968 ( .A(n8385), .B(n8383), .ZN(n11479) );
  NAND2_X1 U10969 ( .A1(n11479), .A2(n8470), .ZN(n8373) );
  INV_X1 U10970 ( .A(SI_21_), .ZN(n11480) );
  OR2_X1 U10971 ( .A1(n12569), .A2(n11480), .ZN(n8372) );
  INV_X1 U10972 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8374) );
  OR2_X1 U10973 ( .A1(n8375), .A2(n8374), .ZN(n8376) );
  NAND2_X1 U10974 ( .A1(n8390), .A2(n8376), .ZN(n13211) );
  NAND2_X1 U10975 ( .A1(n13211), .A2(n8428), .ZN(n8381) );
  INV_X1 U10976 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13210) );
  NAND2_X1 U10977 ( .A1(n8473), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U10978 ( .A1(n8392), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8377) );
  OAI211_X1 U10979 ( .C1(n6534), .C2(n13210), .A(n8378), .B(n8377), .ZN(n8379)
         );
  INV_X1 U10980 ( .A(n8379), .ZN(n8380) );
  AND2_X1 U10981 ( .A1(n13417), .A2(n13222), .ZN(n8382) );
  INV_X1 U10982 ( .A(n8383), .ZN(n8384) );
  NAND2_X1 U10983 ( .A1(n8385), .A2(n8384), .ZN(n8387) );
  NAND2_X1 U10984 ( .A1(n12382), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8386) );
  XNOR2_X1 U10985 ( .A(n8402), .B(P1_DATAO_REG_22__SCAN_IN), .ZN(n8399) );
  XNOR2_X1 U10986 ( .A(n8401), .B(n8399), .ZN(n11579) );
  NAND2_X1 U10987 ( .A1(n11579), .A2(n8470), .ZN(n8389) );
  OR2_X1 U10988 ( .A1(n12569), .A2(n6960), .ZN(n8388) );
  NAND2_X1 U10989 ( .A1(n8390), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10990 ( .A1(n8412), .A2(n8391), .ZN(n13201) );
  NAND2_X1 U10991 ( .A1(n13201), .A2(n8428), .ZN(n8397) );
  INV_X1 U10992 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13200) );
  NAND2_X1 U10993 ( .A1(n8392), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10994 ( .A1(n8473), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8393) );
  OAI211_X1 U10995 ( .C1(n6535), .C2(n13200), .A(n8394), .B(n8393), .ZN(n8395)
         );
  INV_X1 U10996 ( .A(n8395), .ZN(n8396) );
  NOR2_X1 U10997 ( .A1(n13411), .A2(n13208), .ZN(n8398) );
  INV_X1 U10998 ( .A(n8399), .ZN(n8400) );
  NAND2_X1 U10999 ( .A1(n8402), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8403) );
  INV_X1 U11000 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8404) );
  NAND2_X1 U11001 ( .A1(n8404), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8421) );
  INV_X1 U11002 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11928) );
  NAND2_X1 U11003 ( .A1(n11928), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8405) );
  NAND2_X1 U11004 ( .A1(n8421), .A2(n8405), .ZN(n8407) );
  INV_X1 U11005 ( .A(n8407), .ZN(n8406) );
  NAND2_X1 U11006 ( .A1(n8408), .A2(n8407), .ZN(n8409) );
  NAND2_X1 U11007 ( .A1(n8422), .A2(n8409), .ZN(n11869) );
  NAND2_X1 U11008 ( .A1(n11869), .A2(n8470), .ZN(n8411) );
  INV_X1 U11009 ( .A(SI_23_), .ZN(n11871) );
  OR2_X1 U11010 ( .A1(n12569), .A2(n11871), .ZN(n8410) );
  AND2_X1 U11011 ( .A1(n8412), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8413) );
  OR2_X1 U11012 ( .A1(n8426), .A2(n8413), .ZN(n13190) );
  NAND2_X1 U11013 ( .A1(n13190), .A2(n8428), .ZN(n8419) );
  INV_X1 U11014 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n15708) );
  INV_X1 U11015 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n8414) );
  OR2_X1 U11016 ( .A1(n6535), .A2(n8414), .ZN(n8416) );
  INV_X1 U11017 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n15797) );
  OR2_X1 U11018 ( .A1(n12562), .A2(n15797), .ZN(n8415) );
  OAI211_X1 U11019 ( .C1(n12563), .C2(n15708), .A(n8416), .B(n8415), .ZN(n8417) );
  INV_X1 U11020 ( .A(n8417), .ZN(n8418) );
  NAND2_X1 U11021 ( .A1(n13189), .A2(n12913), .ZN(n12621) );
  NAND2_X1 U11022 ( .A1(n13189), .A2(n13198), .ZN(n8420) );
  XNOR2_X1 U11023 ( .A(n8435), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n12170) );
  NAND2_X1 U11024 ( .A1(n12170), .A2(n8470), .ZN(n8424) );
  INV_X1 U11025 ( .A(SI_24_), .ZN(n12173) );
  OR2_X1 U11026 ( .A1(n12569), .A2(n12173), .ZN(n8423) );
  NAND2_X1 U11027 ( .A1(n8424), .A2(n8423), .ZN(n8571) );
  INV_X1 U11028 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8425) );
  OR2_X1 U11029 ( .A1(n8426), .A2(n8425), .ZN(n8427) );
  NAND2_X1 U11030 ( .A1(n8427), .A2(n8443), .ZN(n13173) );
  NAND2_X1 U11031 ( .A1(n13173), .A2(n8428), .ZN(n8434) );
  INV_X1 U11032 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n8431) );
  NAND2_X1 U11033 ( .A1(n6539), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U11034 ( .A1(n8473), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8429) );
  OAI211_X1 U11035 ( .C1(n8431), .C2(n12563), .A(n8430), .B(n8429), .ZN(n8432)
         );
  INV_X1 U11036 ( .A(n8432), .ZN(n8433) );
  AND2_X1 U11037 ( .A1(n8571), .A2(n12965), .ZN(n13149) );
  INV_X1 U11038 ( .A(n8435), .ZN(n8436) );
  NAND2_X1 U11039 ( .A1(n8436), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U11040 ( .A1(n8439), .A2(n8438), .ZN(n8452) );
  XNOR2_X1 U11041 ( .A(n12126), .B(P1_DATAO_REG_25__SCAN_IN), .ZN(n8450) );
  XNOR2_X1 U11042 ( .A(n8452), .B(n8450), .ZN(n12284) );
  NAND2_X1 U11043 ( .A1(n12284), .A2(n8470), .ZN(n8441) );
  OR2_X1 U11044 ( .A1(n12569), .A2(n12285), .ZN(n8440) );
  NAND2_X1 U11045 ( .A1(n6539), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8448) );
  INV_X1 U11046 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n8442) );
  AOI21_X1 U11047 ( .B1(P3_REG3_REG_25__SCAN_IN), .B2(n8443), .A(n8457), .ZN(
        n13161) );
  OR2_X1 U11048 ( .A1(n8510), .A2(n13161), .ZN(n8446) );
  INV_X1 U11049 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n8444) );
  OR2_X1 U11050 ( .A1(n12563), .A2(n8444), .ZN(n8445) );
  AND2_X1 U11051 ( .A1(n13339), .A2(n13168), .ZN(n8462) );
  OR2_X1 U11052 ( .A1(n13149), .A2(n8462), .ZN(n8449) );
  INV_X1 U11053 ( .A(n8450), .ZN(n8451) );
  NAND2_X1 U11054 ( .A1(n8452), .A2(n8451), .ZN(n8454) );
  NAND2_X1 U11055 ( .A1(n12126), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U11056 ( .A1(n8454), .A2(n8453), .ZN(n8468) );
  INV_X1 U11057 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12353) );
  XNOR2_X1 U11058 ( .A(n12353), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8466) );
  XNOR2_X1 U11059 ( .A(n8468), .B(n8466), .ZN(n13491) );
  NAND2_X1 U11060 ( .A1(n13491), .A2(n8470), .ZN(n8456) );
  INV_X1 U11061 ( .A(SI_26_), .ZN(n13492) );
  OR2_X1 U11062 ( .A1(n12569), .A2(n13492), .ZN(n8455) );
  NAND2_X1 U11063 ( .A1(n8473), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8461) );
  INV_X1 U11064 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13401) );
  OR2_X1 U11065 ( .A1(n12563), .A2(n13401), .ZN(n8460) );
  INV_X1 U11066 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n12941) );
  NAND2_X1 U11067 ( .A1(n8457), .A2(n12941), .ZN(n8476) );
  INV_X1 U11068 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n13145) );
  OR2_X1 U11069 ( .A1(n6535), .A2(n13145), .ZN(n8458) );
  OR2_X1 U11070 ( .A1(n8574), .A2(n13129), .ZN(n8463) );
  OR2_X1 U11071 ( .A1(n8571), .A2(n12965), .ZN(n13150) );
  NAND2_X1 U11072 ( .A1(n8574), .A2(n13129), .ZN(n8464) );
  NAND2_X1 U11073 ( .A1(n8465), .A2(n8464), .ZN(n13127) );
  INV_X1 U11074 ( .A(n8466), .ZN(n8467) );
  NAND2_X1 U11075 ( .A1(n15628), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8469) );
  XNOR2_X1 U11076 ( .A(n12379), .B(P1_DATAO_REG_27__SCAN_IN), .ZN(n8482) );
  XNOR2_X1 U11077 ( .A(n8484), .B(n8482), .ZN(n13486) );
  NAND2_X1 U11078 ( .A1(n13486), .A2(n8470), .ZN(n8472) );
  INV_X1 U11079 ( .A(SI_27_), .ZN(n13488) );
  OR2_X1 U11080 ( .A1(n12569), .A2(n13488), .ZN(n8471) );
  NAND2_X1 U11081 ( .A1(n8473), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8481) );
  INV_X1 U11082 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n13133) );
  OR2_X1 U11083 ( .A1(n6534), .A2(n13133), .ZN(n8480) );
  INV_X1 U11084 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U11085 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(n8476), .ZN(n8477) );
  INV_X1 U11086 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13399) );
  OR2_X1 U11087 ( .A1(n12563), .A2(n13399), .ZN(n8478) );
  INV_X1 U11088 ( .A(n13143), .ZN(n12964) );
  OR2_X1 U11089 ( .A1(n13333), .A2(n12964), .ZN(n8503) );
  NAND2_X1 U11090 ( .A1(n8505), .A2(n8503), .ZN(n8498) );
  INV_X1 U11091 ( .A(n8482), .ZN(n8483) );
  NAND2_X1 U11092 ( .A1(n12379), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8485) );
  INV_X1 U11093 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10377) );
  XNOR2_X1 U11094 ( .A(n10377), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8486) );
  XNOR2_X1 U11095 ( .A(n10379), .B(n8486), .ZN(n12385) );
  NAND2_X1 U11096 ( .A1(n12385), .A2(n8470), .ZN(n8488) );
  INV_X1 U11097 ( .A(SI_28_), .ZN(n15723) );
  OR2_X1 U11098 ( .A1(n12569), .A2(n15723), .ZN(n8487) );
  NAND2_X1 U11099 ( .A1(n6539), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8497) );
  INV_X1 U11100 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9423) );
  OR2_X1 U11101 ( .A1(n12562), .A2(n9423), .ZN(n8496) );
  INV_X1 U11102 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U11103 ( .A1(n8490), .A2(n8489), .ZN(n13106) );
  NAND2_X1 U11104 ( .A1(n8491), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8492) );
  AND2_X1 U11105 ( .A1(n13106), .A2(n8492), .ZN(n12463) );
  INV_X1 U11106 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8493) );
  OR2_X1 U11107 ( .A1(n12563), .A2(n8493), .ZN(n8494) );
  NAND2_X1 U11108 ( .A1(n8498), .A2(n7315), .ZN(n8506) );
  NAND2_X1 U11109 ( .A1(n8499), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8500) );
  MUX2_X1 U11110 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8500), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8502) );
  NAND2_X1 U11111 ( .A1(n12766), .A2(n12579), .ZN(n8536) );
  AND2_X1 U11112 ( .A1(n12745), .A2(n8503), .ZN(n8504) );
  NAND3_X1 U11113 ( .A1(n8506), .A2(n13308), .A3(n10395), .ZN(n8516) );
  NAND2_X1 U11114 ( .A1(n7080), .A2(n8507), .ZN(n11256) );
  INV_X1 U11115 ( .A(n11256), .ZN(n8509) );
  INV_X1 U11116 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10398) );
  OR2_X1 U11117 ( .A1(n12562), .A2(n10398), .ZN(n8513) );
  INV_X1 U11118 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n10404) );
  OR2_X1 U11119 ( .A1(n12563), .A2(n10404), .ZN(n8512) );
  INV_X1 U11120 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n15589) );
  OR2_X1 U11121 ( .A1(n6534), .A2(n15589), .ZN(n8511) );
  OAI22_X1 U11122 ( .A1(n13143), .A2(n15492), .B1(n12576), .B2(n15491), .ZN(
        n8514) );
  INV_X1 U11123 ( .A(n8514), .ZN(n8515) );
  NAND2_X1 U11124 ( .A1(n8516), .A2(n8515), .ZN(n13120) );
  INV_X1 U11125 ( .A(P3_B_REG_SCAN_IN), .ZN(n10389) );
  XNOR2_X1 U11126 ( .A(n8517), .B(n10389), .ZN(n8518) );
  NAND2_X1 U11127 ( .A1(n8518), .A2(n12286), .ZN(n8519) );
  OR2_X1 U11128 ( .A1(n8517), .A2(n8520), .ZN(n8521) );
  NAND2_X1 U11129 ( .A1(n12286), .A2(n13493), .ZN(n8523) );
  NAND2_X1 U11130 ( .A1(n13473), .A2(n13471), .ZN(n9418) );
  INV_X1 U11131 ( .A(n9418), .ZN(n8535) );
  NOR2_X1 U11132 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .ZN(
        n15563) );
  NOR4_X1 U11133 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .A3(
        P3_D_REG_8__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n8527) );
  NOR4_X1 U11134 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n8526) );
  NOR4_X1 U11135 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n8525) );
  NAND4_X1 U11136 ( .A1(n15563), .A2(n8527), .A3(n8526), .A4(n8525), .ZN(n8533) );
  NOR4_X1 U11137 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n8531) );
  NOR4_X1 U11138 ( .A1(P3_D_REG_10__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8530) );
  NOR4_X1 U11139 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_4__SCAN_IN), .ZN(n8529) );
  NOR4_X1 U11140 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8528) );
  NAND4_X1 U11141 ( .A1(n8531), .A2(n8530), .A3(n8529), .A4(n8528), .ZN(n8532)
         );
  NOR2_X1 U11142 ( .A1(n8533), .A2(n8532), .ZN(n8534) );
  INV_X1 U11143 ( .A(n11385), .ZN(n9409) );
  NAND2_X1 U11144 ( .A1(n12627), .A2(n9409), .ZN(n12615) );
  NOR2_X1 U11145 ( .A1(n8536), .A2(n12615), .ZN(n11233) );
  AND2_X1 U11146 ( .A1(n11245), .A2(n11233), .ZN(n11248) );
  NOR2_X1 U11147 ( .A1(n12764), .A2(n11248), .ZN(n8537) );
  INV_X1 U11148 ( .A(n9419), .ZN(n8538) );
  NOR2_X1 U11149 ( .A1(n11763), .A2(n9409), .ZN(n8539) );
  XNOR2_X1 U11150 ( .A(n8539), .B(n9408), .ZN(n8541) );
  NAND2_X1 U11151 ( .A1(n12627), .A2(n12613), .ZN(n8540) );
  NAND2_X1 U11152 ( .A1(n8541), .A2(n8540), .ZN(n11244) );
  NAND3_X1 U11153 ( .A1(n11249), .A2(n11245), .A3(n11244), .ZN(n8542) );
  INV_X1 U11154 ( .A(n8544), .ZN(n8582) );
  AND2_X1 U11155 ( .A1(n12634), .A2(n8545), .ZN(n12637) );
  INV_X1 U11156 ( .A(n15502), .ZN(n8547) );
  NAND2_X1 U11157 ( .A1(n12974), .A2(n15513), .ZN(n8546) );
  NAND2_X1 U11158 ( .A1(n8547), .A2(n8546), .ZN(n11263) );
  OR2_X1 U11159 ( .A1(n12974), .A2(n15513), .ZN(n12624) );
  NAND2_X1 U11160 ( .A1(n11263), .A2(n12624), .ZN(n15490) );
  NAND2_X1 U11161 ( .A1(n12637), .A2(n15490), .ZN(n8552) );
  INV_X1 U11162 ( .A(n11644), .ZN(n8550) );
  INV_X1 U11163 ( .A(n8548), .ZN(n8549) );
  NAND2_X1 U11164 ( .A1(n8552), .A2(n8551), .ZN(n11656) );
  XNOR2_X1 U11165 ( .A(n12973), .B(n11436), .ZN(n12641) );
  NAND2_X1 U11166 ( .A1(n11656), .A2(n12641), .ZN(n11762) );
  OR2_X1 U11167 ( .A1(n12973), .A2(n15472), .ZN(n11761) );
  INV_X1 U11168 ( .A(n12647), .ZN(n11815) );
  NAND2_X1 U11169 ( .A1(n11815), .A2(n12651), .ZN(n8554) );
  OAI211_X1 U11170 ( .C1(n12652), .C2(n11761), .A(n12658), .B(n8554), .ZN(
        n8555) );
  INV_X1 U11171 ( .A(n8555), .ZN(n8556) );
  NAND2_X1 U11172 ( .A1(n12219), .A2(n12969), .ZN(n12665) );
  NAND2_X1 U11173 ( .A1(n12970), .A2(n12000), .ZN(n12659) );
  NAND3_X1 U11174 ( .A1(n11846), .A2(n12665), .A3(n12659), .ZN(n8559) );
  NOR2_X1 U11175 ( .A1(n12970), .A2(n12000), .ZN(n12660) );
  NAND2_X1 U11176 ( .A1(n12660), .A2(n12665), .ZN(n8557) );
  OR2_X1 U11177 ( .A1(n12219), .A2(n12969), .ZN(n12666) );
  AND2_X1 U11178 ( .A1(n8557), .A2(n12666), .ZN(n8558) );
  NAND2_X1 U11179 ( .A1(n8559), .A2(n8558), .ZN(n11932) );
  NAND2_X1 U11180 ( .A1(n11932), .A2(n12671), .ZN(n8560) );
  OR2_X1 U11181 ( .A1(n12235), .A2(n13314), .ZN(n12684) );
  NAND2_X1 U11182 ( .A1(n12235), .A2(n13314), .ZN(n12685) );
  NAND2_X1 U11183 ( .A1(n8563), .A2(n12689), .ZN(n13301) );
  NAND2_X1 U11184 ( .A1(n12263), .A2(n13319), .ZN(n12694) );
  XNOR2_X1 U11185 ( .A(n13373), .B(n13283), .ZN(n13270) );
  INV_X1 U11186 ( .A(n13283), .ZN(n12955) );
  NAND2_X1 U11187 ( .A1(n13373), .A2(n12955), .ZN(n12706) );
  NAND2_X1 U11188 ( .A1(n13267), .A2(n12706), .ZN(n13258) );
  OR2_X1 U11189 ( .A1(n13432), .A2(n13243), .ZN(n12718) );
  INV_X1 U11190 ( .A(n12718), .ZN(n8567) );
  OR2_X1 U11191 ( .A1(n13254), .A2(n8567), .ZN(n13215) );
  OR2_X1 U11192 ( .A1(n13215), .A2(n13218), .ZN(n8565) );
  INV_X1 U11193 ( .A(n12722), .ZN(n8568) );
  AND2_X1 U11194 ( .A1(n6591), .A2(n13228), .ZN(n8566) );
  NAND2_X1 U11195 ( .A1(n13417), .A2(n12443), .ZN(n12726) );
  INV_X1 U11196 ( .A(n12617), .ZN(n8570) );
  AOI21_X1 U11197 ( .B1(n13184), .B2(n13178), .A(n8570), .ZN(n13172) );
  OR2_X1 U11198 ( .A1(n8571), .A2(n13181), .ZN(n12618) );
  NAND2_X1 U11199 ( .A1(n8571), .A2(n13181), .ZN(n12620) );
  NAND2_X1 U11200 ( .A1(n13172), .A2(n13171), .ZN(n13170) );
  NAND2_X1 U11201 ( .A1(n13170), .A2(n12620), .ZN(n13160) );
  NAND2_X1 U11202 ( .A1(n13160), .A2(n13159), .ZN(n13158) );
  INV_X1 U11203 ( .A(n13339), .ZN(n13164) );
  NAND2_X2 U11204 ( .A1(n13158), .A2(n8573), .ZN(n13138) );
  NAND2_X1 U11205 ( .A1(n13333), .A2(n13143), .ZN(n12746) );
  XNOR2_X1 U11206 ( .A(n10397), .B(n12745), .ZN(n13124) );
  AND2_X1 U11207 ( .A1(n15512), .A2(n12760), .ZN(n8575) );
  NAND2_X1 U11208 ( .A1(n11244), .A2(n8575), .ZN(n8578) );
  NOR2_X1 U11209 ( .A1(n11385), .A2(n12579), .ZN(n8576) );
  AND2_X1 U11210 ( .A1(n12766), .A2(n8576), .ZN(n9415) );
  INV_X1 U11211 ( .A(n9415), .ZN(n8577) );
  INV_X1 U11212 ( .A(n8579), .ZN(n10383) );
  OAI22_X1 U11213 ( .A1(n13124), .A2(n13461), .B1(n10383), .B2(n13470), .ZN(
        n8580) );
  INV_X1 U11214 ( .A(n8580), .ZN(n8581) );
  NAND3_X1 U11215 ( .A1(n8719), .A2(n8589), .A3(n8732), .ZN(n8708) );
  AND3_X2 U11216 ( .A1(n8591), .A2(n8590), .A3(n6813), .ZN(n8718) );
  XNOR2_X2 U11217 ( .A(n8596), .B(n15152), .ZN(n8603) );
  AND2_X2 U11218 ( .A1(n8603), .A2(n8598), .ZN(n8736) );
  NAND2_X1 U11219 ( .A1(n8736), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8607) );
  INV_X1 U11220 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14736) );
  OR2_X1 U11221 ( .A1(n9257), .A2(n14736), .ZN(n8606) );
  NAND2_X1 U11222 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n8600) );
  NAND2_X1 U11223 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n8601) );
  NOR2_X2 U11224 ( .A1(n8948), .A2(n15815), .ZN(n8963) );
  OR2_X2 U11225 ( .A1(n9073), .A2(n9052), .ZN(n9054) );
  INV_X1 U11226 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8999) );
  OR2_X2 U11227 ( .A1(n9026), .A2(n8999), .ZN(n9001) );
  INV_X1 U11228 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8987) );
  INV_X1 U11229 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14494) );
  INV_X1 U11230 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14384) );
  INV_X1 U11231 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14421) );
  OR2_X2 U11232 ( .A1(n9217), .A2(n14421), .ZN(n9236) );
  INV_X1 U11233 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14527) );
  NAND2_X1 U11234 ( .A1(n9252), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9253) );
  INV_X1 U11235 ( .A(n9253), .ZN(n8602) );
  NAND2_X1 U11236 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n8602), .ZN(n12485) );
  OAI21_X1 U11237 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(n8602), .A(n12485), .ZN(
        n14735) );
  INV_X1 U11238 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10359) );
  OR2_X1 U11239 ( .A1(n9316), .A2(n10359), .ZN(n8604) );
  INV_X1 U11240 ( .A(n10364), .ZN(n14550) );
  INV_X1 U11241 ( .A(SI_2_), .ZN(n8608) );
  NAND3_X1 U11242 ( .A1(n8769), .A2(n8751), .A3(n8753), .ZN(n8617) );
  NAND2_X1 U11243 ( .A1(n8612), .A2(SI_1_), .ZN(n8766) );
  INV_X1 U11244 ( .A(n8766), .ZN(n8613) );
  NAND2_X1 U11245 ( .A1(n8613), .A2(n8769), .ZN(n8616) );
  INV_X1 U11246 ( .A(n8614), .ZN(n8615) );
  NAND2_X1 U11247 ( .A1(n8615), .A2(SI_2_), .ZN(n8768) );
  INV_X1 U11248 ( .A(SI_4_), .ZN(n8618) );
  NAND2_X1 U11249 ( .A1(n6546), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8619) );
  INV_X1 U11250 ( .A(n8624), .ZN(n8621) );
  INV_X1 U11251 ( .A(SI_3_), .ZN(n8620) );
  NAND2_X1 U11252 ( .A1(n8621), .A2(n8620), .ZN(n8790) );
  AND2_X1 U11253 ( .A1(n8816), .A2(n8790), .ZN(n8827) );
  MUX2_X1 U11254 ( .A(n10520), .B(n10493), .S(n6546), .Z(n8629) );
  INV_X1 U11255 ( .A(SI_5_), .ZN(n8623) );
  NAND2_X1 U11256 ( .A1(n8629), .A2(n8623), .ZN(n8833) );
  INV_X1 U11257 ( .A(n8813), .ZN(n8625) );
  NAND2_X1 U11258 ( .A1(n8625), .A2(n8816), .ZN(n8628) );
  INV_X1 U11259 ( .A(n8626), .ZN(n8627) );
  NAND2_X1 U11260 ( .A1(n8627), .A2(SI_4_), .ZN(n8815) );
  NAND2_X1 U11261 ( .A1(n8628), .A2(n8815), .ZN(n8829) );
  INV_X1 U11262 ( .A(n8629), .ZN(n8630) );
  NAND2_X1 U11263 ( .A1(n8630), .A2(SI_5_), .ZN(n8832) );
  INV_X1 U11264 ( .A(n8832), .ZN(n8631) );
  AOI21_X1 U11265 ( .B1(n8829), .B2(n8833), .A(n8631), .ZN(n8632) );
  MUX2_X1 U11266 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n8609), .Z(n8635) );
  INV_X1 U11267 ( .A(n8635), .ZN(n8634) );
  NAND2_X1 U11268 ( .A1(n8634), .A2(n10446), .ZN(n8636) );
  NAND2_X1 U11269 ( .A1(n8635), .A2(SI_6_), .ZN(n8638) );
  INV_X1 U11270 ( .A(n8855), .ZN(n8637) );
  NAND2_X1 U11271 ( .A1(n8854), .A2(n8637), .ZN(n8858) );
  NAND2_X1 U11272 ( .A1(n8858), .A2(n8638), .ZN(n8867) );
  NAND2_X1 U11273 ( .A1(n8639), .A2(SI_7_), .ZN(n8642) );
  INV_X1 U11274 ( .A(n8639), .ZN(n8641) );
  INV_X1 U11275 ( .A(SI_7_), .ZN(n8640) );
  NAND2_X1 U11276 ( .A1(n8867), .A2(n8866), .ZN(n8869) );
  INV_X1 U11277 ( .A(SI_8_), .ZN(n10502) );
  MUX2_X1 U11278 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n9277), .Z(n8644) );
  NAND2_X1 U11279 ( .A1(n8644), .A2(SI_9_), .ZN(n8647) );
  INV_X1 U11280 ( .A(n8644), .ZN(n8645) );
  NAND2_X1 U11281 ( .A1(n8645), .A2(n10496), .ZN(n8646) );
  MUX2_X1 U11282 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n9277), .Z(n8648) );
  INV_X1 U11283 ( .A(n8648), .ZN(n8649) );
  MUX2_X1 U11284 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n9277), .Z(n8955) );
  INV_X1 U11285 ( .A(n8955), .ZN(n8650) );
  INV_X1 U11286 ( .A(n8954), .ZN(n8651) );
  AOI22_X1 U11287 ( .A1(n8651), .A2(n8969), .B1(n8955), .B2(SI_11_), .ZN(n8653) );
  MUX2_X1 U11288 ( .A(n10832), .B(n8652), .S(n9277), .Z(n8656) );
  XNOR2_X1 U11289 ( .A(n8656), .B(SI_12_), .ZN(n8972) );
  MUX2_X1 U11290 ( .A(n10820), .B(n10818), .S(n9277), .Z(n8657) );
  NAND2_X1 U11291 ( .A1(n8657), .A2(n10573), .ZN(n8658) );
  MUX2_X1 U11292 ( .A(n11080), .B(n11060), .S(n9277), .Z(n9060) );
  INV_X1 U11293 ( .A(n9014), .ZN(n8660) );
  INV_X1 U11294 ( .A(n8661), .ZN(n8659) );
  XNOR2_X1 U11295 ( .A(n8661), .B(SI_15_), .ZN(n9047) );
  INV_X1 U11296 ( .A(n9060), .ZN(n8662) );
  NAND2_X1 U11297 ( .A1(n8662), .A2(SI_14_), .ZN(n8663) );
  MUX2_X1 U11298 ( .A(n15748), .B(n15681), .S(n9277), .Z(n8666) );
  XNOR2_X1 U11299 ( .A(n8666), .B(SI_16_), .ZN(n9017) );
  INV_X1 U11300 ( .A(n9017), .ZN(n8664) );
  MUX2_X1 U11301 ( .A(n15707), .B(n15783), .S(n9277), .Z(n9032) );
  MUX2_X1 U11302 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n9277), .Z(n8993) );
  MUX2_X1 U11303 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n9277), .Z(n8668) );
  NAND2_X1 U11304 ( .A1(n8668), .A2(SI_19_), .ZN(n8982) );
  OAI21_X1 U11305 ( .B1(n8979), .B2(n15667), .A(n8982), .ZN(n8672) );
  NAND3_X1 U11306 ( .A1(n8982), .A2(n15667), .A3(n8979), .ZN(n8670) );
  INV_X1 U11307 ( .A(n8668), .ZN(n8669) );
  NAND2_X1 U11308 ( .A1(n8669), .A2(n11163), .ZN(n8981) );
  MUX2_X1 U11309 ( .A(n12380), .B(n11543), .S(n9277), .Z(n9148) );
  NAND2_X1 U11310 ( .A1(n9165), .A2(SI_20_), .ZN(n8673) );
  MUX2_X1 U11311 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n9277), .Z(n8677) );
  XNOR2_X1 U11312 ( .A(n8677), .B(SI_21_), .ZN(n9170) );
  NOR2_X1 U11313 ( .A1(n9165), .A2(SI_20_), .ZN(n8674) );
  NOR2_X1 U11314 ( .A1(n9170), .A2(n8674), .ZN(n8675) );
  NAND2_X1 U11315 ( .A1(n8677), .A2(SI_21_), .ZN(n8678) );
  MUX2_X1 U11316 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n9277), .Z(n9955) );
  NAND2_X1 U11317 ( .A1(n8679), .A2(SI_22_), .ZN(n8680) );
  MUX2_X1 U11318 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n9277), .Z(n9195) );
  INV_X1 U11319 ( .A(n9195), .ZN(n8681) );
  NAND2_X1 U11320 ( .A1(n8681), .A2(n11871), .ZN(n8682) );
  NAND2_X1 U11321 ( .A1(n9195), .A2(SI_23_), .ZN(n8683) );
  MUX2_X1 U11322 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n9277), .Z(n8686) );
  XNOR2_X1 U11323 ( .A(n8686), .B(SI_24_), .ZN(n9210) );
  NAND2_X1 U11324 ( .A1(n8686), .A2(SI_24_), .ZN(n8687) );
  MUX2_X1 U11325 ( .A(n12124), .B(n12126), .S(n9277), .Z(n8689) );
  NAND2_X1 U11326 ( .A1(n8689), .A2(n12285), .ZN(n8692) );
  INV_X1 U11327 ( .A(n8689), .ZN(n8690) );
  NAND2_X1 U11328 ( .A1(n8690), .A2(SI_25_), .ZN(n8691) );
  NAND2_X1 U11329 ( .A1(n8692), .A2(n8691), .ZN(n9224) );
  MUX2_X1 U11330 ( .A(n12353), .B(n15628), .S(n9277), .Z(n9244) );
  INV_X1 U11331 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14361) );
  MUX2_X1 U11332 ( .A(n14361), .B(n12379), .S(n9277), .Z(n9261) );
  INV_X1 U11333 ( .A(n9261), .ZN(n8693) );
  NOR2_X1 U11334 ( .A1(n8693), .A2(SI_27_), .ZN(n8695) );
  NAND2_X1 U11335 ( .A1(n8693), .A2(SI_27_), .ZN(n8694) );
  INV_X1 U11336 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15840) );
  MUX2_X1 U11337 ( .A(n10377), .B(n15840), .S(n9277), .Z(n8696) );
  NAND2_X1 U11338 ( .A1(n8696), .A2(n15723), .ZN(n9275) );
  INV_X1 U11339 ( .A(n8696), .ZN(n8697) );
  NAND2_X1 U11340 ( .A1(n8697), .A2(SI_28_), .ZN(n8698) );
  NAND2_X1 U11341 ( .A1(n9275), .A2(n8698), .ZN(n8699) );
  NAND2_X1 U11342 ( .A1(n8700), .A2(n8699), .ZN(n8701) );
  NAND2_X1 U11343 ( .A1(n14355), .A2(n8870), .ZN(n8714) );
  OR2_X1 U11344 ( .A1(n9324), .A2(n15840), .ZN(n8713) );
  NAND2_X1 U11345 ( .A1(n8721), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8722) );
  MUX2_X1 U11346 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8722), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8723) );
  XNOR2_X1 U11347 ( .A(n9520), .B(n9521), .ZN(n8731) );
  INV_X1 U11348 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8727) );
  INV_X1 U11349 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8728) );
  BUF_X2 U11350 ( .A(n8760), .Z(n9151) );
  MUX2_X1 U11351 ( .A(n14550), .B(n14738), .S(n8760), .Z(n9270) );
  INV_X1 U11352 ( .A(n9270), .ZN(n9274) );
  INV_X1 U11353 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11341) );
  OR2_X1 U11354 ( .A1(n8784), .A2(n11341), .ZN(n8738) );
  INV_X1 U11355 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8735) );
  INV_X2 U11356 ( .A(n8736), .ZN(n8804) );
  INV_X1 U11357 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10125) );
  INV_X1 U11358 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n15239) );
  INV_X1 U11359 ( .A(SI_0_), .ZN(n8739) );
  NOR2_X1 U11360 ( .A1(n6545), .A2(n8739), .ZN(n8740) );
  XNOR2_X1 U11361 ( .A(n8740), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n15166) );
  MUX2_X1 U11362 ( .A(n15239), .B(n15166), .S(n6531), .Z(n11343) );
  INV_X1 U11363 ( .A(n11343), .ZN(n11441) );
  OR2_X1 U11364 ( .A1(n10118), .A2(n11441), .ZN(n8741) );
  NAND2_X1 U11365 ( .A1(n10118), .A2(n11441), .ZN(n11445) );
  INV_X1 U11366 ( .A(n10107), .ZN(n10106) );
  NAND2_X1 U11367 ( .A1(n11347), .A2(n10106), .ZN(n8759) );
  XNOR2_X1 U11368 ( .A(n9480), .B(n9151), .ZN(n8758) );
  NAND2_X1 U11369 ( .A1(n8736), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8747) );
  INV_X1 U11370 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14571) );
  OR2_X1 U11371 ( .A1(n8784), .A2(n14571), .ZN(n8746) );
  INV_X1 U11372 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10747) );
  OR2_X1 U11373 ( .A1(n9257), .A2(n10747), .ZN(n8745) );
  INV_X1 U11374 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n8743) );
  OR2_X1 U11375 ( .A1(n9316), .A2(n8743), .ZN(n8744) );
  AND4_X2 U11376 ( .A1(n8747), .A2(n8746), .A3(n8745), .A4(n8744), .ZN(n9429)
         );
  INV_X1 U11377 ( .A(n9429), .ZN(n8757) );
  NAND2_X1 U11378 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8748) );
  MUX2_X1 U11379 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8748), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8750) );
  INV_X1 U11380 ( .A(n8749), .ZN(n8772) );
  NAND2_X1 U11381 ( .A1(n8750), .A2(n8772), .ZN(n12477) );
  INV_X1 U11382 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n12475) );
  NAND2_X1 U11383 ( .A1(n8751), .A2(n8766), .ZN(n8754) );
  INV_X1 U11384 ( .A(n8754), .ZN(n8752) );
  NAND2_X1 U11385 ( .A1(n8752), .A2(n8753), .ZN(n8767) );
  INV_X1 U11386 ( .A(n8753), .ZN(n8755) );
  NAND2_X1 U11387 ( .A1(n8755), .A2(n8754), .ZN(n8756) );
  NAND2_X1 U11388 ( .A1(n9429), .A2(n15294), .ZN(n9479) );
  INV_X1 U11389 ( .A(n11444), .ZN(n9360) );
  NAND3_X1 U11390 ( .A1(n8759), .A2(n8758), .A3(n9360), .ZN(n8780) );
  INV_X1 U11391 ( .A(n8760), .ZN(n8799) );
  INV_X1 U11392 ( .A(n8799), .ZN(n8822) );
  NAND2_X1 U11393 ( .A1(n8736), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8765) );
  INV_X1 U11394 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11356) );
  OR2_X1 U11395 ( .A1(n8784), .A2(n11356), .ZN(n8764) );
  INV_X1 U11396 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10749) );
  INV_X1 U11397 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n8761) );
  OR2_X1 U11398 ( .A1(n9316), .A2(n8761), .ZN(n8762) );
  NAND2_X1 U11399 ( .A1(n8767), .A2(n8766), .ZN(n8771) );
  NAND2_X1 U11400 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  XNOR2_X1 U11401 ( .A(n8771), .B(n8770), .ZN(n10490) );
  NAND2_X1 U11402 ( .A1(n10490), .A2(n8870), .ZN(n8778) );
  NAND2_X1 U11403 ( .A1(n8772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8774) );
  OR2_X1 U11404 ( .A1(n6531), .A2(n14596), .ZN(n8777) );
  OR2_X1 U11405 ( .A1(n8775), .A2(n10518), .ZN(n8776) );
  OR2_X2 U11406 ( .A1(n9433), .A2(n15306), .ZN(n15274) );
  NAND2_X1 U11407 ( .A1(n9433), .A2(n15306), .ZN(n8781) );
  NAND3_X1 U11408 ( .A1(n8780), .A2(n8779), .A3(n11360), .ZN(n8783) );
  MUX2_X1 U11409 ( .A(n8781), .B(n15274), .S(n8822), .Z(n8782) );
  NAND2_X1 U11410 ( .A1(n8783), .A2(n8782), .ZN(n8798) );
  NAND2_X1 U11411 ( .A1(n9314), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8789) );
  OR2_X1 U11412 ( .A1(n8784), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8788) );
  INV_X1 U11413 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10752) );
  OR2_X1 U11414 ( .A1(n9257), .A2(n10752), .ZN(n8787) );
  INV_X1 U11415 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8785) );
  OR2_X1 U11416 ( .A1(n9316), .A2(n8785), .ZN(n8786) );
  INV_X1 U11417 ( .A(n8828), .ZN(n8791) );
  NAND2_X1 U11418 ( .A1(n8813), .A2(n8790), .ZN(n8792) );
  NAND2_X1 U11419 ( .A1(n8791), .A2(n8792), .ZN(n8794) );
  INV_X1 U11420 ( .A(n8792), .ZN(n8793) );
  NAND2_X1 U11421 ( .A1(n8828), .A2(n8793), .ZN(n8814) );
  NAND2_X1 U11422 ( .A1(n8870), .A2(n10486), .ZN(n8797) );
  INV_X1 U11423 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n15551) );
  OR2_X1 U11424 ( .A1(n6531), .A2(n14612), .ZN(n8795) );
  NAND2_X1 U11425 ( .A1(n14569), .A2(n15315), .ZN(n8800) );
  INV_X1 U11426 ( .A(n15275), .ZN(n9483) );
  NAND2_X1 U11427 ( .A1(n8798), .A2(n9483), .ZN(n8802) );
  INV_X2 U11428 ( .A(n8799), .ZN(n9307) );
  MUX2_X1 U11429 ( .A(n8800), .B(n9485), .S(n9307), .Z(n8801) );
  NAND2_X1 U11430 ( .A1(n8802), .A2(n8801), .ZN(n8824) );
  NAND2_X1 U11431 ( .A1(n8803), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8812) );
  INV_X1 U11432 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10726) );
  OR2_X1 U11433 ( .A1(n8804), .A2(n10726), .ZN(n8811) );
  INV_X1 U11434 ( .A(n8841), .ZN(n8808) );
  INV_X1 U11435 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8806) );
  INV_X1 U11436 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8805) );
  NAND2_X1 U11437 ( .A1(n8806), .A2(n8805), .ZN(n8807) );
  NAND2_X1 U11438 ( .A1(n8808), .A2(n8807), .ZN(n14465) );
  OR2_X1 U11439 ( .A1(n9317), .A2(n14465), .ZN(n8810) );
  INV_X1 U11440 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11305) );
  OR2_X1 U11441 ( .A1(n9257), .A2(n11305), .ZN(n8809) );
  NAND2_X1 U11442 ( .A1(n8814), .A2(n8813), .ZN(n8818) );
  NAND2_X1 U11443 ( .A1(n8816), .A2(n8815), .ZN(n8817) );
  XNOR2_X1 U11444 ( .A(n8818), .B(n8817), .ZN(n10494) );
  NAND2_X1 U11445 ( .A1(n10494), .A2(n8870), .ZN(n8821) );
  NAND2_X1 U11446 ( .A1(n8819), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8820) );
  MUX2_X1 U11447 ( .A(n14568), .B(n14464), .S(n8822), .Z(n8825) );
  MUX2_X1 U11448 ( .A(n14464), .B(n14568), .S(n8822), .Z(n8823) );
  INV_X1 U11449 ( .A(n8825), .ZN(n8826) );
  NAND2_X1 U11450 ( .A1(n8828), .A2(n8827), .ZN(n8831) );
  INV_X1 U11451 ( .A(n8829), .ZN(n8830) );
  NAND2_X1 U11452 ( .A1(n8831), .A2(n8830), .ZN(n8835) );
  NAND2_X1 U11453 ( .A1(n8833), .A2(n8832), .ZN(n8834) );
  XNOR2_X1 U11454 ( .A(n8835), .B(n8834), .ZN(n10492) );
  NAND2_X1 U11455 ( .A1(n10492), .A2(n8870), .ZN(n8839) );
  INV_X1 U11456 ( .A(n8716), .ZN(n8836) );
  NAND2_X1 U11457 ( .A1(n8836), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8837) );
  XNOR2_X1 U11458 ( .A(n8837), .B(P1_IR_REG_5__SCAN_IN), .ZN(n14637) );
  AOI22_X1 U11459 ( .A1(n9088), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10537), 
        .B2(n14637), .ZN(n8838) );
  AND2_X2 U11460 ( .A1(n8839), .A2(n8838), .ZN(n15262) );
  NAND2_X1 U11461 ( .A1(n8803), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8845) );
  INV_X1 U11462 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n8840) );
  OR2_X1 U11463 ( .A1(n8804), .A2(n8840), .ZN(n8844) );
  OAI21_X1 U11464 ( .B1(n8841), .B2(P1_REG3_REG_5__SCAN_IN), .A(n8878), .ZN(
        n15259) );
  OR2_X1 U11465 ( .A1(n9317), .A2(n15259), .ZN(n8843) );
  INV_X1 U11466 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10757) );
  OR2_X1 U11467 ( .A1(n9257), .A2(n10757), .ZN(n8842) );
  NAND4_X1 U11468 ( .A1(n8845), .A2(n8844), .A3(n8843), .A4(n8842), .ZN(n14567) );
  MUX2_X1 U11469 ( .A(n11576), .B(n14567), .S(n9307), .Z(n8848) );
  MUX2_X1 U11470 ( .A(n14567), .B(n11576), .S(n9307), .Z(n8846) );
  NAND2_X1 U11471 ( .A1(n8803), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8853) );
  INV_X1 U11472 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8849) );
  XNOR2_X1 U11473 ( .A(n8878), .B(n8849), .ZN(n11608) );
  OR2_X1 U11474 ( .A1(n9317), .A2(n11608), .ZN(n8852) );
  INV_X1 U11475 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10731) );
  OR2_X1 U11476 ( .A1(n8804), .A2(n10731), .ZN(n8851) );
  INV_X1 U11477 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11456) );
  OR2_X1 U11478 ( .A1(n9257), .A2(n11456), .ZN(n8850) );
  NAND4_X1 U11479 ( .A1(n8853), .A2(n8852), .A3(n8851), .A4(n8850), .ZN(n14566) );
  NAND2_X1 U11480 ( .A1(n8856), .A2(n8855), .ZN(n8857) );
  AND2_X1 U11481 ( .A1(n8858), .A2(n8857), .ZN(n10498) );
  NAND2_X1 U11482 ( .A1(n10498), .A2(n8870), .ZN(n8862) );
  NAND2_X1 U11483 ( .A1(n8859), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8860) );
  XNOR2_X1 U11484 ( .A(n8860), .B(P1_IR_REG_6__SCAN_IN), .ZN(n14656) );
  AOI22_X1 U11485 ( .A1(n9088), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10537), 
        .B2(n14656), .ZN(n8861) );
  NAND2_X1 U11486 ( .A1(n8862), .A2(n8861), .ZN(n11605) );
  MUX2_X1 U11487 ( .A(n14566), .B(n11605), .S(n9307), .Z(n8864) );
  MUX2_X1 U11488 ( .A(n11605), .B(n14566), .S(n9307), .Z(n8863) );
  INV_X1 U11489 ( .A(n8864), .ZN(n8865) );
  OR2_X1 U11490 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  AND2_X1 U11491 ( .A1(n8869), .A2(n8868), .ZN(n10523) );
  NAND2_X1 U11492 ( .A1(n10523), .A2(n9286), .ZN(n8877) );
  NAND2_X1 U11493 ( .A1(n8872), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8871) );
  MUX2_X1 U11494 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8871), .S(
        P1_IR_REG_7__SCAN_IN), .Z(n8875) );
  INV_X1 U11495 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U11496 ( .A1(n8875), .A2(n8910), .ZN(n14671) );
  INV_X1 U11497 ( .A(n14671), .ZN(n10764) );
  AOI22_X1 U11498 ( .A1(n9088), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10537), 
        .B2(n10764), .ZN(n8876) );
  INV_X1 U11499 ( .A(n15251), .ZN(n9489) );
  NAND2_X1 U11500 ( .A1(n8803), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8884) );
  INV_X1 U11501 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10732) );
  OR2_X1 U11502 ( .A1(n8804), .A2(n10732), .ZN(n8883) );
  INV_X1 U11503 ( .A(n8878), .ZN(n8879) );
  AOI21_X1 U11504 ( .B1(n8879), .B2(P1_REG3_REG_6__SCAN_IN), .A(
        P1_REG3_REG_7__SCAN_IN), .ZN(n8880) );
  OR2_X1 U11505 ( .A1(n8880), .A2(n8896), .ZN(n15248) );
  OR2_X1 U11506 ( .A1(n9317), .A2(n15248), .ZN(n8882) );
  INV_X1 U11507 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10761) );
  OR2_X1 U11508 ( .A1(n9257), .A2(n10761), .ZN(n8881) );
  NAND4_X1 U11509 ( .A1(n8884), .A2(n8883), .A3(n8882), .A4(n8881), .ZN(n14565) );
  MUX2_X1 U11510 ( .A(n9489), .B(n14565), .S(n9307), .Z(n8888) );
  MUX2_X1 U11511 ( .A(n9489), .B(n14565), .S(n9330), .Z(n8885) );
  INV_X1 U11512 ( .A(n8887), .ZN(n8890) );
  INV_X1 U11513 ( .A(n8888), .ZN(n8889) );
  NAND2_X1 U11514 ( .A1(n8910), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8894) );
  XNOR2_X1 U11515 ( .A(n8894), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U11516 ( .A1(n9088), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10809), 
        .B2(n10537), .ZN(n8895) );
  NAND2_X1 U11517 ( .A1(n8803), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8901) );
  INV_X1 U11518 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10736) );
  OR2_X1 U11519 ( .A1(n8804), .A2(n10736), .ZN(n8900) );
  OR2_X1 U11520 ( .A1(n8896), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8897) );
  NAND2_X1 U11521 ( .A1(n8927), .A2(n8897), .ZN(n11902) );
  OR2_X1 U11522 ( .A1(n9317), .A2(n11902), .ZN(n8899) );
  INV_X1 U11523 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10765) );
  OR2_X1 U11524 ( .A1(n9257), .A2(n10765), .ZN(n8898) );
  INV_X1 U11525 ( .A(n9151), .ZN(n9091) );
  MUX2_X1 U11526 ( .A(n10177), .B(n14564), .S(n9091), .Z(n8904) );
  MUX2_X1 U11527 ( .A(n10177), .B(n14564), .S(n9307), .Z(n8902) );
  INV_X1 U11528 ( .A(n8904), .ZN(n8905) );
  NAND2_X1 U11529 ( .A1(n8906), .A2(n8909), .ZN(n10549) );
  NAND2_X1 U11530 ( .A1(n8937), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8911) );
  XNOR2_X1 U11531 ( .A(n8911), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U11532 ( .A1(n10537), .A2(n10793), .B1(n9088), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U11533 ( .A1(n9315), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8919) );
  INV_X1 U11534 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n8914) );
  OR2_X1 U11535 ( .A1(n9316), .A2(n8914), .ZN(n8918) );
  INV_X1 U11536 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n8915) );
  OR2_X1 U11537 ( .A1(n8804), .A2(n8915), .ZN(n8917) );
  INV_X1 U11538 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8926) );
  XNOR2_X1 U11539 ( .A(n8927), .B(n8926), .ZN(n12209) );
  OR2_X1 U11540 ( .A1(n9317), .A2(n12209), .ZN(n8916) );
  INV_X1 U11541 ( .A(n11522), .ZN(n14563) );
  MUX2_X1 U11542 ( .A(n11991), .B(n14563), .S(n9307), .Z(n8922) );
  MUX2_X1 U11543 ( .A(n14563), .B(n11991), .S(n9307), .Z(n8920) );
  NAND2_X1 U11544 ( .A1(n8921), .A2(n8920), .ZN(n8924) );
  NAND2_X1 U11545 ( .A1(n8924), .A2(n8923), .ZN(n8944) );
  NAND2_X1 U11546 ( .A1(n8803), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8932) );
  INV_X1 U11547 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15716) );
  OR2_X1 U11548 ( .A1(n8804), .A2(n15716), .ZN(n8931) );
  INV_X1 U11549 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8925) );
  OAI21_X1 U11550 ( .B1(n8927), .B2(n8926), .A(n8925), .ZN(n8928) );
  NAND2_X1 U11551 ( .A1(n8928), .A2(n8948), .ZN(n12296) );
  OR2_X1 U11552 ( .A1(n9317), .A2(n12296), .ZN(n8930) );
  INV_X1 U11553 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10794) );
  OR2_X1 U11554 ( .A1(n9257), .A2(n10794), .ZN(n8929) );
  INV_X1 U11555 ( .A(n12206), .ZN(n14562) );
  OR2_X1 U11556 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  OR2_X1 U11557 ( .A1(n10570), .A2(n9296), .ZN(n8942) );
  INV_X1 U11558 ( .A(n8937), .ZN(n8939) );
  INV_X1 U11559 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U11560 ( .A1(n8939), .A2(n8938), .ZN(n8956) );
  NAND2_X1 U11561 ( .A1(n8956), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8940) );
  XNOR2_X1 U11562 ( .A(n8940), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U11563 ( .A1(n10840), .A2(n10537), .B1(P2_DATAO_REG_10__SCAN_IN), 
        .B2(n9088), .ZN(n8941) );
  NAND2_X2 U11564 ( .A1(n8942), .A2(n8941), .ZN(n15096) );
  MUX2_X1 U11565 ( .A(n14562), .B(n15096), .S(n9307), .Z(n8945) );
  MUX2_X1 U11566 ( .A(n15096), .B(n14562), .S(n9307), .Z(n8943) );
  INV_X1 U11567 ( .A(n8945), .ZN(n8946) );
  NAND2_X1 U11568 ( .A1(n8803), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8953) );
  INV_X1 U11569 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n8947) );
  OR2_X1 U11570 ( .A1(n8804), .A2(n8947), .ZN(n8952) );
  AND2_X1 U11571 ( .A1(n8948), .A2(n15815), .ZN(n8949) );
  OR2_X1 U11572 ( .A1(n8949), .A2(n8963), .ZN(n14505) );
  OR2_X1 U11573 ( .A1(n9317), .A2(n14505), .ZN(n8951) );
  INV_X1 U11574 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11881) );
  OR2_X1 U11575 ( .A1(n9257), .A2(n11881), .ZN(n8950) );
  NAND4_X1 U11576 ( .A1(n8953), .A2(n8952), .A3(n8951), .A4(n8950), .ZN(n14561) );
  XNOR2_X1 U11577 ( .A(n8955), .B(SI_11_), .ZN(n8970) );
  NAND2_X1 U11578 ( .A1(n10697), .A2(n9286), .ZN(n8959) );
  NAND2_X1 U11579 ( .A1(n8957), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8975) );
  XNOR2_X1 U11580 ( .A(n8975), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U11581 ( .A1(n11020), .A2(n10537), .B1(P2_DATAO_REG_11__SCAN_IN), 
        .B2(n9088), .ZN(n8958) );
  MUX2_X1 U11582 ( .A(n14561), .B(n14507), .S(n9091), .Z(n8962) );
  MUX2_X1 U11583 ( .A(n14561), .B(n14507), .S(n9307), .Z(n8960) );
  NAND2_X1 U11584 ( .A1(n8803), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8968) );
  INV_X1 U11585 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n15084) );
  OR2_X1 U11586 ( .A1(n8804), .A2(n15084), .ZN(n8967) );
  INV_X1 U11587 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11019) );
  OR2_X1 U11588 ( .A1(n9257), .A2(n11019), .ZN(n8966) );
  NOR2_X1 U11589 ( .A1(n8963), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8964) );
  OR2_X1 U11590 ( .A1(n9078), .A2(n8964), .ZN(n12059) );
  OR2_X1 U11591 ( .A1(n9317), .A2(n12059), .ZN(n8965) );
  NAND4_X1 U11592 ( .A1(n8968), .A2(n8967), .A3(n8966), .A4(n8965), .ZN(n14560) );
  INV_X1 U11593 ( .A(n14560), .ZN(n10201) );
  NAND2_X1 U11594 ( .A1(n10715), .A2(n9286), .ZN(n8978) );
  INV_X1 U11595 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U11596 ( .A1(n8975), .A2(n8974), .ZN(n8976) );
  NAND2_X1 U11597 ( .A1(n8976), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9065) );
  XNOR2_X1 U11598 ( .A(n9065), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U11599 ( .A1(n11133), .A2(n10537), .B1(n9088), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8977) );
  INV_X1 U11600 ( .A(n14974), .ZN(n15148) );
  MUX2_X1 U11601 ( .A(n10201), .B(n15148), .S(n9307), .Z(n9096) );
  MUX2_X1 U11602 ( .A(n14560), .B(n14974), .S(n9091), .Z(n9095) );
  NAND2_X1 U11603 ( .A1(n9096), .A2(n9095), .ZN(n9099) );
  NAND2_X1 U11604 ( .A1(n8982), .A2(n8981), .ZN(n8983) );
  AOI22_X1 U11605 ( .A1(n14731), .A2(n10537), .B1(n9088), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n8985) );
  AND2_X1 U11606 ( .A1(n9001), .A2(n8987), .ZN(n8988) );
  OR2_X1 U11607 ( .A1(n8988), .A2(n9141), .ZN(n14876) );
  INV_X1 U11608 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14877) );
  NAND2_X1 U11609 ( .A1(n8803), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U11610 ( .A1(n9314), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8989) );
  OAI211_X1 U11611 ( .C1(n14877), .C2(n9257), .A(n8990), .B(n8989), .ZN(n8991)
         );
  INV_X1 U11612 ( .A(n8991), .ZN(n8992) );
  XNOR2_X1 U11613 ( .A(n8994), .B(n8993), .ZN(n11418) );
  NAND2_X1 U11614 ( .A1(n11418), .A2(n8870), .ZN(n8998) );
  XNOR2_X1 U11615 ( .A(n8995), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14703) );
  NOR2_X1 U11616 ( .A1(n9324), .A2(n15666), .ZN(n8996) );
  AOI21_X1 U11617 ( .B1(n14703), .B2(n10537), .A(n8996), .ZN(n8997) );
  NAND2_X1 U11618 ( .A1(n9026), .A2(n8999), .ZN(n9000) );
  AND2_X1 U11619 ( .A1(n9001), .A2(n9000), .ZN(n14892) );
  NAND2_X1 U11620 ( .A1(n14892), .A2(n9238), .ZN(n9007) );
  INV_X1 U11621 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U11622 ( .A1(n8736), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U11623 ( .A1(n8803), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9002) );
  OAI211_X1 U11624 ( .C1(n9004), .C2(n9257), .A(n9003), .B(n9002), .ZN(n9005)
         );
  INV_X1 U11625 ( .A(n9005), .ZN(n9006) );
  OR2_X1 U11626 ( .A1(n15048), .A2(n14558), .ZN(n9461) );
  NAND2_X1 U11627 ( .A1(n15048), .A2(n14558), .ZN(n9462) );
  NAND2_X1 U11628 ( .A1(n9461), .A2(n9462), .ZN(n9008) );
  AND2_X1 U11629 ( .A1(n9054), .A2(n9009), .ZN(n9010) );
  OR2_X1 U11630 ( .A1(n9010), .A2(n9025), .ZN(n14927) );
  AOI22_X1 U11631 ( .A1(n8803), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n9314), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n9012) );
  NAND2_X1 U11632 ( .A1(n9315), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9011) );
  OAI211_X1 U11633 ( .C1(n14927), .C2(n9317), .A(n9012), .B(n9011), .ZN(n14941) );
  NAND2_X1 U11634 ( .A1(n9016), .A2(n9015), .ZN(n9018) );
  NAND2_X1 U11635 ( .A1(n8726), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9020) );
  MUX2_X1 U11636 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9020), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9022) );
  INV_X1 U11637 ( .A(n9021), .ZN(n9034) );
  AOI22_X1 U11638 ( .A1(n9088), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12196), 
        .B2(n10537), .ZN(n9023) );
  OR2_X1 U11639 ( .A1(n9025), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9027) );
  AND2_X1 U11640 ( .A1(n9027), .A2(n9026), .ZN(n14911) );
  NAND2_X1 U11641 ( .A1(n14911), .A2(n9238), .ZN(n9030) );
  AOI22_X1 U11642 ( .A1(n8803), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n8736), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U11643 ( .A1(n9315), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U11644 ( .A1(n9118), .A2(n14925), .ZN(n9038) );
  OR2_X1 U11645 ( .A1(n14941), .A2(n9307), .ZN(n9040) );
  XNOR2_X1 U11646 ( .A(n9032), .B(SI_17_), .ZN(n9033) );
  XNOR2_X1 U11647 ( .A(n9031), .B(n9033), .ZN(n11015) );
  NAND2_X1 U11648 ( .A1(n11015), .A2(n9286), .ZN(n9037) );
  NAND2_X1 U11649 ( .A1(n9034), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9035) );
  XNOR2_X1 U11650 ( .A(n9035), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14685) );
  AOI22_X1 U11651 ( .A1(n14685), .A2(n10537), .B1(n9088), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n9036) );
  AOI21_X1 U11652 ( .B1(n9038), .B2(n9040), .A(n7090), .ZN(n9043) );
  NAND2_X1 U11653 ( .A1(n9118), .A2(n14884), .ZN(n9039) );
  NAND2_X1 U11654 ( .A1(n14925), .A2(n9151), .ZN(n9111) );
  OR2_X1 U11655 ( .A1(n15060), .A2(n9111), .ZN(n9042) );
  INV_X1 U11656 ( .A(n9040), .ZN(n9114) );
  NAND2_X1 U11657 ( .A1(n9114), .A2(n14884), .ZN(n9041) );
  NAND2_X1 U11658 ( .A1(n9042), .A2(n9041), .ZN(n9117) );
  NAND2_X1 U11659 ( .A1(n9044), .A2(n10860), .ZN(n9045) );
  NAND2_X1 U11660 ( .A1(n11175), .A2(n8870), .ZN(n9051) );
  INV_X1 U11661 ( .A(n8724), .ZN(n9048) );
  NAND2_X1 U11662 ( .A1(n9048), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9049) );
  XNOR2_X1 U11663 ( .A(n9049), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U11664 ( .A1(n9088), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n10537), 
        .B2(n11812), .ZN(n9050) );
  NAND2_X2 U11665 ( .A1(n9051), .A2(n9050), .ZN(n9456) );
  NAND2_X1 U11666 ( .A1(n9073), .A2(n9052), .ZN(n9053) );
  AND2_X1 U11667 ( .A1(n9054), .A2(n9053), .ZN(n14946) );
  NAND2_X1 U11668 ( .A1(n14946), .A2(n9238), .ZN(n9057) );
  AOI22_X1 U11669 ( .A1(n8803), .A2(P1_REG0_REG_15__SCAN_IN), .B1(n9314), .B2(
        P1_REG1_REG_15__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U11670 ( .A1(n9315), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U11671 ( .A1(n9456), .A2(n14435), .ZN(n9356) );
  OR2_X2 U11672 ( .A1(n9456), .A2(n14435), .ZN(n9496) );
  MUX2_X1 U11673 ( .A(n9356), .B(n9496), .S(n9091), .Z(n9058) );
  NAND2_X1 U11674 ( .A1(n9061), .A2(n9060), .ZN(n9062) );
  NAND2_X1 U11675 ( .A1(n9065), .A2(n9064), .ZN(n9066) );
  NAND2_X1 U11676 ( .A1(n9066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9087) );
  INV_X1 U11677 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U11678 ( .A1(n9087), .A2(n9067), .ZN(n9068) );
  NAND2_X1 U11679 ( .A1(n9068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9069) );
  AOI22_X1 U11680 ( .A1(n11805), .A2(n10537), .B1(n9088), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U11681 ( .A1(n9080), .A2(n9071), .ZN(n9072) );
  NAND2_X1 U11682 ( .A1(n9073), .A2(n9072), .ZN(n14968) );
  OR2_X1 U11683 ( .A1(n14968), .A2(n9317), .ZN(n9077) );
  INV_X1 U11684 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n15138) );
  OR2_X1 U11685 ( .A1(n9316), .A2(n15138), .ZN(n9076) );
  INV_X1 U11686 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15071) );
  OR2_X1 U11687 ( .A1(n8804), .A2(n15071), .ZN(n9075) );
  INV_X1 U11688 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14969) );
  OR2_X1 U11689 ( .A1(n9257), .A2(n14969), .ZN(n9074) );
  NAND2_X1 U11690 ( .A1(n14957), .A2(n14480), .ZN(n9102) );
  NAND2_X1 U11691 ( .A1(n8803), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9084) );
  OR2_X1 U11692 ( .A1(n9078), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9079) );
  NAND2_X1 U11693 ( .A1(n9080), .A2(n9079), .ZN(n14985) );
  OR2_X1 U11694 ( .A1(n9317), .A2(n14985), .ZN(n9083) );
  INV_X1 U11695 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n15079) );
  OR2_X1 U11696 ( .A1(n8804), .A2(n15079), .ZN(n9082) );
  INV_X1 U11697 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n14986) );
  OR2_X1 U11698 ( .A1(n9257), .A2(n14986), .ZN(n9081) );
  NAND4_X1 U11699 ( .A1(n9084), .A2(n9083), .A3(n9082), .A4(n9081), .ZN(n14559) );
  XNOR2_X1 U11700 ( .A(n9085), .B(n9086), .ZN(n10817) );
  NAND2_X1 U11701 ( .A1(n10817), .A2(n9286), .ZN(n9090) );
  XNOR2_X1 U11702 ( .A(n9087), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U11703 ( .A1(n11205), .A2(n10537), .B1(P2_DATAO_REG_13__SCAN_IN), 
        .B2(n9088), .ZN(n9089) );
  MUX2_X1 U11704 ( .A(n14559), .B(n14984), .S(n9091), .Z(n9105) );
  INV_X1 U11705 ( .A(n9151), .ZN(n9330) );
  NOR2_X1 U11706 ( .A1(n14984), .A2(n9330), .ZN(n9093) );
  NOR2_X1 U11707 ( .A1(n9307), .A2(n14559), .ZN(n9092) );
  OR3_X1 U11708 ( .A1(n9105), .A2(n9093), .A3(n9092), .ZN(n9094) );
  OAI211_X1 U11709 ( .C1(n9096), .C2(n9095), .A(n14967), .B(n9094), .ZN(n9097)
         );
  INV_X1 U11710 ( .A(n9100), .ZN(n9140) );
  NAND2_X1 U11711 ( .A1(n9496), .A2(n9495), .ZN(n9101) );
  NAND2_X1 U11712 ( .A1(n9101), .A2(n9307), .ZN(n9109) );
  NAND2_X1 U11713 ( .A1(n9356), .A2(n9102), .ZN(n9103) );
  NAND2_X1 U11714 ( .A1(n9103), .A2(n9330), .ZN(n9108) );
  INV_X1 U11715 ( .A(n14559), .ZN(n14377) );
  NOR2_X1 U11716 ( .A1(n9151), .A2(n14377), .ZN(n9104) );
  AOI21_X1 U11717 ( .B1(n14984), .B2(n9151), .A(n9104), .ZN(n9106) );
  NAND3_X1 U11718 ( .A1(n14967), .A2(n9106), .A3(n9105), .ZN(n9107) );
  NAND3_X1 U11719 ( .A1(n9109), .A2(n9108), .A3(n9107), .ZN(n9123) );
  INV_X1 U11720 ( .A(n9110), .ZN(n9113) );
  INV_X1 U11721 ( .A(n9111), .ZN(n9112) );
  AOI21_X1 U11722 ( .B1(n9118), .B2(n9113), .A(n9112), .ZN(n9121) );
  NAND2_X1 U11723 ( .A1(n9118), .A2(n9114), .ZN(n9115) );
  OAI21_X1 U11724 ( .B1(n14925), .B2(n9151), .A(n9115), .ZN(n9116) );
  NAND2_X1 U11725 ( .A1(n9116), .A2(n15055), .ZN(n9120) );
  NAND2_X1 U11726 ( .A1(n9118), .A2(n9117), .ZN(n9119) );
  OAI211_X1 U11727 ( .C1(n9121), .C2(n15055), .A(n9120), .B(n9119), .ZN(n9122)
         );
  AND2_X1 U11728 ( .A1(n14910), .A2(n9330), .ZN(n9124) );
  NAND2_X1 U11729 ( .A1(n15048), .A2(n9124), .ZN(n9129) );
  NAND2_X1 U11730 ( .A1(n14875), .A2(n9129), .ZN(n9128) );
  NAND2_X1 U11731 ( .A1(n14558), .A2(n9151), .ZN(n9130) );
  INV_X1 U11732 ( .A(n9130), .ZN(n9125) );
  NAND2_X1 U11733 ( .A1(n9125), .A2(n14557), .ZN(n9126) );
  OAI22_X1 U11734 ( .A1(n15048), .A2(n9126), .B1(n9151), .B2(n14557), .ZN(
        n9127) );
  OR2_X1 U11735 ( .A1(n9128), .A2(n9127), .ZN(n9134) );
  NOR2_X1 U11736 ( .A1(n9129), .A2(n14557), .ZN(n9132) );
  INV_X1 U11737 ( .A(n14557), .ZN(n14885) );
  OAI22_X1 U11738 ( .A1(n15048), .A2(n9130), .B1(n9330), .B2(n14885), .ZN(
        n9131) );
  OR3_X1 U11739 ( .A1(n9132), .A2(n14875), .A3(n9131), .ZN(n9133) );
  NAND2_X1 U11740 ( .A1(n9134), .A2(n9133), .ZN(n9135) );
  OAI21_X1 U11741 ( .B1(n9137), .B2(n9136), .A(n9135), .ZN(n9138) );
  INV_X1 U11742 ( .A(n9138), .ZN(n9139) );
  NOR2_X1 U11743 ( .A1(n9141), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9142) );
  OR2_X1 U11744 ( .A1(n9157), .A2(n9142), .ZN(n14472) );
  INV_X1 U11745 ( .A(n14472), .ZN(n14860) );
  NAND2_X1 U11746 ( .A1(n14860), .A2(n9238), .ZN(n9147) );
  INV_X1 U11747 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14862) );
  NAND2_X1 U11748 ( .A1(n8803), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9144) );
  NAND2_X1 U11749 ( .A1(n8736), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9143) );
  OAI211_X1 U11750 ( .C1(n14862), .C2(n9257), .A(n9144), .B(n9143), .ZN(n9145)
         );
  INV_X1 U11751 ( .A(n9145), .ZN(n9146) );
  XNOR2_X1 U11752 ( .A(n9166), .B(n9148), .ZN(n11542) );
  NAND2_X1 U11753 ( .A1(n11542), .A2(n8870), .ZN(n9150) );
  OR2_X1 U11754 ( .A1(n9324), .A2(n11543), .ZN(n9149) );
  INV_X1 U11755 ( .A(n14858), .ZN(n15036) );
  MUX2_X1 U11756 ( .A(n14401), .B(n15036), .S(n9151), .Z(n9153) );
  INV_X1 U11757 ( .A(n14401), .ZN(n14556) );
  MUX2_X1 U11758 ( .A(n14556), .B(n14858), .S(n9091), .Z(n9152) );
  NAND2_X1 U11759 ( .A1(n9154), .A2(n9153), .ZN(n9155) );
  OR2_X1 U11760 ( .A1(n9157), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9158) );
  AND2_X1 U11761 ( .A1(n9176), .A2(n9158), .ZN(n14836) );
  NAND2_X1 U11762 ( .A1(n14836), .A2(n9238), .ZN(n9164) );
  INV_X1 U11763 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U11764 ( .A1(n8803), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U11765 ( .A1(n9314), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9159) );
  OAI211_X1 U11766 ( .C1(n9161), .C2(n9257), .A(n9160), .B(n9159), .ZN(n9162)
         );
  INV_X1 U11767 ( .A(n9162), .ZN(n9163) );
  NAND2_X1 U11768 ( .A1(n9164), .A2(n9163), .ZN(n14555) );
  NAND2_X1 U11769 ( .A1(n9166), .A2(n9165), .ZN(n9169) );
  OR2_X1 U11770 ( .A1(n9167), .A2(n11384), .ZN(n9168) );
  NAND2_X1 U11771 ( .A1(n9169), .A2(n9168), .ZN(n9171) );
  XNOR2_X1 U11772 ( .A(n9171), .B(n9170), .ZN(n11694) );
  NAND2_X1 U11773 ( .A1(n11694), .A2(n9286), .ZN(n9173) );
  OR2_X1 U11774 ( .A1(n9324), .A2(n12382), .ZN(n9172) );
  MUX2_X1 U11775 ( .A(n14555), .B(n9519), .S(n9330), .Z(n9175) );
  MUX2_X1 U11776 ( .A(n14555), .B(n9519), .S(n9151), .Z(n9174) );
  NAND2_X1 U11777 ( .A1(n9176), .A2(n14494), .ZN(n9177) );
  AND2_X1 U11778 ( .A1(n9189), .A2(n9177), .ZN(n14814) );
  NAND2_X1 U11779 ( .A1(n14814), .A2(n9238), .ZN(n9182) );
  INV_X1 U11780 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n15640) );
  NAND2_X1 U11781 ( .A1(n9315), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9179) );
  INV_X1 U11782 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n15755) );
  OR2_X1 U11783 ( .A1(n8804), .A2(n15755), .ZN(n9178) );
  OAI211_X1 U11784 ( .C1(n9316), .C2(n15640), .A(n9179), .B(n9178), .ZN(n9180)
         );
  INV_X1 U11785 ( .A(n9180), .ZN(n9181) );
  NAND2_X1 U11786 ( .A1(n9182), .A2(n9181), .ZN(n14554) );
  OR2_X1 U11787 ( .A1(n9956), .A2(n6545), .ZN(n9183) );
  XNOR2_X1 U11788 ( .A(n9183), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15164) );
  MUX2_X1 U11789 ( .A(n14554), .B(n7511), .S(n8760), .Z(n9187) );
  INV_X1 U11790 ( .A(n14554), .ZN(n10269) );
  MUX2_X1 U11791 ( .A(n10269), .B(n14817), .S(n9330), .Z(n9185) );
  AOI21_X1 U11792 ( .B1(n9188), .B2(n9187), .A(n9185), .ZN(n9186) );
  AND2_X1 U11793 ( .A1(n9189), .A2(n14384), .ZN(n9190) );
  OR2_X1 U11794 ( .A1(n9190), .A2(n9202), .ZN(n14791) );
  INV_X1 U11795 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14801) );
  NAND2_X1 U11796 ( .A1(n8803), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9192) );
  NAND2_X1 U11797 ( .A1(n8736), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9191) );
  OAI211_X1 U11798 ( .C1(n14801), .C2(n9257), .A(n9192), .B(n9191), .ZN(n9193)
         );
  INV_X1 U11799 ( .A(n9193), .ZN(n9194) );
  OAI21_X2 U11800 ( .B1(n14791), .B2(n9317), .A(n9194), .ZN(n14553) );
  XNOR2_X1 U11801 ( .A(n9195), .B(SI_23_), .ZN(n9196) );
  XNOR2_X1 U11802 ( .A(n9197), .B(n9196), .ZN(n11925) );
  NAND2_X1 U11803 ( .A1(n11925), .A2(n8870), .ZN(n9199) );
  OR2_X1 U11804 ( .A1(n9324), .A2(n11928), .ZN(n9198) );
  MUX2_X1 U11805 ( .A(n14553), .B(n14800), .S(n9330), .Z(n9201) );
  MUX2_X1 U11806 ( .A(n14553), .B(n14800), .S(n8760), .Z(n9200) );
  OR2_X1 U11807 ( .A1(n9202), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U11808 ( .A1(n9217), .A2(n9203), .ZN(n14456) );
  OR2_X1 U11809 ( .A1(n14456), .A2(n9317), .ZN(n9209) );
  INV_X1 U11810 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9206) );
  NAND2_X1 U11811 ( .A1(n8803), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11812 ( .A1(n9314), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9204) );
  OAI211_X1 U11813 ( .C1(n9206), .C2(n9257), .A(n9205), .B(n9204), .ZN(n9207)
         );
  INV_X1 U11814 ( .A(n9207), .ZN(n9208) );
  XNOR2_X1 U11815 ( .A(n9211), .B(n9210), .ZN(n12104) );
  NAND2_X1 U11816 ( .A1(n12104), .A2(n9286), .ZN(n9213) );
  INV_X1 U11817 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12105) );
  OR2_X1 U11818 ( .A1(n9324), .A2(n12105), .ZN(n9212) );
  MUX2_X1 U11819 ( .A(n14552), .B(n15117), .S(n8760), .Z(n9215) );
  MUX2_X1 U11820 ( .A(n14552), .B(n15117), .S(n9091), .Z(n9214) );
  INV_X1 U11821 ( .A(n9215), .ZN(n9216) );
  NAND2_X1 U11822 ( .A1(n9217), .A2(n14421), .ZN(n9218) );
  NAND2_X1 U11823 ( .A1(n9236), .A2(n9218), .ZN(n14767) );
  OR2_X1 U11824 ( .A1(n14767), .A2(n9317), .ZN(n9223) );
  INV_X1 U11825 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n14766) );
  NAND2_X1 U11826 ( .A1(n8803), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U11827 ( .A1(n8736), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9219) );
  OAI211_X1 U11828 ( .C1(n14766), .C2(n9257), .A(n9220), .B(n9219), .ZN(n9221)
         );
  INV_X1 U11829 ( .A(n9221), .ZN(n9222) );
  XNOR2_X1 U11830 ( .A(n9225), .B(n9224), .ZN(n12123) );
  NAND2_X1 U11831 ( .A1(n12123), .A2(n8870), .ZN(n9227) );
  OR2_X1 U11832 ( .A1(n9324), .A2(n12126), .ZN(n9226) );
  MUX2_X1 U11833 ( .A(n14747), .B(n14765), .S(n9330), .Z(n9231) );
  NAND2_X1 U11834 ( .A1(n9230), .A2(n9231), .ZN(n9229) );
  MUX2_X1 U11835 ( .A(n14747), .B(n14765), .S(n8760), .Z(n9228) );
  NAND2_X1 U11836 ( .A1(n9229), .A2(n9228), .ZN(n9235) );
  INV_X1 U11837 ( .A(n9231), .ZN(n9232) );
  NAND2_X1 U11838 ( .A1(n9233), .A2(n9232), .ZN(n9234) );
  AND2_X1 U11839 ( .A1(n9236), .A2(n14527), .ZN(n9237) );
  OR2_X1 U11840 ( .A1(n9252), .A2(n9237), .ZN(n14529) );
  NAND2_X1 U11841 ( .A1(n14749), .A2(n9238), .ZN(n9243) );
  INV_X1 U11842 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n15569) );
  NAND2_X1 U11843 ( .A1(n8803), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9240) );
  NAND2_X1 U11844 ( .A1(n9314), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9239) );
  OAI211_X1 U11845 ( .C1(n15569), .C2(n9257), .A(n9240), .B(n9239), .ZN(n9241)
         );
  INV_X1 U11846 ( .A(n9241), .ZN(n9242) );
  AND2_X2 U11847 ( .A1(n9243), .A2(n9242), .ZN(n10365) );
  XNOR2_X1 U11848 ( .A(n9244), .B(SI_26_), .ZN(n9245) );
  NAND2_X1 U11849 ( .A1(n12351), .A2(n9286), .ZN(n9248) );
  OR2_X1 U11850 ( .A1(n9324), .A2(n15628), .ZN(n9247) );
  MUX2_X1 U11851 ( .A(n14551), .B(n14753), .S(n8760), .Z(n9250) );
  MUX2_X1 U11852 ( .A(n14551), .B(n14753), .S(n9330), .Z(n9249) );
  OR2_X1 U11853 ( .A1(n9252), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U11854 ( .A1(n9254), .A2(n9253), .ZN(n14367) );
  OR2_X1 U11855 ( .A1(n14367), .A2(n9317), .ZN(n9260) );
  INV_X1 U11856 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n12398) );
  NAND2_X1 U11857 ( .A1(n9314), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9256) );
  NAND2_X1 U11858 ( .A1(n8803), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9255) );
  OAI211_X1 U11859 ( .C1(n12398), .C2(n9257), .A(n9256), .B(n9255), .ZN(n9258)
         );
  INV_X1 U11860 ( .A(n9258), .ZN(n9259) );
  XNOR2_X1 U11861 ( .A(n9261), .B(SI_27_), .ZN(n9262) );
  NAND2_X1 U11862 ( .A1(n12378), .A2(n9286), .ZN(n9265) );
  OR2_X1 U11863 ( .A1(n9324), .A2(n12379), .ZN(n9264) );
  MUX2_X1 U11864 ( .A(n14748), .B(n10373), .S(n9330), .Z(n9267) );
  MUX2_X1 U11865 ( .A(n14748), .B(n10373), .S(n9151), .Z(n9266) );
  INV_X1 U11866 ( .A(n9267), .ZN(n9268) );
  INV_X1 U11867 ( .A(n9271), .ZN(n9273) );
  MUX2_X1 U11868 ( .A(n12472), .B(n10364), .S(n8760), .Z(n9269) );
  INV_X1 U11869 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14353) );
  INV_X1 U11870 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15158) );
  MUX2_X1 U11871 ( .A(n14353), .B(n15158), .S(n9277), .Z(n9278) );
  XNOR2_X1 U11872 ( .A(n9278), .B(SI_29_), .ZN(n9322) );
  INV_X1 U11873 ( .A(SI_29_), .ZN(n15777) );
  MUX2_X1 U11874 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6546), .Z(n9279) );
  NAND2_X1 U11875 ( .A1(n9279), .A2(SI_30_), .ZN(n9282) );
  INV_X1 U11876 ( .A(n9279), .ZN(n9280) );
  INV_X1 U11877 ( .A(SI_30_), .ZN(n15606) );
  NAND2_X1 U11878 ( .A1(n9280), .A2(n15606), .ZN(n9281) );
  NAND2_X1 U11879 ( .A1(n9282), .A2(n9281), .ZN(n9292) );
  MUX2_X1 U11880 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6545), .Z(n9283) );
  XNOR2_X1 U11881 ( .A(n9283), .B(SI_31_), .ZN(n9284) );
  NAND2_X1 U11882 ( .A1(n15156), .A2(n9286), .ZN(n9288) );
  INV_X1 U11883 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15682) );
  OR2_X1 U11884 ( .A1(n9324), .A2(n15682), .ZN(n9287) );
  INV_X1 U11885 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n15555) );
  NAND2_X1 U11886 ( .A1(n8736), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9290) );
  INV_X1 U11887 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15782) );
  OR2_X1 U11888 ( .A1(n9316), .A2(n15782), .ZN(n9289) );
  OAI211_X1 U11889 ( .C1(n9257), .C2(n15555), .A(n9290), .B(n9289), .ZN(n14719) );
  XNOR2_X1 U11890 ( .A(n14717), .B(n14719), .ZN(n9353) );
  OR2_X1 U11891 ( .A1(n8984), .A2(n10107), .ZN(n11349) );
  AND2_X1 U11892 ( .A1(n9520), .A2(n11544), .ZN(n9477) );
  OR2_X1 U11893 ( .A1(n10539), .A2(n9477), .ZN(n9291) );
  NAND2_X1 U11894 ( .A1(n11349), .A2(n9291), .ZN(n9332) );
  INV_X1 U11895 ( .A(n9332), .ZN(n9345) );
  NAND2_X1 U11896 ( .A1(n9353), .A2(n9345), .ZN(n9350) );
  NAND2_X1 U11897 ( .A1(n9293), .A2(n9292), .ZN(n9294) );
  INV_X1 U11898 ( .A(n13800), .ZN(n9297) );
  INV_X1 U11899 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12554) );
  OR2_X1 U11900 ( .A1(n9324), .A2(n12554), .ZN(n9298) );
  INV_X1 U11901 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U11902 ( .A1(n8736), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9301) );
  NAND2_X1 U11903 ( .A1(n8803), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9300) );
  OAI211_X1 U11904 ( .C1(n9257), .C2(n9302), .A(n9301), .B(n9300), .ZN(n14548)
         );
  OAI21_X1 U11905 ( .B1(n14719), .B2(n11544), .A(n14548), .ZN(n9303) );
  INV_X1 U11906 ( .A(n14719), .ZN(n9306) );
  OR2_X1 U11907 ( .A1(n9307), .A2(n9306), .ZN(n9331) );
  XNOR2_X1 U11908 ( .A(n8984), .B(n15165), .ZN(n9309) );
  NAND2_X1 U11909 ( .A1(n9309), .A2(n12384), .ZN(n9311) );
  INV_X1 U11910 ( .A(n14548), .ZN(n9310) );
  AOI21_X1 U11911 ( .B1(n9331), .B2(n9311), .A(n9310), .ZN(n9312) );
  AOI21_X1 U11912 ( .B1(n14725), .B2(n8760), .A(n9312), .ZN(n9337) );
  NAND2_X1 U11913 ( .A1(n9314), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9321) );
  NAND2_X1 U11914 ( .A1(n9315), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9320) );
  INV_X1 U11915 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n15693) );
  OR2_X1 U11916 ( .A1(n9316), .A2(n15693), .ZN(n9319) );
  OR2_X1 U11917 ( .A1(n9317), .A2(n12485), .ZN(n9318) );
  NAND4_X1 U11918 ( .A1(n9321), .A2(n9320), .A3(n9319), .A4(n9318), .ZN(n14549) );
  NAND2_X1 U11919 ( .A1(n14352), .A2(n8870), .ZN(n9326) );
  OR2_X1 U11920 ( .A1(n9324), .A2(n15158), .ZN(n9325) );
  MUX2_X1 U11921 ( .A(n14549), .B(n12491), .S(n9151), .Z(n9334) );
  INV_X1 U11922 ( .A(n9334), .ZN(n9327) );
  NAND2_X1 U11923 ( .A1(n9327), .A2(n9333), .ZN(n9328) );
  NAND2_X1 U11924 ( .A1(n12384), .A2(n9521), .ZN(n9375) );
  AND2_X1 U11925 ( .A1(n9332), .A2(n9375), .ZN(n9341) );
  NAND2_X1 U11926 ( .A1(n9338), .A2(n9337), .ZN(n9336) );
  NAND2_X1 U11927 ( .A1(n9336), .A2(n9335), .ZN(n9340) );
  OR2_X1 U11928 ( .A1(n9338), .A2(n9337), .ZN(n9339) );
  NAND2_X1 U11929 ( .A1(n9340), .A2(n9339), .ZN(n9346) );
  INV_X1 U11930 ( .A(n9346), .ZN(n9351) );
  INV_X1 U11931 ( .A(n9341), .ZN(n9342) );
  OAI21_X1 U11932 ( .B1(n9353), .B2(n9342), .A(n9344), .ZN(n9343) );
  OAI21_X1 U11933 ( .B1(n9345), .B2(n9344), .A(n9343), .ZN(n9349) );
  OAI211_X1 U11934 ( .C1(n9351), .C2(n9350), .A(n9349), .B(n9348), .ZN(n9352)
         );
  XNOR2_X1 U11935 ( .A(n14725), .B(n14548), .ZN(n9373) );
  NAND2_X1 U11936 ( .A1(n14738), .A2(n10364), .ZN(n9513) );
  OR2_X1 U11937 ( .A1(n14738), .A2(n10364), .ZN(n9354) );
  NAND2_X1 U11938 ( .A1(n9513), .A2(n9354), .ZN(n10352) );
  XNOR2_X2 U11939 ( .A(n14753), .B(n10365), .ZN(n14744) );
  XNOR2_X1 U11940 ( .A(n15117), .B(n9507), .ZN(n14773) );
  XNOR2_X1 U11941 ( .A(n14800), .B(n14553), .ZN(n14806) );
  INV_X1 U11942 ( .A(n14806), .ZN(n14793) );
  XNOR2_X1 U11943 ( .A(n14817), .B(n14554), .ZN(n14820) );
  XNOR2_X1 U11944 ( .A(n9519), .B(n14555), .ZN(n14827) );
  NAND2_X1 U11945 ( .A1(n14858), .A2(n14401), .ZN(n9355) );
  NAND2_X1 U11946 ( .A1(n15048), .A2(n14910), .ZN(n9502) );
  NAND2_X1 U11947 ( .A1(n14870), .A2(n9502), .ZN(n14895) );
  XNOR2_X1 U11948 ( .A(n14507), .B(n14561), .ZN(n11873) );
  XNOR2_X1 U11949 ( .A(n10177), .B(n11861), .ZN(n11497) );
  CLKBUF_X1 U11950 ( .A(n9357), .Z(n9432) );
  NOR2_X1 U11951 ( .A1(n9432), .A2(n15275), .ZN(n9359) );
  NOR2_X1 U11952 ( .A1(n14568), .A2(n14464), .ZN(n9437) );
  NAND2_X1 U11953 ( .A1(n14568), .A2(n14464), .ZN(n9436) );
  INV_X1 U11954 ( .A(n9436), .ZN(n9358) );
  OR2_X1 U11955 ( .A1(n9437), .A2(n9358), .ZN(n11303) );
  AND4_X1 U11956 ( .A1(n9360), .A2(n9359), .A3(n11303), .A4(n11347), .ZN(n9361) );
  XNOR2_X1 U11957 ( .A(n15251), .B(n11491), .ZN(n11939) );
  XNOR2_X1 U11958 ( .A(n14567), .B(n11576), .ZN(n11587) );
  XNOR2_X1 U11959 ( .A(n11605), .B(n14566), .ZN(n11394) );
  NAND4_X1 U11960 ( .A1(n9361), .A2(n11939), .A3(n11587), .A4(n11394), .ZN(
        n9362) );
  NOR2_X1 U11961 ( .A1(n11497), .A2(n9362), .ZN(n9364) );
  XNOR2_X1 U11962 ( .A(n15096), .B(n12206), .ZN(n11517) );
  INV_X1 U11963 ( .A(n11517), .ZN(n9363) );
  AND4_X1 U11964 ( .A1(n11873), .A2(n9364), .A3(n9363), .A4(n7782), .ZN(n9365)
         );
  XNOR2_X1 U11965 ( .A(n14984), .B(n14559), .ZN(n9494) );
  XNOR2_X1 U11966 ( .A(n14974), .B(n14560), .ZN(n12053) );
  AND4_X1 U11967 ( .A1(n14967), .A2(n9365), .A3(n9494), .A4(n12053), .ZN(n9367) );
  XNOR2_X1 U11968 ( .A(n15055), .B(n14925), .ZN(n14901) );
  OR2_X1 U11969 ( .A1(n15060), .A2(n14941), .ZN(n9458) );
  NAND2_X1 U11970 ( .A1(n15060), .A2(n14941), .ZN(n9366) );
  INV_X1 U11971 ( .A(n14918), .ZN(n14922) );
  NAND4_X1 U11972 ( .A1(n14827), .A2(n14855), .A3(n9369), .A4(n9368), .ZN(
        n9370) );
  NOR4_X1 U11973 ( .A1(n10352), .A2(n14744), .A3(n14761), .A4(n9371), .ZN(
        n9372) );
  XNOR2_X1 U11974 ( .A(n12491), .B(n14549), .ZN(n9515) );
  XNOR2_X1 U11975 ( .A(n9374), .B(n14731), .ZN(n9377) );
  INV_X1 U11976 ( .A(n9375), .ZN(n9376) );
  INV_X1 U11977 ( .A(n9384), .ZN(n9381) );
  NAND2_X1 U11978 ( .A1(n9381), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9382) );
  MUX2_X1 U11979 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9382), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9385) );
  NAND2_X1 U11980 ( .A1(n9385), .A2(n9389), .ZN(n10538) );
  OR2_X1 U11981 ( .A1(n10538), .A2(P1_U3086), .ZN(n11926) );
  NAND2_X1 U11982 ( .A1(n8984), .A2(n11544), .ZN(n9524) );
  NAND2_X1 U11983 ( .A1(n9524), .A2(n10539), .ZN(n9545) );
  NAND2_X1 U11984 ( .A1(n9389), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9388) );
  NAND2_X1 U11985 ( .A1(n9391), .A2(n9390), .ZN(n9397) );
  NAND2_X1 U11986 ( .A1(n8724), .A2(n9395), .ZN(n9399) );
  NAND2_X1 U11987 ( .A1(n9399), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9396) );
  NOR2_X1 U11988 ( .A1(n12106), .A2(n9532), .ZN(n9401) );
  NAND2_X1 U11989 ( .A1(n9397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9398) );
  AND2_X1 U11990 ( .A1(n10409), .A2(n10538), .ZN(n9402) );
  AND2_X1 U11991 ( .A1(n9545), .A2(n9402), .ZN(n10333) );
  NOR2_X1 U11992 ( .A1(n14586), .A2(P1_U3086), .ZN(n9405) );
  NAND3_X1 U11993 ( .A1(n10333), .A2(n14939), .A3(n9405), .ZN(n9406) );
  OAI211_X1 U11994 ( .C1(n15165), .C2(n11926), .A(n9406), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9407) );
  INV_X1 U11995 ( .A(n13120), .ZN(n9428) );
  OAI22_X1 U11996 ( .A1(n15512), .A2(n9409), .B1(n12579), .B2(n9408), .ZN(
        n9410) );
  INV_X1 U11997 ( .A(n12760), .ZN(n9412) );
  NAND2_X1 U11998 ( .A1(n9410), .A2(n9412), .ZN(n9411) );
  NAND2_X1 U11999 ( .A1(n9411), .A2(n12742), .ZN(n9413) );
  AOI21_X1 U12000 ( .B1(n9414), .B2(n9413), .A(n11532), .ZN(n9417) );
  NOR2_X1 U12001 ( .A1(n12752), .A2(n9415), .ZN(n11530) );
  NAND2_X1 U12002 ( .A1(n13471), .A2(n11530), .ZN(n9416) );
  NAND3_X1 U12003 ( .A1(n9418), .A2(n9417), .A3(n9416), .ZN(n9422) );
  AND2_X1 U12004 ( .A1(n9419), .A2(n11245), .ZN(n9420) );
  NAND2_X1 U12005 ( .A1(n9421), .A2(n9420), .ZN(n11531) );
  NOR2_X1 U12006 ( .A1(n15549), .A2(n9423), .ZN(n9424) );
  NAND2_X1 U12007 ( .A1(n11444), .A2(n11445), .ZN(n9431) );
  NAND2_X1 U12008 ( .A1(n9429), .A2(n10117), .ZN(n9430) );
  NAND2_X1 U12009 ( .A1(n9431), .A2(n9430), .ZN(n11351) );
  INV_X1 U12010 ( .A(n9433), .ZN(n10136) );
  NAND2_X1 U12011 ( .A1(n10136), .A2(n15306), .ZN(n9434) );
  INV_X1 U12012 ( .A(n14569), .ZN(n10144) );
  NAND2_X1 U12013 ( .A1(n10144), .A2(n15315), .ZN(n9435) );
  INV_X1 U12014 ( .A(n11584), .ZN(n9439) );
  NAND2_X1 U12015 ( .A1(n11396), .A2(n15262), .ZN(n9440) );
  NAND2_X1 U12016 ( .A1(n11582), .A2(n9440), .ZN(n11387) );
  AOI22_X1 U12017 ( .A1(n10177), .A2(n14564), .B1(n14565), .B2(n9489), .ZN(
        n9447) );
  NAND2_X1 U12018 ( .A1(n11605), .A2(n14566), .ZN(n9441) );
  NOR2_X1 U12019 ( .A1(n11605), .A2(n14566), .ZN(n11484) );
  NAND2_X1 U12020 ( .A1(n15251), .A2(n11491), .ZN(n11486) );
  NAND2_X1 U12021 ( .A1(n11486), .A2(n14564), .ZN(n9443) );
  NAND2_X1 U12022 ( .A1(n15336), .A2(n9443), .ZN(n9445) );
  NAND3_X1 U12023 ( .A1(n15251), .A2(n11491), .A3(n11861), .ZN(n9444) );
  NAND2_X1 U12024 ( .A1(n9445), .A2(n9444), .ZN(n9446) );
  AOI21_X1 U12025 ( .B1(n9447), .B2(n11484), .A(n9446), .ZN(n9448) );
  NAND2_X1 U12026 ( .A1(n12205), .A2(n11522), .ZN(n9450) );
  NAND2_X1 U12027 ( .A1(n12301), .A2(n12206), .ZN(n9451) );
  NAND2_X1 U12028 ( .A1(n11513), .A2(n9451), .ZN(n11879) );
  INV_X1 U12029 ( .A(n11873), .ZN(n11878) );
  NAND2_X1 U12030 ( .A1(n11879), .A2(n11878), .ZN(n11877) );
  OR2_X1 U12031 ( .A1(n14507), .A2(n14561), .ZN(n9452) );
  NAND2_X1 U12032 ( .A1(n11877), .A2(n9452), .ZN(n12057) );
  OR2_X1 U12033 ( .A1(n14974), .A2(n14560), .ZN(n9453) );
  NAND2_X1 U12034 ( .A1(n12056), .A2(n9453), .ZN(n14983) );
  INV_X1 U12035 ( .A(n9494), .ZN(n14982) );
  OR2_X1 U12036 ( .A1(n14984), .A2(n14559), .ZN(n9454) );
  INV_X1 U12037 ( .A(n14952), .ZN(n9457) );
  INV_X1 U12038 ( .A(n14480), .ZN(n14938) );
  NAND2_X1 U12039 ( .A1(n14957), .A2(n14938), .ZN(n9455) );
  INV_X1 U12040 ( .A(n9455), .ZN(n14950) );
  NOR2_X1 U12041 ( .A1(n15055), .A2(n14925), .ZN(n9460) );
  NAND2_X1 U12042 ( .A1(n15055), .A2(n14925), .ZN(n9459) );
  OR2_X1 U12043 ( .A1(n14875), .A2(n14557), .ZN(n14851) );
  INV_X1 U12044 ( .A(n14855), .ZN(n9463) );
  AND2_X1 U12045 ( .A1(n14851), .A2(n9463), .ZN(n9464) );
  NAND2_X1 U12046 ( .A1(n14858), .A2(n14556), .ZN(n9465) );
  OR2_X1 U12047 ( .A1(n9519), .A2(n14555), .ZN(n9466) );
  NAND2_X1 U12048 ( .A1(n14817), .A2(n10269), .ZN(n9467) );
  NAND2_X1 U12049 ( .A1(n14800), .A2(n14553), .ZN(n9468) );
  INV_X1 U12050 ( .A(n14773), .ZN(n14778) );
  OR2_X1 U12051 ( .A1(n15117), .A2(n14552), .ZN(n9469) );
  AND2_X2 U12052 ( .A1(n14781), .A2(n9469), .ZN(n14758) );
  NAND2_X1 U12053 ( .A1(n14765), .A2(n14747), .ZN(n9470) );
  AND2_X1 U12054 ( .A1(n14753), .A2(n14551), .ZN(n9471) );
  OR2_X1 U12055 ( .A1(n10373), .A2(n14748), .ZN(n9472) );
  INV_X1 U12056 ( .A(n10352), .ZN(n10346) );
  XNOR2_X1 U12057 ( .A(n9473), .B(n9515), .ZN(n12498) );
  INV_X1 U12058 ( .A(n12498), .ZN(n9478) );
  NAND2_X1 U12059 ( .A1(n8984), .A2(n15165), .ZN(n9474) );
  NAND2_X1 U12060 ( .A1(n9474), .A2(n10107), .ZN(n10134) );
  OR2_X1 U12062 ( .A1(n10107), .A2(n9520), .ZN(n9475) );
  AND2_X1 U12063 ( .A1(n8984), .A2(n9475), .ZN(n9476) );
  NAND2_X1 U12064 ( .A1(n10270), .A2(n9476), .ZN(n11940) );
  NAND2_X1 U12065 ( .A1(n14731), .A2(n9477), .ZN(n15310) );
  NAND2_X1 U12066 ( .A1(n9478), .A2(n15339), .ZN(n9528) );
  AND2_X1 U12067 ( .A1(n9482), .A2(n9481), .ZN(n11361) );
  NAND2_X1 U12068 ( .A1(n11361), .A2(n11360), .ZN(n11359) );
  NAND2_X1 U12069 ( .A1(n11359), .A2(n15274), .ZN(n9484) );
  NAND2_X1 U12070 ( .A1(n15322), .A2(n14568), .ZN(n9486) );
  NAND2_X1 U12071 ( .A1(n10150), .A2(n14464), .ZN(n11585) );
  INV_X1 U12072 ( .A(n14566), .ZN(n11548) );
  NAND2_X1 U12073 ( .A1(n11548), .A2(n11605), .ZN(n9487) );
  NAND2_X1 U12074 ( .A1(n15251), .A2(n14565), .ZN(n9488) );
  NAND2_X1 U12075 ( .A1(n9489), .A2(n11491), .ZN(n9490) );
  INV_X1 U12076 ( .A(n11497), .ZN(n9491) );
  OR2_X2 U12077 ( .A1(n11518), .A2(n11517), .ZN(n11516) );
  NAND2_X1 U12078 ( .A1(n12301), .A2(n14562), .ZN(n9492) );
  INV_X1 U12079 ( .A(n14561), .ZN(n10200) );
  OR2_X1 U12080 ( .A1(n14507), .A2(n10200), .ZN(n9493) );
  OR2_X1 U12081 ( .A1(n14974), .A2(n10201), .ZN(n14978) );
  OR2_X1 U12082 ( .A1(n14984), .A2(n14377), .ZN(n14960) );
  INV_X1 U12083 ( .A(n14941), .ZN(n14908) );
  NAND2_X1 U12084 ( .A1(n15060), .A2(n14908), .ZN(n9497) );
  NOR2_X1 U12085 ( .A1(n15055), .A2(n14884), .ZN(n14869) );
  NAND2_X1 U12086 ( .A1(n9502), .A2(n14869), .ZN(n9498) );
  AND2_X1 U12087 ( .A1(n9498), .A2(n14870), .ZN(n9499) );
  NAND2_X1 U12088 ( .A1(n15055), .A2(n14884), .ZN(n9501) );
  AND2_X1 U12089 ( .A1(n9502), .A2(n9501), .ZN(n14844) );
  NAND2_X1 U12090 ( .A1(n14875), .A2(n14885), .ZN(n14846) );
  INV_X1 U12091 ( .A(n14555), .ZN(n10264) );
  OR2_X1 U12092 ( .A1(n9519), .A2(n10264), .ZN(n9503) );
  OR2_X1 U12093 ( .A1(n14817), .A2(n14554), .ZN(n9504) );
  INV_X1 U12094 ( .A(n14553), .ZN(n9505) );
  NAND2_X1 U12095 ( .A1(n14800), .A2(n9505), .ZN(n9506) );
  OR2_X1 U12096 ( .A1(n15117), .A2(n9507), .ZN(n9508) );
  NAND2_X1 U12097 ( .A1(n14765), .A2(n9509), .ZN(n9510) );
  AND2_X1 U12098 ( .A1(n14753), .A2(n10365), .ZN(n9512) );
  OR2_X1 U12099 ( .A1(n14753), .A2(n10365), .ZN(n9511) );
  INV_X1 U12100 ( .A(n14748), .ZN(n14532) );
  NAND2_X1 U12101 ( .A1(n10373), .A2(n14532), .ZN(n10351) );
  AOI21_X2 U12102 ( .B1(n10361), .B2(n10351), .A(n10352), .ZN(n10355) );
  INV_X1 U12103 ( .A(n9513), .ZN(n9514) );
  NAND2_X1 U12104 ( .A1(n14731), .A2(n15165), .ZN(n9517) );
  NAND2_X1 U12105 ( .A1(n9308), .A2(n9521), .ZN(n9516) );
  NAND2_X1 U12106 ( .A1(n10117), .A2(n11343), .ZN(n11443) );
  INV_X1 U12107 ( .A(n15306), .ZN(n11362) );
  NAND2_X1 U12108 ( .A1(n11880), .A2(n15087), .ZN(n14975) );
  AND2_X2 U12109 ( .A1(n14856), .A2(n15127), .ZN(n14834) );
  AND2_X2 U12110 ( .A1(n14746), .A2(n15002), .ZN(n10371) );
  AND2_X2 U12111 ( .A1(n10371), .A2(n15110), .ZN(n10372) );
  NAND2_X1 U12112 ( .A1(n9520), .A2(n12384), .ZN(n10863) );
  AOI21_X1 U12113 ( .B1(n12491), .B2(n10350), .A(n15323), .ZN(n9522) );
  NAND2_X1 U12114 ( .A1(n9522), .A2(n14724), .ZN(n12494) );
  INV_X1 U12115 ( .A(n10863), .ZN(n9523) );
  NAND2_X1 U12116 ( .A1(n12491), .A2(n15295), .ZN(n9527) );
  OR2_X1 U12117 ( .A1(n10364), .A2(n14907), .ZN(n12488) );
  INV_X1 U12118 ( .A(n15163), .ZN(n14587) );
  INV_X1 U12119 ( .A(n14586), .ZN(n15236) );
  AND2_X1 U12120 ( .A1(n15236), .A2(P1_B_REG_SCAN_IN), .ZN(n9526) );
  NOR2_X1 U12121 ( .A1(n14909), .A2(n9526), .ZN(n14720) );
  NAND2_X1 U12122 ( .A1(n14720), .A2(n14548), .ZN(n12486) );
  NAND3_X1 U12123 ( .A1(n12128), .A2(P1_B_REG_SCAN_IN), .A3(n12106), .ZN(n9531) );
  OAI21_X1 U12124 ( .B1(n12106), .B2(P1_B_REG_SCAN_IN), .A(n10532), .ZN(n9529)
         );
  INV_X1 U12125 ( .A(n9529), .ZN(n9530) );
  NAND2_X1 U12126 ( .A1(n12128), .A2(n9532), .ZN(n9533) );
  NAND2_X1 U12127 ( .A1(n9534), .A2(n9533), .ZN(n10319) );
  NOR2_X1 U12128 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n15550) );
  NOR4_X1 U12129 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n9537) );
  NOR4_X1 U12130 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9536) );
  NOR4_X1 U12131 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n9535) );
  AND4_X1 U12132 ( .A1(n15550), .A2(n9537), .A3(n9536), .A4(n9535), .ZN(n9543)
         );
  NOR4_X1 U12133 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9541) );
  NOR4_X1 U12134 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9540) );
  NOR4_X1 U12135 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9539) );
  NOR4_X1 U12136 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9538) );
  AND4_X1 U12137 ( .A1(n9541), .A2(n9540), .A3(n9539), .A4(n9538), .ZN(n9542)
         );
  AND2_X1 U12138 ( .A1(n9543), .A2(n9542), .ZN(n9544) );
  NAND2_X1 U12139 ( .A1(n10536), .A2(n9545), .ZN(n10853) );
  NAND2_X1 U12140 ( .A1(n12106), .A2(n9532), .ZN(n10553) );
  NOR2_X1 U12141 ( .A1(n10853), .A2(n11297), .ZN(n9547) );
  NAND2_X1 U12142 ( .A1(n9553), .A2(n15348), .ZN(n9550) );
  NAND2_X1 U12143 ( .A1(n9548), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U12144 ( .A1(n9550), .A2(n9549), .ZN(P1_U3557) );
  INV_X1 U12145 ( .A(n11297), .ZN(n10320) );
  NOR2_X1 U12146 ( .A1(n10320), .A2(n10853), .ZN(n9552) );
  NAND2_X1 U12147 ( .A1(n9553), .A2(n15342), .ZN(n9556) );
  NAND2_X1 U12148 ( .A1(n9554), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9555) );
  NAND2_X1 U12149 ( .A1(n9556), .A2(n9555), .ZN(P1_U3525) );
  INV_X4 U12150 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U12151 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n9557) );
  NAND2_X1 U12152 ( .A1(n9577), .A2(n9557), .ZN(n9561) );
  NAND4_X1 U12153 ( .A1(n9560), .A2(n9559), .A3(n9558), .A4(n9829), .ZN(n9578)
         );
  NOR2_X2 U12154 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n9589) );
  NAND2_X1 U12155 ( .A1(n9601), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9569) );
  MUX2_X1 U12156 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9569), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n9571) );
  INV_X1 U12157 ( .A(n10051), .ZN(n9570) );
  NAND2_X1 U12158 ( .A1(n9603), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9572) );
  XNOR2_X2 U12159 ( .A(n9572), .B(n9584), .ZN(n13833) );
  INV_X1 U12160 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9573) );
  INV_X1 U12161 ( .A(n13643), .ZN(n9581) );
  NAND2_X1 U12162 ( .A1(n9581), .A2(n13884), .ZN(n9575) );
  NAND2_X1 U12163 ( .A1(n13836), .A2(n9575), .ZN(n9580) );
  NAND2_X1 U12164 ( .A1(n9576), .A2(n9577), .ZN(n9794) );
  NAND2_X2 U12165 ( .A1(n9580), .A2(n14152), .ZN(n10685) );
  INV_X1 U12166 ( .A(n12473), .ZN(n9587) );
  INV_X2 U12167 ( .A(n9603), .ZN(n9605) );
  NOR2_X1 U12168 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n9583) );
  NOR2_X1 U12169 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n9582) );
  NAND3_X1 U12170 ( .A1(n9583), .A2(n9582), .A3(n10076), .ZN(n9597) );
  NAND2_X1 U12171 ( .A1(n9584), .A2(n14345), .ZN(n9585) );
  NOR2_X2 U12172 ( .A1(n9597), .A2(n9585), .ZN(n9604) );
  INV_X1 U12173 ( .A(n9604), .ZN(n9608) );
  NOR2_X2 U12174 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n9606) );
  INV_X1 U12175 ( .A(n9606), .ZN(n14347) );
  NAND2_X1 U12176 ( .A1(n9606), .A2(n9573), .ZN(n9586) );
  NAND2_X1 U12177 ( .A1(n9587), .A2(n6544), .ZN(n9594) );
  NAND2_X1 U12178 ( .A1(n9663), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n9593) );
  MUX2_X1 U12179 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9588), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9590) );
  INV_X1 U12180 ( .A(n9589), .ZN(n9630) );
  NAND3_X2 U12181 ( .A1(n9594), .A2(n9593), .A3(n9592), .ZN(n10871) );
  AND2_X4 U12182 ( .A1(n10826), .A2(n13833), .ZN(n14308) );
  NOR2_X1 U12183 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n9595) );
  INV_X1 U12184 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14344) );
  NAND3_X1 U12185 ( .A1(n9606), .A2(n9595), .A3(P2_IR_REG_30__SCAN_IN), .ZN(
        n9598) );
  XNOR2_X1 U12186 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_30__SCAN_IN), .ZN(
        n9596) );
  OAI21_X1 U12187 ( .B1(n9598), .B2(n9597), .A(n9596), .ZN(n9599) );
  NAND3_X1 U12188 ( .A1(n9601), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_30__SCAN_IN), .ZN(n9602) );
  NAND3_X1 U12189 ( .A1(n9603), .A2(P2_IR_REG_31__SCAN_IN), .A3(n14343), .ZN(
        n9613) );
  NAND2_X1 U12190 ( .A1(n9606), .A2(n14343), .ZN(n9607) );
  NOR2_X1 U12191 ( .A1(n9608), .A2(n9607), .ZN(n9610) );
  XNOR2_X1 U12192 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_29__SCAN_IN), .ZN(
        n9609) );
  NAND2_X1 U12193 ( .A1(n9653), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9617) );
  NAND2_X1 U12194 ( .A1(n6548), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U12195 ( .A1(n9674), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9615) );
  AND2_X2 U12196 ( .A1(n12388), .A2(n14354), .ZN(n9655) );
  NAND2_X1 U12197 ( .A1(n9655), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9614) );
  NAND2_X1 U12198 ( .A1(n9652), .A2(n6543), .ZN(n9627) );
  INV_X1 U12199 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10676) );
  OR2_X1 U12200 ( .A1(n6537), .A2(n11717), .ZN(n9625) );
  NAND2_X1 U12201 ( .A1(n6548), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U12202 ( .A1(n9674), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9622) );
  NAND2_X1 U12203 ( .A1(n9652), .A2(n10865), .ZN(n9624) );
  INV_X1 U12204 ( .A(n9626), .ZN(n9628) );
  NAND2_X1 U12205 ( .A1(n9628), .A2(n9627), .ZN(n10992) );
  NAND2_X1 U12206 ( .A1(n10490), .A2(n6544), .ZN(n9636) );
  NAND2_X1 U12207 ( .A1(n9630), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9631) );
  MUX2_X1 U12208 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9631), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n9633) );
  INV_X1 U12209 ( .A(n9632), .ZN(n9647) );
  NAND2_X1 U12210 ( .A1(n9633), .A2(n9647), .ZN(n15350) );
  INV_X1 U12211 ( .A(n15350), .ZN(n10620) );
  AND2_X1 U12212 ( .A1(n9732), .A2(n10620), .ZN(n9634) );
  XNOR2_X1 U12213 ( .A(n6537), .B(n10867), .ZN(n9641) );
  NAND2_X1 U12214 ( .A1(n9653), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U12215 ( .A1(n6548), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9639) );
  NAND2_X1 U12216 ( .A1(n9674), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U12217 ( .A1(n9655), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9637) );
  XNOR2_X1 U12218 ( .A(n9641), .B(n9642), .ZN(n10991) );
  INV_X1 U12219 ( .A(n9641), .ZN(n9643) );
  NAND2_X1 U12220 ( .A1(n9643), .A2(n9642), .ZN(n9644) );
  NAND2_X1 U12221 ( .A1(n10486), .A2(n6544), .ZN(n9651) );
  NAND2_X1 U12222 ( .A1(n9647), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9646) );
  MUX2_X1 U12223 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9646), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9648) );
  AND2_X1 U12224 ( .A1(n9732), .A2(n10649), .ZN(n9649) );
  AOI21_X1 U12225 ( .B1(n9913), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n9649), .ZN(
        n9650) );
  XNOR2_X1 U12226 ( .A(n6537), .B(n13662), .ZN(n9661) );
  BUF_X1 U12227 ( .A(n9652), .Z(n9981) );
  NAND2_X1 U12228 ( .A1(n9653), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9659) );
  INV_X1 U12229 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9685) );
  NAND2_X1 U12230 ( .A1(n9973), .A2(n9685), .ZN(n9658) );
  INV_X1 U12231 ( .A(n9707), .ZN(n10028) );
  NAND2_X1 U12232 ( .A1(n10028), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9657) );
  NAND2_X1 U12233 ( .A1(n9655), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9656) );
  NAND4_X2 U12234 ( .A1(n9659), .A2(n9658), .A3(n9657), .A4(n9656), .ZN(n13905) );
  AND2_X1 U12235 ( .A1(n9652), .A2(n13905), .ZN(n9660) );
  NAND2_X1 U12236 ( .A1(n9661), .A2(n9660), .ZN(n11007) );
  OR2_X1 U12237 ( .A1(n9661), .A2(n9660), .ZN(n9662) );
  NAND2_X1 U12238 ( .A1(n11007), .A2(n9662), .ZN(n11111) );
  NAND2_X1 U12239 ( .A1(n10492), .A2(n6550), .ZN(n9670) );
  INV_X1 U12240 ( .A(n9679), .ZN(n9665) );
  INV_X1 U12241 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9664) );
  NAND2_X1 U12242 ( .A1(n9665), .A2(n9664), .ZN(n9681) );
  NAND2_X1 U12243 ( .A1(n9681), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9666) );
  MUX2_X1 U12244 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9666), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9667) );
  AOI22_X1 U12245 ( .A1(n9913), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10664), 
        .B2(n6540), .ZN(n9669) );
  NAND2_X2 U12246 ( .A1(n9670), .A2(n9669), .ZN(n13676) );
  XNOR2_X1 U12247 ( .A(n6537), .B(n13676), .ZN(n9697) );
  NAND2_X1 U12248 ( .A1(n9653), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9678) );
  INV_X1 U12249 ( .A(n9686), .ZN(n9671) );
  INV_X1 U12250 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U12251 ( .A1(n9686), .A2(n9672), .ZN(n9673) );
  AND2_X1 U12252 ( .A1(n9705), .A2(n9673), .ZN(n11081) );
  NAND2_X1 U12253 ( .A1(n9973), .A2(n11081), .ZN(n9677) );
  INV_X1 U12254 ( .A(n9707), .ZN(n10017) );
  NAND2_X1 U12255 ( .A1(n10017), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9676) );
  NAND2_X1 U12256 ( .A1(n9655), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9675) );
  NAND2_X1 U12257 ( .A1(n9652), .A2(n13903), .ZN(n9698) );
  XNOR2_X1 U12258 ( .A(n9697), .B(n9698), .ZN(n11082) );
  NAND2_X1 U12259 ( .A1(n10494), .A2(n6550), .ZN(n9684) );
  NAND2_X1 U12260 ( .A1(n9679), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9680) );
  MUX2_X1 U12261 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9680), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n9682) );
  NAND2_X1 U12262 ( .A1(n9682), .A2(n9681), .ZN(n15362) );
  INV_X1 U12263 ( .A(n15362), .ZN(n10624) );
  AOI22_X1 U12264 ( .A1(n9913), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10624), 
        .B2(n6540), .ZN(n9683) );
  XNOR2_X1 U12265 ( .A(n6537), .B(n13670), .ZN(n9692) );
  NAND2_X1 U12266 ( .A1(n9653), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9691) );
  INV_X1 U12267 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n15586) );
  NAND2_X1 U12268 ( .A1(n15586), .A2(n9685), .ZN(n9687) );
  AND2_X1 U12269 ( .A1(n9687), .A2(n9686), .ZN(n11669) );
  NAND2_X1 U12270 ( .A1(n9973), .A2(n11669), .ZN(n9690) );
  NAND2_X1 U12271 ( .A1(n10017), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9689) );
  NAND2_X1 U12272 ( .A1(n9655), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9688) );
  NAND4_X2 U12273 ( .A1(n9691), .A2(n9690), .A3(n9689), .A4(n9688), .ZN(n13904) );
  NAND2_X1 U12274 ( .A1(n9652), .A2(n13904), .ZN(n9693) );
  XNOR2_X1 U12275 ( .A(n9692), .B(n9693), .ZN(n11006) );
  AND3_X1 U12276 ( .A1(n11082), .A2(n11006), .A3(n11007), .ZN(n9696) );
  INV_X1 U12277 ( .A(n9692), .ZN(n9694) );
  AND2_X1 U12278 ( .A1(n9694), .A2(n9693), .ZN(n11083) );
  AND2_X1 U12279 ( .A1(n11082), .A2(n11083), .ZN(n9695) );
  INV_X1 U12280 ( .A(n9697), .ZN(n9699) );
  NAND2_X1 U12281 ( .A1(n9699), .A2(n9698), .ZN(n9700) );
  NAND2_X1 U12282 ( .A1(n10498), .A2(n13785), .ZN(n9703) );
  NAND2_X1 U12283 ( .A1(n9716), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9701) );
  AOI22_X1 U12284 ( .A1(n9913), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n15377), 
        .B2(n6540), .ZN(n9702) );
  XNOR2_X1 U12285 ( .A(n6537), .B(n15438), .ZN(n9712) );
  NAND2_X1 U12286 ( .A1(n9653), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9711) );
  INV_X1 U12287 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n15374) );
  NAND2_X1 U12288 ( .A1(n9705), .A2(n15374), .ZN(n9706) );
  AND2_X1 U12289 ( .A1(n9721), .A2(n9706), .ZN(n11118) );
  NAND2_X1 U12290 ( .A1(n9973), .A2(n11118), .ZN(n9710) );
  NAND2_X1 U12291 ( .A1(n9655), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9709) );
  INV_X1 U12292 ( .A(n9707), .ZN(n9974) );
  NAND2_X1 U12293 ( .A1(n9974), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9708) );
  NAND4_X1 U12294 ( .A1(n9711), .A2(n9710), .A3(n9709), .A4(n9708), .ZN(n13902) );
  AND2_X1 U12295 ( .A1(n9981), .A2(n13902), .ZN(n9713) );
  NAND2_X1 U12296 ( .A1(n9712), .A2(n9713), .ZN(n9715) );
  OR2_X1 U12297 ( .A1(n9713), .A2(n9712), .ZN(n9714) );
  AND2_X1 U12298 ( .A1(n9715), .A2(n9714), .ZN(n11120) );
  NAND2_X1 U12299 ( .A1(n10523), .A2(n13785), .ZN(n9719) );
  OAI21_X1 U12300 ( .B1(n9716), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9717) );
  XNOR2_X1 U12301 ( .A(n9717), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U12302 ( .A1(n9913), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n13913), 
        .B2(n6540), .ZN(n9718) );
  NAND2_X1 U12303 ( .A1(n9719), .A2(n9718), .ZN(n13687) );
  XNOR2_X1 U12304 ( .A(n13687), .B(n6537), .ZN(n9728) );
  INV_X1 U12305 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11729) );
  NAND2_X1 U12306 ( .A1(n10028), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9720) );
  NAND2_X1 U12307 ( .A1(n9721), .A2(n15585), .ZN(n9722) );
  NAND2_X1 U12308 ( .A1(n9737), .A2(n9722), .ZN(n11731) );
  NAND2_X1 U12309 ( .A1(n9655), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9723) );
  OAI21_X1 U12310 ( .B1(n11731), .B2(n10089), .A(n9723), .ZN(n9724) );
  INV_X1 U12311 ( .A(n9724), .ZN(n9725) );
  NAND2_X1 U12312 ( .A1(n9652), .A2(n13901), .ZN(n9726) );
  XNOR2_X1 U12313 ( .A(n9728), .B(n9726), .ZN(n11166) );
  NAND2_X1 U12314 ( .A1(n11167), .A2(n11166), .ZN(n11165) );
  INV_X1 U12315 ( .A(n9726), .ZN(n9727) );
  NAND2_X1 U12316 ( .A1(n9728), .A2(n9727), .ZN(n9729) );
  NAND2_X1 U12317 ( .A1(n11165), .A2(n9729), .ZN(n11410) );
  INV_X1 U12318 ( .A(n9576), .ZN(n9730) );
  NAND2_X1 U12319 ( .A1(n9730), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9731) );
  XNOR2_X1 U12320 ( .A(n9731), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U12321 ( .A1(n9913), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10707), 
        .B2(n6540), .ZN(n9733) );
  XNOR2_X1 U12322 ( .A(n14314), .B(n10014), .ZN(n9743) );
  INV_X1 U12323 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11742) );
  NAND2_X1 U12324 ( .A1(n9974), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9735) );
  OAI21_X1 U12325 ( .B1(n11742), .B2(n12536), .A(n9735), .ZN(n9736) );
  INV_X1 U12326 ( .A(n9736), .ZN(n9742) );
  NAND2_X1 U12327 ( .A1(n9737), .A2(n15651), .ZN(n9738) );
  NAND2_X1 U12328 ( .A1(n9767), .A2(n9738), .ZN(n11746) );
  NAND2_X1 U12329 ( .A1(n9655), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9739) );
  OAI21_X1 U12330 ( .B1(n11746), .B2(n10089), .A(n9739), .ZN(n9740) );
  INV_X1 U12331 ( .A(n9740), .ZN(n9741) );
  NAND2_X1 U12332 ( .A1(n9652), .A2(n6832), .ZN(n9744) );
  NAND2_X1 U12333 ( .A1(n9743), .A2(n9744), .ZN(n11409) );
  NAND2_X1 U12334 ( .A1(n11410), .A2(n11409), .ZN(n9747) );
  INV_X1 U12335 ( .A(n9743), .ZN(n9746) );
  INV_X1 U12336 ( .A(n9744), .ZN(n9745) );
  NAND2_X1 U12337 ( .A1(n9746), .A2(n9745), .ZN(n11408) );
  OR2_X1 U12338 ( .A1(n10549), .A2(n9629), .ZN(n9751) );
  INV_X1 U12339 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U12340 ( .A1(n9576), .A2(n9748), .ZN(n9762) );
  NAND2_X1 U12341 ( .A1(n9762), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9749) );
  XNOR2_X1 U12342 ( .A(n9749), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10931) );
  AOI22_X1 U12343 ( .A1(n9913), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10931), 
        .B2(n6540), .ZN(n9750) );
  XNOR2_X1 U12344 ( .A(n14307), .B(n10014), .ZN(n9756) );
  AOI22_X1 U12345 ( .A1(n9653), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n9974), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n9755) );
  INV_X1 U12346 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10637) );
  XNOR2_X1 U12347 ( .A(n9767), .B(n10637), .ZN(n11755) );
  NAND2_X1 U12348 ( .A1(n9655), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9752) );
  OAI21_X1 U12349 ( .B1(n11755), .B2(n10089), .A(n9752), .ZN(n9753) );
  INV_X1 U12350 ( .A(n9753), .ZN(n9754) );
  NAND2_X1 U12351 ( .A1(n9652), .A2(n13900), .ZN(n9757) );
  NAND2_X1 U12352 ( .A1(n9756), .A2(n9757), .ZN(n9761) );
  INV_X1 U12353 ( .A(n9756), .ZN(n9759) );
  INV_X1 U12354 ( .A(n9757), .ZN(n9758) );
  NAND2_X1 U12355 ( .A1(n9759), .A2(n9758), .ZN(n9760) );
  NAND2_X1 U12356 ( .A1(n9761), .A2(n9760), .ZN(n11754) );
  NAND2_X1 U12357 ( .A1(n9777), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9763) );
  XNOR2_X1 U12358 ( .A(n9763), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U12359 ( .A1(n9913), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10946), 
        .B2(n6540), .ZN(n9764) );
  XNOR2_X1 U12360 ( .A(n14302), .B(n10014), .ZN(n9773) );
  NAND2_X1 U12361 ( .A1(n9653), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9772) );
  INV_X1 U12362 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9766) );
  OAI21_X1 U12363 ( .B1(n9767), .B2(n10637), .A(n9766), .ZN(n9768) );
  AND2_X1 U12364 ( .A1(n9783), .A2(n9768), .ZN(n11797) );
  NAND2_X1 U12365 ( .A1(n9973), .A2(n11797), .ZN(n9771) );
  NAND2_X1 U12366 ( .A1(n9655), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9770) );
  NAND2_X1 U12367 ( .A1(n10028), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9769) );
  NAND4_X1 U12368 ( .A1(n9772), .A2(n9771), .A3(n9770), .A4(n9769), .ZN(n13899) );
  NAND2_X1 U12369 ( .A1(n9652), .A2(n13899), .ZN(n9774) );
  XNOR2_X1 U12370 ( .A(n9773), .B(n9774), .ZN(n11774) );
  INV_X1 U12371 ( .A(n9773), .ZN(n9776) );
  INV_X1 U12372 ( .A(n9774), .ZN(n9775) );
  NAND2_X1 U12373 ( .A1(n10697), .A2(n13785), .ZN(n9780) );
  OAI21_X1 U12374 ( .B1(n9777), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9778) );
  XNOR2_X1 U12375 ( .A(n9778), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U12376 ( .A1(n9913), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n11469), 
        .B2(n6540), .ZN(n9779) );
  XNOR2_X1 U12377 ( .A(n13711), .B(n6537), .ZN(n9791) );
  AOI22_X1 U12378 ( .A1(n9653), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10028), 
        .B2(P2_REG1_REG_11__SCAN_IN), .ZN(n9788) );
  INV_X1 U12379 ( .A(n9783), .ZN(n9781) );
  INV_X1 U12380 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9782) );
  NAND2_X1 U12381 ( .A1(n9783), .A2(n9782), .ZN(n9784) );
  NAND2_X1 U12382 ( .A1(n9800), .A2(n9784), .ZN(n12014) );
  NAND2_X1 U12383 ( .A1(n9655), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9785) );
  OAI21_X1 U12384 ( .B1(n12014), .B2(n10089), .A(n9785), .ZN(n9786) );
  INV_X1 U12385 ( .A(n9786), .ZN(n9787) );
  NAND2_X1 U12386 ( .A1(n9652), .A2(n13898), .ZN(n9789) );
  XNOR2_X1 U12387 ( .A(n9791), .B(n9789), .ZN(n12006) );
  NAND2_X1 U12388 ( .A1(n12007), .A2(n12006), .ZN(n9793) );
  INV_X1 U12389 ( .A(n9789), .ZN(n9790) );
  NAND2_X1 U12390 ( .A1(n9791), .A2(n9790), .ZN(n9792) );
  NAND2_X1 U12391 ( .A1(n10715), .A2(n13785), .ZN(n9798) );
  NAND2_X1 U12392 ( .A1(n9794), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9795) );
  MUX2_X1 U12393 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9795), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n9796) );
  AOI22_X1 U12394 ( .A1(n9913), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n11472), 
        .B2(n6540), .ZN(n9797) );
  XNOR2_X1 U12395 ( .A(n13716), .B(n10014), .ZN(n9806) );
  NAND2_X1 U12396 ( .A1(n9800), .A2(n9799), .ZN(n9801) );
  AND2_X1 U12397 ( .A1(n9814), .A2(n9801), .ZN(n12164) );
  NAND2_X1 U12398 ( .A1(n9973), .A2(n12164), .ZN(n9805) );
  NAND2_X1 U12399 ( .A1(n9653), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9804) );
  NAND2_X1 U12400 ( .A1(n10017), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9803) );
  NAND2_X1 U12401 ( .A1(n13788), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9802) );
  NAND4_X1 U12402 ( .A1(n9805), .A2(n9804), .A3(n9803), .A4(n9802), .ZN(n13897) );
  AND2_X1 U12403 ( .A1(n9981), .A2(n13897), .ZN(n9807) );
  AND2_X1 U12404 ( .A1(n9806), .A2(n9807), .ZN(n12159) );
  INV_X1 U12405 ( .A(n9806), .ZN(n9809) );
  INV_X1 U12406 ( .A(n9807), .ZN(n9808) );
  NAND2_X1 U12407 ( .A1(n9809), .A2(n9808), .ZN(n12160) );
  NAND2_X1 U12408 ( .A1(n10817), .A2(n13785), .ZN(n9812) );
  NAND2_X1 U12409 ( .A1(n9828), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9810) );
  XNOR2_X1 U12410 ( .A(n9810), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U12411 ( .A1(n9913), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n11473), 
        .B2(n6540), .ZN(n9811) );
  XNOR2_X1 U12412 ( .A(n14292), .B(n6537), .ZN(n9822) );
  INV_X1 U12413 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U12414 ( .A1(n9814), .A2(n9813), .ZN(n9815) );
  NAND2_X1 U12415 ( .A1(n9835), .A2(n9815), .ZN(n12321) );
  OR2_X1 U12416 ( .A1(n10089), .A2(n12321), .ZN(n9821) );
  INV_X1 U12417 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9818) );
  NAND2_X1 U12418 ( .A1(n9974), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U12419 ( .A1(n13788), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9816) );
  OAI211_X1 U12420 ( .C1(n12536), .C2(n9818), .A(n9817), .B(n9816), .ZN(n9819)
         );
  INV_X1 U12421 ( .A(n9819), .ZN(n9820) );
  AND2_X1 U12422 ( .A1(n13896), .A2(n9981), .ZN(n9823) );
  NAND2_X1 U12423 ( .A1(n9822), .A2(n9823), .ZN(n9827) );
  INV_X1 U12424 ( .A(n9822), .ZN(n9825) );
  INV_X1 U12425 ( .A(n9823), .ZN(n9824) );
  NAND2_X1 U12426 ( .A1(n9825), .A2(n9824), .ZN(n9826) );
  NAND2_X1 U12427 ( .A1(n9827), .A2(n9826), .ZN(n12317) );
  INV_X1 U12428 ( .A(n9828), .ZN(n9830) );
  NAND2_X1 U12429 ( .A1(n9830), .A2(n9829), .ZN(n9846) );
  NAND2_X1 U12430 ( .A1(n9846), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9831) );
  XNOR2_X1 U12431 ( .A(n9831), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U12432 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n9913), .B1(n11977), 
        .B2(n6540), .ZN(n9832) );
  NAND2_X2 U12433 ( .A1(n9833), .A2(n9832), .ZN(n13724) );
  XNOR2_X1 U12434 ( .A(n13724), .B(n10014), .ZN(n9844) );
  NAND2_X1 U12435 ( .A1(n9835), .A2(n9834), .ZN(n9836) );
  AND2_X1 U12436 ( .A1(n9851), .A2(n9836), .ZN(n13507) );
  NAND2_X1 U12437 ( .A1(n13507), .A2(n9973), .ZN(n9842) );
  INV_X1 U12438 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9839) );
  NAND2_X1 U12439 ( .A1(n10017), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U12440 ( .A1(n13788), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9837) );
  OAI211_X1 U12441 ( .C1(n12536), .C2(n9839), .A(n9838), .B(n9837), .ZN(n9840)
         );
  INV_X1 U12442 ( .A(n9840), .ZN(n9841) );
  NAND2_X1 U12443 ( .A1(n9842), .A2(n9841), .ZN(n13895) );
  NAND2_X1 U12444 ( .A1(n13895), .A2(n9981), .ZN(n9843) );
  XNOR2_X1 U12445 ( .A(n9844), .B(n9843), .ZN(n13506) );
  NAND2_X1 U12446 ( .A1(n9844), .A2(n9843), .ZN(n9845) );
  NAND2_X1 U12447 ( .A1(n11175), .A2(n13785), .ZN(n9849) );
  NAND2_X1 U12448 ( .A1(n9859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9847) );
  XNOR2_X1 U12449 ( .A(n9847), .B(P2_IR_REG_15__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U12450 ( .A1(n12136), .A2(n6540), .B1(P1_DATAO_REG_15__SCAN_IN), 
        .B2(n9913), .ZN(n9848) );
  XNOR2_X1 U12451 ( .A(n14280), .B(n10014), .ZN(n13545) );
  OR2_X2 U12452 ( .A1(n9851), .A2(n9850), .ZN(n9870) );
  NAND2_X1 U12453 ( .A1(n9851), .A2(n9850), .ZN(n9852) );
  AND2_X1 U12454 ( .A1(n9870), .A2(n9852), .ZN(n14168) );
  NAND2_X1 U12455 ( .A1(n14168), .A2(n9973), .ZN(n9858) );
  INV_X1 U12456 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U12457 ( .A1(n9974), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9854) );
  NAND2_X1 U12458 ( .A1(n13788), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9853) );
  OAI211_X1 U12459 ( .C1(n12536), .C2(n9855), .A(n9854), .B(n9853), .ZN(n9856)
         );
  INV_X1 U12460 ( .A(n9856), .ZN(n9857) );
  NAND2_X1 U12461 ( .A1(n9858), .A2(n9857), .ZN(n13894) );
  AND2_X1 U12462 ( .A1(n13894), .A2(n9981), .ZN(n13629) );
  NAND2_X1 U12463 ( .A1(n11005), .A2(n13785), .ZN(n9867) );
  INV_X1 U12464 ( .A(n9859), .ZN(n9861) );
  INV_X1 U12465 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U12466 ( .A1(n9861), .A2(n9860), .ZN(n9863) );
  NAND2_X1 U12467 ( .A1(n9863), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9862) );
  MUX2_X1 U12468 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9862), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n9864) );
  NOR2_X1 U12469 ( .A1(n9878), .A2(n15748), .ZN(n9865) );
  AOI21_X1 U12470 ( .B1(n12141), .B2(n6540), .A(n9865), .ZN(n9866) );
  XNOR2_X1 U12471 ( .A(n14274), .B(n10014), .ZN(n13544) );
  INV_X1 U12472 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U12473 ( .A1(n9870), .A2(n9869), .ZN(n9871) );
  NAND2_X1 U12474 ( .A1(n9883), .A2(n9871), .ZN(n14147) );
  OR2_X1 U12475 ( .A1(n14147), .A2(n10089), .ZN(n9876) );
  INV_X1 U12476 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12140) );
  NAND2_X1 U12477 ( .A1(n10017), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U12478 ( .A1(n13788), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9872) );
  OAI211_X1 U12479 ( .C1(n12536), .C2(n12140), .A(n9873), .B(n9872), .ZN(n9874) );
  INV_X1 U12480 ( .A(n9874), .ZN(n9875) );
  NAND2_X1 U12481 ( .A1(n9876), .A2(n9875), .ZN(n13893) );
  NAND2_X1 U12482 ( .A1(n13893), .A2(n9981), .ZN(n13543) );
  NAND2_X1 U12483 ( .A1(n13544), .A2(n13543), .ZN(n13556) );
  OAI21_X1 U12484 ( .B1(n13545), .B2(n13629), .A(n13556), .ZN(n9893) );
  NAND2_X1 U12485 ( .A1(n11015), .A2(n13785), .ZN(n9881) );
  NAND2_X1 U12486 ( .A1(n9898), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9877) );
  XNOR2_X1 U12487 ( .A(n9877), .B(P2_IR_REG_17__SCAN_IN), .ZN(n12410) );
  NOR2_X1 U12488 ( .A1(n9878), .A2(n15707), .ZN(n9879) );
  AOI21_X1 U12489 ( .B1(n12410), .B2(n6540), .A(n9879), .ZN(n9880) );
  XNOR2_X1 U12490 ( .A(n13742), .B(n10014), .ZN(n9894) );
  NAND2_X1 U12491 ( .A1(n9883), .A2(n9882), .ZN(n9884) );
  AND2_X1 U12492 ( .A1(n9918), .A2(n9884), .ZN(n14132) );
  NAND2_X1 U12493 ( .A1(n14132), .A2(n9973), .ZN(n9889) );
  INV_X1 U12494 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14134) );
  NAND2_X1 U12495 ( .A1(n10028), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9886) );
  NAND2_X1 U12496 ( .A1(n13788), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9885) );
  OAI211_X1 U12497 ( .C1(n12536), .C2(n14134), .A(n9886), .B(n9885), .ZN(n9887) );
  INV_X1 U12498 ( .A(n9887), .ZN(n9888) );
  NAND2_X1 U12499 ( .A1(n9889), .A2(n9888), .ZN(n14107) );
  NAND2_X1 U12500 ( .A1(n14107), .A2(n9981), .ZN(n9895) );
  XNOR2_X1 U12501 ( .A(n9894), .B(n9895), .ZN(n13557) );
  NAND3_X1 U12502 ( .A1(n13545), .A2(n13629), .A3(n13556), .ZN(n9890) );
  OAI211_X1 U12503 ( .C1(n13544), .C2(n13543), .A(n13557), .B(n9890), .ZN(
        n9891) );
  INV_X1 U12504 ( .A(n9891), .ZN(n9892) );
  INV_X1 U12505 ( .A(n9894), .ZN(n9896) );
  NAND2_X1 U12506 ( .A1(n9896), .A2(n9895), .ZN(n9897) );
  OAI21_X1 U12507 ( .B1(n9898), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9899) );
  XNOR2_X1 U12508 ( .A(n9899), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U12509 ( .A1(n12413), .A2(n6540), .B1(P1_DATAO_REG_18__SCAN_IN), 
        .B2(n9913), .ZN(n9900) );
  XNOR2_X1 U12510 ( .A(n14115), .B(n6537), .ZN(n9907) );
  XNOR2_X1 U12511 ( .A(n9918), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n14113) );
  NAND2_X1 U12512 ( .A1(n14113), .A2(n9973), .ZN(n9906) );
  INV_X1 U12513 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9903) );
  NAND2_X1 U12514 ( .A1(n10017), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U12515 ( .A1(n13788), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9901) );
  OAI211_X1 U12516 ( .C1(n12536), .C2(n9903), .A(n9902), .B(n9901), .ZN(n9904)
         );
  INV_X1 U12517 ( .A(n9904), .ZN(n9905) );
  NAND2_X1 U12518 ( .A1(n13892), .A2(n9981), .ZN(n9908) );
  XNOR2_X1 U12519 ( .A(n9907), .B(n9908), .ZN(n13611) );
  INV_X1 U12520 ( .A(n9907), .ZN(n9910) );
  INV_X1 U12521 ( .A(n9908), .ZN(n9909) );
  NAND2_X1 U12522 ( .A1(n9910), .A2(n9909), .ZN(n9911) );
  NAND2_X1 U12523 ( .A1(n11511), .A2(n6550), .ZN(n9915) );
  AOI22_X1 U12524 ( .A1(n9913), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9912), 
        .B2(n6540), .ZN(n9914) );
  XNOR2_X1 U12525 ( .A(n14257), .B(n10014), .ZN(n9926) );
  INV_X1 U12526 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9917) );
  INV_X1 U12527 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9916) );
  OAI21_X1 U12528 ( .B1(n9918), .B2(n9917), .A(n9916), .ZN(n9920) );
  AND2_X1 U12529 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n9919) );
  NAND2_X1 U12530 ( .A1(n9920), .A2(n9932), .ZN(n14099) );
  OR2_X1 U12531 ( .A1(n14099), .A2(n10089), .ZN(n9925) );
  INV_X1 U12532 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14100) );
  NAND2_X1 U12533 ( .A1(n10028), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U12534 ( .A1(n13788), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9921) );
  OAI211_X1 U12535 ( .C1(n12536), .C2(n14100), .A(n9922), .B(n9921), .ZN(n9923) );
  INV_X1 U12536 ( .A(n9923), .ZN(n9924) );
  NAND2_X1 U12537 ( .A1(n14109), .A2(n9981), .ZN(n9927) );
  NAND2_X1 U12538 ( .A1(n9926), .A2(n9927), .ZN(n13520) );
  INV_X1 U12539 ( .A(n9926), .ZN(n9929) );
  INV_X1 U12540 ( .A(n9927), .ZN(n9928) );
  NAND2_X1 U12541 ( .A1(n9929), .A2(n9928), .ZN(n13519) );
  NAND2_X1 U12542 ( .A1(n11542), .A2(n13785), .ZN(n9931) );
  NAND2_X1 U12543 ( .A1(n9913), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9930) );
  XNOR2_X1 U12544 ( .A(n14252), .B(n10014), .ZN(n9940) );
  NAND2_X1 U12545 ( .A1(n9932), .A2(n13587), .ZN(n9933) );
  NAND2_X1 U12546 ( .A1(n9946), .A2(n9933), .ZN(n14072) );
  OR2_X1 U12547 ( .A1(n14072), .A2(n10089), .ZN(n9939) );
  INV_X1 U12548 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9936) );
  NAND2_X1 U12549 ( .A1(n13788), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9935) );
  NAND2_X1 U12550 ( .A1(n10017), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9934) );
  OAI211_X1 U12551 ( .C1(n12536), .C2(n9936), .A(n9935), .B(n9934), .ZN(n9937)
         );
  INV_X1 U12552 ( .A(n9937), .ZN(n9938) );
  NAND2_X1 U12553 ( .A1(n14057), .A2(n9981), .ZN(n9941) );
  NAND2_X1 U12554 ( .A1(n9940), .A2(n9941), .ZN(n9945) );
  INV_X1 U12555 ( .A(n9940), .ZN(n9943) );
  INV_X1 U12556 ( .A(n9941), .ZN(n9942) );
  NAND2_X1 U12557 ( .A1(n9943), .A2(n9942), .ZN(n9944) );
  NAND2_X1 U12558 ( .A1(n9945), .A2(n9944), .ZN(n13586) );
  XNOR2_X1 U12559 ( .A(n14064), .B(n6537), .ZN(n9954) );
  INV_X1 U12560 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13530) );
  NAND2_X1 U12561 ( .A1(n9946), .A2(n13530), .ZN(n9947) );
  NAND2_X1 U12562 ( .A1(n9959), .A2(n9947), .ZN(n14061) );
  INV_X1 U12563 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U12564 ( .A1(n10017), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U12565 ( .A1(n13788), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9948) );
  OAI211_X1 U12566 ( .C1(n12536), .C2(n9950), .A(n9949), .B(n9948), .ZN(n9951)
         );
  INV_X1 U12567 ( .A(n9951), .ZN(n9952) );
  NAND2_X1 U12568 ( .A1(n14081), .A2(n9981), .ZN(n9953) );
  XNOR2_X1 U12569 ( .A(n9954), .B(n9953), .ZN(n13528) );
  NAND2_X1 U12570 ( .A1(n11922), .A2(n13785), .ZN(n9958) );
  NAND2_X1 U12571 ( .A1(n9913), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9957) );
  XNOR2_X1 U12572 ( .A(n14049), .B(n6537), .ZN(n13592) );
  INV_X1 U12573 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13596) );
  NAND2_X1 U12574 ( .A1(n9959), .A2(n13596), .ZN(n9960) );
  AND2_X1 U12575 ( .A1(n9984), .A2(n9960), .ZN(n14048) );
  NAND2_X1 U12576 ( .A1(n14048), .A2(n6548), .ZN(n9966) );
  INV_X1 U12577 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9963) );
  NAND2_X1 U12578 ( .A1(n9974), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9962) );
  NAND2_X1 U12579 ( .A1(n13788), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9961) );
  OAI211_X1 U12580 ( .C1(n12536), .C2(n9963), .A(n9962), .B(n9961), .ZN(n9964)
         );
  INV_X1 U12581 ( .A(n9964), .ZN(n9965) );
  AND2_X1 U12582 ( .A1(n14058), .A2(n9981), .ZN(n13593) );
  NAND2_X1 U12583 ( .A1(n13595), .A2(n13592), .ZN(n9967) );
  NAND2_X1 U12584 ( .A1(n12104), .A2(n13785), .ZN(n9970) );
  NAND2_X1 U12585 ( .A1(n9663), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9969) );
  XOR2_X1 U12586 ( .A(n6537), .B(n14230), .Z(n13574) );
  INV_X1 U12587 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13577) );
  OR2_X2 U12588 ( .A1(n9986), .A2(n13577), .ZN(n9999) );
  NAND2_X1 U12589 ( .A1(n9986), .A2(n13577), .ZN(n9972) );
  AND2_X1 U12590 ( .A1(n9999), .A2(n9972), .ZN(n14015) );
  NAND2_X1 U12591 ( .A1(n14015), .A2(n6548), .ZN(n9980) );
  INV_X1 U12592 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9977) );
  NAND2_X1 U12593 ( .A1(n9974), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U12594 ( .A1(n13788), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9975) );
  OAI211_X1 U12595 ( .C1(n12536), .C2(n9977), .A(n9976), .B(n9975), .ZN(n9978)
         );
  INV_X1 U12596 ( .A(n9978), .ZN(n9979) );
  AND2_X1 U12597 ( .A1(n13998), .A2(n9981), .ZN(n13573) );
  INV_X1 U12598 ( .A(n13573), .ZN(n9992) );
  NAND2_X1 U12599 ( .A1(n11925), .A2(n6550), .ZN(n9983) );
  NAND2_X1 U12600 ( .A1(n9913), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9982) );
  XNOR2_X1 U12601 ( .A(n14034), .B(n6537), .ZN(n13513) );
  INV_X1 U12602 ( .A(n13513), .ZN(n13569) );
  INV_X1 U12603 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13514) );
  NAND2_X1 U12604 ( .A1(n9984), .A2(n13514), .ZN(n9985) );
  NAND2_X1 U12605 ( .A1(n9986), .A2(n9985), .ZN(n14031) );
  INV_X1 U12606 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14032) );
  NAND2_X1 U12607 ( .A1(n10028), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U12608 ( .A1(n13788), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9987) );
  OAI211_X1 U12609 ( .C1(n12536), .C2(n14032), .A(n9988), .B(n9987), .ZN(n9989) );
  INV_X1 U12610 ( .A(n9989), .ZN(n9990) );
  NAND2_X1 U12611 ( .A1(n14041), .A2(n9981), .ZN(n13571) );
  OAI22_X1 U12612 ( .A1(n13574), .A2(n9992), .B1(n13569), .B2(n13571), .ZN(
        n9996) );
  OAI21_X1 U12613 ( .B1(n13513), .B2(n14041), .A(n13573), .ZN(n9994) );
  OAI21_X1 U12614 ( .B1(n13998), .B2(n14041), .A(n9652), .ZN(n9993) );
  AOI22_X1 U12615 ( .A1(n13574), .A2(n9994), .B1(n13569), .B2(n9993), .ZN(
        n9995) );
  INV_X1 U12616 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U12617 ( .A1(n9999), .A2(n9998), .ZN(n10000) );
  NAND2_X1 U12618 ( .A1(n10015), .A2(n10000), .ZN(n13989) );
  INV_X1 U12619 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n10003) );
  NAND2_X1 U12620 ( .A1(n9974), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U12621 ( .A1(n13788), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n10001) );
  OAI211_X1 U12622 ( .C1(n12536), .C2(n10003), .A(n10002), .B(n10001), .ZN(
        n10004) );
  INV_X1 U12623 ( .A(n10004), .ZN(n10005) );
  NAND2_X1 U12624 ( .A1(n14007), .A2(n9981), .ZN(n10010) );
  NAND2_X1 U12625 ( .A1(n12123), .A2(n6550), .ZN(n10008) );
  NAND2_X1 U12626 ( .A1(n9663), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n10007) );
  XNOR2_X1 U12627 ( .A(n14225), .B(n6537), .ZN(n10009) );
  XOR2_X1 U12628 ( .A(n10010), .B(n10009), .Z(n13535) );
  INV_X1 U12629 ( .A(n10009), .ZN(n10011) );
  NAND2_X1 U12630 ( .A1(n12351), .A2(n13785), .ZN(n10013) );
  NAND2_X1 U12631 ( .A1(n9913), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n10012) );
  XNOR2_X1 U12632 ( .A(n14220), .B(n10014), .ZN(n10024) );
  INV_X1 U12633 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n15702) );
  OR2_X2 U12634 ( .A1(n10015), .A2(n15702), .ZN(n10040) );
  NAND2_X1 U12635 ( .A1(n10015), .A2(n15702), .ZN(n10016) );
  NAND2_X1 U12636 ( .A1(n13979), .A2(n6548), .ZN(n10022) );
  INV_X1 U12637 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n15583) );
  NAND2_X1 U12638 ( .A1(n10017), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n10019) );
  NAND2_X1 U12639 ( .A1(n13788), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n10018) );
  OAI211_X1 U12640 ( .C1(n12536), .C2(n15583), .A(n10019), .B(n10018), .ZN(
        n10020) );
  INV_X1 U12641 ( .A(n10020), .ZN(n10021) );
  NAND2_X1 U12642 ( .A1(n13999), .A2(n9981), .ZN(n10023) );
  NAND2_X1 U12643 ( .A1(n10024), .A2(n10023), .ZN(n10025) );
  OAI21_X1 U12644 ( .B1(n10024), .B2(n10023), .A(n10025), .ZN(n13616) );
  NAND2_X1 U12645 ( .A1(n12378), .A2(n13785), .ZN(n10027) );
  NAND2_X1 U12646 ( .A1(n9913), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n10026) );
  XNOR2_X1 U12647 ( .A(n14211), .B(n6537), .ZN(n10036) );
  XNOR2_X1 U12648 ( .A(n10040), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13966) );
  NAND2_X1 U12649 ( .A1(n13966), .A2(n6548), .ZN(n10034) );
  INV_X1 U12650 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n10031) );
  NAND2_X1 U12651 ( .A1(n10028), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n10030) );
  NAND2_X1 U12652 ( .A1(n13788), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n10029) );
  OAI211_X1 U12653 ( .C1(n12536), .C2(n10031), .A(n10030), .B(n10029), .ZN(
        n10032) );
  INV_X1 U12654 ( .A(n10032), .ZN(n10033) );
  NAND2_X1 U12655 ( .A1(n13891), .A2(n9981), .ZN(n10035) );
  XNOR2_X1 U12656 ( .A(n10036), .B(n10035), .ZN(n13496) );
  INV_X1 U12657 ( .A(n10035), .ZN(n10037) );
  NAND2_X1 U12658 ( .A1(n14355), .A2(n6550), .ZN(n10039) );
  NAND2_X1 U12659 ( .A1(n9913), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n10038) );
  INV_X1 U12660 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13497) );
  INV_X1 U12661 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n15703) );
  OAI21_X1 U12662 ( .B1(n10040), .B2(n13497), .A(n15703), .ZN(n10043) );
  INV_X1 U12663 ( .A(n10040), .ZN(n10042) );
  AND2_X1 U12664 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(P2_REG3_REG_27__SCAN_IN), 
        .ZN(n10041) );
  NAND2_X1 U12665 ( .A1(n10042), .A2(n10041), .ZN(n12545) );
  NAND2_X1 U12666 ( .A1(n10043), .A2(n12545), .ZN(n13950) );
  INV_X1 U12667 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13949) );
  NAND2_X1 U12668 ( .A1(n10017), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n10045) );
  NAND2_X1 U12669 ( .A1(n13788), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n10044) );
  OAI211_X1 U12670 ( .C1(n12536), .C2(n13949), .A(n10045), .B(n10044), .ZN(
        n10046) );
  INV_X1 U12671 ( .A(n10046), .ZN(n10047) );
  NAND2_X1 U12672 ( .A1(n13961), .A2(n9981), .ZN(n10049) );
  XNOR2_X1 U12673 ( .A(n10049), .B(n6537), .ZN(n10050) );
  NAND2_X1 U12674 ( .A1(n10051), .A2(n15600), .ZN(n10075) );
  NAND2_X1 U12675 ( .A1(n10054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10053) );
  XNOR2_X1 U12676 ( .A(n12109), .B(P2_B_REG_SCAN_IN), .ZN(n10057) );
  INV_X1 U12677 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U12678 ( .A1(n10057), .A2(n12125), .ZN(n10061) );
  NAND2_X1 U12679 ( .A1(n10059), .A2(n10058), .ZN(n14348) );
  NAND2_X1 U12680 ( .A1(n14348), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10060) );
  INV_X1 U12681 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15430) );
  NAND2_X1 U12682 ( .A1(n15427), .A2(n15430), .ZN(n10063) );
  NAND2_X1 U12683 ( .A1(n12109), .A2(n12354), .ZN(n10062) );
  INV_X1 U12684 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15435) );
  NAND2_X1 U12685 ( .A1(n15427), .A2(n15435), .ZN(n10065) );
  NAND2_X1 U12686 ( .A1(n12125), .A2(n12354), .ZN(n10064) );
  NAND2_X1 U12687 ( .A1(n10065), .A2(n10064), .ZN(n10681) );
  INV_X1 U12688 ( .A(n10681), .ZN(n11326) );
  NOR4_X1 U12689 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n10069) );
  NOR4_X1 U12690 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n10068) );
  NOR4_X1 U12691 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n10067) );
  NOR4_X1 U12692 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n10066) );
  NAND4_X1 U12693 ( .A1(n10069), .A2(n10068), .A3(n10067), .A4(n10066), .ZN(
        n10074) );
  NOR2_X1 U12694 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .ZN(
        n15564) );
  NOR4_X1 U12695 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n10072) );
  NOR4_X1 U12696 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n10071) );
  NOR4_X1 U12697 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n10070) );
  NAND4_X1 U12698 ( .A1(n15564), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n10073) );
  OAI21_X1 U12699 ( .B1(n10074), .B2(n10073), .A(n15427), .ZN(n11325) );
  NAND3_X1 U12700 ( .A1(n10684), .A2(n11326), .A3(n11325), .ZN(n10096) );
  NAND2_X1 U12701 ( .A1(n10075), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10077) );
  XNOR2_X1 U12702 ( .A(n10077), .B(n10076), .ZN(n11907) );
  INV_X1 U12703 ( .A(n10574), .ZN(n10078) );
  NAND2_X1 U12704 ( .A1(n14152), .A2(n13833), .ZN(n13835) );
  NAND3_X1 U12705 ( .A1(n15432), .A2(n10078), .A3(n15451), .ZN(n10079) );
  AND2_X1 U12706 ( .A1(n10826), .A2(n10080), .ZN(n11329) );
  NAND2_X1 U12707 ( .A1(n15432), .A2(n11329), .ZN(n10081) );
  OR2_X1 U12708 ( .A1(n10096), .A2(n10081), .ZN(n10082) );
  NAND2_X1 U12709 ( .A1(n14308), .A2(n9912), .ZN(n10682) );
  NAND2_X1 U12710 ( .A1(n14207), .A2(n13623), .ZN(n10103) );
  NAND2_X1 U12711 ( .A1(n10083), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10581) );
  INV_X1 U12712 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n10084) );
  NAND2_X1 U12713 ( .A1(n10581), .A2(n10084), .ZN(n10085) );
  NAND2_X1 U12714 ( .A1(n10085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10087) );
  INV_X1 U12715 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n10086) );
  XNOR2_X1 U12716 ( .A(n10087), .B(n10086), .ZN(n10580) );
  INV_X1 U12717 ( .A(n10580), .ZN(n10088) );
  OR2_X1 U12718 ( .A1(n12545), .A2(n10089), .ZN(n10094) );
  INV_X1 U12719 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n12544) );
  NAND2_X1 U12720 ( .A1(n13788), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U12721 ( .A1(n9974), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n10090) );
  OAI211_X1 U12722 ( .C1(n12536), .C2(n12544), .A(n10091), .B(n10090), .ZN(
        n10092) );
  INV_X1 U12723 ( .A(n10092), .ZN(n10093) );
  OAI22_X1 U12724 ( .A1(n13978), .A2(n14092), .B1(n13799), .B2(n14094), .ZN(
        n13945) );
  NOR2_X1 U12725 ( .A1(n15434), .A2(n13835), .ZN(n13882) );
  INV_X1 U12726 ( .A(n13882), .ZN(n10095) );
  NAND2_X1 U12727 ( .A1(n10096), .A2(n10682), .ZN(n10100) );
  NAND2_X1 U12728 ( .A1(n10574), .A2(n13835), .ZN(n11327) );
  INV_X1 U12729 ( .A(n11327), .ZN(n10097) );
  NOR2_X1 U12730 ( .A1(n10098), .A2(n10097), .ZN(n10099) );
  NAND2_X1 U12731 ( .A1(n10100), .A2(n10099), .ZN(n10962) );
  OAI22_X1 U12732 ( .A1(n13950), .A2(n13599), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15703), .ZN(n10101) );
  AOI21_X1 U12733 ( .B1(n13945), .B2(n13550), .A(n10101), .ZN(n10102) );
  OAI21_X1 U12734 ( .B1(n10105), .B2(n13625), .A(n10104), .ZN(P2_U3192) );
  INV_X2 U12735 ( .A(n10109), .ZN(n10110) );
  OR2_X4 U12736 ( .A1(n10115), .A2(n10110), .ZN(n10314) );
  AND2_X1 U12737 ( .A1(n14557), .A2(n10305), .ZN(n10111) );
  AOI21_X1 U12738 ( .B1(n14875), .B2(n10316), .A(n10111), .ZN(n10256) );
  INV_X1 U12739 ( .A(n10256), .ZN(n10258) );
  NAND2_X1 U12740 ( .A1(n14875), .A2(n10309), .ZN(n10113) );
  NAND2_X1 U12741 ( .A1(n14557), .A2(n10307), .ZN(n10112) );
  NAND2_X1 U12742 ( .A1(n10113), .A2(n10112), .ZN(n10114) );
  XNOR2_X1 U12743 ( .A(n10114), .B(n10270), .ZN(n10257) );
  OAI22_X1 U12744 ( .A1(n9429), .A2(n10133), .B1(n10115), .B2(n10117), .ZN(
        n10116) );
  OAI22_X1 U12745 ( .A1(n10314), .A2(n9429), .B1(n10117), .B2(n10133), .ZN(
        n10128) );
  XNOR2_X1 U12746 ( .A(n10129), .B(n10128), .ZN(n12389) );
  INV_X1 U12747 ( .A(n10314), .ZN(n10119) );
  NAND2_X1 U12748 ( .A1(n10119), .A2(n12392), .ZN(n10122) );
  INV_X1 U12749 ( .A(n10409), .ZN(n10120) );
  AOI22_X1 U12750 ( .A1(n10307), .A2(n11441), .B1(n10120), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n10121) );
  OR2_X1 U12751 ( .A1(n10115), .A2(n11343), .ZN(n10123) );
  OAI211_X1 U12752 ( .C1(n10125), .C2(n10409), .A(n10124), .B(n10123), .ZN(
        n10851) );
  NAND2_X1 U12753 ( .A1(n10852), .A2(n10851), .ZN(n10850) );
  INV_X1 U12754 ( .A(n10851), .ZN(n10126) );
  NAND2_X1 U12755 ( .A1(n10850), .A2(n10127), .ZN(n12391) );
  NAND2_X1 U12756 ( .A1(n12389), .A2(n12391), .ZN(n10132) );
  INV_X1 U12757 ( .A(n10128), .ZN(n10130) );
  NAND2_X1 U12758 ( .A1(n10130), .A2(n10129), .ZN(n10131) );
  NAND2_X1 U12759 ( .A1(n10132), .A2(n10131), .ZN(n12478) );
  OAI22_X1 U12760 ( .A1(n10136), .A2(n10133), .B1(n10115), .B2(n15306), .ZN(
        n10135) );
  XNOR2_X1 U12761 ( .A(n10135), .B(n10190), .ZN(n10138) );
  OAI22_X1 U12762 ( .A1(n10314), .A2(n10136), .B1(n15306), .B2(n10310), .ZN(
        n10137) );
  XNOR2_X1 U12763 ( .A(n10138), .B(n10137), .ZN(n12480) );
  NAND2_X1 U12764 ( .A1(n12478), .A2(n12480), .ZN(n10141) );
  INV_X1 U12765 ( .A(n10137), .ZN(n10139) );
  NAND2_X1 U12766 ( .A1(n10139), .A2(n10138), .ZN(n10140) );
  NAND2_X1 U12767 ( .A1(n10141), .A2(n10140), .ZN(n10429) );
  INV_X1 U12768 ( .A(n10429), .ZN(n10146) );
  OR2_X1 U12769 ( .A1(n10310), .A2(n10144), .ZN(n10142) );
  OAI21_X1 U12770 ( .B1(n10115), .B2(n15315), .A(n10142), .ZN(n10143) );
  XNOR2_X1 U12771 ( .A(n10143), .B(n10270), .ZN(n10148) );
  OAI22_X1 U12772 ( .A1(n10314), .A2(n10144), .B1(n15315), .B2(n10310), .ZN(
        n10147) );
  XNOR2_X1 U12773 ( .A(n10148), .B(n10147), .ZN(n10432) );
  NAND2_X1 U12774 ( .A1(n10148), .A2(n10147), .ZN(n10149) );
  OAI22_X1 U12775 ( .A1(n10314), .A2(n10150), .B1(n15322), .B2(n10310), .ZN(
        n11566) );
  OAI21_X1 U12776 ( .B1(n10115), .B2(n15322), .A(n10151), .ZN(n10152) );
  OR2_X1 U12777 ( .A1(n10115), .A2(n15262), .ZN(n10153) );
  OAI21_X1 U12778 ( .B1(n10310), .B2(n11396), .A(n10153), .ZN(n10154) );
  XNOR2_X1 U12779 ( .A(n10154), .B(n10270), .ZN(n11568) );
  OAI22_X1 U12780 ( .A1(n10314), .A2(n11396), .B1(n15262), .B2(n10310), .ZN(
        n10157) );
  AOI22_X1 U12781 ( .A1(n11566), .A2(n14462), .B1(n11568), .B2(n10157), .ZN(
        n10155) );
  INV_X1 U12782 ( .A(n11568), .ZN(n10160) );
  NAND2_X1 U12783 ( .A1(n10156), .A2(n10157), .ZN(n10159) );
  INV_X1 U12784 ( .A(n10156), .ZN(n10158) );
  INV_X1 U12785 ( .A(n10157), .ZN(n11569) );
  AOI22_X1 U12786 ( .A1(n10160), .A2(n10159), .B1(n10158), .B2(n11569), .ZN(
        n10161) );
  INV_X1 U12787 ( .A(n11603), .ZN(n10165) );
  INV_X1 U12788 ( .A(n11605), .ZN(n11457) );
  OR2_X1 U12789 ( .A1(n10310), .A2(n11548), .ZN(n10162) );
  OAI21_X1 U12790 ( .B1(n10115), .B2(n11457), .A(n10162), .ZN(n10163) );
  XNOR2_X1 U12791 ( .A(n10163), .B(n10270), .ZN(n10167) );
  OAI22_X1 U12792 ( .A1(n10314), .A2(n11548), .B1(n11457), .B2(n10310), .ZN(
        n10166) );
  XNOR2_X1 U12793 ( .A(n10167), .B(n10166), .ZN(n11604) );
  NAND2_X1 U12794 ( .A1(n10167), .A2(n10166), .ZN(n10168) );
  NAND2_X1 U12795 ( .A1(n11601), .A2(n10168), .ZN(n11547) );
  OAI22_X1 U12796 ( .A1(n15251), .A2(n10115), .B1(n11491), .B2(n10310), .ZN(
        n10169) );
  XNOR2_X1 U12797 ( .A(n10169), .B(n10190), .ZN(n10170) );
  OAI22_X1 U12798 ( .A1(n11491), .A2(n10314), .B1(n15251), .B2(n10310), .ZN(
        n10171) );
  XNOR2_X1 U12799 ( .A(n10170), .B(n10171), .ZN(n11546) );
  NAND2_X1 U12800 ( .A1(n11547), .A2(n11546), .ZN(n11545) );
  INV_X1 U12801 ( .A(n10170), .ZN(n10172) );
  NAND2_X1 U12802 ( .A1(n10172), .A2(n10171), .ZN(n10173) );
  NAND2_X1 U12803 ( .A1(n10177), .A2(n10309), .ZN(n10175) );
  OR2_X1 U12804 ( .A1(n10310), .A2(n11861), .ZN(n10174) );
  NAND2_X1 U12805 ( .A1(n10175), .A2(n10174), .ZN(n10176) );
  XNOR2_X1 U12806 ( .A(n10176), .B(n10190), .ZN(n10182) );
  NAND2_X1 U12807 ( .A1(n10177), .A2(n10307), .ZN(n10179) );
  NAND2_X1 U12808 ( .A1(n10305), .A2(n14564), .ZN(n10178) );
  NAND2_X1 U12809 ( .A1(n10179), .A2(n10178), .ZN(n10180) );
  XNOR2_X1 U12810 ( .A(n10182), .B(n10180), .ZN(n11900) );
  INV_X1 U12811 ( .A(n10180), .ZN(n10181) );
  NAND2_X1 U12812 ( .A1(n10182), .A2(n10181), .ZN(n10183) );
  OAI22_X1 U12813 ( .A1(n12301), .A2(n10115), .B1(n12206), .B2(n10310), .ZN(
        n10184) );
  NOR2_X1 U12814 ( .A1(n10314), .A2(n12206), .ZN(n10185) );
  AOI21_X1 U12815 ( .B1(n15096), .B2(n10316), .A(n10185), .ZN(n12293) );
  NAND2_X1 U12816 ( .A1(n11991), .A2(n10316), .ZN(n10187) );
  NAND2_X1 U12817 ( .A1(n10305), .A2(n14563), .ZN(n10186) );
  NAND2_X1 U12818 ( .A1(n10187), .A2(n10186), .ZN(n12288) );
  INV_X1 U12819 ( .A(n12288), .ZN(n10193) );
  NAND2_X1 U12820 ( .A1(n11991), .A2(n10309), .ZN(n10189) );
  OR2_X1 U12821 ( .A1(n10310), .A2(n11522), .ZN(n10188) );
  NAND2_X1 U12822 ( .A1(n10189), .A2(n10188), .ZN(n10191) );
  XNOR2_X1 U12823 ( .A(n10191), .B(n10303), .ZN(n12290) );
  INV_X1 U12824 ( .A(n12290), .ZN(n10192) );
  AOI22_X1 U12825 ( .A1(n12292), .A2(n12293), .B1(n10193), .B2(n10192), .ZN(
        n10197) );
  NAND2_X1 U12826 ( .A1(n12290), .A2(n12288), .ZN(n10194) );
  AOI21_X1 U12827 ( .B1(n12293), .B2(n10194), .A(n12292), .ZN(n10196) );
  NOR2_X1 U12828 ( .A1(n10194), .A2(n12293), .ZN(n10195) );
  NOR2_X1 U12829 ( .A1(n10310), .A2(n10200), .ZN(n10198) );
  AOI21_X1 U12830 ( .B1(n14507), .B2(n10309), .A(n10198), .ZN(n10199) );
  XNOR2_X1 U12831 ( .A(n10199), .B(n10303), .ZN(n10207) );
  OAI22_X1 U12832 ( .A1(n15087), .A2(n10310), .B1(n10200), .B2(n10314), .ZN(
        n10205) );
  XNOR2_X1 U12833 ( .A(n10207), .B(n10205), .ZN(n14502) );
  NAND2_X1 U12834 ( .A1(n14501), .A2(n14502), .ZN(n14409) );
  OAI22_X1 U12835 ( .A1(n15148), .A2(n10310), .B1(n10201), .B2(n10314), .ZN(
        n10209) );
  NAND2_X1 U12836 ( .A1(n14974), .A2(n10309), .ZN(n10203) );
  NAND2_X1 U12837 ( .A1(n10316), .A2(n14560), .ZN(n10202) );
  NAND2_X1 U12838 ( .A1(n10203), .A2(n10202), .ZN(n10204) );
  XNOR2_X1 U12839 ( .A(n10204), .B(n10303), .ZN(n10208) );
  XOR2_X1 U12840 ( .A(n10209), .B(n10208), .Z(n14412) );
  INV_X1 U12841 ( .A(n10205), .ZN(n10206) );
  NAND2_X1 U12842 ( .A1(n10207), .A2(n10206), .ZN(n14410) );
  NAND3_X1 U12843 ( .A1(n14409), .A2(n14412), .A3(n14410), .ZN(n14411) );
  NOR2_X1 U12844 ( .A1(n10314), .A2(n14377), .ZN(n10211) );
  AOI21_X1 U12845 ( .B1(n14984), .B2(n10316), .A(n10211), .ZN(n10214) );
  AOI22_X1 U12846 ( .A1(n14984), .A2(n10309), .B1(n10316), .B2(n14559), .ZN(
        n10212) );
  XNOR2_X1 U12847 ( .A(n10212), .B(n10303), .ZN(n10213) );
  XOR2_X1 U12848 ( .A(n10214), .B(n10213), .Z(n14478) );
  INV_X1 U12849 ( .A(n10213), .ZN(n10216) );
  INV_X1 U12850 ( .A(n10214), .ZN(n10215) );
  NAND2_X1 U12851 ( .A1(n10316), .A2(n14938), .ZN(n10218) );
  XNOR2_X1 U12852 ( .A(n10219), .B(n10190), .ZN(n10229) );
  INV_X1 U12853 ( .A(n10229), .ZN(n10222) );
  NOR2_X1 U12854 ( .A1(n10314), .A2(n14480), .ZN(n10220) );
  AOI21_X1 U12855 ( .B1(n14957), .B2(n10316), .A(n10220), .ZN(n10228) );
  INV_X1 U12856 ( .A(n10228), .ZN(n10221) );
  NAND2_X1 U12857 ( .A1(n9456), .A2(n10309), .ZN(n10224) );
  INV_X1 U12858 ( .A(n14435), .ZN(n14924) );
  NAND2_X1 U12859 ( .A1(n14924), .A2(n10316), .ZN(n10223) );
  NAND2_X1 U12860 ( .A1(n10224), .A2(n10223), .ZN(n10225) );
  XNOR2_X1 U12861 ( .A(n10225), .B(n10303), .ZN(n14428) );
  NAND2_X1 U12862 ( .A1(n9456), .A2(n10316), .ZN(n10227) );
  NAND2_X1 U12863 ( .A1(n10305), .A2(n14924), .ZN(n10226) );
  NAND2_X1 U12864 ( .A1(n10227), .A2(n10226), .ZN(n14536) );
  NOR2_X1 U12865 ( .A1(n10229), .A2(n10228), .ZN(n14373) );
  NAND2_X1 U12866 ( .A1(n15060), .A2(n10309), .ZN(n10231) );
  NAND2_X1 U12867 ( .A1(n14941), .A2(n10316), .ZN(n10230) );
  NAND2_X1 U12868 ( .A1(n10231), .A2(n10230), .ZN(n10232) );
  XNOR2_X1 U12869 ( .A(n10232), .B(n10190), .ZN(n10238) );
  AND2_X1 U12870 ( .A1(n10305), .A2(n14941), .ZN(n10233) );
  AOI21_X1 U12871 ( .B1(n15060), .B2(n10316), .A(n10233), .ZN(n10237) );
  NOR2_X1 U12872 ( .A1(n10238), .A2(n10237), .ZN(n10235) );
  AOI211_X1 U12873 ( .C1(n14428), .C2(n14536), .A(n14373), .B(n10235), .ZN(
        n10234) );
  INV_X1 U12874 ( .A(n10235), .ZN(n14431) );
  INV_X1 U12875 ( .A(n14536), .ZN(n10236) );
  NAND2_X1 U12876 ( .A1(n14431), .A2(n10236), .ZN(n10239) );
  NAND2_X1 U12877 ( .A1(n10238), .A2(n10237), .ZN(n14430) );
  NAND2_X1 U12878 ( .A1(n15055), .A2(n10309), .ZN(n10242) );
  NAND2_X1 U12879 ( .A1(n14925), .A2(n10316), .ZN(n10241) );
  NAND2_X1 U12880 ( .A1(n10242), .A2(n10241), .ZN(n10243) );
  XNOR2_X1 U12881 ( .A(n10243), .B(n10303), .ZN(n10246) );
  NAND2_X1 U12882 ( .A1(n15055), .A2(n10316), .ZN(n10245) );
  NAND2_X1 U12883 ( .A1(n14925), .A2(n10305), .ZN(n10244) );
  NAND2_X1 U12884 ( .A1(n10245), .A2(n10244), .ZN(n10247) );
  NAND2_X1 U12885 ( .A1(n10246), .A2(n10247), .ZN(n14444) );
  INV_X1 U12886 ( .A(n10246), .ZN(n10249) );
  INV_X1 U12887 ( .A(n10247), .ZN(n10248) );
  NAND2_X1 U12888 ( .A1(n10249), .A2(n10248), .ZN(n14443) );
  NAND2_X1 U12889 ( .A1(n14441), .A2(n14443), .ZN(n14513) );
  OAI22_X1 U12890 ( .A1(n14894), .A2(n10310), .B1(n14910), .B2(n10314), .ZN(
        n10253) );
  NAND2_X1 U12891 ( .A1(n15048), .A2(n10309), .ZN(n10251) );
  NAND2_X1 U12892 ( .A1(n14558), .A2(n10316), .ZN(n10250) );
  NAND2_X1 U12893 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  XNOR2_X1 U12894 ( .A(n10252), .B(n10303), .ZN(n10254) );
  XOR2_X1 U12895 ( .A(n10253), .B(n10254), .Z(n14514) );
  NAND2_X1 U12896 ( .A1(n14513), .A2(n14514), .ZN(n14512) );
  OR2_X1 U12897 ( .A1(n10254), .A2(n10253), .ZN(n10255) );
  XOR2_X1 U12898 ( .A(n10256), .B(n10257), .Z(n14393) );
  NAND2_X1 U12899 ( .A1(n14858), .A2(n10309), .ZN(n10260) );
  OR2_X1 U12900 ( .A1(n14401), .A2(n10310), .ZN(n10259) );
  NAND2_X1 U12901 ( .A1(n10260), .A2(n10259), .ZN(n10261) );
  XNOR2_X1 U12902 ( .A(n10261), .B(n10270), .ZN(n10263) );
  OAI22_X1 U12903 ( .A1(n15036), .A2(n10310), .B1(n14401), .B2(n10314), .ZN(
        n10262) );
  XNOR2_X1 U12904 ( .A(n10263), .B(n10262), .ZN(n14473) );
  OAI22_X1 U12905 ( .A1(n15127), .A2(n10310), .B1(n10264), .B2(n10314), .ZN(
        n10266) );
  OAI22_X1 U12906 ( .A1(n15127), .A2(n10115), .B1(n10264), .B2(n10310), .ZN(
        n10265) );
  XNOR2_X1 U12907 ( .A(n10265), .B(n10270), .ZN(n10267) );
  XOR2_X1 U12908 ( .A(n10266), .B(n10267), .Z(n14399) );
  NAND2_X1 U12909 ( .A1(n14398), .A2(n14399), .ZN(n14397) );
  OR2_X1 U12910 ( .A1(n10267), .A2(n10266), .ZN(n10268) );
  NAND2_X1 U12911 ( .A1(n14397), .A2(n10268), .ZN(n14489) );
  OAI22_X1 U12912 ( .A1(n14817), .A2(n10310), .B1(n10269), .B2(n10314), .ZN(
        n10272) );
  OAI22_X1 U12913 ( .A1(n14817), .A2(n10115), .B1(n10269), .B2(n10310), .ZN(
        n10271) );
  XNOR2_X1 U12914 ( .A(n10271), .B(n10270), .ZN(n10273) );
  XOR2_X1 U12915 ( .A(n10272), .B(n10273), .Z(n14490) );
  NAND2_X1 U12916 ( .A1(n14489), .A2(n14490), .ZN(n14488) );
  NAND2_X1 U12917 ( .A1(n14800), .A2(n10309), .ZN(n10276) );
  NAND2_X1 U12918 ( .A1(n14553), .A2(n10316), .ZN(n10275) );
  NAND2_X1 U12919 ( .A1(n10276), .A2(n10275), .ZN(n10277) );
  XNOR2_X1 U12920 ( .A(n10277), .B(n10303), .ZN(n10278) );
  AOI22_X1 U12921 ( .A1(n14800), .A2(n10316), .B1(n10305), .B2(n14553), .ZN(
        n10279) );
  XNOR2_X1 U12922 ( .A(n10278), .B(n10279), .ZN(n14383) );
  INV_X1 U12923 ( .A(n10278), .ZN(n10280) );
  AOI22_X1 U12924 ( .A1(n15117), .A2(n10316), .B1(n10305), .B2(n14552), .ZN(
        n10284) );
  NAND2_X1 U12925 ( .A1(n15117), .A2(n10309), .ZN(n10282) );
  NAND2_X1 U12926 ( .A1(n14552), .A2(n10307), .ZN(n10281) );
  NAND2_X1 U12927 ( .A1(n10282), .A2(n10281), .ZN(n10283) );
  XNOR2_X1 U12928 ( .A(n10283), .B(n10303), .ZN(n10286) );
  XOR2_X1 U12929 ( .A(n10284), .B(n10286), .Z(n14454) );
  INV_X1 U12930 ( .A(n10284), .ZN(n10285) );
  NAND2_X1 U12931 ( .A1(n14765), .A2(n10309), .ZN(n10289) );
  NAND2_X1 U12932 ( .A1(n14747), .A2(n10307), .ZN(n10288) );
  NAND2_X1 U12933 ( .A1(n10289), .A2(n10288), .ZN(n10290) );
  XNOR2_X1 U12934 ( .A(n10290), .B(n10303), .ZN(n10291) );
  AOI22_X1 U12935 ( .A1(n14765), .A2(n10316), .B1(n10305), .B2(n14747), .ZN(
        n10292) );
  XNOR2_X1 U12936 ( .A(n10291), .B(n10292), .ZN(n14420) );
  INV_X1 U12937 ( .A(n10291), .ZN(n10293) );
  NAND2_X1 U12938 ( .A1(n10293), .A2(n10292), .ZN(n10294) );
  OAI22_X1 U12939 ( .A1(n15002), .A2(n10310), .B1(n10365), .B2(n10314), .ZN(
        n10298) );
  NAND2_X1 U12940 ( .A1(n14753), .A2(n10309), .ZN(n10296) );
  OR2_X1 U12941 ( .A1(n10365), .A2(n10310), .ZN(n10295) );
  NAND2_X1 U12942 ( .A1(n10296), .A2(n10295), .ZN(n10297) );
  XNOR2_X1 U12943 ( .A(n10297), .B(n10303), .ZN(n10299) );
  XOR2_X1 U12944 ( .A(n10298), .B(n10299), .Z(n14526) );
  NOR2_X1 U12945 ( .A1(n10299), .A2(n10298), .ZN(n10300) );
  INV_X1 U12946 ( .A(n14365), .ZN(n10308) );
  NAND2_X1 U12947 ( .A1(n10373), .A2(n10309), .ZN(n10302) );
  NAND2_X1 U12948 ( .A1(n14748), .A2(n10316), .ZN(n10301) );
  NAND2_X1 U12949 ( .A1(n10302), .A2(n10301), .ZN(n10304) );
  XNOR2_X1 U12950 ( .A(n10304), .B(n10303), .ZN(n10325) );
  AND2_X1 U12951 ( .A1(n14748), .A2(n10305), .ZN(n10306) );
  AOI21_X1 U12952 ( .B1(n10373), .B2(n10307), .A(n10306), .ZN(n10323) );
  XNOR2_X1 U12953 ( .A(n10325), .B(n10323), .ZN(n14364) );
  NAND2_X1 U12954 ( .A1(n10308), .A2(n14364), .ZN(n10345) );
  NAND2_X1 U12955 ( .A1(n14738), .A2(n10309), .ZN(n10312) );
  OR2_X1 U12956 ( .A1(n10310), .A2(n10364), .ZN(n10311) );
  NAND2_X1 U12957 ( .A1(n10312), .A2(n10311), .ZN(n10313) );
  XNOR2_X1 U12958 ( .A(n10313), .B(n10190), .ZN(n10318) );
  NOR2_X1 U12959 ( .A1(n10314), .A2(n10364), .ZN(n10315) );
  AOI21_X1 U12960 ( .B1(n14738), .B2(n10316), .A(n10315), .ZN(n10317) );
  XNOR2_X1 U12961 ( .A(n10318), .B(n10317), .ZN(n10339) );
  INV_X1 U12962 ( .A(n10339), .ZN(n10322) );
  INV_X1 U12963 ( .A(n10319), .ZN(n11298) );
  NAND2_X1 U12964 ( .A1(n10331), .A2(n10536), .ZN(n10328) );
  OR2_X1 U12965 ( .A1(n15295), .A2(n10539), .ZN(n10321) );
  NAND2_X1 U12966 ( .A1(n10322), .A2(n14515), .ZN(n10344) );
  INV_X1 U12967 ( .A(n10323), .ZN(n10324) );
  OR2_X1 U12968 ( .A1(n10325), .A2(n10324), .ZN(n10338) );
  AND2_X1 U12969 ( .A1(n10339), .A2(n10326), .ZN(n10327) );
  NAND2_X1 U12970 ( .A1(n10345), .A2(n10327), .ZN(n10343) );
  OR2_X1 U12971 ( .A1(n10863), .A2(n11544), .ZN(n11306) );
  OR2_X1 U12972 ( .A1(n10328), .A2(n11306), .ZN(n10330) );
  INV_X1 U12973 ( .A(n10331), .ZN(n10335) );
  NAND2_X1 U12974 ( .A1(n10335), .A2(n10332), .ZN(n10854) );
  NAND2_X1 U12975 ( .A1(n10854), .A2(n10333), .ZN(n10334) );
  NAND2_X1 U12976 ( .A1(n14748), .A2(n14538), .ZN(n10337) );
  AOI22_X1 U12977 ( .A1(n14521), .A2(n14549), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10336) );
  OAI211_X1 U12978 ( .C1(n14528), .C2(n14735), .A(n10337), .B(n10336), .ZN(
        n10341) );
  NOR3_X1 U12979 ( .A1(n10339), .A2(n14546), .A3(n10338), .ZN(n10340) );
  AOI211_X1 U12980 ( .C1(n14738), .C2(n14544), .A(n10341), .B(n10340), .ZN(
        n10342) );
  OAI211_X1 U12981 ( .C1(n10345), .C2(n10344), .A(n10343), .B(n10342), .ZN(
        P1_U3220) );
  INV_X1 U12982 ( .A(n10348), .ZN(n10349) );
  NAND2_X1 U12983 ( .A1(n6652), .A2(n10349), .ZN(n14741) );
  OAI211_X1 U12984 ( .C1(n12472), .C2(n10372), .A(n10110), .B(n10350), .ZN(
        n14732) );
  OAI21_X1 U12985 ( .B1(n14741), .B2(n15100), .A(n14732), .ZN(n10358) );
  AND2_X1 U12986 ( .A1(n10352), .A2(n10351), .ZN(n10353) );
  AND2_X1 U12987 ( .A1(n10361), .A2(n10353), .ZN(n10354) );
  OAI21_X1 U12988 ( .B1(n10355), .B2(n10354), .A(n15331), .ZN(n10357) );
  AOI22_X1 U12989 ( .A1(n14748), .A2(n14939), .B1(n14940), .B2(n14549), .ZN(
        n10356) );
  NAND2_X1 U12990 ( .A1(n10357), .A2(n10356), .ZN(n14734) );
  NOR2_X1 U12991 ( .A1(n10358), .A2(n14734), .ZN(n12469) );
  MUX2_X1 U12992 ( .A(n10359), .B(n12469), .S(n15342), .Z(n10360) );
  NAND2_X1 U12993 ( .A1(n10360), .A2(n7838), .ZN(P1_U3524) );
  INV_X1 U12994 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10376) );
  OAI21_X1 U12995 ( .B1(n10363), .B2(n10362), .A(n10361), .ZN(n10366) );
  OAI22_X1 U12996 ( .A1(n10365), .A2(n14907), .B1(n10364), .B2(n14909), .ZN(
        n14370) );
  AOI21_X1 U12997 ( .B1(n10366), .B2(n15331), .A(n14370), .ZN(n10370) );
  INV_X1 U12998 ( .A(n15310), .ZN(n15320) );
  INV_X1 U12999 ( .A(n10371), .ZN(n14745) );
  AOI211_X1 U13000 ( .C1(n10373), .C2(n14745), .A(n15323), .B(n10372), .ZN(
        n12401) );
  NAND2_X1 U13001 ( .A1(n10377), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n10378) );
  XNOR2_X1 U13002 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .ZN(n12551) );
  XNOR2_X1 U13003 ( .A(n12553), .B(n12551), .ZN(n13483) );
  NAND2_X1 U13004 ( .A1(n13483), .A2(n8470), .ZN(n10381) );
  OR2_X1 U13005 ( .A1(n12569), .A2(n15777), .ZN(n10380) );
  INV_X1 U13006 ( .A(n12550), .ZN(n12754) );
  INV_X1 U13007 ( .A(n12611), .ZN(n10382) );
  INV_X1 U13008 ( .A(n10391), .ZN(n13128) );
  AOI211_X1 U13009 ( .C1(n13128), .C2(n8579), .A(n15508), .B(n10382), .ZN(
        n10394) );
  NOR4_X1 U13010 ( .A1(n12611), .A2(n10383), .A3(n10391), .A4(n15508), .ZN(
        n10393) );
  INV_X1 U13011 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n15807) );
  OR2_X1 U13012 ( .A1(n6534), .A2(n15807), .ZN(n10388) );
  INV_X1 U13013 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n10384) );
  OR2_X1 U13014 ( .A1(n12562), .A2(n10384), .ZN(n10387) );
  INV_X1 U13015 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n10385) );
  OR2_X1 U13016 ( .A1(n12563), .A2(n10385), .ZN(n10386) );
  OR2_X1 U13017 ( .A1(n7986), .A2(n10389), .ZN(n10390) );
  NAND2_X1 U13018 ( .A1(n13320), .A2(n10390), .ZN(n13107) );
  OAI22_X1 U13019 ( .A1(n10391), .A2(n15492), .B1(n12584), .B2(n13107), .ZN(
        n10392) );
  INV_X1 U13020 ( .A(n10396), .ZN(n12577) );
  NOR2_X1 U13021 ( .A1(n12577), .A2(n15512), .ZN(n13115) );
  OR2_X1 U13022 ( .A1(n10403), .A2(n15546), .ZN(n10402) );
  XNOR2_X1 U13023 ( .A(n12591), .B(n12611), .ZN(n13119) );
  OR2_X1 U13024 ( .A1(n15549), .A2(n10398), .ZN(n10399) );
  NAND2_X1 U13025 ( .A1(n10402), .A2(n10401), .ZN(P3_U3488) );
  OAI22_X1 U13026 ( .A1(n13119), .A2(n13461), .B1(n15540), .B2(n10404), .ZN(
        n10405) );
  INV_X1 U13027 ( .A(n10405), .ZN(n10406) );
  NAND2_X1 U13028 ( .A1(n10407), .A2(n10406), .ZN(P3_U3456) );
  INV_X1 U13029 ( .A(n10408), .ZN(n10552) );
  OR2_X2 U13030 ( .A1(n10409), .A2(n10552), .ZN(n14570) );
  INV_X1 U13031 ( .A(n10410), .ZN(n10413) );
  AND2_X1 U13032 ( .A1(n11907), .A2(n10411), .ZN(n10412) );
  NAND2_X1 U13033 ( .A1(n10413), .A2(n10412), .ZN(n10577) );
  AOI211_X1 U13034 ( .C1(n10415), .C2(n10414), .A(n13030), .B(n6702), .ZN(
        n10428) );
  OR3_X1 U13035 ( .A1(n12983), .A2(n10417), .A3(n10416), .ZN(n10418) );
  AOI21_X1 U13036 ( .B1(n10419), .B2(n10418), .A(n13046), .ZN(n10427) );
  NAND3_X1 U13037 ( .A1(n12978), .A2(n6718), .A3(n10420), .ZN(n10421) );
  AOI21_X1 U13038 ( .B1(n10422), .B2(n10421), .A(n13077), .ZN(n10426) );
  NAND2_X1 U13039 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n12334)
         );
  INV_X1 U13040 ( .A(n12334), .ZN(n10423) );
  AOI21_X1 U13041 ( .B1(n15467), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n10423), 
        .ZN(n10424) );
  OAI21_X1 U13042 ( .B1(n13088), .B2(n10567), .A(n10424), .ZN(n10425) );
  INV_X1 U13043 ( .A(n10430), .ZN(n10431) );
  AOI211_X1 U13044 ( .C1(n10432), .C2(n10429), .A(n14546), .B(n10431), .ZN(
        n10437) );
  MUX2_X1 U13045 ( .A(n14539), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n10436) );
  NAND2_X1 U13046 ( .A1(n14939), .A2(n9433), .ZN(n10434) );
  NAND2_X1 U13047 ( .A1(n14940), .A2(n14568), .ZN(n10433) );
  AND2_X1 U13048 ( .A1(n10434), .A2(n10433), .ZN(n15272) );
  OAI22_X1 U13049 ( .A1(n14524), .A2(n15315), .B1(n15272), .B2(n14458), .ZN(
        n10435) );
  OR3_X1 U13050 ( .A1(n10437), .A2(n10436), .A3(n10435), .ZN(P1_U3218) );
  NAND2_X1 U13051 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_STATE_REG_SCAN_IN), .ZN(
        n10438) );
  OAI21_X1 U13052 ( .B1(n10439), .B2(P3_STATE_REG_SCAN_IN), .A(n10438), .ZN(
        P3_U3295) );
  NOR2_X1 U13053 ( .A1(n6545), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13480) );
  OAI222_X1 U13054 ( .A1(n13495), .A2(n10441), .B1(n11197), .B2(P3_U3151), 
        .C1(n10440), .C2(n13487), .ZN(P3_U3294) );
  INV_X1 U13055 ( .A(n13487), .ZN(n10973) );
  AOI222_X1 U13056 ( .A1(n10442), .A2(n13480), .B1(SI_2_), .B2(n10973), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n11161), .ZN(n10443) );
  INV_X1 U13057 ( .A(n10443), .ZN(P3_U3293) );
  OAI222_X1 U13058 ( .A1(n13487), .A2(n10446), .B1(n10445), .B2(P3_U3151), 
        .C1(n13495), .C2(n10444), .ZN(P3_U3289) );
  AOI222_X1 U13059 ( .A1(n10447), .A2(n13480), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11215), .C1(SI_5_), .C2(n10973), .ZN(n10448) );
  INV_X1 U13060 ( .A(n10448), .ZN(P3_U3290) );
  AOI222_X1 U13061 ( .A1(n10449), .A2(n13480), .B1(n11106), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n10973), .ZN(n10450) );
  INV_X1 U13062 ( .A(n10450), .ZN(P3_U3291) );
  AOI222_X1 U13063 ( .A1(n10452), .A2(n13480), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10451), .C1(SI_3_), .C2(n10973), .ZN(n10453) );
  INV_X1 U13064 ( .A(n10453), .ZN(P3_U3292) );
  AOI222_X1 U13065 ( .A1(n10455), .A2(n13480), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10454), .C1(SI_7_), .C2(n10973), .ZN(n10456) );
  INV_X1 U13066 ( .A(n10456), .ZN(P3_U3288) );
  NAND2_X1 U13067 ( .A1(n14572), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10457) );
  NAND2_X1 U13068 ( .A1(n15554), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10460) );
  INV_X1 U13069 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U13070 ( .A1(n10458), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10459) );
  NAND2_X1 U13071 ( .A1(n10469), .A2(n10468), .ZN(n10461) );
  INV_X1 U13072 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10462) );
  XNOR2_X1 U13073 ( .A(n10504), .B(n10463), .ZN(n10464) );
  NAND2_X1 U13074 ( .A1(n10464), .A2(n15556), .ZN(n10506) );
  OR2_X1 U13075 ( .A1(n10464), .A2(n15556), .ZN(n10465) );
  INV_X1 U13076 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10466) );
  XNOR2_X1 U13077 ( .A(n10467), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n10478) );
  XNOR2_X1 U13078 ( .A(n10469), .B(n10468), .ZN(n15234) );
  NAND2_X1 U13079 ( .A1(n15234), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10475) );
  XNOR2_X1 U13080 ( .A(n10470), .B(n10471), .ZN(n10474) );
  INV_X1 U13081 ( .A(n10471), .ZN(n10472) );
  OAI21_X1 U13082 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n10473), .A(n10472), .ZN(
        n15168) );
  NAND2_X1 U13083 ( .A1(n15168), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n15867) );
  XNOR2_X1 U13084 ( .A(n10474), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(n15866) );
  NOR2_X1 U13085 ( .A1(n15867), .A2(n15866), .ZN(n15865) );
  AOI21_X1 U13086 ( .B1(n10474), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n15865), .ZN(
        n15233) );
  NAND2_X1 U13087 ( .A1(n10475), .A2(n15233), .ZN(n10477) );
  OR2_X1 U13088 ( .A1(n15234), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n10476) );
  NAND2_X1 U13089 ( .A1(n10477), .A2(n10476), .ZN(n10479) );
  NAND2_X1 U13090 ( .A1(n10478), .A2(n10479), .ZN(n15862) );
  NAND2_X1 U13091 ( .A1(n15862), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n10482) );
  INV_X1 U13092 ( .A(n10478), .ZN(n10481) );
  INV_X1 U13093 ( .A(n10479), .ZN(n10480) );
  NAND2_X1 U13094 ( .A1(n10481), .A2(n10480), .ZN(n15863) );
  NAND2_X1 U13095 ( .A1(n10482), .A2(n15863), .ZN(n10483) );
  NAND2_X1 U13096 ( .A1(n10484), .A2(n10483), .ZN(n10511) );
  OAI21_X1 U13097 ( .B1(n10484), .B2(n10483), .A(n10511), .ZN(n10485) );
  INV_X1 U13098 ( .A(n10485), .ZN(SUB_1596_U59) );
  INV_X1 U13099 ( .A(n10649), .ZN(n10657) );
  NOR2_X1 U13100 ( .A1(n6546), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14356) );
  INV_X2 U13101 ( .A(n14356), .ZN(n14362) );
  INV_X1 U13102 ( .A(n10486), .ZN(n10488) );
  OAI222_X1 U13103 ( .A1(P2_U3088), .A2(n10657), .B1(n14362), .B2(n10487), 
        .C1(n14360), .C2(n10488), .ZN(P2_U3324) );
  NAND2_X1 U13104 ( .A1(n6546), .A2(P1_U3086), .ZN(n12476) );
  NOR2_X1 U13105 ( .A1(n6545), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15155) );
  INV_X2 U13106 ( .A(n15155), .ZN(n12474) );
  OAI222_X1 U13107 ( .A1(n14612), .A2(P1_U3086), .B1(n12476), .B2(n10489), 
        .C1(n12474), .C2(n10488), .ZN(P1_U3352) );
  INV_X1 U13108 ( .A(n10490), .ZN(n10519) );
  OAI222_X1 U13109 ( .A1(n15350), .A2(P2_U3088), .B1(n14360), .B2(n10519), 
        .C1(n10491), .C2(n14362), .ZN(P2_U3325) );
  INV_X1 U13110 ( .A(n10664), .ZN(n10672) );
  INV_X1 U13111 ( .A(n10492), .ZN(n10521) );
  OAI222_X1 U13112 ( .A1(n10672), .A2(P2_U3088), .B1(n14360), .B2(n10521), 
        .C1(n10493), .C2(n14362), .ZN(P2_U3322) );
  INV_X1 U13113 ( .A(n10494), .ZN(n10516) );
  OAI222_X1 U13114 ( .A1(n15362), .A2(P2_U3088), .B1(n14360), .B2(n10516), 
        .C1(n10495), .C2(n14362), .ZN(P2_U3323) );
  OAI222_X1 U13115 ( .A1(n13495), .A2(n10497), .B1(n12028), .B2(P3_U3151), 
        .C1(n10496), .C2(n13487), .ZN(P3_U3286) );
  INV_X1 U13116 ( .A(n10498), .ZN(n10512) );
  AOI22_X1 U13117 ( .A1(n15377), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n14356), .ZN(n10499) );
  OAI21_X1 U13118 ( .B1(n10512), .B2(n14360), .A(n10499), .ZN(P2_U3321) );
  INV_X1 U13119 ( .A(n10500), .ZN(n10501) );
  OAI222_X1 U13120 ( .A1(n13487), .A2(n10502), .B1(n7489), .B2(P3_U3151), .C1(
        n13495), .C2(n10501), .ZN(P3_U3287) );
  OAI222_X1 U13121 ( .A1(n14362), .A2(n10503), .B1(n14360), .B2(n12473), .C1(
        n10597), .C2(P2_U3088), .ZN(P2_U3326) );
  NAND2_X1 U13122 ( .A1(n10504), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10505) );
  NAND2_X1 U13123 ( .A1(n10506), .A2(n10505), .ZN(n10507) );
  NAND2_X1 U13124 ( .A1(n10507), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10560) );
  INV_X1 U13125 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14635) );
  NAND2_X1 U13126 ( .A1(n10509), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n10510) );
  INV_X1 U13127 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10663) );
  XNOR2_X1 U13128 ( .A(n10555), .B(n10663), .ZN(SUB_1596_U58) );
  INV_X1 U13129 ( .A(n14656), .ZN(n10514) );
  OAI222_X1 U13130 ( .A1(n10514), .A2(P1_U3086), .B1(n12476), .B2(n10513), 
        .C1(n12474), .C2(n10512), .ZN(P1_U3349) );
  INV_X1 U13131 ( .A(n14625), .ZN(n10517) );
  INV_X1 U13132 ( .A(n12476), .ZN(n10716) );
  INV_X1 U13133 ( .A(n10716), .ZN(n15161) );
  OAI222_X1 U13134 ( .A1(P1_U3086), .A2(n10517), .B1(n12474), .B2(n10516), 
        .C1(n10515), .C2(n15161), .ZN(P1_U3351) );
  OAI222_X1 U13135 ( .A1(P1_U3086), .A2(n14596), .B1(n12474), .B2(n10519), 
        .C1(n10518), .C2(n15161), .ZN(P1_U3353) );
  INV_X1 U13136 ( .A(n14637), .ZN(n10522) );
  OAI222_X1 U13137 ( .A1(P1_U3086), .A2(n10522), .B1(n12474), .B2(n10521), 
        .C1(n10520), .C2(n15161), .ZN(P1_U3350) );
  INV_X1 U13138 ( .A(n10523), .ZN(n10525) );
  OAI222_X1 U13139 ( .A1(n14671), .A2(P1_U3086), .B1(n15161), .B2(n10524), 
        .C1(n12474), .C2(n10525), .ZN(P1_U3348) );
  INV_X1 U13140 ( .A(n13913), .ZN(n10527) );
  OAI222_X1 U13141 ( .A1(P2_U3088), .A2(n10527), .B1(n14362), .B2(n10526), 
        .C1(n14360), .C2(n10525), .ZN(P2_U3320) );
  OAI222_X1 U13142 ( .A1(n13495), .A2(n10530), .B1(n10529), .B2(P3_U3151), 
        .C1(n10528), .C2(n13487), .ZN(P3_U3285) );
  INV_X1 U13143 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10535) );
  NOR3_X1 U13144 ( .A1(n10533), .A2(n10532), .A3(n10552), .ZN(n10534) );
  AOI21_X1 U13145 ( .B1(n15859), .B2(n10535), .A(n10534), .ZN(P1_U3446) );
  OR2_X1 U13146 ( .A1(n10536), .A2(n9386), .ZN(n10743) );
  INV_X1 U13147 ( .A(n10743), .ZN(n10540) );
  AOI21_X1 U13148 ( .B1(n10539), .B2(n10538), .A(n10537), .ZN(n10742) );
  NOR2_X1 U13149 ( .A1(n15244), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U13150 ( .A(n10809), .ZN(n10542) );
  OAI222_X1 U13151 ( .A1(n10542), .A2(P1_U3086), .B1(n15161), .B2(n10541), 
        .C1(n12474), .C2(n6896), .ZN(P1_U3347) );
  INV_X1 U13152 ( .A(n10707), .ZN(n10714) );
  OAI222_X1 U13153 ( .A1(P2_U3088), .A2(n10714), .B1(n14362), .B2(n10543), 
        .C1(n14360), .C2(n6896), .ZN(P2_U3319) );
  NAND2_X1 U13154 ( .A1(P1_U4016), .A2(n12392), .ZN(n10544) );
  OAI21_X1 U13155 ( .B1(P1_U4016), .B2(n10545), .A(n10544), .ZN(P1_U3560) );
  OAI222_X1 U13156 ( .A1(n13495), .A2(n10547), .B1(n12982), .B2(P3_U3151), 
        .C1(n10546), .C2(n13487), .ZN(P3_U3284) );
  INV_X1 U13157 ( .A(n10931), .ZN(n10639) );
  OAI222_X1 U13158 ( .A1(P2_U3088), .A2(n10639), .B1(n14362), .B2(n10548), 
        .C1(n14360), .C2(n10549), .ZN(P2_U3318) );
  INV_X1 U13159 ( .A(n10793), .ZN(n10551) );
  OAI222_X1 U13160 ( .A1(n10551), .A2(P1_U3086), .B1(n15161), .B2(n10550), 
        .C1(n12474), .C2(n10549), .ZN(P1_U3346) );
  INV_X1 U13161 ( .A(n15859), .ZN(n15293) );
  OAI22_X1 U13162 ( .A1(n15293), .A2(P1_D_REG_0__SCAN_IN), .B1(n10553), .B2(
        n10552), .ZN(n10554) );
  INV_X1 U13163 ( .A(n10554), .ZN(P1_U3445) );
  INV_X1 U13164 ( .A(n10556), .ZN(n10558) );
  NAND2_X1 U13165 ( .A1(n10558), .A2(n10557), .ZN(n10559) );
  OAI21_X1 U13166 ( .B1(n10561), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10560), .ZN(
        n10778) );
  XNOR2_X1 U13167 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n10562) );
  XNOR2_X1 U13168 ( .A(n10778), .B(n10562), .ZN(n10563) );
  OAI21_X1 U13169 ( .B1(n10564), .B2(n10563), .A(n10783), .ZN(n10565) );
  INV_X1 U13170 ( .A(n10565), .ZN(SUB_1596_U57) );
  OAI222_X1 U13171 ( .A1(n13487), .A2(n10568), .B1(n10567), .B2(P3_U3151), 
        .C1(n13495), .C2(n10566), .ZN(P3_U3283) );
  INV_X1 U13172 ( .A(n10840), .ZN(n10791) );
  OAI222_X1 U13173 ( .A1(n10791), .A2(P1_U3086), .B1(n15161), .B2(n10569), 
        .C1(n12474), .C2(n10570), .ZN(P1_U3345) );
  INV_X1 U13174 ( .A(n10946), .ZN(n10940) );
  OAI222_X1 U13175 ( .A1(P2_U3088), .A2(n10940), .B1(n14362), .B2(n10571), 
        .C1(n14360), .C2(n10570), .ZN(P2_U3317) );
  OAI222_X1 U13176 ( .A1(n13487), .A2(n10573), .B1(n12998), .B2(P3_U3151), 
        .C1(n13495), .C2(n10572), .ZN(P3_U3282) );
  NAND2_X1 U13177 ( .A1(n10574), .A2(n11907), .ZN(n10575) );
  NAND2_X1 U13178 ( .A1(n10575), .A2(n7247), .ZN(n10576) );
  AND2_X1 U13179 ( .A1(n10577), .A2(n10576), .ZN(n10578) );
  NAND2_X1 U13180 ( .A1(n10589), .A2(n10580), .ZN(n15349) );
  INV_X1 U13181 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11073) );
  AND2_X1 U13182 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10584) );
  INV_X1 U13183 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11508) );
  MUX2_X1 U13184 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n11508), .S(n10597), .Z(
        n10579) );
  INV_X1 U13185 ( .A(n10579), .ZN(n10583) );
  OR2_X1 U13186 ( .A1(n10580), .A2(P2_U3088), .ZN(n14357) );
  XNOR2_X1 U13187 ( .A(n10581), .B(P2_IR_REG_27__SCAN_IN), .ZN(n13881) );
  INV_X1 U13188 ( .A(n13881), .ZN(n14363) );
  NOR2_X1 U13189 ( .A1(n14357), .A2(n14363), .ZN(n10582) );
  OAI211_X1 U13190 ( .C1(n10584), .C2(n10583), .A(n15394), .B(n10619), .ZN(
        n10585) );
  OAI21_X1 U13191 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n11073), .A(n10585), .ZN(
        n10594) );
  AND2_X1 U13192 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10586) );
  INV_X1 U13193 ( .A(n10586), .ZN(n10592) );
  INV_X1 U13194 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10696) );
  MUX2_X1 U13195 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n10696), .S(n10597), .Z(
        n10591) );
  MUX2_X1 U13196 ( .A(n10696), .B(P2_REG1_REG_1__SCAN_IN), .S(n10597), .Z(
        n10587) );
  NAND2_X1 U13197 ( .A1(n10587), .A2(n10586), .ZN(n10599) );
  INV_X1 U13198 ( .A(n10599), .ZN(n10590) );
  NOR2_X1 U13199 ( .A1(n14357), .A2(n13881), .ZN(n10588) );
  NAND2_X1 U13200 ( .A1(n10589), .A2(n10588), .ZN(n15420) );
  AOI211_X1 U13201 ( .C1(n10592), .C2(n10591), .A(n10590), .B(n15420), .ZN(
        n10593) );
  AOI211_X1 U13202 ( .C1(n15408), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n10594), .B(
        n10593), .ZN(n10595) );
  OAI21_X1 U13203 ( .B1(n10597), .B2(n15412), .A(n10595), .ZN(P2_U3215) );
  XNOR2_X1 U13204 ( .A(n10931), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n10929) );
  INV_X1 U13205 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10596) );
  MUX2_X1 U13206 ( .A(n10596), .B(P2_REG1_REG_2__SCAN_IN), .S(n15350), .Z(
        n15354) );
  NAND2_X1 U13207 ( .A1(n9591), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10598) );
  NAND2_X1 U13208 ( .A1(n10599), .A2(n10598), .ZN(n15353) );
  NAND2_X1 U13209 ( .A1(n10620), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10644) );
  NAND2_X1 U13210 ( .A1(n15352), .A2(n10644), .ZN(n10602) );
  INV_X1 U13211 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10600) );
  MUX2_X1 U13212 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10600), .S(n10649), .Z(
        n10601) );
  NAND2_X1 U13213 ( .A1(n10602), .A2(n10601), .ZN(n10647) );
  NAND2_X1 U13214 ( .A1(n10649), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10603) );
  NAND2_X1 U13215 ( .A1(n10647), .A2(n10603), .ZN(n15365) );
  INV_X1 U13216 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10604) );
  MUX2_X1 U13217 ( .A(n10604), .B(P2_REG1_REG_4__SCAN_IN), .S(n15362), .Z(
        n15366) );
  NAND2_X1 U13218 ( .A1(n10624), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10658) );
  NAND2_X1 U13219 ( .A1(n15364), .A2(n10658), .ZN(n10607) );
  INV_X1 U13220 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10605) );
  MUX2_X1 U13221 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10605), .S(n10664), .Z(
        n10606) );
  NAND2_X1 U13222 ( .A1(n10607), .A2(n10606), .ZN(n10661) );
  NAND2_X1 U13223 ( .A1(n10664), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10608) );
  NAND2_X1 U13224 ( .A1(n10661), .A2(n10608), .ZN(n15379) );
  INV_X1 U13225 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10609) );
  MUX2_X1 U13226 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10609), .S(n15377), .Z(
        n15380) );
  NAND2_X1 U13227 ( .A1(n15377), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n13915) );
  NAND2_X1 U13228 ( .A1(n15378), .A2(n13915), .ZN(n10612) );
  INV_X1 U13229 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10610) );
  MUX2_X1 U13230 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10610), .S(n13913), .Z(
        n10611) );
  NAND2_X1 U13231 ( .A1(n10612), .A2(n10611), .ZN(n13917) );
  NAND2_X1 U13232 ( .A1(n13913), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10613) );
  NAND2_X1 U13233 ( .A1(n13917), .A2(n10613), .ZN(n10702) );
  INV_X1 U13234 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10614) );
  XNOR2_X1 U13235 ( .A(n10707), .B(n10614), .ZN(n10703) );
  NAND2_X1 U13236 ( .A1(n10702), .A2(n10703), .ZN(n10616) );
  NAND2_X1 U13237 ( .A1(n10707), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10615) );
  NAND2_X1 U13238 ( .A1(n10616), .A2(n10615), .ZN(n10930) );
  XOR2_X1 U13239 ( .A(n10929), .B(n10930), .Z(n10643) );
  INV_X1 U13240 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10617) );
  MUX2_X1 U13241 ( .A(n10617), .B(P2_REG2_REG_2__SCAN_IN), .S(n15350), .Z(
        n15357) );
  NAND2_X1 U13242 ( .A1(n9591), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10618) );
  NAND2_X1 U13243 ( .A1(n10619), .A2(n10618), .ZN(n15356) );
  NAND2_X1 U13244 ( .A1(n10620), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10650) );
  NAND2_X1 U13245 ( .A1(n15355), .A2(n10650), .ZN(n10622) );
  INV_X1 U13246 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11681) );
  MUX2_X1 U13247 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11681), .S(n10649), .Z(
        n10621) );
  NAND2_X1 U13248 ( .A1(n10622), .A2(n10621), .ZN(n10653) );
  NAND2_X1 U13249 ( .A1(n10649), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10623) );
  NAND2_X1 U13250 ( .A1(n10653), .A2(n10623), .ZN(n15368) );
  INV_X1 U13251 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11674) );
  MUX2_X1 U13252 ( .A(n11674), .B(P2_REG2_REG_4__SCAN_IN), .S(n15362), .Z(
        n15369) );
  NAND2_X1 U13253 ( .A1(n10624), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10666) );
  NAND2_X1 U13254 ( .A1(n15367), .A2(n10666), .ZN(n10626) );
  INV_X1 U13255 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11690) );
  MUX2_X1 U13256 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n11690), .S(n10664), .Z(
        n10625) );
  NAND2_X1 U13257 ( .A1(n10626), .A2(n10625), .ZN(n10668) );
  NAND2_X1 U13258 ( .A1(n10664), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10627) );
  NAND2_X1 U13259 ( .A1(n10668), .A2(n10627), .ZN(n15382) );
  INV_X1 U13260 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11705) );
  MUX2_X1 U13261 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11705), .S(n15377), .Z(
        n15383) );
  NAND2_X1 U13262 ( .A1(n15377), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n13910) );
  NAND2_X1 U13263 ( .A1(n15381), .A2(n13910), .ZN(n10629) );
  MUX2_X1 U13264 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11729), .S(n13913), .Z(
        n10628) );
  NAND2_X1 U13265 ( .A1(n10629), .A2(n10628), .ZN(n13912) );
  NAND2_X1 U13266 ( .A1(n13913), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10709) );
  NAND2_X1 U13267 ( .A1(n13912), .A2(n10709), .ZN(n10631) );
  MUX2_X1 U13268 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11742), .S(n10707), .Z(
        n10630) );
  NAND2_X1 U13269 ( .A1(n10631), .A2(n10630), .ZN(n10711) );
  NAND2_X1 U13270 ( .A1(n10707), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10632) );
  NAND2_X1 U13271 ( .A1(n10711), .A2(n10632), .ZN(n10634) );
  INV_X1 U13272 ( .A(n10634), .ZN(n10636) );
  MUX2_X1 U13273 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11626), .S(n10931), .Z(
        n10635) );
  INV_X1 U13274 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11626) );
  MUX2_X1 U13275 ( .A(n11626), .B(P2_REG2_REG_9__SCAN_IN), .S(n10931), .Z(
        n10633) );
  OAI21_X1 U13276 ( .B1(n10636), .B2(n10635), .A(n10924), .ZN(n10641) );
  NOR2_X1 U13277 ( .A1(n10637), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11757) );
  AOI21_X1 U13278 ( .B1(n15408), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n11757), .ZN(
        n10638) );
  OAI21_X1 U13279 ( .B1(n10639), .B2(n15412), .A(n10638), .ZN(n10640) );
  AOI21_X1 U13280 ( .B1(n15394), .B2(n10641), .A(n10640), .ZN(n10642) );
  OAI21_X1 U13281 ( .B1(n10643), .B2(n15420), .A(n10642), .ZN(P2_U3223) );
  MUX2_X1 U13282 ( .A(n10600), .B(P2_REG1_REG_3__SCAN_IN), .S(n10649), .Z(
        n10645) );
  NAND3_X1 U13283 ( .A1(n15352), .A2(n10645), .A3(n10644), .ZN(n10646) );
  AND3_X1 U13284 ( .A1(n15398), .A2(n10647), .A3(n10646), .ZN(n10648) );
  AOI21_X1 U13285 ( .B1(n15408), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n10648), .ZN(
        n10656) );
  MUX2_X1 U13286 ( .A(n11681), .B(P2_REG2_REG_3__SCAN_IN), .S(n10649), .Z(
        n10651) );
  NAND3_X1 U13287 ( .A1(n10651), .A2(n15355), .A3(n10650), .ZN(n10652) );
  AND3_X1 U13288 ( .A1(n15394), .A2(n10653), .A3(n10652), .ZN(n10654) );
  AOI21_X1 U13289 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_U3088), .A(n10654), 
        .ZN(n10655) );
  OAI211_X1 U13290 ( .C1(n10657), .C2(n15412), .A(n10656), .B(n10655), .ZN(
        P2_U3217) );
  INV_X1 U13291 ( .A(n15408), .ZN(n15406) );
  MUX2_X1 U13292 ( .A(n10605), .B(P2_REG1_REG_5__SCAN_IN), .S(n10664), .Z(
        n10659) );
  NAND3_X1 U13293 ( .A1(n15364), .A2(n10659), .A3(n10658), .ZN(n10660) );
  NAND3_X1 U13294 ( .A1(n15398), .A2(n10661), .A3(n10660), .ZN(n10662) );
  OAI21_X1 U13295 ( .B1(n15406), .B2(n10663), .A(n10662), .ZN(n10670) );
  AND2_X1 U13296 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n11087) );
  MUX2_X1 U13297 ( .A(n11690), .B(P2_REG2_REG_5__SCAN_IN), .S(n10664), .Z(
        n10665) );
  NAND3_X1 U13298 ( .A1(n15367), .A2(n10666), .A3(n10665), .ZN(n10667) );
  AND3_X1 U13299 ( .A1(n15394), .A2(n10668), .A3(n10667), .ZN(n10669) );
  NOR3_X1 U13300 ( .A1(n10670), .A2(n11087), .A3(n10669), .ZN(n10671) );
  OAI21_X1 U13301 ( .B1(n10672), .B2(n15412), .A(n10671), .ZN(P2_U3219) );
  INV_X1 U13302 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10673) );
  NAND2_X1 U13303 ( .A1(n15394), .A2(n10673), .ZN(n10674) );
  OAI211_X1 U13304 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15420), .A(n10674), .B(
        n15412), .ZN(n10675) );
  INV_X1 U13305 ( .A(n10675), .ZN(n10678) );
  AOI22_X1 U13306 ( .A1(n15398), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15394), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10677) );
  MUX2_X1 U13307 ( .A(n10678), .B(n10677), .S(n10676), .Z(n10680) );
  AOI22_X1 U13308 ( .A1(n15408), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10679) );
  NAND2_X1 U13309 ( .A1(n10680), .A2(n10679), .ZN(P2_U3214) );
  AND2_X1 U13310 ( .A1(n15432), .A2(n10681), .ZN(n15433) );
  AND3_X1 U13311 ( .A1(n11325), .A2(n10682), .A3(n11327), .ZN(n10683) );
  XNOR2_X1 U13312 ( .A(n10822), .B(n10871), .ZN(n10687) );
  XOR2_X1 U13313 ( .A(n10865), .B(n13846), .Z(n11503) );
  NAND2_X1 U13314 ( .A1(n11924), .A2(n9912), .ZN(n13642) );
  NAND2_X1 U13315 ( .A1(n10687), .A2(n13641), .ZN(n10873) );
  OAI21_X1 U13316 ( .B1(n13641), .B2(n13846), .A(n10873), .ZN(n10689) );
  NAND2_X1 U13317 ( .A1(n13884), .A2(n9912), .ZN(n13803) );
  NAND2_X1 U13318 ( .A1(n13877), .A2(n10080), .ZN(n10688) );
  NAND2_X1 U13319 ( .A1(n10689), .A2(n14180), .ZN(n10691) );
  AOI22_X1 U13320 ( .A1(n14108), .A2(n13906), .B1(n14106), .B2(n10686), .ZN(
        n10690) );
  NAND2_X1 U13321 ( .A1(n10691), .A2(n10690), .ZN(n11505) );
  INV_X1 U13322 ( .A(n11505), .ZN(n10694) );
  AND2_X1 U13323 ( .A1(n10871), .A2(n11717), .ZN(n10692) );
  NOR2_X1 U13324 ( .A1(n10869), .A2(n10692), .ZN(n11504) );
  AOI22_X1 U13325 ( .A1(n11504), .A2(n14308), .B1(n14315), .B2(n10871), .ZN(
        n10693) );
  OAI211_X1 U13326 ( .C1(n11503), .C2(n14319), .A(n10694), .B(n10693), .ZN(
        n10969) );
  NAND2_X1 U13327 ( .A1(n15466), .A2(n10969), .ZN(n10695) );
  OAI21_X1 U13328 ( .B1(n15466), .B2(n10696), .A(n10695), .ZN(P2_U3500) );
  INV_X1 U13329 ( .A(n11020), .ZN(n10699) );
  INV_X1 U13330 ( .A(n10697), .ZN(n10701) );
  OAI222_X1 U13331 ( .A1(P1_U3086), .A2(n10699), .B1(n12474), .B2(n10701), 
        .C1(n10698), .C2(n15161), .ZN(P1_U3344) );
  INV_X1 U13332 ( .A(n11469), .ZN(n10953) );
  OAI222_X1 U13333 ( .A1(n10953), .A2(P2_U3088), .B1(n14360), .B2(n10701), 
        .C1(n10700), .C2(n14362), .ZN(P2_U3316) );
  NAND2_X1 U13334 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n11412) );
  XOR2_X1 U13335 ( .A(n10702), .B(n10703), .Z(n10704) );
  NAND2_X1 U13336 ( .A1(n15398), .A2(n10704), .ZN(n10705) );
  NAND2_X1 U13337 ( .A1(n11412), .A2(n10705), .ZN(n10706) );
  AOI21_X1 U13338 ( .B1(n15408), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n10706), .ZN(
        n10713) );
  MUX2_X1 U13339 ( .A(n11742), .B(P2_REG2_REG_8__SCAN_IN), .S(n10707), .Z(
        n10708) );
  NAND3_X1 U13340 ( .A1(n13912), .A2(n10709), .A3(n10708), .ZN(n10710) );
  NAND3_X1 U13341 ( .A1(n15394), .A2(n10711), .A3(n10710), .ZN(n10712) );
  OAI211_X1 U13342 ( .C1(n15412), .C2(n10714), .A(n10713), .B(n10712), .ZN(
        P2_U3222) );
  INV_X1 U13343 ( .A(n10715), .ZN(n10831) );
  AOI22_X1 U13344 ( .A1(n11133), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10716), .ZN(n10717) );
  OAI21_X1 U13345 ( .B1(n10831), .B2(n12474), .A(n10717), .ZN(P1_U3343) );
  MUX2_X1 U13346 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n8915), .S(n10793), .Z(
        n10738) );
  OR2_X1 U13347 ( .A1(n10809), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10737) );
  INV_X1 U13348 ( .A(n10737), .ZN(n10718) );
  NOR2_X1 U13349 ( .A1(n10738), .A2(n10718), .ZN(n10741) );
  INV_X1 U13350 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10719) );
  MUX2_X1 U13351 ( .A(n10719), .B(P1_REG1_REG_1__SCAN_IN), .S(n12477), .Z(
        n14575) );
  AND2_X1 U13352 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n14576) );
  NAND2_X1 U13353 ( .A1(n14575), .A2(n14576), .ZN(n14598) );
  INV_X1 U13354 ( .A(n12477), .ZN(n14574) );
  NAND2_X1 U13355 ( .A1(n14574), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n14597) );
  NAND2_X1 U13356 ( .A1(n14598), .A2(n14597), .ZN(n10722) );
  INV_X1 U13357 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10720) );
  MUX2_X1 U13358 ( .A(n10720), .B(P1_REG1_REG_2__SCAN_IN), .S(n14596), .Z(
        n10721) );
  NAND2_X1 U13359 ( .A1(n10722), .A2(n10721), .ZN(n14606) );
  OR2_X1 U13360 ( .A1(n14596), .A2(n10720), .ZN(n14605) );
  NAND2_X1 U13361 ( .A1(n14606), .A2(n14605), .ZN(n10725) );
  INV_X1 U13362 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10723) );
  MUX2_X1 U13363 ( .A(n10723), .B(P1_REG1_REG_3__SCAN_IN), .S(n14612), .Z(
        n10724) );
  OR2_X1 U13364 ( .A1(n14612), .A2(n10723), .ZN(n14620) );
  NAND2_X1 U13365 ( .A1(n14622), .A2(n14620), .ZN(n10728) );
  MUX2_X1 U13366 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10726), .S(n14625), .Z(
        n10727) );
  NAND2_X1 U13367 ( .A1(n10728), .A2(n10727), .ZN(n14624) );
  NAND2_X1 U13368 ( .A1(n14625), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10729) );
  MUX2_X1 U13369 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n8840), .S(n14637), .Z(
        n14644) );
  NAND2_X1 U13370 ( .A1(n14643), .A2(n14644), .ZN(n14642) );
  OR2_X1 U13371 ( .A1(n14637), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n10730) );
  AND2_X1 U13372 ( .A1(n14642), .A2(n10730), .ZN(n14655) );
  MUX2_X1 U13373 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10731), .S(n14656), .Z(
        n14654) );
  NAND2_X1 U13374 ( .A1(n14656), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n14667) );
  NAND2_X1 U13375 ( .A1(n14668), .A2(n14667), .ZN(n10734) );
  MUX2_X1 U13376 ( .A(n10732), .B(P1_REG1_REG_7__SCAN_IN), .S(n14671), .Z(
        n10733) );
  NAND2_X1 U13377 ( .A1(n10734), .A2(n10733), .ZN(n14670) );
  NAND2_X1 U13378 ( .A1(n10764), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10735) );
  NAND2_X1 U13379 ( .A1(n14670), .A2(n10735), .ZN(n10806) );
  MUX2_X1 U13380 ( .A(n10736), .B(P1_REG1_REG_8__SCAN_IN), .S(n10809), .Z(
        n10807) );
  NAND2_X1 U13381 ( .A1(n10804), .A2(n10737), .ZN(n10739) );
  NAND2_X1 U13382 ( .A1(n10739), .A2(n10738), .ZN(n10790) );
  INV_X1 U13383 ( .A(n10790), .ZN(n10740) );
  AOI21_X1 U13384 ( .B1(n10741), .B2(n10804), .A(n10740), .ZN(n10776) );
  NAND2_X1 U13385 ( .A1(n10743), .A2(n10742), .ZN(n15247) );
  INV_X1 U13386 ( .A(n15247), .ZN(n10746) );
  NAND2_X1 U13387 ( .A1(n10746), .A2(n14586), .ZN(n14714) );
  NAND2_X1 U13388 ( .A1(n10746), .A2(n15163), .ZN(n14709) );
  INV_X1 U13389 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n11322) );
  NAND2_X1 U13390 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n12207) );
  OAI21_X1 U13391 ( .B1(n14650), .B2(n11322), .A(n12207), .ZN(n10744) );
  AOI21_X1 U13392 ( .B1(n10793), .B2(n14653), .A(n10744), .ZN(n10775) );
  NOR2_X1 U13393 ( .A1(n14586), .A2(n15163), .ZN(n10745) );
  NAND2_X1 U13394 ( .A1(n10746), .A2(n10745), .ZN(n14712) );
  MUX2_X1 U13395 ( .A(n10747), .B(P1_REG2_REG_1__SCAN_IN), .S(n12477), .Z(
        n14577) );
  AND2_X1 U13396 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10748) );
  NAND2_X1 U13397 ( .A1(n14577), .A2(n10748), .ZN(n14593) );
  NAND2_X1 U13398 ( .A1(n14574), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n14592) );
  NAND2_X1 U13399 ( .A1(n14593), .A2(n14592), .ZN(n10751) );
  MUX2_X1 U13400 ( .A(n10749), .B(P1_REG2_REG_2__SCAN_IN), .S(n14596), .Z(
        n10750) );
  NAND2_X1 U13401 ( .A1(n10751), .A2(n10750), .ZN(n14610) );
  OR2_X1 U13402 ( .A1(n14596), .A2(n10749), .ZN(n14609) );
  NAND2_X1 U13403 ( .A1(n14610), .A2(n14609), .ZN(n10754) );
  MUX2_X1 U13404 ( .A(n10752), .B(P1_REG2_REG_3__SCAN_IN), .S(n14612), .Z(
        n10753) );
  NAND2_X1 U13405 ( .A1(n10754), .A2(n10753), .ZN(n14628) );
  OR2_X1 U13406 ( .A1(n14612), .A2(n10752), .ZN(n14626) );
  NAND2_X1 U13407 ( .A1(n14628), .A2(n14626), .ZN(n10756) );
  MUX2_X1 U13408 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11305), .S(n14625), .Z(
        n10755) );
  NAND2_X1 U13409 ( .A1(n14625), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14639) );
  NAND2_X1 U13410 ( .A1(n14640), .A2(n14639), .ZN(n10759) );
  MUX2_X1 U13411 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10757), .S(n14637), .Z(
        n10758) );
  NAND2_X1 U13412 ( .A1(n14637), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n14658) );
  MUX2_X1 U13413 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11456), .S(n14656), .Z(
        n10760) );
  NAND2_X1 U13414 ( .A1(n14656), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n14673) );
  MUX2_X1 U13415 ( .A(n10761), .B(P1_REG2_REG_7__SCAN_IN), .S(n14671), .Z(
        n10762) );
  NAND2_X1 U13416 ( .A1(n10763), .A2(n10762), .ZN(n14676) );
  NAND2_X1 U13417 ( .A1(n10764), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10811) );
  NAND2_X1 U13418 ( .A1(n14676), .A2(n10811), .ZN(n10767) );
  MUX2_X1 U13419 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10765), .S(n10809), .Z(
        n10766) );
  NAND2_X1 U13420 ( .A1(n10809), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10772) );
  NAND2_X1 U13421 ( .A1(n10813), .A2(n10772), .ZN(n10769) );
  MUX2_X1 U13422 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10770), .S(n10793), .Z(
        n10768) );
  INV_X1 U13423 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10770) );
  MUX2_X1 U13424 ( .A(n10770), .B(P1_REG2_REG_9__SCAN_IN), .S(n10793), .Z(
        n10771) );
  NAND3_X1 U13425 ( .A1(n10813), .A2(n10772), .A3(n10771), .ZN(n10773) );
  NAND3_X1 U13426 ( .A1(n14677), .A2(n10798), .A3(n10773), .ZN(n10774) );
  OAI211_X1 U13427 ( .C1(n10776), .C2(n14714), .A(n10775), .B(n10774), .ZN(
        P1_U3252) );
  INV_X1 U13428 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10780) );
  INV_X1 U13429 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14649) );
  NAND2_X1 U13430 ( .A1(n10778), .A2(n10777), .ZN(n10779) );
  INV_X1 U13431 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10781) );
  XNOR2_X1 U13432 ( .A(n11002), .B(n10781), .ZN(n11001) );
  INV_X1 U13433 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n15779) );
  XNOR2_X1 U13434 ( .A(n11001), .B(n15779), .ZN(n10786) );
  NAND2_X1 U13435 ( .A1(n6645), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10782) );
  INV_X1 U13436 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10784) );
  OR2_X1 U13437 ( .A1(n10793), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10787) );
  XNOR2_X1 U13438 ( .A(n10840), .B(n15716), .ZN(n10788) );
  AOI21_X1 U13439 ( .B1(n10790), .B2(n10787), .A(n10788), .ZN(n10803) );
  AND2_X1 U13440 ( .A1(n10788), .A2(n10787), .ZN(n10789) );
  NAND2_X1 U13441 ( .A1(n10790), .A2(n10789), .ZN(n10834) );
  NAND2_X1 U13442 ( .A1(n10834), .A2(n14708), .ZN(n10802) );
  AND2_X1 U13443 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n12298) );
  NOR2_X1 U13444 ( .A1(n14709), .A2(n10791), .ZN(n10792) );
  AOI211_X1 U13445 ( .C1(n15244), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n12298), 
        .B(n10792), .ZN(n10801) );
  NAND2_X1 U13446 ( .A1(n10793), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10797) );
  MUX2_X1 U13447 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10794), .S(n10840), .Z(
        n10795) );
  MUX2_X1 U13448 ( .A(n10794), .B(P1_REG2_REG_10__SCAN_IN), .S(n10840), .Z(
        n10796) );
  NAND3_X1 U13449 ( .A1(n10798), .A2(n10797), .A3(n10796), .ZN(n10799) );
  NAND3_X1 U13450 ( .A1(n14677), .A2(n10845), .A3(n10799), .ZN(n10800) );
  OAI211_X1 U13451 ( .C1(n10803), .C2(n10802), .A(n10801), .B(n10800), .ZN(
        P1_U3253) );
  INV_X1 U13452 ( .A(n10804), .ZN(n10805) );
  AOI21_X1 U13453 ( .B1(n10807), .B2(n10806), .A(n10805), .ZN(n10816) );
  AND2_X1 U13454 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11904) );
  INV_X1 U13455 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15735) );
  NOR2_X1 U13456 ( .A1(n14650), .A2(n15735), .ZN(n10808) );
  AOI211_X1 U13457 ( .C1(n14653), .C2(n10809), .A(n11904), .B(n10808), .ZN(
        n10815) );
  MUX2_X1 U13458 ( .A(n10765), .B(P1_REG2_REG_8__SCAN_IN), .S(n10809), .Z(
        n10810) );
  NAND3_X1 U13459 ( .A1(n14676), .A2(n10811), .A3(n10810), .ZN(n10812) );
  NAND3_X1 U13460 ( .A1(n14677), .A2(n10813), .A3(n10812), .ZN(n10814) );
  OAI211_X1 U13461 ( .C1(n10816), .C2(n14714), .A(n10815), .B(n10814), .ZN(
        P1_U3251) );
  INV_X1 U13462 ( .A(n11205), .ZN(n11143) );
  INV_X1 U13463 ( .A(n10817), .ZN(n10819) );
  OAI222_X1 U13464 ( .A1(n11143), .A2(P1_U3086), .B1(n12476), .B2(n10818), 
        .C1(n12474), .C2(n10819), .ZN(P1_U3342) );
  INV_X1 U13465 ( .A(n11473), .ZN(n15411) );
  OAI222_X1 U13466 ( .A1(P2_U3088), .A2(n15411), .B1(n14362), .B2(n10820), 
        .C1(n14360), .C2(n10819), .ZN(P2_U3314) );
  INV_X1 U13467 ( .A(n15466), .ZN(n15464) );
  NOR2_X1 U13468 ( .A1(n10686), .A2(n11717), .ZN(n10821) );
  OR2_X1 U13469 ( .A1(n10865), .A2(n10821), .ZN(n13847) );
  INV_X1 U13470 ( .A(n13847), .ZN(n10825) );
  NAND2_X1 U13471 ( .A1(n10685), .A2(n14162), .ZN(n10824) );
  INV_X1 U13472 ( .A(n6543), .ZN(n13639) );
  NOR2_X1 U13473 ( .A1(n13639), .A2(n14094), .ZN(n10823) );
  AOI21_X1 U13474 ( .B1(n10825), .B2(n10824), .A(n10823), .ZN(n11715) );
  INV_X1 U13475 ( .A(n10826), .ZN(n10827) );
  OAI22_X1 U13476 ( .A1(n13847), .A2(n14301), .B1(n13640), .B2(n10827), .ZN(
        n10828) );
  INV_X1 U13477 ( .A(n10828), .ZN(n10829) );
  AND2_X1 U13478 ( .A1(n11715), .A2(n10829), .ZN(n15437) );
  NAND2_X1 U13479 ( .A1(n15464), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10830) );
  OAI21_X1 U13480 ( .B1(n15464), .B2(n15437), .A(n10830), .ZN(P2_U3499) );
  INV_X1 U13481 ( .A(n11472), .ZN(n15402) );
  OAI222_X1 U13482 ( .A1(P2_U3088), .A2(n15402), .B1(n14362), .B2(n10832), 
        .C1(n14360), .C2(n10831), .ZN(P2_U3315) );
  NAND2_X1 U13483 ( .A1(n10840), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10833) );
  NAND2_X1 U13484 ( .A1(n10834), .A2(n10833), .ZN(n10838) );
  OR2_X1 U13485 ( .A1(n11020), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U13486 ( .A1(n11020), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10835) );
  NAND2_X1 U13487 ( .A1(n11028), .A2(n10835), .ZN(n10837) );
  INV_X1 U13488 ( .A(n11029), .ZN(n10836) );
  AOI21_X1 U13489 ( .B1(n10838), .B2(n10837), .A(n10836), .ZN(n10849) );
  AND2_X1 U13490 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n14504) );
  INV_X1 U13491 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15705) );
  NOR2_X1 U13492 ( .A1(n14650), .A2(n15705), .ZN(n10839) );
  AOI211_X1 U13493 ( .C1(n14653), .C2(n11020), .A(n14504), .B(n10839), .ZN(
        n10848) );
  NAND2_X1 U13494 ( .A1(n10840), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10844) );
  MUX2_X1 U13495 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11881), .S(n11020), .Z(
        n10841) );
  NAND2_X1 U13496 ( .A1(n10842), .A2(n10841), .ZN(n11022) );
  MUX2_X1 U13497 ( .A(n11881), .B(P1_REG2_REG_11__SCAN_IN), .S(n11020), .Z(
        n10843) );
  NAND3_X1 U13498 ( .A1(n10845), .A2(n10844), .A3(n10843), .ZN(n10846) );
  NAND3_X1 U13499 ( .A1(n11022), .A2(n14677), .A3(n10846), .ZN(n10847) );
  OAI211_X1 U13500 ( .C1(n10849), .C2(n14714), .A(n10848), .B(n10847), .ZN(
        P1_U3254) );
  AOI22_X1 U13501 ( .A1(n14544), .A2(n11441), .B1(n14521), .B2(n8757), .ZN(
        n10856) );
  OAI21_X1 U13502 ( .B1(n10852), .B2(n10851), .A(n10850), .ZN(n14582) );
  INV_X1 U13503 ( .A(n10853), .ZN(n11299) );
  NAND2_X1 U13504 ( .A1(n10854), .A2(n11299), .ZN(n12482) );
  AOI22_X1 U13505 ( .A1(n14515), .A2(n14582), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n12482), .ZN(n10855) );
  NAND2_X1 U13506 ( .A1(n10856), .A2(n10855), .ZN(P1_U3232) );
  INV_X1 U13507 ( .A(n10857), .ZN(n10859) );
  OAI222_X1 U13508 ( .A1(n13487), .A2(n10860), .B1(n13495), .B2(n10859), .C1(
        P3_U3151), .C2(n10858), .ZN(P3_U3281) );
  INV_X1 U13509 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15625) );
  INV_X1 U13510 ( .A(n11347), .ZN(n10861) );
  OAI21_X1 U13511 ( .B1(n15339), .B2(n15331), .A(n10861), .ZN(n10862) );
  OR2_X1 U13512 ( .A1(n9429), .A2(n14909), .ZN(n11342) );
  OAI211_X1 U13513 ( .C1(n10863), .C2(n11343), .A(n10862), .B(n11342), .ZN(
        n15101) );
  NAND2_X1 U13514 ( .A1(n15101), .A2(n15342), .ZN(n10864) );
  OAI21_X1 U13515 ( .B1(n15342), .B2(n15625), .A(n10864), .ZN(P1_U3459) );
  INV_X1 U13516 ( .A(n14301), .ZN(n15443) );
  OR2_X1 U13517 ( .A1(n6543), .A2(n10871), .ZN(n10866) );
  NOR2_X1 U13518 ( .A1(n10869), .A2(n11340), .ZN(n10870) );
  OR2_X1 U13519 ( .A1(n6728), .A2(n10870), .ZN(n11332) );
  OAI22_X1 U13520 ( .A1(n11332), .A2(n15453), .B1(n11340), .B2(n15451), .ZN(
        n10877) );
  INV_X1 U13521 ( .A(n10871), .ZN(n11068) );
  NAND2_X1 U13522 ( .A1(n10873), .A2(n10872), .ZN(n10914) );
  XNOR2_X1 U13523 ( .A(n10914), .B(n13848), .ZN(n10876) );
  INV_X1 U13524 ( .A(n10685), .ZN(n15444) );
  INV_X1 U13525 ( .A(n13905), .ZN(n13660) );
  OAI22_X1 U13526 ( .A1(n14092), .A2(n13639), .B1(n13660), .B2(n14094), .ZN(
        n10874) );
  AOI21_X1 U13527 ( .B1(n11336), .B2(n15444), .A(n10874), .ZN(n10875) );
  OAI21_X1 U13528 ( .B1(n14162), .B2(n10876), .A(n10875), .ZN(n11335) );
  AOI211_X1 U13529 ( .C1(n15443), .C2(n11336), .A(n10877), .B(n11335), .ZN(
        n10959) );
  NAND2_X1 U13530 ( .A1(n15464), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10878) );
  OAI21_X1 U13531 ( .B1(n10959), .B2(n15464), .A(n10878), .ZN(P2_U3501) );
  INV_X1 U13532 ( .A(n10879), .ZN(n10880) );
  CLKBUF_X1 U13533 ( .A(n10887), .Z(n10909) );
  INV_X1 U13534 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10881) );
  NOR2_X1 U13535 ( .A1(n10909), .A2(n10881), .ZN(P3_U3246) );
  INV_X1 U13536 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10882) );
  NOR2_X1 U13537 ( .A1(n10909), .A2(n10882), .ZN(P3_U3261) );
  INV_X1 U13538 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10883) );
  NOR2_X1 U13539 ( .A1(n10909), .A2(n10883), .ZN(P3_U3251) );
  INV_X1 U13540 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10884) );
  NOR2_X1 U13541 ( .A1(n10909), .A2(n10884), .ZN(P3_U3253) );
  INV_X1 U13542 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10885) );
  NOR2_X1 U13543 ( .A1(n10909), .A2(n10885), .ZN(P3_U3255) );
  INV_X1 U13544 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10886) );
  NOR2_X1 U13545 ( .A1(n10909), .A2(n10886), .ZN(P3_U3256) );
  INV_X1 U13546 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n15762) );
  NOR2_X1 U13547 ( .A1(n10909), .A2(n15762), .ZN(P3_U3257) );
  INV_X1 U13548 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10888) );
  NOR2_X1 U13549 ( .A1(n10909), .A2(n10888), .ZN(P3_U3245) );
  INV_X1 U13550 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10889) );
  NOR2_X1 U13551 ( .A1(n10909), .A2(n10889), .ZN(P3_U3254) );
  INV_X1 U13552 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10890) );
  NOR2_X1 U13553 ( .A1(n10887), .A2(n10890), .ZN(P3_U3242) );
  INV_X1 U13554 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10891) );
  NOR2_X1 U13555 ( .A1(n10909), .A2(n10891), .ZN(P3_U3247) );
  INV_X1 U13556 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10892) );
  NOR2_X1 U13557 ( .A1(n10909), .A2(n10892), .ZN(P3_U3248) );
  INV_X1 U13558 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10893) );
  NOR2_X1 U13559 ( .A1(n10909), .A2(n10893), .ZN(P3_U3252) );
  INV_X1 U13560 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10894) );
  NOR2_X1 U13561 ( .A1(n10909), .A2(n10894), .ZN(P3_U3250) );
  INV_X1 U13562 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10895) );
  NOR2_X1 U13563 ( .A1(n10887), .A2(n10895), .ZN(P3_U3240) );
  INV_X1 U13564 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10896) );
  NOR2_X1 U13565 ( .A1(n10887), .A2(n10896), .ZN(P3_U3239) );
  INV_X1 U13566 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10897) );
  NOR2_X1 U13567 ( .A1(n10887), .A2(n10897), .ZN(P3_U3238) );
  INV_X1 U13568 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10898) );
  NOR2_X1 U13569 ( .A1(n10887), .A2(n10898), .ZN(P3_U3237) );
  INV_X1 U13570 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10899) );
  NOR2_X1 U13571 ( .A1(n10887), .A2(n10899), .ZN(P3_U3236) );
  INV_X1 U13572 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10900) );
  NOR2_X1 U13573 ( .A1(n10909), .A2(n10900), .ZN(P3_U3259) );
  INV_X1 U13574 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10901) );
  NOR2_X1 U13575 ( .A1(n10887), .A2(n10901), .ZN(P3_U3234) );
  INV_X1 U13576 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10902) );
  NOR2_X1 U13577 ( .A1(n10887), .A2(n10902), .ZN(P3_U3258) );
  INV_X1 U13578 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10903) );
  NOR2_X1 U13579 ( .A1(n10887), .A2(n10903), .ZN(P3_U3243) );
  INV_X1 U13580 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10904) );
  NOR2_X1 U13581 ( .A1(n10887), .A2(n10904), .ZN(P3_U3260) );
  INV_X1 U13582 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n15637) );
  NOR2_X1 U13583 ( .A1(n10887), .A2(n15637), .ZN(P3_U3244) );
  INV_X1 U13584 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10905) );
  NOR2_X1 U13585 ( .A1(n10909), .A2(n10905), .ZN(P3_U3262) );
  INV_X1 U13586 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10906) );
  NOR2_X1 U13587 ( .A1(n10909), .A2(n10906), .ZN(P3_U3263) );
  INV_X1 U13588 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10907) );
  NOR2_X1 U13589 ( .A1(n10909), .A2(n10907), .ZN(P3_U3241) );
  INV_X1 U13590 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n15749) );
  NOR2_X1 U13591 ( .A1(n10909), .A2(n15749), .ZN(P3_U3235) );
  INV_X1 U13592 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10908) );
  NOR2_X1 U13593 ( .A1(n10909), .A2(n10908), .ZN(P3_U3249) );
  OR2_X1 U13594 ( .A1(n13906), .A2(n10867), .ZN(n10910) );
  XNOR2_X2 U13595 ( .A(n13662), .B(n13905), .ZN(n13845) );
  INV_X1 U13596 ( .A(n13845), .ZN(n10911) );
  NAND2_X1 U13597 ( .A1(n10912), .A2(n10911), .ZN(n10977) );
  OAI21_X1 U13598 ( .B1(n10912), .B2(n10911), .A(n10977), .ZN(n10913) );
  INV_X1 U13599 ( .A(n10913), .ZN(n11684) );
  NAND2_X1 U13600 ( .A1(n10914), .A2(n13650), .ZN(n10916) );
  INV_X1 U13601 ( .A(n13906), .ZN(n11115) );
  NAND2_X1 U13602 ( .A1(n11115), .A2(n10867), .ZN(n10915) );
  NAND2_X1 U13603 ( .A1(n10916), .A2(n10915), .ZN(n10981) );
  XNOR2_X1 U13604 ( .A(n13845), .B(n10981), .ZN(n10917) );
  AOI222_X1 U13605 ( .A1(n14180), .A2(n10917), .B1(n13904), .B2(n14108), .C1(
        n13906), .C2(n14106), .ZN(n11680) );
  OAI21_X1 U13606 ( .B1(n6728), .B2(n13659), .A(n10985), .ZN(n11678) );
  INV_X1 U13607 ( .A(n11678), .ZN(n10918) );
  AOI22_X1 U13608 ( .A1(n10918), .A2(n14308), .B1(n14315), .B2(n13662), .ZN(
        n10919) );
  OAI211_X1 U13609 ( .C1(n14319), .C2(n11684), .A(n11680), .B(n10919), .ZN(
        n11016) );
  NAND2_X1 U13610 ( .A1(n11016), .A2(n15466), .ZN(n10920) );
  OAI21_X1 U13611 ( .B1(n15466), .B2(n10600), .A(n10920), .ZN(P2_U3502) );
  INV_X1 U13612 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n15650) );
  NAND2_X1 U13613 ( .A1(P3_U3897), .A2(n11659), .ZN(n10921) );
  OAI21_X1 U13614 ( .B1(P3_U3897), .B2(n15650), .A(n10921), .ZN(P3_U3494) );
  INV_X1 U13615 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n15734) );
  NAND2_X1 U13616 ( .A1(P3_U3897), .A2(n13319), .ZN(n10922) );
  OAI21_X1 U13617 ( .B1(P3_U3897), .B2(n15734), .A(n10922), .ZN(P3_U3504) );
  OR2_X1 U13618 ( .A1(n10931), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10923) );
  INV_X1 U13619 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10925) );
  MUX2_X1 U13620 ( .A(n10925), .B(P2_REG2_REG_10__SCAN_IN), .S(n10946), .Z(
        n10926) );
  AOI21_X1 U13621 ( .B1(n10927), .B2(n10926), .A(n15414), .ZN(n10928) );
  NAND2_X1 U13622 ( .A1(n10928), .A2(n10948), .ZN(n10939) );
  NAND2_X1 U13623 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11776)
         );
  XNOR2_X1 U13624 ( .A(n10946), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n10933) );
  OR2_X1 U13625 ( .A1(n10931), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10932) );
  NAND2_X1 U13626 ( .A1(n6624), .A2(n10932), .ZN(n10934) );
  AOI21_X1 U13627 ( .B1(n10933), .B2(n10934), .A(n15420), .ZN(n10935) );
  NAND2_X1 U13628 ( .A1(n10935), .A2(n10944), .ZN(n10936) );
  NAND2_X1 U13629 ( .A1(n11776), .A2(n10936), .ZN(n10937) );
  AOI21_X1 U13630 ( .B1(n15408), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10937), 
        .ZN(n10938) );
  OAI211_X1 U13631 ( .C1(n15412), .C2(n10940), .A(n10939), .B(n10938), .ZN(
        P2_U3224) );
  INV_X1 U13632 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n15649) );
  NAND2_X1 U13633 ( .A1(n12857), .A2(P3_U3897), .ZN(n10941) );
  OAI21_X1 U13634 ( .B1(P3_U3897), .B2(n15649), .A(n10941), .ZN(P3_U3508) );
  INV_X1 U13635 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n15629) );
  NAND2_X1 U13636 ( .A1(n13305), .A2(P3_U3897), .ZN(n10942) );
  OAI21_X1 U13637 ( .B1(P3_U3897), .B2(n15629), .A(n10942), .ZN(P3_U3505) );
  NAND2_X1 U13638 ( .A1(n10946), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10943) );
  NAND2_X1 U13639 ( .A1(n10944), .A2(n10943), .ZN(n11468) );
  INV_X1 U13640 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10945) );
  XNOR2_X1 U13641 ( .A(n11469), .B(n10945), .ZN(n11467) );
  XNOR2_X1 U13642 ( .A(n11468), .B(n11467), .ZN(n10957) );
  NAND2_X1 U13643 ( .A1(n10946), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10947) );
  INV_X1 U13644 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10949) );
  MUX2_X1 U13645 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10949), .S(n11469), .Z(
        n10950) );
  NAND2_X1 U13646 ( .A1(n10951), .A2(n10950), .ZN(n15391) );
  OAI21_X1 U13647 ( .B1(n10951), .B2(n10950), .A(n15391), .ZN(n10955) );
  NAND2_X1 U13648 ( .A1(n15408), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n10952) );
  NAND2_X1 U13649 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12010)
         );
  OAI211_X1 U13650 ( .C1(n15412), .C2(n10953), .A(n10952), .B(n12010), .ZN(
        n10954) );
  AOI21_X1 U13651 ( .B1(n10955), .B2(n15394), .A(n10954), .ZN(n10956) );
  OAI21_X1 U13652 ( .B1(n10957), .B2(n15420), .A(n10956), .ZN(P2_U3225) );
  INV_X2 U13653 ( .A(n15460), .ZN(n15462) );
  INV_X1 U13654 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10961) );
  OR2_X1 U13655 ( .A1(n10959), .A2(n15460), .ZN(n10960) );
  OAI21_X1 U13656 ( .B1(n15462), .B2(n10961), .A(n10960), .ZN(P2_U3436) );
  NOR2_X1 U13657 ( .A1(n10962), .A2(P2_U3088), .ZN(n11074) );
  INV_X1 U13658 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11714) );
  NAND2_X1 U13659 ( .A1(n9652), .A2(n10686), .ZN(n10963) );
  AOI21_X1 U13660 ( .B1(n13627), .B2(n10963), .A(n13623), .ZN(n10966) );
  INV_X1 U13661 ( .A(n10963), .ZN(n10964) );
  NAND2_X1 U13662 ( .A1(n13627), .A2(n10964), .ZN(n10965) );
  MUX2_X1 U13663 ( .A(n10966), .B(n10965), .S(n13640), .Z(n10968) );
  INV_X1 U13664 ( .A(n13621), .ZN(n13537) );
  NAND2_X1 U13665 ( .A1(n13537), .A2(n6543), .ZN(n10967) );
  OAI211_X1 U13666 ( .C1(n11074), .C2(n11714), .A(n10968), .B(n10967), .ZN(
        P2_U3204) );
  INV_X1 U13667 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10971) );
  NAND2_X1 U13668 ( .A1(n15462), .A2(n10969), .ZN(n10970) );
  OAI21_X1 U13669 ( .B1(n15462), .B2(n10971), .A(n10970), .ZN(P2_U3433) );
  INV_X1 U13670 ( .A(n10972), .ZN(n10975) );
  AOI222_X1 U13671 ( .A1(n13035), .A2(P3_STATE_REG_SCAN_IN), .B1(n10975), .B2(
        n13480), .C1(n10974), .C2(n10973), .ZN(P3_U3280) );
  INV_X1 U13672 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10990) );
  OR2_X1 U13673 ( .A1(n13905), .A2(n13662), .ZN(n10976) );
  XNOR2_X1 U13674 ( .A(n13670), .B(n13904), .ZN(n13853) );
  INV_X1 U13675 ( .A(n13853), .ZN(n10978) );
  NAND2_X1 U13676 ( .A1(n10979), .A2(n10978), .ZN(n11050) );
  OAI21_X1 U13677 ( .B1(n10979), .B2(n10978), .A(n11050), .ZN(n10980) );
  INV_X1 U13678 ( .A(n10980), .ZN(n11677) );
  NAND2_X1 U13679 ( .A1(n10981), .A2(n13845), .ZN(n10983) );
  NAND2_X1 U13680 ( .A1(n13660), .A2(n13662), .ZN(n10982) );
  NAND2_X1 U13681 ( .A1(n10983), .A2(n10982), .ZN(n11051) );
  XNOR2_X1 U13682 ( .A(n11051), .B(n13853), .ZN(n10984) );
  OAI22_X1 U13683 ( .A1(n14092), .A2(n13660), .B1(n13675), .B2(n14094), .ZN(
        n11010) );
  AOI21_X1 U13684 ( .B1(n10984), .B2(n14180), .A(n11010), .ZN(n11673) );
  INV_X1 U13685 ( .A(n10985), .ZN(n10986) );
  OAI211_X1 U13686 ( .C1(n10986), .C2(n7575), .A(n14308), .B(n11056), .ZN(
        n11671) );
  INV_X1 U13687 ( .A(n11671), .ZN(n10987) );
  AOI21_X1 U13688 ( .B1(n14315), .B2(n13670), .A(n10987), .ZN(n10988) );
  OAI211_X1 U13689 ( .C1(n11677), .C2(n14319), .A(n11673), .B(n10988), .ZN(
        n14320) );
  NAND2_X1 U13690 ( .A1(n14320), .A2(n15462), .ZN(n10989) );
  OAI21_X1 U13691 ( .B1(n15462), .B2(n10990), .A(n10989), .ZN(P2_U3442) );
  INV_X1 U13692 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11331) );
  NAND2_X1 U13693 ( .A1(n13550), .A2(n14106), .ZN(n13618) );
  OAI22_X1 U13694 ( .A1(n11074), .A2(n11331), .B1(n13618), .B2(n13639), .ZN(
        n10998) );
  OAI22_X1 U13695 ( .A1(n13621), .A2(n13660), .B1(n13637), .B2(n11340), .ZN(
        n10997) );
  INV_X1 U13696 ( .A(n10991), .ZN(n10993) );
  NAND3_X1 U13697 ( .A1(n11065), .A2(n10993), .A3(n10992), .ZN(n10994) );
  AOI21_X1 U13698 ( .B1(n10995), .B2(n10994), .A(n13625), .ZN(n10996) );
  OR3_X1 U13699 ( .A1(n10998), .A2(n10997), .A3(n10996), .ZN(P2_U3209) );
  NAND2_X1 U13700 ( .A1(n10999), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n11000) );
  NAND2_X1 U13701 ( .A1(n11001), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n11004) );
  XNOR2_X1 U13702 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n11318) );
  XNOR2_X1 U13703 ( .A(n11319), .B(n11318), .ZN(n11313) );
  INV_X1 U13704 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n11311) );
  XNOR2_X1 U13705 ( .A(n11312), .B(n11311), .ZN(SUB_1596_U55) );
  INV_X1 U13706 ( .A(n12196), .ZN(n11966) );
  INV_X1 U13707 ( .A(n11005), .ZN(n11064) );
  OAI222_X1 U13708 ( .A1(P1_U3086), .A2(n11966), .B1(n12474), .B2(n11064), 
        .C1(n15681), .C2(n15161), .ZN(P1_U3339) );
  INV_X1 U13709 ( .A(n11006), .ZN(n11009) );
  NAND2_X1 U13710 ( .A1(n11109), .A2(n11007), .ZN(n11008) );
  NOR2_X1 U13711 ( .A1(n11008), .A2(n11009), .ZN(n11084) );
  AOI21_X1 U13712 ( .B1(n11009), .B2(n11008), .A(n11084), .ZN(n11014) );
  AOI22_X1 U13713 ( .A1(n13550), .A2(n11010), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11011) );
  OAI21_X1 U13714 ( .B1(n7575), .B2(n13637), .A(n11011), .ZN(n11012) );
  AOI21_X1 U13715 ( .B1(n11669), .B2(n13634), .A(n11012), .ZN(n11013) );
  OAI21_X1 U13716 ( .B1(n11014), .B2(n13625), .A(n11013), .ZN(P2_U3202) );
  INV_X1 U13717 ( .A(n11015), .ZN(n11078) );
  INV_X1 U13718 ( .A(n14685), .ZN(n12204) );
  OAI222_X1 U13719 ( .A1(n12476), .A2(n15783), .B1(n12474), .B2(n11078), .C1(
        P1_U3086), .C2(n12204), .ZN(P1_U3338) );
  INV_X1 U13720 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11018) );
  NAND2_X1 U13721 ( .A1(n11016), .A2(n15462), .ZN(n11017) );
  OAI21_X1 U13722 ( .B1(n15462), .B2(n11018), .A(n11017), .ZN(P2_U3439) );
  MUX2_X1 U13723 ( .A(n11019), .B(P1_REG2_REG_12__SCAN_IN), .S(n11133), .Z(
        n11025) );
  NAND2_X1 U13724 ( .A1(n11020), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11021) );
  INV_X1 U13725 ( .A(n11135), .ZN(n11023) );
  AOI21_X1 U13726 ( .B1(n11025), .B2(n11024), .A(n11023), .ZN(n11035) );
  INV_X1 U13727 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11026) );
  NOR2_X1 U13728 ( .A1(n11026), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14414) );
  INV_X1 U13729 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n12359) );
  NOR2_X1 U13730 ( .A1(n14650), .A2(n12359), .ZN(n11027) );
  AOI211_X1 U13731 ( .C1(n14653), .C2(n11133), .A(n14414), .B(n11027), .ZN(
        n11034) );
  XNOR2_X1 U13732 ( .A(n11133), .B(n15084), .ZN(n11031) );
  NAND2_X1 U13733 ( .A1(n11030), .A2(n11031), .ZN(n11130) );
  OAI21_X1 U13734 ( .B1(n11031), .B2(n11030), .A(n11130), .ZN(n11032) );
  NAND2_X1 U13735 ( .A1(n11032), .A2(n14708), .ZN(n11033) );
  OAI211_X1 U13736 ( .C1(n11035), .C2(n14712), .A(n11034), .B(n11033), .ZN(
        P1_U3255) );
  OAI21_X1 U13737 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n11036), .A(n11095), .ZN(
        n11041) );
  INV_X1 U13738 ( .A(n11099), .ZN(n11037) );
  AOI21_X1 U13739 ( .B1(n15480), .B2(n6733), .A(n11037), .ZN(n11039) );
  INV_X1 U13740 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15768) );
  NOR2_X1 U13741 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15768), .ZN(n12816) );
  AOI21_X1 U13742 ( .B1(n15467), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n12816), .ZN(
        n11038) );
  OAI21_X1 U13743 ( .B1(n13077), .B2(n11039), .A(n11038), .ZN(n11040) );
  AOI21_X1 U13744 ( .B1(n13100), .B2(n11041), .A(n11040), .ZN(n11047) );
  AND3_X1 U13745 ( .A1(n11152), .A2(n11043), .A3(n11042), .ZN(n11044) );
  OAI21_X1 U13746 ( .B1(n11045), .B2(n11044), .A(n13095), .ZN(n11046) );
  OAI211_X1 U13747 ( .C1(n13088), .C2(n11048), .A(n11047), .B(n11046), .ZN(
        P3_U3185) );
  OR2_X1 U13748 ( .A1(n13670), .A2(n13904), .ZN(n11049) );
  NAND2_X1 U13749 ( .A1(n11050), .A2(n11049), .ZN(n11616) );
  XNOR2_X2 U13750 ( .A(n13676), .B(n13903), .ZN(n13852) );
  XNOR2_X1 U13751 ( .A(n11616), .B(n13852), .ZN(n11693) );
  INV_X1 U13752 ( .A(n13904), .ZN(n11053) );
  NAND2_X1 U13753 ( .A1(n13670), .A2(n11053), .ZN(n11052) );
  XNOR2_X1 U13754 ( .A(n11621), .B(n13852), .ZN(n11054) );
  INV_X1 U13755 ( .A(n13902), .ZN(n11623) );
  OAI22_X1 U13756 ( .A1(n14092), .A2(n11053), .B1(n11623), .B2(n14094), .ZN(
        n11088) );
  AOI21_X1 U13757 ( .B1(n11054), .B2(n14180), .A(n11088), .ZN(n11689) );
  INV_X1 U13758 ( .A(n11706), .ZN(n11055) );
  AOI21_X1 U13759 ( .B1(n13676), .B2(n11056), .A(n11055), .ZN(n11685) );
  AOI22_X1 U13760 ( .A1(n11685), .A2(n14308), .B1(n14315), .B2(n13676), .ZN(
        n11057) );
  OAI211_X1 U13761 ( .C1(n11693), .C2(n14319), .A(n11689), .B(n11057), .ZN(
        n11061) );
  NAND2_X1 U13762 ( .A1(n11061), .A2(n15466), .ZN(n11058) );
  OAI21_X1 U13763 ( .B1(n15466), .B2(n10605), .A(n11058), .ZN(P2_U3504) );
  INV_X1 U13764 ( .A(n11805), .ZN(n11203) );
  OAI222_X1 U13765 ( .A1(P1_U3086), .A2(n11203), .B1(n12474), .B2(n11059), 
        .C1(n11060), .C2(n15161), .ZN(P1_U3341) );
  INV_X1 U13766 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11063) );
  NAND2_X1 U13767 ( .A1(n11061), .A2(n15462), .ZN(n11062) );
  OAI21_X1 U13768 ( .B1(n15462), .B2(n11063), .A(n11062), .ZN(P2_U3445) );
  INV_X1 U13769 ( .A(n12141), .ZN(n12248) );
  OAI222_X1 U13770 ( .A1(P2_U3088), .A2(n12248), .B1(n14362), .B2(n15748), 
        .C1(n14360), .C2(n11064), .ZN(P2_U3311) );
  OAI21_X1 U13771 ( .B1(n11067), .B2(n11066), .A(n11065), .ZN(n11070) );
  OAI22_X1 U13772 ( .A1(n13621), .A2(n11115), .B1(n13637), .B2(n11068), .ZN(
        n11069) );
  AOI21_X1 U13773 ( .B1(n13627), .B2(n11070), .A(n11069), .ZN(n11072) );
  INV_X1 U13774 ( .A(n13618), .ZN(n13605) );
  NAND2_X1 U13775 ( .A1(n13605), .A2(n10686), .ZN(n11071) );
  OAI211_X1 U13776 ( .C1(n11074), .C2(n11073), .A(n11072), .B(n11071), .ZN(
        P2_U3194) );
  INV_X1 U13777 ( .A(n11075), .ZN(n11076) );
  OAI222_X1 U13778 ( .A1(n13487), .A2(n11077), .B1(n13061), .B2(P3_U3151), 
        .C1(n13495), .C2(n11076), .ZN(P3_U3279) );
  INV_X1 U13779 ( .A(n12410), .ZN(n11079) );
  OAI222_X1 U13780 ( .A1(P2_U3088), .A2(n11079), .B1(n14362), .B2(n15707), 
        .C1(n14360), .C2(n11078), .ZN(P2_U3310) );
  INV_X1 U13781 ( .A(n11977), .ZN(n11981) );
  OAI222_X1 U13782 ( .A1(P2_U3088), .A2(n11981), .B1(n14362), .B2(n11080), 
        .C1(n14360), .C2(n11059), .ZN(P2_U3313) );
  INV_X1 U13783 ( .A(n11081), .ZN(n11686) );
  NOR3_X1 U13784 ( .A1(n11084), .A2(n11083), .A3(n11082), .ZN(n11085) );
  OAI21_X1 U13785 ( .B1(n11085), .B2(n6727), .A(n13627), .ZN(n11090) );
  INV_X1 U13786 ( .A(n13676), .ZN(n13674) );
  NOR2_X1 U13787 ( .A1(n13637), .A2(n13674), .ZN(n11086) );
  AOI211_X1 U13788 ( .C1(n13550), .C2(n11088), .A(n11087), .B(n11086), .ZN(
        n11089) );
  OAI211_X1 U13789 ( .C1(n13599), .C2(n11686), .A(n11090), .B(n11089), .ZN(
        P2_U3199) );
  AOI21_X1 U13790 ( .B1(n11092), .B2(n11091), .A(n6723), .ZN(n11108) );
  INV_X1 U13791 ( .A(n13088), .ZN(n13014) );
  AND3_X1 U13792 ( .A1(n11095), .A2(n11094), .A3(n11093), .ZN(n11096) );
  OAI21_X1 U13793 ( .B1(n11097), .B2(n11096), .A(n13100), .ZN(n11104) );
  AND3_X1 U13794 ( .A1(n11099), .A2(n11098), .A3(n7970), .ZN(n11100) );
  OAI21_X1 U13795 ( .B1(n11101), .B2(n11100), .A(n13090), .ZN(n11103) );
  INV_X1 U13796 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15798) );
  NOR2_X1 U13797 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15798), .ZN(n11435) );
  AOI21_X1 U13798 ( .B1(n15467), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11435), .ZN(
        n11102) );
  NAND3_X1 U13799 ( .A1(n11104), .A2(n11103), .A3(n11102), .ZN(n11105) );
  AOI21_X1 U13800 ( .B1(n11106), .B2(n13014), .A(n11105), .ZN(n11107) );
  OAI21_X1 U13801 ( .B1(n11108), .B2(n13030), .A(n11107), .ZN(P3_U3186) );
  INV_X1 U13802 ( .A(n11109), .ZN(n11110) );
  AOI211_X1 U13803 ( .C1(n11112), .C2(n11111), .A(n13625), .B(n11110), .ZN(
        n11117) );
  AOI22_X1 U13804 ( .A1(n13537), .A2(n13904), .B1(n13662), .B2(n13623), .ZN(
        n11114) );
  MUX2_X1 U13805 ( .A(n13599), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n11113) );
  OAI211_X1 U13806 ( .C1(n11115), .C2(n13618), .A(n11114), .B(n11113), .ZN(
        n11116) );
  OR2_X1 U13807 ( .A1(n11117), .A2(n11116), .ZN(P2_U3190) );
  INV_X1 U13808 ( .A(n11118), .ZN(n11709) );
  OAI211_X1 U13809 ( .C1(n11121), .C2(n11120), .A(n11119), .B(n13627), .ZN(
        n11124) );
  AOI22_X1 U13810 ( .A1(n13901), .A2(n14108), .B1(n14106), .B2(n13903), .ZN(
        n11702) );
  OAI22_X1 U13811 ( .A1(n13632), .A2(n11702), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15374), .ZN(n11122) );
  AOI21_X1 U13812 ( .B1(n15438), .B2(n13623), .A(n11122), .ZN(n11123) );
  OAI211_X1 U13813 ( .C1(n13599), .C2(n11709), .A(n11124), .B(n11123), .ZN(
        P2_U3211) );
  INV_X1 U13814 ( .A(SI_17_), .ZN(n11127) );
  INV_X1 U13815 ( .A(n11125), .ZN(n11126) );
  OAI222_X1 U13816 ( .A1(n13487), .A2(n11127), .B1(n13073), .B2(P3_U3151), 
        .C1(n13495), .C2(n11126), .ZN(P3_U3278) );
  OR2_X1 U13817 ( .A1(n11133), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11128) );
  AND2_X1 U13818 ( .A1(n11130), .A2(n11128), .ZN(n11132) );
  XNOR2_X1 U13819 ( .A(n11205), .B(n15079), .ZN(n11131) );
  AND2_X1 U13820 ( .A1(n11131), .A2(n11128), .ZN(n11129) );
  NAND2_X1 U13821 ( .A1(n11130), .A2(n11129), .ZN(n11199) );
  OAI211_X1 U13822 ( .C1(n11132), .C2(n11131), .A(n14708), .B(n11199), .ZN(
        n11142) );
  NAND2_X1 U13823 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14484)
         );
  MUX2_X1 U13824 ( .A(n14986), .B(P1_REG2_REG_13__SCAN_IN), .S(n11205), .Z(
        n11136) );
  OR2_X1 U13825 ( .A1(n11133), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11134) );
  AOI21_X1 U13826 ( .B1(n11136), .B2(n11137), .A(n14712), .ZN(n11138) );
  NAND2_X1 U13827 ( .A1(n11138), .A2(n11210), .ZN(n11139) );
  NAND2_X1 U13828 ( .A1(n14484), .A2(n11139), .ZN(n11140) );
  AOI21_X1 U13829 ( .B1(n15244), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11140), 
        .ZN(n11141) );
  OAI211_X1 U13830 ( .C1(n14709), .C2(n11143), .A(n11142), .B(n11141), .ZN(
        P1_U3256) );
  AOI21_X1 U13831 ( .B1(n11146), .B2(n11145), .A(n11144), .ZN(n11148) );
  AOI22_X1 U13832 ( .A1(n15467), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n11147) );
  OAI21_X1 U13833 ( .B1(n13077), .B2(n11148), .A(n11147), .ZN(n11160) );
  AOI21_X1 U13834 ( .B1(n11151), .B2(n11150), .A(n11149), .ZN(n11158) );
  INV_X1 U13835 ( .A(n11152), .ZN(n11156) );
  NOR3_X1 U13836 ( .A1(n11183), .A2(n11154), .A3(n11153), .ZN(n11155) );
  OAI21_X1 U13837 ( .B1(n11156), .B2(n11155), .A(n13095), .ZN(n11157) );
  OAI21_X1 U13838 ( .B1(n13046), .B2(n11158), .A(n11157), .ZN(n11159) );
  AOI211_X1 U13839 ( .C1(n11161), .C2(n13014), .A(n11160), .B(n11159), .ZN(
        n11162) );
  INV_X1 U13840 ( .A(n11162), .ZN(P3_U3184) );
  OAI222_X1 U13841 ( .A1(n13495), .A2(n11164), .B1(n12613), .B2(P3_U3151), 
        .C1(n11163), .C2(n13487), .ZN(P3_U3276) );
  OAI211_X1 U13842 ( .C1(n11167), .C2(n11166), .A(n11165), .B(n13627), .ZN(
        n11172) );
  INV_X1 U13843 ( .A(n11731), .ZN(n11170) );
  INV_X1 U13844 ( .A(n13687), .ZN(n15452) );
  OAI22_X1 U13845 ( .A1(n13637), .A2(n15452), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15585), .ZN(n11169) );
  OAI22_X1 U13846 ( .A1(n13692), .A2(n13621), .B1(n13618), .B2(n11623), .ZN(
        n11168) );
  AOI211_X1 U13847 ( .C1(n11170), .C2(n13634), .A(n11169), .B(n11168), .ZN(
        n11171) );
  NAND2_X1 U13848 ( .A1(n11172), .A2(n11171), .ZN(P2_U3185) );
  INV_X1 U13849 ( .A(n11173), .ZN(n11174) );
  OAI222_X1 U13850 ( .A1(n13487), .A2(n15667), .B1(n13087), .B2(P3_U3151), 
        .C1(n13495), .C2(n11174), .ZN(P3_U3277) );
  INV_X1 U13851 ( .A(n12136), .ZN(n11985) );
  INV_X1 U13852 ( .A(n11175), .ZN(n11177) );
  INV_X1 U13853 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11176) );
  OAI222_X1 U13854 ( .A1(n11985), .A2(P2_U3088), .B1(n14360), .B2(n11177), 
        .C1(n11176), .C2(n14362), .ZN(P2_U3312) );
  INV_X1 U13855 ( .A(n11812), .ZN(n11955) );
  OAI222_X1 U13856 ( .A1(n12476), .A2(n11178), .B1(n12474), .B2(n11177), .C1(
        n11955), .C2(P1_U3086), .ZN(P1_U3340) );
  AND2_X1 U13857 ( .A1(n15505), .A2(n11483), .ZN(n12626) );
  INV_X1 U13858 ( .A(n12626), .ZN(n12628) );
  AND2_X1 U13859 ( .A1(n15502), .A2(n12628), .ZN(n12598) );
  NOR3_X1 U13860 ( .A1(n12598), .A2(n13374), .A3(n11179), .ZN(n11180) );
  AOI21_X1 U13861 ( .B1(n13320), .B2(n12974), .A(n11180), .ZN(n11538) );
  MUX2_X1 U13862 ( .A(n11538), .B(n11181), .S(n15546), .Z(n11182) );
  OAI21_X1 U13863 ( .B1(n11483), .B2(n13391), .A(n11182), .ZN(P3_U3459) );
  AOI21_X1 U13864 ( .B1(n11185), .B2(n11184), .A(n11183), .ZN(n11186) );
  OAI22_X1 U13865 ( .A1(n13030), .A2(n11186), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11284), .ZN(n11195) );
  AOI21_X1 U13866 ( .B1(n11189), .B2(n11188), .A(n11187), .ZN(n11193) );
  AOI21_X1 U13867 ( .B1(n15541), .B2(n11191), .A(n11190), .ZN(n11192) );
  OAI22_X1 U13868 ( .A1(n11193), .A2(n13077), .B1(n13046), .B2(n11192), .ZN(
        n11194) );
  AOI211_X1 U13869 ( .C1(P3_ADDR_REG_1__SCAN_IN), .C2(n15467), .A(n11195), .B(
        n11194), .ZN(n11196) );
  OAI21_X1 U13870 ( .B1(n11197), .B2(n13088), .A(n11196), .ZN(P3_U3183) );
  XNOR2_X1 U13871 ( .A(n11805), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n11202) );
  NAND2_X1 U13872 ( .A1(n11205), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11198) );
  NAND2_X1 U13873 ( .A1(n11199), .A2(n11198), .ZN(n11201) );
  INV_X1 U13874 ( .A(n11804), .ZN(n11200) );
  AOI21_X1 U13875 ( .B1(n11202), .B2(n11201), .A(n11200), .ZN(n11214) );
  AND2_X1 U13876 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14379) );
  NOR2_X1 U13877 ( .A1(n14709), .A2(n11203), .ZN(n11204) );
  AOI211_X1 U13878 ( .C1(n15244), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n14379), 
        .B(n11204), .ZN(n11213) );
  NAND2_X1 U13879 ( .A1(n11205), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11209) );
  NAND2_X1 U13880 ( .A1(n11210), .A2(n11209), .ZN(n11207) );
  MUX2_X1 U13881 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n14969), .S(n11805), .Z(
        n11206) );
  NAND2_X1 U13882 ( .A1(n11207), .A2(n11206), .ZN(n11807) );
  MUX2_X1 U13883 ( .A(n14969), .B(P1_REG2_REG_14__SCAN_IN), .S(n11805), .Z(
        n11208) );
  NAND3_X1 U13884 ( .A1(n11210), .A2(n11209), .A3(n11208), .ZN(n11211) );
  NAND3_X1 U13885 ( .A1(n11807), .A2(n14677), .A3(n11211), .ZN(n11212) );
  OAI211_X1 U13886 ( .C1(n11214), .C2(n14714), .A(n11213), .B(n11212), .ZN(
        P1_U3257) );
  OAI21_X1 U13887 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n11216), .A(n11375), .ZN(
        n11222) );
  INV_X1 U13888 ( .A(n11217), .ZN(n11218) );
  AOI21_X1 U13889 ( .B1(n15795), .B2(n6719), .A(n11218), .ZN(n11220) );
  AND2_X1 U13890 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n12867) );
  AOI21_X1 U13891 ( .B1(n15467), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n12867), .ZN(
        n11219) );
  OAI21_X1 U13892 ( .B1(n11220), .B2(n13077), .A(n11219), .ZN(n11221) );
  AOI21_X1 U13893 ( .B1(n13100), .B2(n11222), .A(n11221), .ZN(n11231) );
  INV_X1 U13894 ( .A(n11223), .ZN(n11228) );
  OAI21_X1 U13895 ( .B1(n11227), .B2(n11225), .A(n11224), .ZN(n11226) );
  OAI21_X1 U13896 ( .B1(n11228), .B2(n11227), .A(n11226), .ZN(n11229) );
  NAND2_X1 U13897 ( .A1(n11229), .A2(n13095), .ZN(n11230) );
  OAI211_X1 U13898 ( .C1(n13088), .C2(n6911), .A(n11231), .B(n11230), .ZN(
        P3_U3187) );
  NAND2_X1 U13899 ( .A1(n11247), .A2(n11244), .ZN(n11238) );
  NOR2_X1 U13900 ( .A1(n11532), .A2(n11232), .ZN(n11237) );
  INV_X1 U13901 ( .A(n11233), .ZN(n11234) );
  OR2_X1 U13902 ( .A1(n11249), .A2(n11234), .ZN(n11236) );
  NAND4_X1 U13903 ( .A1(n11238), .A2(n11237), .A3(n11236), .A4(n11235), .ZN(
        n11239) );
  NAND2_X1 U13904 ( .A1(n11239), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11242) );
  INV_X1 U13905 ( .A(n12764), .ZN(n11240) );
  OR2_X1 U13906 ( .A1(n11249), .A2(n11240), .ZN(n11241) );
  NOR2_X1 U13907 ( .A1(n12952), .A2(P3_U3151), .ZN(n11285) );
  AND2_X1 U13908 ( .A1(n11249), .A2(n12764), .ZN(n11255) );
  NAND2_X1 U13909 ( .A1(n11247), .A2(n15514), .ZN(n11243) );
  NAND3_X1 U13910 ( .A1(n11245), .A2(n15512), .A3(n11244), .ZN(n11246) );
  NAND2_X1 U13911 ( .A1(n11249), .A2(n11248), .ZN(n11250) );
  OAI22_X1 U13912 ( .A1(n12926), .A2(n11483), .B1(n12960), .B2(n12598), .ZN(
        n11252) );
  AOI21_X1 U13913 ( .B1(n12933), .B2(n12974), .A(n11252), .ZN(n11253) );
  OAI21_X1 U13914 ( .B1(n11285), .B2(n11254), .A(n11253), .ZN(P3_U3172) );
  INV_X1 U13915 ( .A(n12974), .ZN(n15493) );
  INV_X1 U13916 ( .A(n11255), .ZN(n11257) );
  OAI22_X1 U13917 ( .A1(n12926), .A2(n15497), .B1(n15493), .B2(n12922), .ZN(
        n11258) );
  AOI21_X1 U13918 ( .B1(n12933), .B2(n11659), .A(n11258), .ZN(n11273) );
  INV_X1 U13919 ( .A(n12615), .ZN(n11259) );
  OAI21_X1 U13920 ( .B1(n11763), .B2(n12613), .A(n11385), .ZN(n11260) );
  XNOR2_X1 U13921 ( .A(n11421), .B(n11262), .ZN(n11422) );
  INV_X1 U13922 ( .A(n11279), .ZN(n15503) );
  OAI21_X1 U13923 ( .B1(n11421), .B2(n15503), .A(n11263), .ZN(n11266) );
  NAND2_X1 U13924 ( .A1(n11421), .A2(n12624), .ZN(n11264) );
  NAND2_X1 U13925 ( .A1(n11266), .A2(n11280), .ZN(n11278) );
  XNOR2_X1 U13926 ( .A(n11421), .B(n11267), .ZN(n11268) );
  NAND2_X1 U13927 ( .A1(n11268), .A2(n15493), .ZN(n11269) );
  NAND2_X1 U13928 ( .A1(n11278), .A2(n11269), .ZN(n11270) );
  NAND2_X1 U13929 ( .A1(n11271), .A2(n7163), .ZN(n11272) );
  OAI211_X1 U13930 ( .C1(n11285), .C2(n11274), .A(n11273), .B(n11272), .ZN(
        P3_U3177) );
  OAI22_X1 U13931 ( .A1(n12926), .A2(n15513), .B1(n6869), .B2(n12922), .ZN(
        n11275) );
  AOI21_X1 U13932 ( .B1(n12933), .B2(n15506), .A(n11275), .ZN(n11283) );
  INV_X2 U13933 ( .A(n12462), .ZN(n12447) );
  NAND3_X1 U13934 ( .A1(n12447), .A2(n15502), .A3(n11276), .ZN(n11277) );
  OAI211_X1 U13935 ( .C1(n11280), .C2(n11279), .A(n11278), .B(n11277), .ZN(
        n11281) );
  NAND2_X1 U13936 ( .A1(n11281), .A2(n7163), .ZN(n11282) );
  OAI211_X1 U13937 ( .C1(n11285), .C2(n11284), .A(n11283), .B(n11282), .ZN(
        P3_U3162) );
  OR2_X1 U13938 ( .A1(n13100), .A2(n13095), .ZN(n11289) );
  INV_X1 U13939 ( .A(n11288), .ZN(n11286) );
  NAND2_X1 U13940 ( .A1(n11289), .A2(n11286), .ZN(n11287) );
  OAI21_X1 U13941 ( .B1(n13077), .B2(n11539), .A(n11287), .ZN(n11292) );
  OAI21_X1 U13942 ( .B1(n11289), .B2(n13090), .A(n11288), .ZN(n11290) );
  NAND2_X1 U13943 ( .A1(n11290), .A2(n13088), .ZN(n11291) );
  MUX2_X1 U13944 ( .A(n11292), .B(n11291), .S(P3_IR_REG_0__SCAN_IN), .Z(n11295) );
  INV_X1 U13945 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n11293) );
  OAI22_X1 U13946 ( .A1(n13007), .A2(n11293), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11254), .ZN(n11294) );
  OR2_X1 U13947 ( .A1(n11295), .A2(n11294), .ZN(P3_U3182) );
  NAND4_X1 U13948 ( .A1(n11299), .A2(n11298), .A3(n11297), .A4(n11296), .ZN(
        n12487) );
  AND2_X1 U13949 ( .A1(n11940), .A2(n11349), .ZN(n11300) );
  XNOR2_X1 U13950 ( .A(n11301), .B(n11303), .ZN(n15321) );
  XNOR2_X1 U13951 ( .A(n11302), .B(n11303), .ZN(n11304) );
  AOI222_X1 U13952 ( .A1(n15331), .A2(n11304), .B1(n14567), .B2(n14940), .C1(
        n14569), .C2(n14939), .ZN(n15325) );
  MUX2_X1 U13953 ( .A(n11305), .B(n15325), .S(n14987), .Z(n11310) );
  OR2_X2 U13954 ( .A1(n6538), .A2(n11306), .ZN(n15283) );
  NOR2_X1 U13955 ( .A1(n15265), .A2(n15323), .ZN(n14727) );
  INV_X1 U13956 ( .A(n14727), .ZN(n11993) );
  NAND2_X1 U13957 ( .A1(n15286), .A2(n14464), .ZN(n11307) );
  NAND2_X1 U13958 ( .A1(n11592), .A2(n11307), .ZN(n15324) );
  OAI22_X1 U13959 ( .A1(n11993), .A2(n15324), .B1(n14465), .B2(n15280), .ZN(
        n11308) );
  AOI21_X1 U13960 ( .B1(n14752), .B2(n14464), .A(n11308), .ZN(n11309) );
  OAI211_X1 U13961 ( .C1(n14953), .C2(n15321), .A(n11310), .B(n11309), .ZN(
        P1_U3289) );
  NAND2_X1 U13962 ( .A1(n11312), .A2(n11311), .ZN(n11317) );
  INV_X1 U13963 ( .A(n11313), .ZN(n11314) );
  OR2_X1 U13964 ( .A1(n11315), .A2(n11314), .ZN(n11316) );
  INV_X1 U13965 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11830) );
  NAND2_X1 U13966 ( .A1(n11830), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n11320) );
  NAND2_X1 U13967 ( .A1(n11322), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11559) );
  INV_X1 U13968 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n11323) );
  NAND2_X1 U13969 ( .A1(n11323), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U13970 ( .A1(n11559), .A2(n11324), .ZN(n11557) );
  XNOR2_X1 U13971 ( .A(n11558), .B(n11557), .ZN(n11553) );
  NAND4_X1 U13972 ( .A1(n11326), .A2(n15432), .A3(n11325), .A4(n15431), .ZN(
        n11330) );
  INV_X1 U13973 ( .A(n11330), .ZN(n11328) );
  NAND2_X1 U13974 ( .A1(n11328), .A2(n11327), .ZN(n11667) );
  NOR2_X1 U13975 ( .A1(n11330), .A2(n9652), .ZN(n14122) );
  INV_X1 U13976 ( .A(n14122), .ZN(n14052) );
  OAI22_X1 U13977 ( .A1(n14052), .A2(n11332), .B1(n11331), .B2(n14146), .ZN(
        n11333) );
  AOI21_X1 U13978 ( .B1(n14186), .B2(P2_REG2_REG_2__SCAN_IN), .A(n11333), .ZN(
        n11339) );
  NAND2_X1 U13979 ( .A1(n13643), .A2(n9912), .ZN(n11501) );
  INV_X1 U13980 ( .A(n11501), .ZN(n11334) );
  NAND2_X1 U13981 ( .A1(n14135), .A2(n11334), .ZN(n12047) );
  INV_X1 U13982 ( .A(n12047), .ZN(n11337) );
  AOI22_X1 U13983 ( .A1(n11337), .A2(n11336), .B1(n14135), .B2(n11335), .ZN(
        n11338) );
  OAI211_X1 U13984 ( .C1(n11340), .C2(n14188), .A(n11339), .B(n11338), .ZN(
        P2_U3263) );
  NOR2_X1 U13985 ( .A1(n14905), .A2(n14990), .ZN(n11348) );
  OAI22_X1 U13986 ( .A1(n6538), .A2(n11342), .B1(n11341), .B2(n15280), .ZN(
        n11345) );
  AOI21_X1 U13987 ( .B1(n11993), .B2(n15283), .A(n11343), .ZN(n11344) );
  AOI211_X1 U13988 ( .C1(n6538), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11345), .B(
        n11344), .ZN(n11346) );
  OAI21_X1 U13989 ( .B1(n11348), .B2(n11347), .A(n11346), .ZN(P1_U3293) );
  INV_X1 U13990 ( .A(n11349), .ZN(n11350) );
  NAND2_X1 U13991 ( .A1(n14987), .A2(n11350), .ZN(n15285) );
  OAI21_X1 U13992 ( .B1(n6538), .B2(n11940), .A(n15285), .ZN(n14789) );
  INV_X1 U13993 ( .A(n14789), .ZN(n14897) );
  XNOR2_X1 U13994 ( .A(n11351), .B(n11360), .ZN(n15311) );
  NAND2_X1 U13995 ( .A1(n14940), .A2(n14569), .ZN(n11353) );
  OR2_X1 U13996 ( .A1(n9429), .A2(n14907), .ZN(n11352) );
  NAND2_X1 U13997 ( .A1(n11353), .A2(n11352), .ZN(n15303) );
  INV_X1 U13998 ( .A(n11443), .ZN(n11355) );
  INV_X1 U13999 ( .A(n15287), .ZN(n11354) );
  OAI211_X1 U14000 ( .C1(n15306), .C2(n11355), .A(n11354), .B(n10110), .ZN(
        n15305) );
  OAI22_X1 U14001 ( .A1(n15265), .A2(n15305), .B1(n11356), .B2(n15280), .ZN(
        n11358) );
  NOR2_X1 U14002 ( .A1(n14987), .A2(n10749), .ZN(n11357) );
  AOI211_X1 U14003 ( .C1(n14987), .C2(n15303), .A(n11358), .B(n11357), .ZN(
        n11364) );
  OAI21_X1 U14004 ( .B1(n11361), .B2(n11360), .A(n11359), .ZN(n15308) );
  AOI22_X1 U14005 ( .A1(n14905), .A2(n15308), .B1(n14752), .B2(n11362), .ZN(
        n11363) );
  OAI211_X1 U14006 ( .C1(n14897), .C2(n15311), .A(n11364), .B(n11363), .ZN(
        P1_U3291) );
  AOI21_X1 U14007 ( .B1(n11367), .B2(n11366), .A(n11365), .ZN(n11382) );
  AND2_X1 U14008 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n12931) );
  INV_X1 U14009 ( .A(n11368), .ZN(n11371) );
  NAND3_X1 U14010 ( .A1(n11217), .A2(n11369), .A3(n6910), .ZN(n11370) );
  AOI21_X1 U14011 ( .B1(n11371), .B2(n11370), .A(n13077), .ZN(n11372) );
  AOI211_X1 U14012 ( .C1(n15467), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n12931), .B(
        n11372), .ZN(n11381) );
  INV_X1 U14013 ( .A(n11373), .ZN(n11377) );
  NAND3_X1 U14014 ( .A1(n11375), .A2(n11374), .A3(n7908), .ZN(n11376) );
  AOI21_X1 U14015 ( .B1(n11377), .B2(n11376), .A(n13046), .ZN(n11378) );
  AOI21_X1 U14016 ( .B1(n13014), .B2(n11379), .A(n11378), .ZN(n11380) );
  OAI211_X1 U14017 ( .C1(n11382), .C2(n13030), .A(n11381), .B(n11380), .ZN(
        P3_U3188) );
  INV_X1 U14018 ( .A(n11383), .ZN(n11386) );
  OAI222_X1 U14019 ( .A1(n13495), .A2(n11386), .B1(n11385), .B2(P3_U3151), 
        .C1(n11384), .C2(n13487), .ZN(P3_U3275) );
  INV_X1 U14020 ( .A(n11394), .ZN(n11388) );
  AND2_X1 U14021 ( .A1(n11387), .A2(n11388), .ZN(n11485) );
  INV_X1 U14022 ( .A(n11485), .ZN(n11391) );
  INV_X1 U14023 ( .A(n11387), .ZN(n11389) );
  NAND2_X1 U14024 ( .A1(n11389), .A2(n11394), .ZN(n11390) );
  NAND2_X1 U14025 ( .A1(n11391), .A2(n11390), .ZN(n11392) );
  INV_X1 U14026 ( .A(n11392), .ZN(n11462) );
  NAND2_X1 U14027 ( .A1(n11392), .A2(n10368), .ZN(n11400) );
  OAI21_X1 U14028 ( .B1(n11395), .B2(n11394), .A(n11393), .ZN(n11398) );
  OAI22_X1 U14029 ( .A1(n11396), .A2(n14907), .B1(n11491), .B2(n14909), .ZN(
        n11397) );
  AOI21_X1 U14030 ( .B1(n11398), .B2(n15331), .A(n11397), .ZN(n11399) );
  AND2_X1 U14031 ( .A1(n11400), .A2(n11399), .ZN(n11455) );
  AOI211_X1 U14032 ( .C1(n11605), .C2(n11593), .A(n15323), .B(n11944), .ZN(
        n11459) );
  INV_X1 U14033 ( .A(n11459), .ZN(n11401) );
  OAI211_X1 U14034 ( .C1(n11462), .C2(n15310), .A(n11455), .B(n11401), .ZN(
        n11406) );
  OAI22_X1 U14035 ( .A1(n15086), .A2(n11457), .B1(n15348), .B2(n10731), .ZN(
        n11402) );
  AOI21_X1 U14036 ( .B1(n11406), .B2(n15348), .A(n11402), .ZN(n11403) );
  INV_X1 U14037 ( .A(n11403), .ZN(P1_U3534) );
  INV_X1 U14038 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11404) );
  OAI22_X1 U14039 ( .A1(n15147), .A2(n11457), .B1(n15342), .B2(n11404), .ZN(
        n11405) );
  AOI21_X1 U14040 ( .B1(n11406), .B2(n15342), .A(n11405), .ZN(n11407) );
  INV_X1 U14041 ( .A(n11407), .ZN(P1_U3477) );
  NAND2_X1 U14042 ( .A1(n11409), .A2(n11408), .ZN(n11411) );
  XOR2_X1 U14043 ( .A(n11411), .B(n11410), .Z(n11417) );
  INV_X1 U14044 ( .A(n11746), .ZN(n11415) );
  OAI21_X1 U14045 ( .B1(n13637), .B2(n6833), .A(n11412), .ZN(n11414) );
  OAI22_X1 U14046 ( .A1(n11736), .A2(n13618), .B1(n13621), .B2(n11788), .ZN(
        n11413) );
  AOI211_X1 U14047 ( .C1(n11415), .C2(n13634), .A(n11414), .B(n11413), .ZN(
        n11416) );
  OAI21_X1 U14048 ( .B1(n11417), .B2(n13625), .A(n11416), .ZN(P2_U3193) );
  INV_X1 U14049 ( .A(n12413), .ZN(n13928) );
  INV_X1 U14050 ( .A(n11418), .ZN(n11420) );
  OAI222_X1 U14051 ( .A1(n13928), .A2(P2_U3088), .B1(n14360), .B2(n11420), 
        .C1(n11419), .C2(n14362), .ZN(P2_U3309) );
  INV_X1 U14052 ( .A(n14703), .ZN(n14691) );
  OAI222_X1 U14053 ( .A1(n12476), .A2(n15666), .B1(n12474), .B2(n11420), .C1(
        n14691), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U14054 ( .A(n15506), .ZN(n11649) );
  NAND2_X1 U14055 ( .A1(n11422), .A2(n11649), .ZN(n12811) );
  INV_X1 U14056 ( .A(n11423), .ZN(n11424) );
  NAND2_X1 U14057 ( .A1(n11424), .A2(n11659), .ZN(n11425) );
  NAND2_X1 U14058 ( .A1(n12813), .A2(n11425), .ZN(n11433) );
  XNOR2_X1 U14059 ( .A(n11421), .B(n11436), .ZN(n11426) );
  INV_X1 U14060 ( .A(n12973), .ZN(n11648) );
  NAND2_X1 U14061 ( .A1(n11426), .A2(n11648), .ZN(n12214) );
  INV_X1 U14062 ( .A(n11426), .ZN(n11427) );
  NAND2_X1 U14063 ( .A1(n11427), .A2(n12973), .ZN(n11428) );
  NAND2_X1 U14064 ( .A1(n12214), .A2(n11428), .ZN(n11432) );
  INV_X1 U14065 ( .A(n11433), .ZN(n11430) );
  NAND2_X1 U14066 ( .A1(n11430), .A2(n11429), .ZN(n12215) );
  INV_X1 U14067 ( .A(n12215), .ZN(n11431) );
  AOI21_X1 U14068 ( .B1(n11433), .B2(n11432), .A(n11431), .ZN(n11440) );
  INV_X1 U14069 ( .A(n12933), .ZN(n12956) );
  INV_X1 U14070 ( .A(n12972), .ZN(n12217) );
  OAI22_X1 U14071 ( .A1(n12956), .A2(n12217), .B1(n7381), .B2(n12922), .ZN(
        n11434) );
  AOI211_X1 U14072 ( .C1(n12958), .C2(n11436), .A(n11435), .B(n11434), .ZN(
        n11439) );
  INV_X1 U14073 ( .A(n15470), .ZN(n11437) );
  NAND2_X1 U14074 ( .A1(n12952), .A2(n11437), .ZN(n11438) );
  OAI211_X1 U14075 ( .C1(n11440), .C2(n12960), .A(n11439), .B(n11438), .ZN(
        P3_U3170) );
  NAND2_X1 U14076 ( .A1(n11441), .A2(n15294), .ZN(n11442) );
  NAND2_X1 U14077 ( .A1(n11443), .A2(n11442), .ZN(n15298) );
  XNOR2_X1 U14078 ( .A(n11444), .B(n11445), .ZN(n15302) );
  AOI22_X1 U14079 ( .A1(n14990), .A2(n15302), .B1(n14752), .B2(n15294), .ZN(
        n11447) );
  INV_X1 U14080 ( .A(n15280), .ZN(n14945) );
  NAND2_X1 U14081 ( .A1(n14945), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n11446) );
  OAI211_X1 U14082 ( .C1(n15298), .C2(n11993), .A(n11447), .B(n11446), .ZN(
        n11454) );
  OAI21_X1 U14083 ( .B1(n11444), .B2(n8742), .A(n15331), .ZN(n11448) );
  NAND2_X1 U14084 ( .A1(n11448), .A2(n14907), .ZN(n11451) );
  XNOR2_X1 U14085 ( .A(n15298), .B(n9429), .ZN(n11449) );
  OAI21_X1 U14086 ( .B1(n11449), .B2(n15276), .A(n8742), .ZN(n11450) );
  NAND2_X1 U14087 ( .A1(n11451), .A2(n11450), .ZN(n15299) );
  NAND2_X1 U14088 ( .A1(n14940), .A2(n9433), .ZN(n15296) );
  NAND2_X1 U14089 ( .A1(n15299), .A2(n15296), .ZN(n11452) );
  MUX2_X1 U14090 ( .A(n11452), .B(P1_REG2_REG_1__SCAN_IN), .S(n6538), .Z(
        n11453) );
  OR2_X1 U14091 ( .A1(n11454), .A2(n11453), .ZN(P1_U3292) );
  MUX2_X1 U14092 ( .A(n11456), .B(n11455), .S(n14987), .Z(n11461) );
  OAI22_X1 U14093 ( .A1(n15283), .A2(n11457), .B1(n15280), .B2(n11608), .ZN(
        n11458) );
  AOI21_X1 U14094 ( .B1(n11459), .B2(n15289), .A(n11458), .ZN(n11460) );
  OAI211_X1 U14095 ( .C1(n11462), .C2(n15285), .A(n11461), .B(n11460), .ZN(
        P1_U3287) );
  OR2_X1 U14096 ( .A1(n11469), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n15389) );
  NAND2_X1 U14097 ( .A1(n15391), .A2(n15389), .ZN(n11463) );
  INV_X1 U14098 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11464) );
  MUX2_X1 U14099 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11464), .S(n11472), .Z(
        n15388) );
  NAND2_X1 U14100 ( .A1(n11463), .A2(n15388), .ZN(n15393) );
  NAND2_X1 U14101 ( .A1(n15402), .A2(n11464), .ZN(n11465) );
  MUX2_X1 U14102 ( .A(n9818), .B(P2_REG2_REG_13__SCAN_IN), .S(n11473), .Z(
        n15415) );
  NAND2_X1 U14103 ( .A1(n11473), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11466) );
  NAND2_X1 U14104 ( .A1(n15417), .A2(n11466), .ZN(n11978) );
  XNOR2_X1 U14105 ( .A(n11976), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n11478) );
  XNOR2_X1 U14106 ( .A(n11977), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11982) );
  NAND2_X1 U14107 ( .A1(n11468), .A2(n11467), .ZN(n11471) );
  NAND2_X1 U14108 ( .A1(n11469), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11470) );
  NAND2_X1 U14109 ( .A1(n11471), .A2(n11470), .ZN(n15397) );
  XNOR2_X1 U14110 ( .A(n11472), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n15396) );
  XNOR2_X1 U14111 ( .A(n11473), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n15422) );
  NOR2_X1 U14112 ( .A1(n15421), .A2(n15422), .ZN(n15419) );
  XOR2_X1 U14113 ( .A(n11982), .B(n11983), .Z(n11476) );
  NAND2_X1 U14114 ( .A1(n15408), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n11474) );
  NAND2_X1 U14115 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n13508)
         );
  OAI211_X1 U14116 ( .C1(n15412), .C2(n11981), .A(n11474), .B(n13508), .ZN(
        n11475) );
  AOI21_X1 U14117 ( .B1(n11476), .B2(n15398), .A(n11475), .ZN(n11477) );
  OAI21_X1 U14118 ( .B1(n11478), .B2(n15414), .A(n11477), .ZN(P2_U3228) );
  INV_X1 U14119 ( .A(n11479), .ZN(n11481) );
  OAI222_X1 U14120 ( .A1(n13495), .A2(n11481), .B1(n12627), .B2(P3_U3151), 
        .C1(n11480), .C2(n13487), .ZN(P3_U3274) );
  MUX2_X1 U14121 ( .A(n11538), .B(n8065), .S(n15539), .Z(n11482) );
  OAI21_X1 U14122 ( .B1(n13470), .B2(n11483), .A(n11482), .ZN(P3_U3390) );
  NOR2_X1 U14123 ( .A1(n11485), .A2(n11484), .ZN(n11937) );
  NOR2_X1 U14124 ( .A1(n11937), .A2(n11939), .ZN(n11936) );
  INV_X1 U14125 ( .A(n11936), .ZN(n11487) );
  NAND2_X1 U14126 ( .A1(n11487), .A2(n11486), .ZN(n11488) );
  XNOR2_X1 U14127 ( .A(n11488), .B(n11497), .ZN(n15340) );
  INV_X1 U14128 ( .A(n15340), .ZN(n11500) );
  INV_X1 U14129 ( .A(n11489), .ZN(n11490) );
  OAI211_X1 U14130 ( .C1(n11490), .C2(n15336), .A(n10110), .B(n11857), .ZN(
        n15334) );
  INV_X1 U14131 ( .A(n15334), .ZN(n11494) );
  OAI22_X1 U14132 ( .A1(n11491), .A2(n14907), .B1(n11522), .B2(n14909), .ZN(
        n15332) );
  MUX2_X1 U14133 ( .A(n15332), .B(P1_REG2_REG_8__SCAN_IN), .S(n6538), .Z(
        n11493) );
  OAI22_X1 U14134 ( .A1(n15283), .A2(n15336), .B1(n15280), .B2(n11902), .ZN(
        n11492) );
  AOI211_X1 U14135 ( .C1(n11494), .C2(n15289), .A(n11493), .B(n11492), .ZN(
        n11499) );
  NAND2_X1 U14136 ( .A1(n11496), .A2(n11497), .ZN(n15330) );
  NAND3_X1 U14137 ( .A1(n11495), .A2(n15330), .A3(n14905), .ZN(n11498) );
  OAI211_X1 U14138 ( .C1(n11500), .C2(n14953), .A(n11499), .B(n11498), .ZN(
        P1_U3285) );
  NAND2_X1 U14139 ( .A1(n10685), .A2(n11501), .ZN(n11502) );
  OAI22_X1 U14140 ( .A1(n11068), .A2(n14188), .B1(n14191), .B2(n11503), .ZN(
        n11510) );
  INV_X1 U14141 ( .A(n14146), .ZN(n14184) );
  AOI22_X1 U14142 ( .A1(n14122), .A2(n11504), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n14184), .ZN(n11507) );
  NAND2_X1 U14143 ( .A1(n14135), .A2(n11505), .ZN(n11506) );
  OAI211_X1 U14144 ( .C1(n11508), .C2(n14135), .A(n11507), .B(n11506), .ZN(
        n11509) );
  OR2_X1 U14145 ( .A1(n11510), .A2(n11509), .ZN(P2_U3264) );
  INV_X1 U14146 ( .A(n11511), .ZN(n11655) );
  INV_X1 U14147 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11512) );
  OAI222_X1 U14148 ( .A1(P2_U3088), .A2(n14152), .B1(n14360), .B2(n11655), 
        .C1(n11512), .C2(n14362), .ZN(P2_U3308) );
  OAI21_X1 U14149 ( .B1(n11514), .B2(n11517), .A(n11513), .ZN(n11515) );
  INV_X1 U14150 ( .A(n11515), .ZN(n15099) );
  NAND2_X1 U14151 ( .A1(n11518), .A2(n11517), .ZN(n15093) );
  NAND3_X1 U14152 ( .A1(n11516), .A2(n15093), .A3(n14905), .ZN(n11527) );
  OAI21_X1 U14153 ( .B1(n11858), .B2(n12301), .A(n10110), .ZN(n11519) );
  OR2_X1 U14154 ( .A1(n11880), .A2(n11519), .ZN(n11521) );
  NAND2_X1 U14155 ( .A1(n14940), .A2(n14561), .ZN(n11520) );
  NAND2_X1 U14156 ( .A1(n11521), .A2(n11520), .ZN(n15094) );
  NOR2_X1 U14157 ( .A1(n11522), .A2(n14907), .ZN(n15095) );
  OAI22_X1 U14158 ( .A1(n14987), .A2(n10794), .B1(n12296), .B2(n15280), .ZN(
        n11523) );
  AOI21_X1 U14159 ( .B1(n15095), .B2(n14987), .A(n11523), .ZN(n11524) );
  OAI21_X1 U14160 ( .B1(n12301), .B2(n15283), .A(n11524), .ZN(n11525) );
  AOI21_X1 U14161 ( .B1(n15094), .B2(n15289), .A(n11525), .ZN(n11526) );
  OAI211_X1 U14162 ( .C1(n15099), .C2(n14953), .A(n11527), .B(n11526), .ZN(
        P1_U3283) );
  NAND2_X1 U14163 ( .A1(n11528), .A2(n11530), .ZN(n11529) );
  OAI21_X1 U14164 ( .B1(n13471), .B2(n11530), .A(n11529), .ZN(n11535) );
  INV_X1 U14165 ( .A(n11531), .ZN(n11534) );
  INV_X1 U14166 ( .A(n11532), .ZN(n11533) );
  NAND3_X1 U14167 ( .A1(n11535), .A2(n11534), .A3(n11533), .ZN(n11537) );
  AOI22_X1 U14168 ( .A1(n6529), .A2(n6872), .B1(n15516), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n11541) );
  MUX2_X1 U14169 ( .A(n11539), .B(n11538), .S(n15500), .Z(n11540) );
  NAND2_X1 U14170 ( .A1(n11541), .A2(n11540), .ZN(P3_U3233) );
  INV_X1 U14171 ( .A(n11542), .ZN(n12381) );
  OAI222_X1 U14172 ( .A1(n11544), .A2(P1_U3086), .B1(n12474), .B2(n12381), 
        .C1(n11543), .C2(n15161), .ZN(P1_U3335) );
  OAI211_X1 U14173 ( .C1(n11547), .C2(n11546), .A(n11545), .B(n14515), .ZN(
        n11551) );
  OAI22_X1 U14174 ( .A1(n11548), .A2(n14907), .B1(n11861), .B2(n14909), .ZN(
        n11942) );
  AND2_X1 U14175 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14665) );
  NOR2_X1 U14176 ( .A1(n14528), .A2(n15248), .ZN(n11549) );
  AOI211_X1 U14177 ( .C1(n14497), .C2(n11942), .A(n14665), .B(n11549), .ZN(
        n11550) );
  OAI211_X1 U14178 ( .C1(n15251), .C2(n14524), .A(n11551), .B(n11550), .ZN(
        P1_U3213) );
  INV_X1 U14179 ( .A(n11552), .ZN(n11554) );
  NAND2_X1 U14180 ( .A1(n11554), .A2(n11553), .ZN(n11555) );
  INV_X1 U14181 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n11561) );
  XNOR2_X1 U14182 ( .A(n11561), .B(P3_ADDR_REG_10__SCAN_IN), .ZN(n11562) );
  NAND2_X1 U14183 ( .A1(n11563), .A2(n11562), .ZN(n11564) );
  NAND2_X1 U14184 ( .A1(n11910), .A2(n11911), .ZN(n11565) );
  XNOR2_X1 U14185 ( .A(n11565), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  INV_X1 U14186 ( .A(n11566), .ZN(n11567) );
  XNOR2_X1 U14187 ( .A(n6700), .B(n11566), .ZN(n14463) );
  NAND2_X1 U14188 ( .A1(n14463), .A2(n14462), .ZN(n14461) );
  OAI21_X1 U14189 ( .B1(n6700), .B2(n11567), .A(n14461), .ZN(n11571) );
  XNOR2_X1 U14190 ( .A(n11569), .B(n11568), .ZN(n11570) );
  XNOR2_X1 U14191 ( .A(n11571), .B(n11570), .ZN(n11578) );
  NAND2_X1 U14192 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n14634) );
  NAND2_X1 U14193 ( .A1(n14939), .A2(n14568), .ZN(n11573) );
  NAND2_X1 U14194 ( .A1(n14940), .A2(n14566), .ZN(n11572) );
  NAND2_X1 U14195 ( .A1(n11573), .A2(n11572), .ZN(n11590) );
  NAND2_X1 U14196 ( .A1(n14497), .A2(n11590), .ZN(n11574) );
  OAI211_X1 U14197 ( .C1(n14528), .C2(n15259), .A(n14634), .B(n11574), .ZN(
        n11575) );
  AOI21_X1 U14198 ( .B1(n11576), .B2(n14544), .A(n11575), .ZN(n11577) );
  OAI21_X1 U14199 ( .B1(n11578), .B2(n14546), .A(n11577), .ZN(P1_U3227) );
  INV_X1 U14200 ( .A(n11579), .ZN(n11581) );
  OAI22_X1 U14201 ( .A1(n12766), .A2(P3_U3151), .B1(SI_22_), .B2(n13487), .ZN(
        n11580) );
  AOI21_X1 U14202 ( .B1(n11581), .B2(n13480), .A(n11580), .ZN(P3_U3273) );
  INV_X1 U14203 ( .A(n11582), .ZN(n11583) );
  AOI21_X1 U14204 ( .B1(n11587), .B2(n11584), .A(n11583), .ZN(n15266) );
  NAND2_X1 U14205 ( .A1(n11586), .A2(n11585), .ZN(n11588) );
  XNOR2_X1 U14206 ( .A(n11588), .B(n11587), .ZN(n11591) );
  NOR2_X1 U14207 ( .A1(n15266), .A2(n11940), .ZN(n11589) );
  AOI211_X1 U14208 ( .C1(n15331), .C2(n11591), .A(n11590), .B(n11589), .ZN(
        n15270) );
  INV_X1 U14209 ( .A(n11592), .ZN(n11594) );
  OAI211_X1 U14210 ( .C1(n11594), .C2(n15262), .A(n10110), .B(n11593), .ZN(
        n15264) );
  OAI211_X1 U14211 ( .C1(n15266), .C2(n15310), .A(n15270), .B(n15264), .ZN(
        n11599) );
  OAI22_X1 U14212 ( .A1(n15086), .A2(n15262), .B1(n15348), .B2(n8840), .ZN(
        n11595) );
  AOI21_X1 U14213 ( .B1(n11599), .B2(n15348), .A(n11595), .ZN(n11596) );
  INV_X1 U14214 ( .A(n11596), .ZN(P1_U3533) );
  INV_X1 U14215 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n11597) );
  OAI22_X1 U14216 ( .A1(n15147), .A2(n15262), .B1(n15342), .B2(n11597), .ZN(
        n11598) );
  AOI21_X1 U14217 ( .B1(n11599), .B2(n15342), .A(n11598), .ZN(n11600) );
  INV_X1 U14218 ( .A(n11600), .ZN(P1_U3474) );
  INV_X1 U14219 ( .A(n11601), .ZN(n11602) );
  AOI211_X1 U14220 ( .C1(n11604), .C2(n11603), .A(n14546), .B(n11602), .ZN(
        n11610) );
  AOI22_X1 U14221 ( .A1(n14544), .A2(n11605), .B1(n14538), .B2(n14567), .ZN(
        n11607) );
  NOR2_X1 U14222 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8849), .ZN(n14652) );
  AOI21_X1 U14223 ( .B1(n14521), .B2(n14565), .A(n14652), .ZN(n11606) );
  OAI211_X1 U14224 ( .C1(n11608), .C2(n14528), .A(n11607), .B(n11606), .ZN(
        n11609) );
  OR2_X1 U14225 ( .A1(n11610), .A2(n11609), .ZN(P1_U3239) );
  OAI22_X1 U14226 ( .A1(n15438), .A2(n13902), .B1(n13676), .B2(n13903), .ZN(
        n11615) );
  NAND2_X1 U14227 ( .A1(n13676), .A2(n13903), .ZN(n11611) );
  NAND2_X1 U14228 ( .A1(n11611), .A2(n11623), .ZN(n11613) );
  AND2_X1 U14229 ( .A1(n13903), .A2(n13902), .ZN(n11612) );
  AOI22_X1 U14230 ( .A1(n11613), .A2(n15438), .B1(n11612), .B2(n13676), .ZN(
        n11614) );
  NAND2_X1 U14231 ( .A1(n11617), .A2(n11723), .ZN(n11620) );
  AND2_X1 U14232 ( .A1(n13687), .A2(n13901), .ZN(n11618) );
  AOI22_X1 U14233 ( .A1(n11738), .A2(n11618), .B1(n14314), .B2(n6832), .ZN(
        n11619) );
  XNOR2_X1 U14234 ( .A(n14307), .B(n11788), .ZN(n13856) );
  XNOR2_X1 U14235 ( .A(n11782), .B(n13856), .ZN(n14312) );
  NAND2_X1 U14236 ( .A1(n13676), .A2(n13675), .ZN(n11622) );
  XNOR2_X1 U14237 ( .A(n15438), .B(n13902), .ZN(n13680) );
  NAND2_X1 U14238 ( .A1(n13687), .A2(n11736), .ZN(n11724) );
  INV_X1 U14239 ( .A(n11738), .ZN(n13854) );
  NAND2_X1 U14240 ( .A1(n11786), .A2(n13854), .ZN(n11740) );
  NAND2_X1 U14241 ( .A1(n11740), .A2(n11789), .ZN(n11624) );
  XOR2_X1 U14242 ( .A(n13856), .B(n11624), .Z(n11625) );
  AOI222_X1 U14243 ( .A1(n14180), .A2(n11625), .B1(n13899), .B2(n14108), .C1(
        n6832), .C2(n14106), .ZN(n14311) );
  MUX2_X1 U14244 ( .A(n11626), .B(n14311), .S(n14135), .Z(n11630) );
  AOI21_X1 U14245 ( .B1(n14307), .B2(n11743), .A(n11795), .ZN(n14309) );
  INV_X1 U14246 ( .A(n14307), .ZN(n11627) );
  OAI22_X1 U14247 ( .A1(n14188), .A2(n11627), .B1(n11755), .B2(n14146), .ZN(
        n11628) );
  AOI21_X1 U14248 ( .B1(n14309), .B2(n14122), .A(n11628), .ZN(n11629) );
  OAI211_X1 U14249 ( .C1(n14312), .C2(n14191), .A(n11630), .B(n11629), .ZN(
        P2_U3256) );
  XOR2_X1 U14250 ( .A(n11632), .B(n11631), .Z(n11642) );
  INV_X1 U14251 ( .A(n11833), .ZN(n11633) );
  OAI21_X1 U14252 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n6726), .A(n11633), .ZN(
        n11640) );
  AOI21_X1 U14253 ( .B1(n15571), .B2(n11634), .A(n11840), .ZN(n11635) );
  NOR2_X1 U14254 ( .A1(n11635), .A2(n13046), .ZN(n11639) );
  INV_X1 U14255 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11636) );
  NOR2_X1 U14256 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11636), .ZN(n12776) );
  AOI21_X1 U14257 ( .B1(n15467), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12776), .ZN(
        n11637) );
  OAI21_X1 U14258 ( .B1(n13088), .B2(n6938), .A(n11637), .ZN(n11638) );
  AOI211_X1 U14259 ( .C1(n11640), .C2(n13090), .A(n11639), .B(n11638), .ZN(
        n11641) );
  OAI21_X1 U14260 ( .B1(n11642), .B2(n13030), .A(n11641), .ZN(P3_U3189) );
  NAND2_X1 U14261 ( .A1(n15490), .A2(n15489), .ZN(n15488) );
  NAND2_X1 U14262 ( .A1(n15488), .A2(n11644), .ZN(n11646) );
  XNOR2_X1 U14263 ( .A(n11646), .B(n12595), .ZN(n15478) );
  AOI211_X1 U14264 ( .C1(n12595), .C2(n11647), .A(n15508), .B(n6696), .ZN(
        n11651) );
  OAI22_X1 U14265 ( .A1(n11649), .A2(n15492), .B1(n11648), .B2(n15491), .ZN(
        n11650) );
  OR2_X1 U14266 ( .A1(n11651), .A2(n11650), .ZN(n15476) );
  AOI21_X1 U14267 ( .B1(n15478), .B2(n15537), .A(n15476), .ZN(n11666) );
  MUX2_X1 U14268 ( .A(n11652), .B(n11666), .S(n15549), .Z(n11653) );
  OAI21_X1 U14269 ( .B1(n13391), .B2(n15482), .A(n11653), .ZN(P3_U3462) );
  OAI222_X1 U14270 ( .A1(P1_U3086), .A2(n8984), .B1(n12474), .B2(n11655), .C1(
        n11654), .C2(n15161), .ZN(P1_U3336) );
  OAI21_X1 U14271 ( .B1(n11656), .B2(n12641), .A(n11762), .ZN(n15469) );
  NOR2_X1 U14272 ( .A1(n6696), .A2(n11657), .ZN(n11658) );
  XNOR2_X1 U14273 ( .A(n11658), .B(n12641), .ZN(n11661) );
  AOI22_X1 U14274 ( .A1(n13320), .A2(n12972), .B1(n11659), .B2(n15504), .ZN(
        n11660) );
  OAI21_X1 U14275 ( .B1(n11661), .B2(n15508), .A(n11660), .ZN(n15468) );
  AOI21_X1 U14276 ( .B1(n15537), .B2(n15469), .A(n15468), .ZN(n11720) );
  OAI22_X1 U14277 ( .A1(n13470), .A2(n15472), .B1(n8102), .B2(n15540), .ZN(
        n11662) );
  INV_X1 U14278 ( .A(n11662), .ZN(n11663) );
  OAI21_X1 U14279 ( .B1(n11720), .B2(n15539), .A(n11663), .ZN(P3_U3402) );
  OAI22_X1 U14280 ( .A1(n13470), .A2(n15482), .B1(n8088), .B2(n15540), .ZN(
        n11664) );
  INV_X1 U14281 ( .A(n11664), .ZN(n11665) );
  OAI21_X1 U14282 ( .B1(n11666), .B2(n15539), .A(n11665), .ZN(P3_U3399) );
  INV_X1 U14283 ( .A(n11667), .ZN(n11668) );
  INV_X1 U14284 ( .A(n14194), .ZN(n14173) );
  INV_X1 U14285 ( .A(n11669), .ZN(n11670) );
  OAI22_X1 U14286 ( .A1(n14173), .A2(n11671), .B1(n11670), .B2(n14146), .ZN(
        n11672) );
  AOI21_X1 U14287 ( .B1(n14169), .B2(n13670), .A(n11672), .ZN(n11676) );
  MUX2_X1 U14288 ( .A(n11674), .B(n11673), .S(n14135), .Z(n11675) );
  OAI211_X1 U14289 ( .C1(n14191), .C2(n11677), .A(n11676), .B(n11675), .ZN(
        P2_U3261) );
  OAI22_X1 U14290 ( .A1(n14052), .A2(n11678), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14146), .ZN(n11679) );
  AOI21_X1 U14291 ( .B1(n14169), .B2(n13662), .A(n11679), .ZN(n11683) );
  MUX2_X1 U14292 ( .A(n11681), .B(n11680), .S(n14135), .Z(n11682) );
  OAI211_X1 U14293 ( .C1(n11684), .C2(n14191), .A(n11683), .B(n11682), .ZN(
        P2_U3262) );
  INV_X1 U14294 ( .A(n11685), .ZN(n11687) );
  OAI22_X1 U14295 ( .A1(n14052), .A2(n11687), .B1(n11686), .B2(n14146), .ZN(
        n11688) );
  AOI21_X1 U14296 ( .B1(n14169), .B2(n13676), .A(n11688), .ZN(n11692) );
  MUX2_X1 U14297 ( .A(n11690), .B(n11689), .S(n14135), .Z(n11691) );
  OAI211_X1 U14298 ( .C1(n14191), .C2(n11693), .A(n11692), .B(n11691), .ZN(
        P2_U3260) );
  INV_X1 U14299 ( .A(n11694), .ZN(n12383) );
  INV_X1 U14300 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11695) );
  OAI222_X1 U14301 ( .A1(P2_U3088), .A2(n11696), .B1(n14360), .B2(n12383), 
        .C1(n11695), .C2(n14362), .ZN(P2_U3306) );
  OAI21_X1 U14302 ( .B1(n11616), .B2(n13675), .A(n13674), .ZN(n11698) );
  NAND2_X1 U14303 ( .A1(n11616), .A2(n13675), .ZN(n11697) );
  NAND2_X1 U14304 ( .A1(n11698), .A2(n11697), .ZN(n11699) );
  INV_X1 U14305 ( .A(n13680), .ZN(n13850) );
  XNOR2_X1 U14306 ( .A(n11699), .B(n13850), .ZN(n15445) );
  INV_X1 U14307 ( .A(n15445), .ZN(n11713) );
  XNOR2_X1 U14308 ( .A(n11700), .B(n13680), .ZN(n11701) );
  NAND2_X1 U14309 ( .A1(n11701), .A2(n14180), .ZN(n11703) );
  NAND2_X1 U14310 ( .A1(n11703), .A2(n11702), .ZN(n15442) );
  INV_X1 U14311 ( .A(n15442), .ZN(n11704) );
  MUX2_X1 U14312 ( .A(n11705), .B(n11704), .S(n14135), .Z(n11712) );
  INV_X1 U14313 ( .A(n11730), .ZN(n11708) );
  AOI21_X1 U14314 ( .B1(n11706), .B2(n15438), .A(n15453), .ZN(n11707) );
  NAND2_X1 U14315 ( .A1(n11708), .A2(n11707), .ZN(n15439) );
  OAI22_X1 U14316 ( .A1(n14173), .A2(n15439), .B1(n11709), .B2(n14146), .ZN(
        n11710) );
  AOI21_X1 U14317 ( .B1(n14169), .B2(n15438), .A(n11710), .ZN(n11711) );
  OAI211_X1 U14318 ( .C1(n14191), .C2(n11713), .A(n11712), .B(n11711), .ZN(
        P2_U3259) );
  OAI22_X1 U14319 ( .A1(n14186), .A2(n11715), .B1(n11714), .B2(n14146), .ZN(
        n11716) );
  AOI21_X1 U14320 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n14186), .A(n11716), .ZN(
        n11719) );
  OAI21_X1 U14321 ( .B1(n14169), .B2(n14122), .A(n11717), .ZN(n11718) );
  OAI211_X1 U14322 ( .C1(n12047), .C2(n13847), .A(n11719), .B(n11718), .ZN(
        P2_U3265) );
  INV_X1 U14323 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11721) );
  MUX2_X1 U14324 ( .A(n11721), .B(n11720), .S(n15549), .Z(n11722) );
  OAI21_X1 U14325 ( .B1(n13391), .B2(n15472), .A(n11722), .ZN(P3_U3463) );
  INV_X1 U14326 ( .A(n11724), .ZN(n11726) );
  OR2_X1 U14327 ( .A1(n11726), .A2(n11725), .ZN(n13851) );
  XNOR2_X1 U14328 ( .A(n11723), .B(n13851), .ZN(n15450) );
  XNOR2_X1 U14329 ( .A(n11727), .B(n13851), .ZN(n11728) );
  AOI222_X1 U14330 ( .A1(n14180), .A2(n11728), .B1(n13902), .B2(n14106), .C1(
        n6832), .C2(n14108), .ZN(n15455) );
  MUX2_X1 U14331 ( .A(n11729), .B(n15455), .S(n14135), .Z(n11734) );
  OAI21_X1 U14332 ( .B1(n11730), .B2(n15452), .A(n11745), .ZN(n15454) );
  OAI22_X1 U14333 ( .A1(n14052), .A2(n15454), .B1(n11731), .B2(n14146), .ZN(
        n11732) );
  AOI21_X1 U14334 ( .B1(n14169), .B2(n13687), .A(n11732), .ZN(n11733) );
  OAI211_X1 U14335 ( .C1(n14191), .C2(n15450), .A(n11734), .B(n11733), .ZN(
        P2_U3258) );
  INV_X1 U14336 ( .A(n11723), .ZN(n11737) );
  OAI21_X1 U14337 ( .B1(n11723), .B2(n13901), .A(n13687), .ZN(n11735) );
  OAI21_X1 U14338 ( .B1(n11737), .B2(n11736), .A(n11735), .ZN(n11739) );
  XNOR2_X1 U14339 ( .A(n11739), .B(n11738), .ZN(n14318) );
  OAI21_X1 U14340 ( .B1(n13854), .B2(n11786), .A(n11740), .ZN(n11741) );
  AOI222_X1 U14341 ( .A1(n14180), .A2(n11741), .B1(n13900), .B2(n14108), .C1(
        n13901), .C2(n14106), .ZN(n14317) );
  MUX2_X1 U14342 ( .A(n11742), .B(n14317), .S(n14135), .Z(n11750) );
  INV_X1 U14343 ( .A(n11743), .ZN(n11744) );
  AOI211_X1 U14344 ( .C1(n14314), .C2(n11745), .A(n15453), .B(n11744), .ZN(
        n14313) );
  INV_X1 U14345 ( .A(n14313), .ZN(n11747) );
  OAI22_X1 U14346 ( .A1(n11747), .A2(n14173), .B1(n11746), .B2(n14146), .ZN(
        n11748) );
  AOI21_X1 U14347 ( .B1(n14169), .B2(n14314), .A(n11748), .ZN(n11749) );
  OAI211_X1 U14348 ( .C1(n14191), .C2(n14318), .A(n11750), .B(n11749), .ZN(
        P2_U3257) );
  INV_X1 U14349 ( .A(n11751), .ZN(n11752) );
  AOI21_X1 U14350 ( .B1(n11754), .B2(n11753), .A(n11752), .ZN(n11760) );
  AOI22_X1 U14351 ( .A1(n13605), .A2(n6832), .B1(n13537), .B2(n13899), .ZN(
        n11759) );
  NOR2_X1 U14352 ( .A1(n13599), .A2(n11755), .ZN(n11756) );
  AOI211_X1 U14353 ( .C1(n14307), .C2(n13623), .A(n11757), .B(n11756), .ZN(
        n11758) );
  OAI211_X1 U14354 ( .C1(n11760), .C2(n13625), .A(n11759), .B(n11758), .ZN(
        P2_U3203) );
  NAND2_X1 U14355 ( .A1(n11762), .A2(n11761), .ZN(n11816) );
  XNOR2_X1 U14356 ( .A(n11816), .B(n12645), .ZN(n15528) );
  AND2_X1 U14357 ( .A1(n11763), .A2(n12761), .ZN(n15515) );
  NAND2_X1 U14358 ( .A1(n15500), .A2(n15515), .ZN(n13188) );
  INV_X1 U14359 ( .A(n15511), .ZN(n12120) );
  INV_X1 U14360 ( .A(n12645), .ZN(n12596) );
  NOR2_X1 U14361 ( .A1(n11764), .A2(n12596), .ZN(n11820) );
  AND2_X1 U14362 ( .A1(n11764), .A2(n12596), .ZN(n11765) );
  OAI21_X1 U14363 ( .B1(n11820), .B2(n11765), .A(n13308), .ZN(n11767) );
  AOI22_X1 U14364 ( .A1(n13320), .A2(n12971), .B1(n12973), .B2(n15504), .ZN(
        n11766) );
  OAI211_X1 U14365 ( .C1(n12120), .C2(n15528), .A(n11767), .B(n11766), .ZN(
        n15529) );
  MUX2_X1 U14366 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n15529), .S(n15500), .Z(
        n11768) );
  INV_X1 U14367 ( .A(n11768), .ZN(n11773) );
  INV_X1 U14368 ( .A(n11769), .ZN(n13252) );
  NOR2_X1 U14369 ( .A1(n11770), .A2(n15512), .ZN(n15530) );
  INV_X1 U14370 ( .A(n11771), .ZN(n12869) );
  AOI22_X1 U14371 ( .A1(n13252), .A2(n15530), .B1(n15516), .B2(n12869), .ZN(
        n11772) );
  OAI211_X1 U14372 ( .C1(n15528), .C2(n13188), .A(n11773), .B(n11772), .ZN(
        P3_U3228) );
  XNOR2_X1 U14373 ( .A(n11775), .B(n11774), .ZN(n11781) );
  NAND2_X1 U14374 ( .A1(n13623), .A2(n14302), .ZN(n11777) );
  NAND2_X1 U14375 ( .A1(n11777), .A2(n11776), .ZN(n11779) );
  OAI22_X1 U14376 ( .A1(n11788), .A2(n13618), .B1(n13621), .B2(n13709), .ZN(
        n11778) );
  AOI211_X1 U14377 ( .C1(n11797), .C2(n13634), .A(n11779), .B(n11778), .ZN(
        n11780) );
  OAI21_X1 U14378 ( .B1(n11781), .B2(n13625), .A(n11780), .ZN(P2_U3189) );
  NAND2_X1 U14379 ( .A1(n14307), .A2(n13900), .ZN(n11783) );
  INV_X1 U14380 ( .A(n13858), .ZN(n11887) );
  NAND3_X1 U14381 ( .A1(n11786), .A2(n11785), .A3(n11784), .ZN(n11793) );
  OAI21_X1 U14382 ( .B1(n11788), .B2(n11787), .A(n14307), .ZN(n11791) );
  XNOR2_X1 U14383 ( .A(n13858), .B(n11890), .ZN(n11794) );
  AOI222_X1 U14384 ( .A1(n14180), .A2(n11794), .B1(n13898), .B2(n14108), .C1(
        n13900), .C2(n14106), .ZN(n14305) );
  MUX2_X1 U14385 ( .A(n10925), .B(n14305), .S(n14135), .Z(n11802) );
  INV_X1 U14386 ( .A(n11795), .ZN(n11796) );
  INV_X1 U14387 ( .A(n14302), .ZN(n11799) );
  AOI21_X1 U14388 ( .B1(n14302), .B2(n11796), .A(n11889), .ZN(n14303) );
  INV_X1 U14389 ( .A(n11797), .ZN(n11798) );
  OAI22_X1 U14390 ( .A1(n14188), .A2(n11799), .B1(n14146), .B2(n11798), .ZN(
        n11800) );
  AOI21_X1 U14391 ( .B1(n14303), .B2(n14122), .A(n11800), .ZN(n11801) );
  OAI211_X1 U14392 ( .C1(n14306), .C2(n14191), .A(n11802), .B(n11801), .ZN(
        P2_U3255) );
  OR2_X1 U14393 ( .A1(n11805), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11803) );
  NAND2_X1 U14394 ( .A1(n11804), .A2(n11803), .ZN(n11956) );
  XNOR2_X1 U14395 ( .A(n11956), .B(n11812), .ZN(n11954) );
  XNOR2_X1 U14396 ( .A(n11954), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n11814) );
  INV_X1 U14397 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15185) );
  NAND2_X1 U14398 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14540)
         );
  OAI21_X1 U14399 ( .B1(n14650), .B2(n15185), .A(n14540), .ZN(n11811) );
  NAND2_X1 U14400 ( .A1(n11805), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11806) );
  NAND2_X1 U14401 ( .A1(n11808), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11809) );
  AOI21_X1 U14402 ( .B1(n11950), .B2(n11809), .A(n14712), .ZN(n11810) );
  AOI211_X1 U14403 ( .C1(n14653), .C2(n11812), .A(n11811), .B(n11810), .ZN(
        n11813) );
  OAI21_X1 U14404 ( .B1(n14714), .B2(n11814), .A(n11813), .ZN(P1_U3258) );
  OR2_X1 U14405 ( .A1(n15511), .A2(n15515), .ZN(n15477) );
  AOI21_X1 U14406 ( .B1(n11816), .B2(n12596), .A(n11815), .ZN(n11818) );
  XNOR2_X1 U14407 ( .A(n11818), .B(n12597), .ZN(n15533) );
  NOR2_X1 U14408 ( .A1(n11820), .A2(n11819), .ZN(n11821) );
  XNOR2_X1 U14409 ( .A(n11821), .B(n12597), .ZN(n11823) );
  INV_X1 U14410 ( .A(n12970), .ZN(n12222) );
  OAI22_X1 U14411 ( .A1(n12222), .A2(n15491), .B1(n12217), .B2(n15492), .ZN(
        n11822) );
  AOI21_X1 U14412 ( .B1(n11823), .B2(n13308), .A(n11822), .ZN(n15534) );
  MUX2_X1 U14413 ( .A(n6903), .B(n15534), .S(n15500), .Z(n11826) );
  NOR2_X1 U14414 ( .A1(n12216), .A2(n15512), .ZN(n15536) );
  INV_X1 U14415 ( .A(n11824), .ZN(n12934) );
  AOI22_X1 U14416 ( .A1(n13252), .A2(n15536), .B1(n15516), .B2(n12934), .ZN(
        n11825) );
  OAI211_X1 U14417 ( .C1(n13327), .C2(n15533), .A(n11826), .B(n11825), .ZN(
        P3_U3227) );
  XOR2_X1 U14418 ( .A(n11828), .B(n11827), .Z(n11845) );
  AND2_X1 U14419 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n12834) );
  INV_X1 U14420 ( .A(n12834), .ZN(n11829) );
  OAI21_X1 U14421 ( .B1(n13007), .B2(n11830), .A(n11829), .ZN(n11837) );
  OR3_X1 U14422 ( .A1(n11833), .A2(n11832), .A3(n11831), .ZN(n11834) );
  AOI21_X1 U14423 ( .B1(n11835), .B2(n11834), .A(n13077), .ZN(n11836) );
  AOI211_X1 U14424 ( .C1(n13014), .C2(n11838), .A(n11837), .B(n11836), .ZN(
        n11844) );
  NOR3_X1 U14425 ( .A1(n11841), .A2(n11840), .A3(n11839), .ZN(n11842) );
  OAI21_X1 U14426 ( .B1(n6721), .B2(n11842), .A(n13100), .ZN(n11843) );
  OAI211_X1 U14427 ( .C1(n11845), .C2(n13030), .A(n11844), .B(n11843), .ZN(
        P3_U3190) );
  NAND2_X1 U14428 ( .A1(n11847), .A2(n12656), .ZN(n11968) );
  OAI21_X1 U14429 ( .B1(n11847), .B2(n12656), .A(n11968), .ZN(n12004) );
  OAI211_X1 U14430 ( .C1(n11850), .C2(n11849), .A(n11848), .B(n13308), .ZN(
        n11852) );
  AOI22_X1 U14431 ( .A1(n15504), .A2(n12971), .B1(n12969), .B2(n13320), .ZN(
        n11851) );
  NAND2_X1 U14432 ( .A1(n11852), .A2(n11851), .ZN(n12001) );
  AOI21_X1 U14433 ( .B1(n15537), .B2(n12004), .A(n12001), .ZN(n11867) );
  AOI22_X1 U14434 ( .A1(n13458), .A2(n12777), .B1(P3_REG0_REG_7__SCAN_IN), 
        .B2(n15539), .ZN(n11853) );
  OAI21_X1 U14435 ( .B1(n11867), .B2(n15539), .A(n11853), .ZN(P3_U3411) );
  OAI21_X1 U14436 ( .B1(n11856), .B2(n11855), .A(n11854), .ZN(n11998) );
  INV_X1 U14437 ( .A(n11857), .ZN(n11859) );
  OAI21_X1 U14438 ( .B1(n12205), .B2(n11859), .A(n7503), .ZN(n11994) );
  OAI22_X1 U14439 ( .A1(n11994), .A2(n15323), .B1(n12205), .B2(n15335), .ZN(
        n11863) );
  XNOR2_X1 U14440 ( .A(n11860), .B(n7782), .ZN(n11862) );
  OAI222_X1 U14441 ( .A1(n14909), .A2(n12206), .B1(n11862), .B2(n15276), .C1(
        n14907), .C2(n11861), .ZN(n11995) );
  AOI211_X1 U14442 ( .C1(n15339), .C2(n11998), .A(n11863), .B(n11995), .ZN(
        n11866) );
  NAND2_X1 U14443 ( .A1(n9548), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n11864) );
  OAI21_X1 U14444 ( .B1(n11866), .B2(n9548), .A(n11864), .ZN(P1_U3537) );
  NAND2_X1 U14445 ( .A1(n9554), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n11865) );
  OAI21_X1 U14446 ( .B1(n11866), .B2(n9554), .A(n11865), .ZN(P1_U3486) );
  MUX2_X1 U14447 ( .A(n15571), .B(n11867), .S(n15549), .Z(n11868) );
  OAI21_X1 U14448 ( .B1(n13391), .B2(n12000), .A(n11868), .ZN(P3_U3466) );
  NAND2_X1 U14449 ( .A1(n11869), .A2(n13480), .ZN(n11870) );
  OAI211_X1 U14450 ( .C1(n11871), .C2(n13487), .A(n11870), .B(n12768), .ZN(
        P3_U3272) );
  OAI211_X1 U14451 ( .C1(n11874), .C2(n11873), .A(n11872), .B(n15331), .ZN(
        n11876) );
  AOI22_X1 U14452 ( .A1(n14562), .A2(n14939), .B1(n14940), .B2(n14560), .ZN(
        n11875) );
  NAND2_X1 U14453 ( .A1(n11876), .A2(n11875), .ZN(n15089) );
  INV_X1 U14454 ( .A(n15089), .ZN(n11886) );
  OAI21_X1 U14455 ( .B1(n11879), .B2(n11878), .A(n11877), .ZN(n15091) );
  OAI21_X1 U14456 ( .B1(n11880), .B2(n15087), .A(n14975), .ZN(n15088) );
  OAI22_X1 U14457 ( .A1(n14987), .A2(n11881), .B1(n14505), .B2(n15280), .ZN(
        n11882) );
  AOI21_X1 U14458 ( .B1(n14752), .B2(n14507), .A(n11882), .ZN(n11883) );
  OAI21_X1 U14459 ( .B1(n15088), .B2(n11993), .A(n11883), .ZN(n11884) );
  AOI21_X1 U14460 ( .B1(n15091), .B2(n14990), .A(n11884), .ZN(n11885) );
  OAI21_X1 U14461 ( .B1(n11886), .B2(n6538), .A(n11885), .ZN(P1_U3282) );
  NAND2_X1 U14462 ( .A1(n14302), .A2(n13899), .ZN(n11888) );
  XNOR2_X1 U14463 ( .A(n13711), .B(n13709), .ZN(n13862) );
  INV_X1 U14464 ( .A(n13862), .ZN(n13706) );
  XNOR2_X1 U14465 ( .A(n12041), .B(n13706), .ZN(n12021) );
  INV_X1 U14466 ( .A(n13711), .ZN(n12036) );
  OAI211_X1 U14467 ( .C1(n11889), .C2(n12036), .A(n14308), .B(n12045), .ZN(
        n12017) );
  OAI21_X1 U14468 ( .B1(n12036), .B2(n15451), .A(n12017), .ZN(n11894) );
  INV_X1 U14469 ( .A(n13899), .ZN(n11891) );
  XNOR2_X1 U14470 ( .A(n12037), .B(n13706), .ZN(n11893) );
  INV_X1 U14471 ( .A(n13897), .ZN(n13717) );
  OAI22_X1 U14472 ( .A1(n14092), .A2(n11891), .B1(n13717), .B2(n14094), .ZN(
        n12008) );
  INV_X1 U14473 ( .A(n12008), .ZN(n11892) );
  OAI21_X1 U14474 ( .B1(n11893), .B2(n14162), .A(n11892), .ZN(n12018) );
  AOI211_X1 U14475 ( .C1(n15458), .C2(n12021), .A(n11894), .B(n12018), .ZN(
        n11897) );
  NAND2_X1 U14476 ( .A1(n15460), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n11895) );
  OAI21_X1 U14477 ( .B1(n11897), .B2(n15460), .A(n11895), .ZN(P2_U3463) );
  NAND2_X1 U14478 ( .A1(n15464), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11896) );
  OAI21_X1 U14479 ( .B1(n11897), .B2(n15464), .A(n11896), .ZN(P2_U3510) );
  OAI21_X1 U14480 ( .B1(n11900), .B2(n11899), .A(n11898), .ZN(n11901) );
  NAND2_X1 U14481 ( .A1(n11901), .A2(n14515), .ZN(n11906) );
  NOR2_X1 U14482 ( .A1(n14528), .A2(n11902), .ZN(n11903) );
  AOI211_X1 U14483 ( .C1(n14497), .C2(n15332), .A(n11904), .B(n11903), .ZN(
        n11905) );
  OAI211_X1 U14484 ( .C1(n15336), .C2(n14524), .A(n11906), .B(n11905), .ZN(
        P1_U3221) );
  INV_X1 U14485 ( .A(n11925), .ZN(n11909) );
  NAND2_X1 U14486 ( .A1(n14356), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11908) );
  OR2_X1 U14487 ( .A1(n11907), .A2(P2_U3088), .ZN(n13887) );
  OAI211_X1 U14488 ( .C1(n11909), .C2(n14360), .A(n11908), .B(n13887), .ZN(
        P2_U3304) );
  INV_X1 U14489 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n12086) );
  NAND2_X1 U14490 ( .A1(n12086), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n11912) );
  NAND2_X1 U14491 ( .A1(n11913), .A2(n11912), .ZN(n11917) );
  INV_X1 U14492 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11914) );
  NAND2_X1 U14493 ( .A1(n11914), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n12152) );
  NAND2_X1 U14494 ( .A1(n15705), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n11915) );
  AND2_X1 U14495 ( .A1(n12152), .A2(n11915), .ZN(n11916) );
  NAND2_X1 U14496 ( .A1(n11917), .A2(n11916), .ZN(n12153) );
  OR2_X1 U14497 ( .A1(n11917), .A2(n11916), .ZN(n11918) );
  AND2_X1 U14498 ( .A1(n12153), .A2(n11918), .ZN(n11919) );
  NAND2_X1 U14499 ( .A1(n12149), .A2(n12150), .ZN(n11921) );
  XNOR2_X1 U14500 ( .A(n11921), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  INV_X1 U14501 ( .A(n11922), .ZN(n11923) );
  INV_X1 U14502 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n15764) );
  OAI222_X1 U14503 ( .A1(P2_U3088), .A2(n11924), .B1(n14360), .B2(n11923), 
        .C1(n15764), .C2(n14362), .ZN(P2_U3305) );
  NAND2_X1 U14504 ( .A1(n11925), .A2(n15155), .ZN(n11927) );
  OAI211_X1 U14505 ( .C1(n11928), .C2(n12476), .A(n11927), .B(n11926), .ZN(
        P1_U3332) );
  XNOR2_X1 U14506 ( .A(n11930), .B(n12594), .ZN(n11931) );
  AOI222_X1 U14507 ( .A1(n13308), .A2(n11931), .B1(n12967), .B2(n13320), .C1(
        n12969), .C2(n15504), .ZN(n12077) );
  INV_X1 U14508 ( .A(n13461), .ZN(n13465) );
  XNOR2_X1 U14509 ( .A(n11932), .B(n12594), .ZN(n12076) );
  OAI22_X1 U14510 ( .A1(n13470), .A2(n12228), .B1(n11933), .B2(n15540), .ZN(
        n11934) );
  AOI21_X1 U14511 ( .B1(n13465), .B2(n12076), .A(n11934), .ZN(n11935) );
  OAI21_X1 U14512 ( .B1(n12077), .B2(n15539), .A(n11935), .ZN(P3_U3417) );
  AOI21_X1 U14513 ( .B1(n11937), .B2(n11939), .A(n11936), .ZN(n15254) );
  XNOR2_X1 U14514 ( .A(n11938), .B(n11939), .ZN(n11943) );
  NOR2_X1 U14515 ( .A1(n15254), .A2(n11940), .ZN(n11941) );
  AOI211_X1 U14516 ( .C1(n15331), .C2(n11943), .A(n11942), .B(n11941), .ZN(
        n15258) );
  OAI211_X1 U14517 ( .C1(n11944), .C2(n15251), .A(n11489), .B(n10110), .ZN(
        n15253) );
  OAI211_X1 U14518 ( .C1(n15254), .C2(n15310), .A(n15258), .B(n15253), .ZN(
        n11948) );
  OAI22_X1 U14519 ( .A1(n15086), .A2(n15251), .B1(n15348), .B2(n10732), .ZN(
        n11945) );
  AOI21_X1 U14520 ( .B1(n11948), .B2(n15348), .A(n11945), .ZN(n11946) );
  INV_X1 U14521 ( .A(n11946), .ZN(P1_U3535) );
  INV_X1 U14522 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15691) );
  OAI22_X1 U14523 ( .A1(n15147), .A2(n15251), .B1(n15342), .B2(n15691), .ZN(
        n11947) );
  AOI21_X1 U14524 ( .B1(n11948), .B2(n15342), .A(n11947), .ZN(n11949) );
  INV_X1 U14525 ( .A(n11949), .ZN(P1_U3480) );
  INV_X1 U14526 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14932) );
  MUX2_X1 U14527 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n14932), .S(n12196), .Z(
        n11951) );
  OAI211_X1 U14528 ( .C1(n11952), .C2(n11951), .A(n12193), .B(n14677), .ZN(
        n11965) );
  NAND2_X1 U14529 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14434)
         );
  XNOR2_X1 U14530 ( .A(n12196), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11959) );
  INV_X1 U14531 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11953) );
  NAND2_X1 U14532 ( .A1(n11954), .A2(n11953), .ZN(n11958) );
  NAND2_X1 U14533 ( .A1(n11956), .A2(n11955), .ZN(n11957) );
  NAND2_X1 U14534 ( .A1(n11958), .A2(n11957), .ZN(n11960) );
  AOI21_X1 U14535 ( .B1(n11959), .B2(n11960), .A(n14714), .ZN(n11961) );
  NAND2_X1 U14536 ( .A1(n11961), .A2(n12198), .ZN(n11962) );
  NAND2_X1 U14537 ( .A1(n14434), .A2(n11962), .ZN(n11963) );
  AOI21_X1 U14538 ( .B1(n15244), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11963), 
        .ZN(n11964) );
  OAI211_X1 U14539 ( .C1(n14709), .C2(n11966), .A(n11965), .B(n11964), .ZN(
        P1_U3259) );
  INV_X1 U14540 ( .A(n12660), .ZN(n11967) );
  NAND2_X1 U14541 ( .A1(n11968), .A2(n11967), .ZN(n11969) );
  NAND2_X1 U14542 ( .A1(n12666), .A2(n12665), .ZN(n12662) );
  XNOR2_X1 U14543 ( .A(n11969), .B(n12662), .ZN(n12075) );
  INV_X1 U14544 ( .A(n12075), .ZN(n11974) );
  XOR2_X1 U14545 ( .A(n12662), .B(n11970), .Z(n11971) );
  NAND2_X1 U14546 ( .A1(n11971), .A2(n13308), .ZN(n11973) );
  AOI22_X1 U14547 ( .A1(n15504), .A2(n12970), .B1(n12968), .B2(n13320), .ZN(
        n11972) );
  OAI211_X1 U14548 ( .C1(n12120), .C2(n12075), .A(n11973), .B(n11972), .ZN(
        n12070) );
  AOI21_X1 U14549 ( .B1(n6716), .B2(n11974), .A(n12070), .ZN(n12110) );
  AOI22_X1 U14550 ( .A1(n13458), .A2(n7141), .B1(P3_REG0_REG_8__SCAN_IN), .B2(
        n15539), .ZN(n11975) );
  OAI21_X1 U14551 ( .B1(n12110), .B2(n15539), .A(n11975), .ZN(P3_U3414) );
  NAND2_X1 U14552 ( .A1(n11976), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11980) );
  NAND2_X1 U14553 ( .A1(n11978), .A2(n11977), .ZN(n11979) );
  NAND2_X1 U14554 ( .A1(n11980), .A2(n11979), .ZN(n12137) );
  XNOR2_X1 U14555 ( .A(n12137), .B(n11985), .ZN(n12135) );
  XNOR2_X1 U14556 ( .A(n12135), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n11989) );
  INV_X1 U14557 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n15725) );
  OAI22_X1 U14558 ( .A1(n11983), .A2(n11982), .B1(n11981), .B2(n15725), .ZN(
        n12129) );
  XOR2_X1 U14559 ( .A(n12136), .B(n12129), .Z(n12130) );
  XOR2_X1 U14560 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n12130), .Z(n11987) );
  NAND2_X1 U14561 ( .A1(n15408), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n11984) );
  NAND2_X1 U14562 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n13631)
         );
  OAI211_X1 U14563 ( .C1(n15412), .C2(n11985), .A(n11984), .B(n13631), .ZN(
        n11986) );
  AOI21_X1 U14564 ( .B1(n11987), .B2(n15398), .A(n11986), .ZN(n11988) );
  OAI21_X1 U14565 ( .B1(n11989), .B2(n15414), .A(n11988), .ZN(P2_U3229) );
  INV_X1 U14566 ( .A(n12209), .ZN(n11990) );
  AOI22_X1 U14567 ( .A1(n14752), .A2(n11991), .B1(n11990), .B2(n14945), .ZN(
        n11992) );
  OAI21_X1 U14568 ( .B1(n11994), .B2(n11993), .A(n11992), .ZN(n11997) );
  MUX2_X1 U14569 ( .A(n11995), .B(P1_REG2_REG_9__SCAN_IN), .S(n6538), .Z(
        n11996) );
  AOI211_X1 U14570 ( .C1(n14990), .C2(n11998), .A(n11997), .B(n11996), .ZN(
        n11999) );
  INV_X1 U14571 ( .A(n11999), .ZN(P1_U3284) );
  INV_X1 U14572 ( .A(n13327), .ZN(n13255) );
  OAI22_X1 U14573 ( .A1(n15483), .A2(n12000), .B1(n12778), .B2(n15486), .ZN(
        n12003) );
  MUX2_X1 U14574 ( .A(n12001), .B(P3_REG2_REG_7__SCAN_IN), .S(n15519), .Z(
        n12002) );
  AOI211_X1 U14575 ( .C1(n12004), .C2(n13255), .A(n12003), .B(n12002), .ZN(
        n12005) );
  INV_X1 U14576 ( .A(n12005), .ZN(P3_U3226) );
  XNOR2_X1 U14577 ( .A(n12007), .B(n12006), .ZN(n12013) );
  NAND2_X1 U14578 ( .A1(n13550), .A2(n12008), .ZN(n12009) );
  OAI211_X1 U14579 ( .C1(n13599), .C2(n12014), .A(n12010), .B(n12009), .ZN(
        n12011) );
  AOI21_X1 U14580 ( .B1(n13711), .B2(n13623), .A(n12011), .ZN(n12012) );
  OAI21_X1 U14581 ( .B1(n12013), .B2(n13625), .A(n12012), .ZN(P2_U3208) );
  INV_X1 U14582 ( .A(n14191), .ZN(n14019) );
  INV_X1 U14583 ( .A(n12014), .ZN(n12015) );
  AOI22_X1 U14584 ( .A1(n14169), .A2(n13711), .B1(n12015), .B2(n14184), .ZN(
        n12016) );
  OAI21_X1 U14585 ( .B1(n12017), .B2(n14173), .A(n12016), .ZN(n12020) );
  MUX2_X1 U14586 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n12018), .S(n14135), .Z(
        n12019) );
  AOI211_X1 U14587 ( .C1(n14019), .C2(n12021), .A(n12020), .B(n12019), .ZN(
        n12022) );
  INV_X1 U14588 ( .A(n12022), .ZN(P2_U3254) );
  XOR2_X1 U14589 ( .A(n12024), .B(n12023), .Z(n12035) );
  OAI21_X1 U14590 ( .B1(n6720), .B2(P3_REG2_REG_9__SCAN_IN), .A(n12025), .ZN(
        n12033) );
  NOR2_X1 U14591 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12026), .ZN(n12895) );
  AOI21_X1 U14592 ( .B1(n15467), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12895), .ZN(
        n12027) );
  OAI21_X1 U14593 ( .B1(n13088), .B2(n12028), .A(n12027), .ZN(n12032) );
  AOI21_X1 U14594 ( .B1(n12066), .B2(n12029), .A(n12098), .ZN(n12030) );
  NOR2_X1 U14595 ( .A1(n12030), .A2(n13046), .ZN(n12031) );
  AOI211_X1 U14596 ( .C1(n13090), .C2(n12033), .A(n12032), .B(n12031), .ZN(
        n12034) );
  OAI21_X1 U14597 ( .B1(n12035), .B2(n13030), .A(n12034), .ZN(P3_U3191) );
  NOR2_X1 U14598 ( .A1(n14297), .A2(n13897), .ZN(n12178) );
  NAND2_X1 U14599 ( .A1(n14297), .A2(n13897), .ZN(n12177) );
  INV_X1 U14600 ( .A(n12177), .ZN(n12038) );
  OR2_X1 U14601 ( .A1(n12178), .A2(n12038), .ZN(n13860) );
  XNOR2_X1 U14602 ( .A(n12175), .B(n13860), .ZN(n12044) );
  AND2_X1 U14603 ( .A1(n13711), .A2(n13898), .ZN(n12040) );
  OR2_X1 U14604 ( .A1(n13711), .A2(n13898), .ZN(n12039) );
  XNOR2_X1 U14605 ( .A(n12179), .B(n13860), .ZN(n14300) );
  NOR2_X1 U14606 ( .A1(n14300), .A2(n10685), .ZN(n12043) );
  OAI22_X1 U14607 ( .A1(n14092), .A2(n13709), .B1(n13720), .B2(n14094), .ZN(
        n12042) );
  AOI211_X1 U14608 ( .C1(n12044), .C2(n14180), .A(n12043), .B(n12042), .ZN(
        n14299) );
  AOI211_X1 U14609 ( .C1(n14297), .C2(n12045), .A(n15453), .B(n7006), .ZN(
        n14296) );
  AOI22_X1 U14610 ( .A1(n14186), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12164), 
        .B2(n14184), .ZN(n12046) );
  OAI21_X1 U14611 ( .B1(n13716), .B2(n14188), .A(n12046), .ZN(n12049) );
  NOR2_X1 U14612 ( .A1(n14300), .A2(n12047), .ZN(n12048) );
  AOI211_X1 U14613 ( .C1(n14296), .C2(n14194), .A(n12049), .B(n12048), .ZN(
        n12050) );
  OAI21_X1 U14614 ( .B1(n14299), .B2(n14186), .A(n12050), .ZN(P2_U3253) );
  OAI211_X1 U14615 ( .C1(n12053), .C2(n12052), .A(n12051), .B(n15331), .ZN(
        n12055) );
  AOI22_X1 U14616 ( .A1(n14939), .A2(n14561), .B1(n14940), .B2(n14559), .ZN(
        n12054) );
  NAND2_X1 U14617 ( .A1(n12055), .A2(n12054), .ZN(n15081) );
  INV_X1 U14618 ( .A(n15081), .ZN(n12064) );
  OAI21_X1 U14619 ( .B1(n12057), .B2(n7748), .A(n12056), .ZN(n15083) );
  XNOR2_X1 U14620 ( .A(n14975), .B(n14974), .ZN(n12058) );
  NOR2_X1 U14621 ( .A1(n12058), .A2(n15323), .ZN(n15082) );
  NAND2_X1 U14622 ( .A1(n15082), .A2(n15289), .ZN(n12061) );
  INV_X1 U14623 ( .A(n12059), .ZN(n14415) );
  AOI22_X1 U14624 ( .A1(n6538), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n14415), 
        .B2(n14945), .ZN(n12060) );
  OAI211_X1 U14625 ( .C1(n15148), .C2(n15283), .A(n12061), .B(n12060), .ZN(
        n12062) );
  AOI21_X1 U14626 ( .B1(n15083), .B2(n14789), .A(n12062), .ZN(n12063) );
  OAI21_X1 U14627 ( .B1(n12064), .B2(n6538), .A(n12063), .ZN(P1_U3281) );
  NAND2_X1 U14628 ( .A1(n12966), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n12065) );
  OAI21_X1 U14629 ( .B1(n12966), .B2(n12584), .A(n12065), .ZN(P3_U3521) );
  MUX2_X1 U14630 ( .A(n12066), .B(n12077), .S(n15549), .Z(n12068) );
  INV_X1 U14631 ( .A(n13386), .ZN(n13388) );
  INV_X1 U14632 ( .A(n12228), .ZN(n12896) );
  AOI22_X1 U14633 ( .A1(n12076), .A2(n13388), .B1(n12896), .B2(n13383), .ZN(
        n12067) );
  NAND2_X1 U14634 ( .A1(n12068), .A2(n12067), .ZN(P3_U3468) );
  INV_X1 U14635 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n15639) );
  NAND2_X1 U14636 ( .A1(n13129), .A2(P3_U3897), .ZN(n12069) );
  OAI21_X1 U14637 ( .B1(P3_U3897), .B2(n15639), .A(n12069), .ZN(P3_U3517) );
  INV_X1 U14638 ( .A(n12070), .ZN(n12072) );
  MUX2_X1 U14639 ( .A(n12072), .B(n12071), .S(n15519), .Z(n12074) );
  AOI22_X1 U14640 ( .A1(n6529), .A2(n7141), .B1(n15516), .B2(n12835), .ZN(
        n12073) );
  OAI211_X1 U14641 ( .C1(n12075), .C2(n13188), .A(n12074), .B(n12073), .ZN(
        P3_U3225) );
  INV_X1 U14642 ( .A(n12076), .ZN(n12082) );
  MUX2_X1 U14643 ( .A(n12078), .B(n12077), .S(n15500), .Z(n12081) );
  INV_X1 U14644 ( .A(n12079), .ZN(n12897) );
  AOI22_X1 U14645 ( .A1(n6529), .A2(n12896), .B1(n15516), .B2(n12897), .ZN(
        n12080) );
  OAI211_X1 U14646 ( .C1(n12082), .C2(n13327), .A(n12081), .B(n12080), .ZN(
        P3_U3224) );
  XOR2_X1 U14647 ( .A(n12084), .B(n12083), .Z(n12103) );
  AND2_X1 U14648 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n12804) );
  INV_X1 U14649 ( .A(n12804), .ZN(n12085) );
  OAI21_X1 U14650 ( .B1(n13007), .B2(n12086), .A(n12085), .ZN(n12093) );
  INV_X1 U14651 ( .A(n12087), .ZN(n12089) );
  NAND3_X1 U14652 ( .A1(n12025), .A2(n12089), .A3(n12088), .ZN(n12090) );
  AOI21_X1 U14653 ( .B1(n12091), .B2(n12090), .A(n13077), .ZN(n12092) );
  AOI211_X1 U14654 ( .C1(n13014), .C2(n12094), .A(n12093), .B(n12092), .ZN(
        n12102) );
  INV_X1 U14655 ( .A(n12095), .ZN(n12100) );
  NOR3_X1 U14656 ( .A1(n12098), .A2(n12097), .A3(n12096), .ZN(n12099) );
  OAI21_X1 U14657 ( .B1(n12100), .B2(n12099), .A(n13100), .ZN(n12101) );
  OAI211_X1 U14658 ( .C1(n12103), .C2(n13030), .A(n12102), .B(n12101), .ZN(
        P3_U3192) );
  INV_X1 U14659 ( .A(n12104), .ZN(n12108) );
  OAI222_X1 U14660 ( .A1(P1_U3086), .A2(n12106), .B1(n12474), .B2(n12108), 
        .C1(n12105), .C2(n15161), .ZN(P1_U3331) );
  INV_X1 U14661 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12107) );
  OAI222_X1 U14662 ( .A1(n12109), .A2(P2_U3088), .B1(n14360), .B2(n12108), 
        .C1(n12107), .C2(n14362), .ZN(P2_U3303) );
  MUX2_X1 U14663 ( .A(n12111), .B(n12110), .S(n15549), .Z(n12112) );
  OAI21_X1 U14664 ( .B1(n12219), .B2(n13391), .A(n12112), .ZN(P3_U3467) );
  NAND2_X1 U14665 ( .A1(n12113), .A2(n12680), .ZN(n12114) );
  NAND2_X1 U14666 ( .A1(n12115), .A2(n12114), .ZN(n12274) );
  INV_X1 U14667 ( .A(n12274), .ZN(n12121) );
  XNOR2_X1 U14668 ( .A(n12116), .B(n8561), .ZN(n12117) );
  NAND2_X1 U14669 ( .A1(n12117), .A2(n13308), .ZN(n12119) );
  AOI22_X1 U14670 ( .A1(n13320), .A2(n13314), .B1(n12968), .B2(n15504), .ZN(
        n12118) );
  OAI211_X1 U14671 ( .C1(n12120), .C2(n12274), .A(n12119), .B(n12118), .ZN(
        n12268) );
  AOI21_X1 U14672 ( .B1(n6716), .B2(n12121), .A(n12268), .ZN(n12305) );
  INV_X1 U14673 ( .A(n12308), .ZN(n12805) );
  AOI22_X1 U14674 ( .A1(n13458), .A2(n12805), .B1(P3_REG0_REG_10__SCAN_IN), 
        .B2(n15539), .ZN(n12122) );
  OAI21_X1 U14675 ( .B1(n12305), .B2(n15539), .A(n12122), .ZN(P3_U3420) );
  INV_X1 U14676 ( .A(n12123), .ZN(n12127) );
  OAI222_X1 U14677 ( .A1(n12125), .A2(P2_U3088), .B1(n14360), .B2(n12127), 
        .C1(n12124), .C2(n14362), .ZN(P2_U3302) );
  OAI222_X1 U14678 ( .A1(P1_U3086), .A2(n12128), .B1(n12474), .B2(n12127), 
        .C1(n12126), .C2(n15161), .ZN(P1_U3330) );
  AOI22_X1 U14679 ( .A1(n12130), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n12136), 
        .B2(n12129), .ZN(n12245) );
  XNOR2_X1 U14680 ( .A(n12141), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n12244) );
  INV_X1 U14681 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n12131) );
  OAI22_X1 U14682 ( .A1(n12245), .A2(n12244), .B1(n12131), .B2(n12248), .ZN(
        n12406) );
  INV_X1 U14683 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n12132) );
  XNOR2_X1 U14684 ( .A(n12410), .B(n12132), .ZN(n12405) );
  XNOR2_X1 U14685 ( .A(n12406), .B(n12405), .ZN(n12148) );
  INV_X1 U14686 ( .A(n15412), .ZN(n13908) );
  INV_X1 U14687 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n12133) );
  NAND2_X1 U14688 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13564)
         );
  OAI21_X1 U14689 ( .B1(n15406), .B2(n12133), .A(n13564), .ZN(n12134) );
  AOI21_X1 U14690 ( .B1(n12410), .B2(n13908), .A(n12134), .ZN(n12147) );
  NAND2_X1 U14691 ( .A1(n12135), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n12139) );
  NAND2_X1 U14692 ( .A1(n12137), .A2(n12136), .ZN(n12138) );
  NAND2_X1 U14693 ( .A1(n12139), .A2(n12138), .ZN(n12243) );
  XNOR2_X1 U14694 ( .A(n12141), .B(n12140), .ZN(n12242) );
  NAND2_X1 U14695 ( .A1(n12243), .A2(n12242), .ZN(n12143) );
  NAND2_X1 U14696 ( .A1(n12141), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n12142) );
  NAND2_X1 U14697 ( .A1(n12143), .A2(n12142), .ZN(n12145) );
  MUX2_X1 U14698 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n14134), .S(n12410), .Z(
        n12144) );
  NAND2_X1 U14699 ( .A1(n12145), .A2(n12144), .ZN(n12412) );
  OAI211_X1 U14700 ( .C1(n12145), .C2(n12144), .A(n12412), .B(n15394), .ZN(
        n12146) );
  OAI211_X1 U14701 ( .C1(n12148), .C2(n15420), .A(n12147), .B(n12146), .ZN(
        P2_U3231) );
  NAND2_X1 U14702 ( .A1(n12153), .A2(n12152), .ZN(n12358) );
  INV_X1 U14703 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n12154) );
  XNOR2_X1 U14704 ( .A(n12154), .B(P1_ADDR_REG_12__SCAN_IN), .ZN(n12357) );
  XNOR2_X1 U14705 ( .A(n12358), .B(n12357), .ZN(n12155) );
  NAND2_X1 U14706 ( .A1(n12156), .A2(n12155), .ZN(n12356) );
  NAND2_X1 U14707 ( .A1(n12355), .A2(n12356), .ZN(n12157) );
  XNOR2_X1 U14708 ( .A(n12157), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  INV_X1 U14709 ( .A(n12159), .ZN(n12161) );
  NAND2_X1 U14710 ( .A1(n12161), .A2(n12160), .ZN(n12162) );
  XNOR2_X1 U14711 ( .A(n12158), .B(n12162), .ZN(n12163) );
  NAND2_X1 U14712 ( .A1(n12163), .A2(n13627), .ZN(n12169) );
  INV_X1 U14713 ( .A(n12164), .ZN(n12165) );
  OAI22_X1 U14714 ( .A1(n13621), .A2(n13720), .B1(n13599), .B2(n12165), .ZN(
        n12167) );
  NAND2_X1 U14715 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n15404)
         );
  OAI21_X1 U14716 ( .B1(n13618), .B2(n13709), .A(n15404), .ZN(n12166) );
  NOR2_X1 U14717 ( .A1(n12167), .A2(n12166), .ZN(n12168) );
  OAI211_X1 U14718 ( .C1(n13716), .C2(n13637), .A(n12169), .B(n12168), .ZN(
        P2_U3196) );
  INV_X1 U14719 ( .A(n12170), .ZN(n12172) );
  INV_X1 U14720 ( .A(n8517), .ZN(n12171) );
  OAI222_X1 U14721 ( .A1(n13487), .A2(n12173), .B1(n13495), .B2(n12172), .C1(
        n12171), .C2(P3_U3151), .ZN(P3_U3271) );
  NOR2_X1 U14722 ( .A1(n13716), .A2(n13897), .ZN(n12174) );
  NOR2_X1 U14723 ( .A1(n14292), .A2(n13720), .ZN(n13861) );
  XNOR2_X1 U14724 ( .A(n13724), .B(n13895), .ZN(n13866) );
  XNOR2_X1 U14725 ( .A(n12520), .B(n13866), .ZN(n12176) );
  AOI222_X1 U14726 ( .A1(n14180), .A2(n12176), .B1(n13894), .B2(n14108), .C1(
        n13896), .C2(n14106), .ZN(n14289) );
  INV_X1 U14727 ( .A(n13866), .ZN(n12180) );
  NAND2_X1 U14728 ( .A1(n12181), .A2(n13866), .ZN(n12182) );
  NAND2_X1 U14729 ( .A1(n12500), .A2(n12182), .ZN(n14290) );
  INV_X1 U14730 ( .A(n14290), .ZN(n12187) );
  INV_X1 U14731 ( .A(n13724), .ZN(n14285) );
  NOR2_X1 U14732 ( .A1(n14182), .A2(n14285), .ZN(n12183) );
  OR2_X1 U14733 ( .A1(n14167), .A2(n12183), .ZN(n14286) );
  AOI22_X1 U14734 ( .A1(n14186), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n13507), 
        .B2(n14184), .ZN(n12185) );
  NAND2_X1 U14735 ( .A1(n13724), .A2(n14169), .ZN(n12184) );
  OAI211_X1 U14736 ( .C1(n14286), .C2(n14052), .A(n12185), .B(n12184), .ZN(
        n12186) );
  AOI21_X1 U14737 ( .B1(n12187), .B2(n14019), .A(n12186), .ZN(n12188) );
  OAI21_X1 U14738 ( .B1(n14289), .B2(n14186), .A(n12188), .ZN(P2_U3251) );
  NAND2_X1 U14739 ( .A1(n12196), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n12192) );
  INV_X1 U14740 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n12189) );
  MUX2_X1 U14741 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n12189), .S(n14685), .Z(
        n12190) );
  MUX2_X1 U14742 ( .A(n12189), .B(P1_REG2_REG_17__SCAN_IN), .S(n14685), .Z(
        n12191) );
  NAND3_X1 U14743 ( .A1(n12193), .A2(n12192), .A3(n12191), .ZN(n12194) );
  NAND3_X1 U14744 ( .A1(n14682), .A2(n14677), .A3(n12194), .ZN(n12203) );
  NAND2_X1 U14745 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14447)
         );
  INV_X1 U14746 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n12195) );
  XNOR2_X1 U14747 ( .A(n14685), .B(n12195), .ZN(n14683) );
  NAND2_X1 U14748 ( .A1(n12196), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n12197) );
  NAND2_X1 U14749 ( .A1(n12198), .A2(n12197), .ZN(n14684) );
  XOR2_X1 U14750 ( .A(n14683), .B(n14684), .Z(n12199) );
  NAND2_X1 U14751 ( .A1(n14708), .A2(n12199), .ZN(n12200) );
  NAND2_X1 U14752 ( .A1(n14447), .A2(n12200), .ZN(n12201) );
  AOI21_X1 U14753 ( .B1(n15244), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n12201), 
        .ZN(n12202) );
  OAI211_X1 U14754 ( .C1(n14709), .C2(n12204), .A(n12203), .B(n12202), .ZN(
        P1_U3260) );
  XNOR2_X1 U14755 ( .A(n12289), .B(n12288), .ZN(n12291) );
  XNOR2_X1 U14756 ( .A(n12291), .B(n12290), .ZN(n12212) );
  INV_X1 U14757 ( .A(n14521), .ZN(n14542) );
  OAI22_X1 U14758 ( .A1(n12206), .A2(n14542), .B1(n14524), .B2(n12205), .ZN(
        n12211) );
  NAND2_X1 U14759 ( .A1(n14538), .A2(n14564), .ZN(n12208) );
  OAI211_X1 U14760 ( .C1(n14528), .C2(n12209), .A(n12208), .B(n12207), .ZN(
        n12210) );
  AOI211_X1 U14761 ( .C1(n12212), .C2(n14515), .A(n12211), .B(n12210), .ZN(
        n12213) );
  INV_X1 U14762 ( .A(n12213), .ZN(P1_U3231) );
  XNOR2_X1 U14763 ( .A(n12447), .B(n12868), .ZN(n12218) );
  XNOR2_X1 U14764 ( .A(n12218), .B(n12972), .ZN(n12865) );
  NAND2_X1 U14765 ( .A1(n12864), .A2(n12865), .ZN(n12863) );
  XNOR2_X1 U14766 ( .A(n12447), .B(n12216), .ZN(n12773) );
  NAND2_X1 U14767 ( .A1(n12218), .A2(n12217), .ZN(n12772) );
  XNOR2_X1 U14768 ( .A(n12447), .B(n12656), .ZN(n12223) );
  OAI211_X1 U14769 ( .C1(n12773), .C2(n12971), .A(n12772), .B(n12223), .ZN(
        n12220) );
  INV_X1 U14770 ( .A(n12223), .ZN(n12829) );
  OAI21_X1 U14771 ( .B1(n12831), .B2(n12222), .A(n12829), .ZN(n12226) );
  NAND2_X1 U14772 ( .A1(n12773), .A2(n12971), .ZN(n12774) );
  AOI22_X1 U14773 ( .A1(n12226), .A2(n12225), .B1(n12224), .B2(n12969), .ZN(
        n12227) );
  XNOR2_X1 U14774 ( .A(n12447), .B(n12228), .ZN(n12229) );
  XNOR2_X1 U14775 ( .A(n12229), .B(n12968), .ZN(n12893) );
  XNOR2_X1 U14776 ( .A(n12447), .B(n12308), .ZN(n12233) );
  XNOR2_X1 U14777 ( .A(n12233), .B(n12237), .ZN(n12802) );
  INV_X1 U14778 ( .A(n12229), .ZN(n12231) );
  NAND2_X1 U14779 ( .A1(n12231), .A2(n12230), .ZN(n12800) );
  AND2_X1 U14780 ( .A1(n12802), .A2(n12800), .ZN(n12232) );
  NAND2_X1 U14781 ( .A1(n12233), .A2(n12967), .ZN(n12234) );
  XNOR2_X1 U14782 ( .A(n12235), .B(n12462), .ZN(n12325) );
  XNOR2_X1 U14783 ( .A(n12327), .B(n12325), .ZN(n12328) );
  XNOR2_X1 U14784 ( .A(n12328), .B(n13314), .ZN(n12241) );
  INV_X1 U14785 ( .A(n12235), .ZN(n12313) );
  NAND2_X1 U14786 ( .A1(n12933), .A2(n13306), .ZN(n12236) );
  NAND2_X1 U14787 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12979)
         );
  OAI211_X1 U14788 ( .C1(n12237), .C2(n12922), .A(n12236), .B(n12979), .ZN(
        n12239) );
  INV_X1 U14789 ( .A(n12952), .ZN(n12944) );
  NOR2_X1 U14790 ( .A1(n12944), .A2(n12311), .ZN(n12238) );
  AOI211_X1 U14791 ( .C1(n12958), .C2(n12313), .A(n12239), .B(n12238), .ZN(
        n12240) );
  OAI21_X1 U14792 ( .B1(n12241), .B2(n12960), .A(n12240), .ZN(P3_U3176) );
  XNOR2_X1 U14793 ( .A(n12243), .B(n12242), .ZN(n12252) );
  NAND2_X1 U14794 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13552)
         );
  XOR2_X1 U14795 ( .A(n12245), .B(n12244), .Z(n12246) );
  NAND2_X1 U14796 ( .A1(n15398), .A2(n12246), .ZN(n12247) );
  NAND2_X1 U14797 ( .A1(n13552), .A2(n12247), .ZN(n12250) );
  NOR2_X1 U14798 ( .A1(n15412), .A2(n12248), .ZN(n12249) );
  AOI211_X1 U14799 ( .C1(n15408), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n12250), 
        .B(n12249), .ZN(n12251) );
  OAI21_X1 U14800 ( .B1(n12252), .B2(n15414), .A(n12251), .ZN(P2_U3230) );
  XNOR2_X1 U14801 ( .A(n13469), .B(n12447), .ZN(n12253) );
  NAND2_X1 U14802 ( .A1(n12253), .A2(n13306), .ZN(n12330) );
  OAI21_X1 U14803 ( .B1(n12336), .B2(n12325), .A(n12330), .ZN(n12257) );
  NAND3_X1 U14804 ( .A1(n12330), .A2(n12336), .A3(n12325), .ZN(n12255) );
  INV_X1 U14805 ( .A(n12253), .ZN(n12254) );
  NAND2_X1 U14806 ( .A1(n12254), .A2(n12262), .ZN(n12329) );
  AND2_X1 U14807 ( .A1(n12255), .A2(n12329), .ZN(n12256) );
  XNOR2_X1 U14808 ( .A(n12263), .B(n12462), .ZN(n12258) );
  INV_X1 U14809 ( .A(n12258), .ZN(n12259) );
  NAND2_X1 U14810 ( .A1(n12259), .A2(n13319), .ZN(n12341) );
  NAND2_X1 U14811 ( .A1(n6722), .A2(n12341), .ZN(n12260) );
  XNOR2_X1 U14812 ( .A(n12342), .B(n12260), .ZN(n12267) );
  NAND2_X1 U14813 ( .A1(n12933), .A2(n13305), .ZN(n12261) );
  NAND2_X1 U14814 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12997)
         );
  OAI211_X1 U14815 ( .C1(n12262), .C2(n12922), .A(n12261), .B(n12997), .ZN(
        n12265) );
  NOR2_X1 U14816 ( .A1(n12926), .A2(n12263), .ZN(n12264) );
  AOI211_X1 U14817 ( .C1(n13310), .C2(n12952), .A(n12265), .B(n12264), .ZN(
        n12266) );
  OAI21_X1 U14818 ( .B1(n12267), .B2(n12960), .A(n12266), .ZN(P3_U3174) );
  INV_X1 U14819 ( .A(n12268), .ZN(n12269) );
  MUX2_X1 U14820 ( .A(n12270), .B(n12269), .S(n15500), .Z(n12273) );
  INV_X1 U14821 ( .A(n12271), .ZN(n12806) );
  AOI22_X1 U14822 ( .A1(n6529), .A2(n12805), .B1(n15516), .B2(n12806), .ZN(
        n12272) );
  OAI211_X1 U14823 ( .C1(n12274), .C2(n13188), .A(n12273), .B(n12272), .ZN(
        P3_U3223) );
  XNOR2_X1 U14824 ( .A(n12276), .B(n12679), .ZN(n12277) );
  AOI222_X1 U14825 ( .A1(n13308), .A2(n12277), .B1(n12967), .B2(n15504), .C1(
        n13306), .C2(n13320), .ZN(n12310) );
  MUX2_X1 U14826 ( .A(n15739), .B(n12310), .S(n15549), .Z(n12280) );
  OAI21_X1 U14827 ( .B1(n6712), .B2(n12679), .A(n12278), .ZN(n12309) );
  AOI22_X1 U14828 ( .A1(n12309), .A2(n13388), .B1(n12313), .B2(n13383), .ZN(
        n12279) );
  NAND2_X1 U14829 ( .A1(n12280), .A2(n12279), .ZN(P3_U3470) );
  MUX2_X1 U14830 ( .A(n12281), .B(n12310), .S(n15540), .Z(n12283) );
  AOI22_X1 U14831 ( .A1(n12309), .A2(n13465), .B1(n12313), .B2(n13458), .ZN(
        n12282) );
  NAND2_X1 U14832 ( .A1(n12283), .A2(n12282), .ZN(P3_U3423) );
  INV_X1 U14833 ( .A(n12284), .ZN(n12287) );
  OAI222_X1 U14834 ( .A1(n13495), .A2(n12287), .B1(P3_U3151), .B2(n12286), 
        .C1(n12285), .C2(n13487), .ZN(P3_U3270) );
  OAI22_X1 U14835 ( .A1(n12291), .A2(n12290), .B1(n12289), .B2(n12288), .ZN(
        n12295) );
  XOR2_X1 U14836 ( .A(n12293), .B(n12292), .Z(n12294) );
  XNOR2_X1 U14837 ( .A(n12295), .B(n12294), .ZN(n12303) );
  INV_X1 U14838 ( .A(n12296), .ZN(n12297) );
  AOI22_X1 U14839 ( .A1(n14539), .A2(n12297), .B1(n14521), .B2(n14561), .ZN(
        n12300) );
  AOI21_X1 U14840 ( .B1(n14538), .B2(n14563), .A(n12298), .ZN(n12299) );
  OAI211_X1 U14841 ( .C1(n12301), .C2(n14524), .A(n12300), .B(n12299), .ZN(
        n12302) );
  AOI21_X1 U14842 ( .B1(n12303), .B2(n14515), .A(n12302), .ZN(n12304) );
  INV_X1 U14843 ( .A(n12304), .ZN(P1_U3217) );
  MUX2_X1 U14844 ( .A(n12306), .B(n12305), .S(n15549), .Z(n12307) );
  OAI21_X1 U14845 ( .B1(n13391), .B2(n12308), .A(n12307), .ZN(P3_U3469) );
  INV_X1 U14846 ( .A(n12309), .ZN(n12316) );
  MUX2_X1 U14847 ( .A(n7465), .B(n12310), .S(n15500), .Z(n12315) );
  INV_X1 U14848 ( .A(n12311), .ZN(n12312) );
  AOI22_X1 U14849 ( .A1(n6529), .A2(n12313), .B1(n15516), .B2(n12312), .ZN(
        n12314) );
  OAI211_X1 U14850 ( .C1(n12316), .C2(n13327), .A(n12315), .B(n12314), .ZN(
        P3_U3222) );
  AOI21_X1 U14851 ( .B1(n12318), .B2(n12317), .A(n13625), .ZN(n12320) );
  NAND2_X1 U14852 ( .A1(n12320), .A2(n12319), .ZN(n12324) );
  INV_X1 U14853 ( .A(n12321), .ZN(n14185) );
  AOI22_X1 U14854 ( .A1(n13895), .A2(n14108), .B1(n14106), .B2(n13897), .ZN(
        n14178) );
  NAND2_X1 U14855 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n15410)
         );
  OAI21_X1 U14856 ( .B1(n13632), .B2(n14178), .A(n15410), .ZN(n12322) );
  AOI21_X1 U14857 ( .B1(n13634), .B2(n14185), .A(n12322), .ZN(n12323) );
  OAI211_X1 U14858 ( .C1(n7578), .C2(n13637), .A(n12324), .B(n12323), .ZN(
        P2_U3206) );
  INV_X1 U14859 ( .A(n12325), .ZN(n12326) );
  AOI22_X1 U14860 ( .A1(n12328), .A2(n13314), .B1(n12327), .B2(n12326), .ZN(
        n12332) );
  NAND2_X1 U14861 ( .A1(n12330), .A2(n12329), .ZN(n12331) );
  XNOR2_X1 U14862 ( .A(n12332), .B(n12331), .ZN(n12340) );
  INV_X1 U14863 ( .A(n12333), .ZN(n13322) );
  NAND2_X1 U14864 ( .A1(n12933), .A2(n13319), .ZN(n12335) );
  OAI211_X1 U14865 ( .C1(n12336), .C2(n12922), .A(n12335), .B(n12334), .ZN(
        n12338) );
  NOR2_X1 U14866 ( .A1(n12926), .A2(n13469), .ZN(n12337) );
  AOI211_X1 U14867 ( .C1(n13322), .C2(n12952), .A(n12338), .B(n12337), .ZN(
        n12339) );
  OAI21_X1 U14868 ( .B1(n12340), .B2(n12960), .A(n12339), .ZN(P3_U3164) );
  INV_X1 U14869 ( .A(n13452), .ZN(n12350) );
  XNOR2_X1 U14870 ( .A(n13452), .B(n12447), .ZN(n12425) );
  XNOR2_X1 U14871 ( .A(n12425), .B(n13305), .ZN(n12343) );
  OAI211_X1 U14872 ( .C1(n12344), .C2(n12343), .A(n12428), .B(n7163), .ZN(
        n12349) );
  NAND2_X1 U14873 ( .A1(n12933), .A2(n13295), .ZN(n12345) );
  NAND2_X1 U14874 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13006)
         );
  OAI211_X1 U14875 ( .C1(n12346), .C2(n12922), .A(n12345), .B(n13006), .ZN(
        n12347) );
  AOI21_X1 U14876 ( .B1(n13298), .B2(n12952), .A(n12347), .ZN(n12348) );
  OAI211_X1 U14877 ( .C1(n12350), .C2(n12926), .A(n12349), .B(n12348), .ZN(
        P3_U3155) );
  INV_X1 U14878 ( .A(n12351), .ZN(n12352) );
  OAI222_X1 U14879 ( .A1(n9532), .A2(P1_U3086), .B1(n12474), .B2(n12352), .C1(
        n15628), .C2(n15161), .ZN(P1_U3329) );
  OAI222_X1 U14880 ( .A1(P2_U3088), .A2(n12354), .B1(n14362), .B2(n12353), 
        .C1(n14360), .C2(n12352), .ZN(P2_U3301) );
  NAND2_X1 U14881 ( .A1(n12359), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n12360) );
  XNOR2_X1 U14882 ( .A(P1_ADDR_REG_13__SCAN_IN), .B(P3_ADDR_REG_13__SCAN_IN), 
        .ZN(n12362) );
  XNOR2_X1 U14883 ( .A(n12371), .B(n12362), .ZN(n12363) );
  NAND2_X1 U14884 ( .A1(n12366), .A2(n12367), .ZN(n12365) );
  XNOR2_X1 U14885 ( .A(n12365), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  INV_X1 U14886 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n12369) );
  NAND2_X1 U14887 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n12369), .ZN(n12370) );
  NAND2_X1 U14888 ( .A1(n12371), .A2(n12370), .ZN(n12374) );
  INV_X1 U14889 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n12372) );
  NAND2_X1 U14890 ( .A1(n12372), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n12373) );
  NAND2_X1 U14891 ( .A1(n12374), .A2(n12373), .ZN(n15174) );
  INV_X1 U14892 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n12375) );
  XNOR2_X1 U14893 ( .A(n12375), .B(P3_ADDR_REG_14__SCAN_IN), .ZN(n15173) );
  INV_X1 U14894 ( .A(n15173), .ZN(n12376) );
  XNOR2_X1 U14895 ( .A(n15174), .B(n12376), .ZN(n15170) );
  XNOR2_X1 U14896 ( .A(n15170), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(n12377) );
  XNOR2_X1 U14897 ( .A(n15169), .B(n12377), .ZN(SUB_1596_U66) );
  INV_X1 U14898 ( .A(n12378), .ZN(n14359) );
  OAI222_X1 U14899 ( .A1(P1_U3086), .A2(n14586), .B1(n12474), .B2(n14359), 
        .C1(n12379), .C2(n15161), .ZN(P1_U3328) );
  OAI222_X1 U14900 ( .A1(n14360), .A2(n12381), .B1(n14362), .B2(n12380), .C1(
        P2_U3088), .C2(n13833), .ZN(P2_U3307) );
  OAI222_X1 U14901 ( .A1(P1_U3086), .A2(n12384), .B1(n12474), .B2(n12383), 
        .C1(n12382), .C2(n15161), .ZN(P1_U3334) );
  INV_X1 U14902 ( .A(n12385), .ZN(n12386) );
  OAI222_X1 U14903 ( .A1(n13495), .A2(n12386), .B1(n7986), .B2(P3_U3151), .C1(
        n15723), .C2(n13487), .ZN(P3_U3267) );
  OAI222_X1 U14904 ( .A1(n12474), .A2(n13800), .B1(n8603), .B2(P1_U3086), .C1(
        n12554), .C2(n15161), .ZN(P1_U3325) );
  INV_X1 U14905 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12387) );
  OAI222_X1 U14906 ( .A1(n12388), .A2(P2_U3088), .B1(n14362), .B2(n12387), 
        .C1(n14360), .C2(n13800), .ZN(P2_U3297) );
  XOR2_X1 U14907 ( .A(n12391), .B(n12389), .Z(n12395) );
  AOI22_X1 U14908 ( .A1(n14544), .A2(n15294), .B1(n14538), .B2(n12392), .ZN(
        n12394) );
  AOI22_X1 U14909 ( .A1(n14521), .A2(n9433), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n12482), .ZN(n12393) );
  OAI211_X1 U14910 ( .C1(n12395), .C2(n14546), .A(n12394), .B(n12393), .ZN(
        P1_U3222) );
  INV_X1 U14911 ( .A(n12396), .ZN(n12404) );
  NAND2_X1 U14912 ( .A1(n12397), .A2(n14987), .ZN(n12403) );
  NOR2_X1 U14913 ( .A1(n15110), .A2(n15283), .ZN(n12400) );
  OAI22_X1 U14914 ( .A1(n14367), .A2(n15280), .B1(n12398), .B2(n14987), .ZN(
        n12399) );
  AOI211_X1 U14915 ( .C1(n12401), .C2(n15289), .A(n12400), .B(n12399), .ZN(
        n12402) );
  OAI211_X1 U14916 ( .C1(n12404), .C2(n15285), .A(n12403), .B(n12402), .ZN(
        P1_U3266) );
  XNOR2_X1 U14917 ( .A(n12407), .B(n12413), .ZN(n13925) );
  INV_X1 U14918 ( .A(n12407), .ZN(n12408) );
  AOI22_X1 U14919 ( .A1(n13925), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n12413), 
        .B2(n12408), .ZN(n12409) );
  XNOR2_X1 U14920 ( .A(n12409), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n12419) );
  NAND2_X1 U14921 ( .A1(n12410), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12411) );
  NAND2_X1 U14922 ( .A1(n12412), .A2(n12411), .ZN(n12414) );
  NAND2_X1 U14923 ( .A1(n12414), .A2(n12413), .ZN(n12415) );
  NAND2_X1 U14924 ( .A1(n12416), .A2(n12415), .ZN(n13924) );
  OR2_X2 U14925 ( .A1(n13924), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13922) );
  NAND2_X1 U14926 ( .A1(n13922), .A2(n12416), .ZN(n12417) );
  XNOR2_X1 U14927 ( .A(n12417), .B(n14100), .ZN(n12421) );
  INV_X1 U14928 ( .A(n12421), .ZN(n12418) );
  OAI21_X1 U14929 ( .B1(n12419), .B2(n15420), .A(n15412), .ZN(n12420) );
  NAND2_X1 U14930 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13523)
         );
  OAI211_X1 U14931 ( .C1(n12424), .C2(n15406), .A(n12423), .B(n13523), .ZN(
        P2_U3233) );
  XNOR2_X1 U14932 ( .A(n13411), .B(n12462), .ZN(n12791) );
  INV_X1 U14933 ( .A(n12425), .ZN(n12426) );
  NAND2_X1 U14934 ( .A1(n12426), .A2(n13305), .ZN(n12427) );
  XNOR2_X1 U14935 ( .A(n13446), .B(n12462), .ZN(n12948) );
  OAI21_X1 U14936 ( .B1(n12950), .B2(n12948), .A(n13295), .ZN(n12430) );
  NAND2_X1 U14937 ( .A1(n12950), .A2(n12948), .ZN(n12429) );
  XNOR2_X1 U14938 ( .A(n13373), .B(n12462), .ZN(n12854) );
  AND2_X1 U14939 ( .A1(n12854), .A2(n13283), .ZN(n12431) );
  INV_X1 U14940 ( .A(n12854), .ZN(n12432) );
  NAND2_X1 U14941 ( .A1(n12432), .A2(n12955), .ZN(n12433) );
  XNOR2_X1 U14942 ( .A(n13436), .B(n11421), .ZN(n12435) );
  XNOR2_X1 U14943 ( .A(n12435), .B(n13273), .ZN(n12874) );
  INV_X1 U14944 ( .A(n12874), .ZN(n12434) );
  INV_X1 U14945 ( .A(n12435), .ZN(n12436) );
  XNOR2_X1 U14946 ( .A(n13247), .B(n12447), .ZN(n12437) );
  XNOR2_X1 U14947 ( .A(n12437), .B(n13261), .ZN(n12918) );
  INV_X1 U14948 ( .A(n12437), .ZN(n12438) );
  NAND2_X1 U14949 ( .A1(n12438), .A2(n13261), .ZN(n12439) );
  XNOR2_X1 U14950 ( .A(n13432), .B(n12447), .ZN(n12440) );
  XNOR2_X1 U14951 ( .A(n12440), .B(n12906), .ZN(n12822) );
  NAND2_X1 U14952 ( .A1(n12440), .A2(n13243), .ZN(n12441) );
  XNOR2_X1 U14953 ( .A(n13423), .B(n12447), .ZN(n12442) );
  XNOR2_X1 U14954 ( .A(n12442), .B(n13233), .ZN(n12903) );
  XNOR2_X1 U14955 ( .A(n13417), .B(n12447), .ZN(n12444) );
  XNOR2_X1 U14956 ( .A(n12444), .B(n13222), .ZN(n12841) );
  NAND2_X1 U14957 ( .A1(n12444), .A2(n12443), .ZN(n12445) );
  XNOR2_X1 U14958 ( .A(n8571), .B(n11421), .ZN(n12886) );
  XNOR2_X1 U14959 ( .A(n13189), .B(n12447), .ZN(n12451) );
  INV_X1 U14960 ( .A(n12451), .ZN(n12884) );
  AOI22_X1 U14961 ( .A1(n12884), .A2(n13198), .B1(n12791), .B2(n13208), .ZN(
        n12448) );
  OAI21_X1 U14962 ( .B1(n12886), .B2(n13181), .A(n12448), .ZN(n12449) );
  INV_X1 U14963 ( .A(n12449), .ZN(n12450) );
  INV_X1 U14964 ( .A(n12886), .ZN(n12454) );
  AOI21_X1 U14965 ( .B1(n12451), .B2(n12913), .A(n13181), .ZN(n12453) );
  NAND3_X1 U14966 ( .A1(n12451), .A2(n12913), .A3(n13181), .ZN(n12452) );
  NAND2_X1 U14967 ( .A1(n12457), .A2(n12456), .ZN(n12847) );
  XNOR2_X1 U14968 ( .A(n13339), .B(n12447), .ZN(n12458) );
  XNOR2_X1 U14969 ( .A(n12458), .B(n13168), .ZN(n12848) );
  XNOR2_X1 U14970 ( .A(n8574), .B(n12462), .ZN(n12459) );
  XNOR2_X1 U14971 ( .A(n12459), .B(n13129), .ZN(n12940) );
  XNOR2_X1 U14972 ( .A(n13333), .B(n12462), .ZN(n12460) );
  XNOR2_X1 U14973 ( .A(n12460), .B(n13143), .ZN(n12785) );
  INV_X1 U14974 ( .A(n12460), .ZN(n12461) );
  AOI22_X1 U14975 ( .A1(n12951), .A2(n12964), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12465) );
  INV_X1 U14976 ( .A(n12463), .ZN(n13121) );
  NAND2_X1 U14977 ( .A1(n12952), .A2(n13121), .ZN(n12464) );
  OAI211_X1 U14978 ( .C1(n12576), .C2(n12956), .A(n12465), .B(n12464), .ZN(
        n12466) );
  AOI21_X1 U14979 ( .B1(n8579), .B2(n12958), .A(n12466), .ZN(n12467) );
  OAI21_X1 U14980 ( .B1(n12468), .B2(n12960), .A(n12467), .ZN(P3_U3160) );
  INV_X1 U14981 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n12470) );
  OAI21_X1 U14982 ( .B1(n12472), .B2(n15086), .A(n12471), .ZN(P1_U3556) );
  OAI222_X1 U14983 ( .A1(n12477), .A2(P1_U3086), .B1(n12476), .B2(n12475), 
        .C1(n12474), .C2(n12473), .ZN(P1_U3354) );
  XNOR2_X1 U14984 ( .A(n12480), .B(n12479), .ZN(n12481) );
  NAND2_X1 U14985 ( .A1(n12481), .A2(n14515), .ZN(n12484) );
  AOI22_X1 U14986 ( .A1(n14497), .A2(n15303), .B1(n12482), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n12483) );
  OAI211_X1 U14987 ( .C1(n15306), .C2(n14524), .A(n12484), .B(n12483), .ZN(
        P1_U3237) );
  OAI22_X1 U14988 ( .A1(n12487), .A2(n12486), .B1(n12485), .B2(n15280), .ZN(
        n12490) );
  NOR2_X1 U14989 ( .A1(n6538), .A2(n12488), .ZN(n12489) );
  AOI211_X1 U14990 ( .C1(n6538), .C2(P1_REG2_REG_29__SCAN_IN), .A(n12490), .B(
        n12489), .ZN(n12493) );
  NAND2_X1 U14991 ( .A1(n12491), .A2(n14752), .ZN(n12492) );
  OAI211_X1 U14992 ( .C1(n12494), .C2(n15265), .A(n12493), .B(n12492), .ZN(
        n12495) );
  AOI21_X1 U14993 ( .B1(n12496), .B2(n14905), .A(n12495), .ZN(n12497) );
  OAI21_X1 U14994 ( .B1(n12498), .B2(n14953), .A(n12497), .ZN(P1_U3356) );
  NAND2_X1 U14995 ( .A1(n13724), .A2(n13895), .ZN(n12499) );
  XNOR2_X1 U14996 ( .A(n14170), .B(n13733), .ZN(n14165) );
  OR2_X1 U14997 ( .A1(n14170), .A2(n13894), .ZN(n12501) );
  XNOR2_X1 U14998 ( .A(n14274), .B(n13893), .ZN(n13864) );
  NAND2_X1 U14999 ( .A1(n14274), .A2(n13893), .ZN(n12502) );
  INV_X1 U15000 ( .A(n14107), .ZN(n13743) );
  XNOR2_X1 U15001 ( .A(n14268), .B(n13743), .ZN(n14130) );
  NAND2_X1 U15002 ( .A1(n14268), .A2(n14107), .ZN(n12503) );
  XNOR2_X1 U15003 ( .A(n14262), .B(n13892), .ZN(n14119) );
  OR2_X1 U15004 ( .A1(n14262), .A2(n13892), .ZN(n12505) );
  AND2_X1 U15005 ( .A1(n14252), .A2(n14057), .ZN(n12506) );
  OR2_X1 U15006 ( .A1(n14252), .A2(n14057), .ZN(n12507) );
  INV_X1 U15007 ( .A(n14081), .ZN(n13600) );
  XNOR2_X1 U15008 ( .A(n14246), .B(n13600), .ZN(n13844) );
  INV_X1 U15009 ( .A(n14044), .ZN(n12508) );
  XNOR2_X1 U15010 ( .A(n14034), .B(n13597), .ZN(n14029) );
  NAND2_X1 U15011 ( .A1(n14049), .A2(n14058), .ZN(n14027) );
  AND2_X1 U15012 ( .A1(n14029), .A2(n14027), .ZN(n12509) );
  XNOR2_X1 U15013 ( .A(n14230), .B(n13998), .ZN(n14005) );
  INV_X1 U15014 ( .A(n14005), .ZN(n14012) );
  OR2_X1 U15015 ( .A1(n14034), .A2(n14041), .ZN(n14009) );
  AND2_X1 U15016 ( .A1(n14012), .A2(n14009), .ZN(n12510) );
  NAND2_X1 U15017 ( .A1(n14230), .A2(n13998), .ZN(n12511) );
  OR2_X1 U15018 ( .A1(n14225), .A2(n14007), .ZN(n12513) );
  AND2_X1 U15019 ( .A1(n14225), .A2(n14007), .ZN(n12512) );
  NAND2_X1 U15020 ( .A1(n14220), .A2(n13999), .ZN(n12514) );
  INV_X1 U15021 ( .A(n13959), .ZN(n13970) );
  INV_X1 U15022 ( .A(n12515), .ZN(n12516) );
  NAND2_X1 U15023 ( .A1(n13954), .A2(n12516), .ZN(n12519) );
  NAND2_X1 U15024 ( .A1(n14352), .A2(n13785), .ZN(n12518) );
  NAND2_X1 U15025 ( .A1(n9663), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12517) );
  INV_X1 U15026 ( .A(n14058), .ZN(n14024) );
  INV_X1 U15027 ( .A(n13895), .ZN(n12521) );
  NAND2_X1 U15028 ( .A1(n13724), .A2(n12521), .ZN(n12522) );
  INV_X1 U15029 ( .A(n14274), .ZN(n12524) );
  NAND2_X1 U15030 ( .A1(n13742), .A2(n14107), .ZN(n12525) );
  INV_X1 U15031 ( .A(n13892), .ZN(n14091) );
  NAND2_X1 U15032 ( .A1(n14257), .A2(n13607), .ZN(n14077) );
  OR2_X1 U15033 ( .A1(n14257), .A2(n13607), .ZN(n12527) );
  NAND2_X1 U15034 ( .A1(n14077), .A2(n12527), .ZN(n14089) );
  INV_X1 U15035 ( .A(n14077), .ZN(n12528) );
  XNOR2_X1 U15036 ( .A(n14252), .B(n14057), .ZN(n14076) );
  INV_X1 U15037 ( .A(n14252), .ZN(n14075) );
  NAND2_X1 U15038 ( .A1(n14064), .A2(n14081), .ZN(n12529) );
  NOR2_X1 U15039 ( .A1(n14034), .A2(n13597), .ZN(n12530) );
  INV_X1 U15040 ( .A(n13998), .ZN(n14025) );
  NAND2_X1 U15041 ( .A1(n14230), .A2(n14025), .ZN(n13995) );
  XNOR2_X1 U15042 ( .A(n14225), .B(n14007), .ZN(n13994) );
  INV_X1 U15043 ( .A(n14007), .ZN(n13977) );
  NAND2_X1 U15044 ( .A1(n14225), .A2(n13977), .ZN(n12531) );
  OR2_X1 U15045 ( .A1(n14220), .A2(n13782), .ZN(n13843) );
  NAND2_X1 U15046 ( .A1(n13975), .A2(n13843), .ZN(n12532) );
  NAND2_X1 U15047 ( .A1(n14220), .A2(n13782), .ZN(n13842) );
  NAND2_X1 U15048 ( .A1(n14211), .A2(n13978), .ZN(n12533) );
  AOI211_X1 U15049 ( .C1(n13953), .C2(n13961), .A(n14162), .B(n13872), .ZN(
        n12541) );
  NAND3_X1 U15050 ( .A1(n13953), .A2(n13961), .A3(n14180), .ZN(n12538) );
  AOI21_X1 U15051 ( .B1(n13881), .B2(P2_B_REG_SCAN_IN), .A(n14094), .ZN(n13934) );
  INV_X1 U15052 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n13939) );
  NAND2_X1 U15053 ( .A1(n9974), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n12535) );
  NAND2_X1 U15054 ( .A1(n13788), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n12534) );
  OAI211_X1 U15055 ( .C1(n12536), .C2(n13939), .A(n12535), .B(n12534), .ZN(
        n13889) );
  AOI22_X1 U15056 ( .A1(n13961), .A2(n14106), .B1(n13934), .B2(n13889), .ZN(
        n12537) );
  OAI21_X1 U15057 ( .B1(n12539), .B2(n12538), .A(n12537), .ZN(n12540) );
  NAND2_X1 U15058 ( .A1(n6653), .A2(n14135), .ZN(n12549) );
  NAND2_X1 U15059 ( .A1(n14112), .A2(n14098), .ZN(n14095) );
  INV_X1 U15060 ( .A(n14049), .ZN(n14241) );
  INV_X1 U15061 ( .A(n14034), .ZN(n14235) );
  INV_X1 U15062 ( .A(n14220), .ZN(n13781) );
  AND2_X2 U15063 ( .A1(n13988), .A2(n13781), .ZN(n13973) );
  INV_X1 U15064 ( .A(n14203), .ZN(n13798) );
  NOR2_X1 U15065 ( .A1(n13798), .A2(n14188), .ZN(n12547) );
  OAI22_X1 U15066 ( .A1(n12545), .A2(n14146), .B1(n12544), .B2(n14135), .ZN(
        n12546) );
  AOI211_X1 U15067 ( .C1(n14202), .C2(n14194), .A(n12547), .B(n12546), .ZN(
        n12548) );
  OAI211_X1 U15068 ( .C1(n14205), .C2(n14191), .A(n12549), .B(n12548), .ZN(
        P2_U3236) );
  NOR3_X1 U15069 ( .A1(n12591), .A2(n12550), .A3(n12613), .ZN(n12575) );
  NOR3_X1 U15070 ( .A1(n10396), .A2(n12576), .A3(n12613), .ZN(n12574) );
  INV_X1 U15071 ( .A(n12551), .ZN(n12552) );
  NAND2_X1 U15072 ( .A1(n12554), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12555) );
  INV_X1 U15073 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12557) );
  XNOR2_X1 U15074 ( .A(n12557), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12558) );
  NAND2_X1 U15075 ( .A1(n13481), .A2(n8470), .ZN(n12561) );
  INV_X1 U15076 ( .A(SI_31_), .ZN(n13476) );
  OR2_X1 U15077 ( .A1(n12569), .A2(n13476), .ZN(n12560) );
  INV_X1 U15078 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n13110) );
  OR2_X1 U15079 ( .A1(n6535), .A2(n13110), .ZN(n12566) );
  INV_X1 U15080 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13330) );
  OR2_X1 U15081 ( .A1(n12562), .A2(n13330), .ZN(n12565) );
  INV_X1 U15082 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13394) );
  OR2_X1 U15083 ( .A1(n12563), .A2(n13394), .ZN(n12564) );
  XNOR2_X1 U15084 ( .A(n12568), .B(n6731), .ZN(n12769) );
  NAND2_X1 U15085 ( .A1(n12769), .A2(n8470), .ZN(n12571) );
  OR2_X1 U15086 ( .A1(n12569), .A2(n15606), .ZN(n12570) );
  NAND2_X1 U15087 ( .A1(n13395), .A2(n12584), .ZN(n12572) );
  AND2_X1 U15088 ( .A1(n13395), .A2(n13108), .ZN(n12578) );
  NOR2_X1 U15089 ( .A1(n12583), .A2(n12578), .ZN(n12573) );
  INV_X1 U15090 ( .A(n12576), .ZN(n12963) );
  NOR3_X1 U15091 ( .A1(n12577), .A2(n12579), .A3(n12963), .ZN(n12582) );
  INV_X1 U15092 ( .A(n12578), .ZN(n12580) );
  NOR2_X1 U15093 ( .A1(n12580), .A2(n12579), .ZN(n12581) );
  AOI211_X1 U15094 ( .C1(n12613), .C2(n12583), .A(n12582), .B(n12581), .ZN(
        n12589) );
  NAND2_X1 U15095 ( .A1(n12587), .A2(n13108), .ZN(n12586) );
  OR2_X1 U15096 ( .A1(n13395), .A2(n12584), .ZN(n12585) );
  NAND2_X1 U15097 ( .A1(n12586), .A2(n12585), .ZN(n12592) );
  NAND2_X1 U15098 ( .A1(n12592), .A2(n12587), .ZN(n12756) );
  INV_X1 U15099 ( .A(n12756), .ZN(n12588) );
  OR2_X1 U15100 ( .A1(n12589), .A2(n12588), .ZN(n12590) );
  INV_X1 U15101 ( .A(n12592), .ZN(n12757) );
  XNOR2_X1 U15102 ( .A(n13432), .B(n13243), .ZN(n13230) );
  AND2_X1 U15103 ( .A1(n12693), .A2(n12694), .ZN(n12691) );
  NAND2_X1 U15104 ( .A1(n8561), .A2(n12594), .ZN(n12670) );
  INV_X1 U15105 ( .A(n12670), .ZN(n12603) );
  INV_X1 U15106 ( .A(n12641), .ZN(n12601) );
  NAND3_X1 U15107 ( .A1(n12597), .A2(n12596), .A3(n12595), .ZN(n12600) );
  NAND3_X1 U15108 ( .A1(n11265), .A2(n15489), .A3(n12598), .ZN(n12599) );
  NOR4_X1 U15109 ( .A1(n12662), .A2(n12601), .A3(n12600), .A4(n12599), .ZN(
        n12602) );
  NAND4_X1 U15110 ( .A1(n12679), .A2(n12656), .A3(n12603), .A4(n12602), .ZN(
        n12604) );
  NOR4_X1 U15111 ( .A1(n12695), .A2(n13303), .A3(n12605), .A4(n12604), .ZN(
        n12606) );
  NAND4_X1 U15112 ( .A1(n13259), .A2(n13281), .A3(n12606), .A4(n13270), .ZN(
        n12607) );
  NOR4_X1 U15113 ( .A1(n13218), .A2(n13230), .A3(n13254), .A4(n12607), .ZN(
        n12609) );
  INV_X1 U15114 ( .A(n12608), .ZN(n12729) );
  XNOR2_X1 U15115 ( .A(n13417), .B(n13222), .ZN(n13205) );
  NOR4_X1 U15116 ( .A1(n12611), .A2(n12745), .A3(n13125), .A4(n12610), .ZN(
        n12612) );
  NAND3_X1 U15117 ( .A1(n12755), .A2(n12757), .A3(n12612), .ZN(n12614) );
  XNOR2_X1 U15118 ( .A(n12614), .B(n12613), .ZN(n12616) );
  NOR2_X1 U15119 ( .A1(n12616), .A2(n12615), .ZN(n12762) );
  NAND2_X1 U15120 ( .A1(n12618), .A2(n12617), .ZN(n12619) );
  AND2_X1 U15121 ( .A1(n12619), .A2(n12620), .ZN(n12623) );
  OAI21_X1 U15122 ( .B1(n12731), .B2(n12621), .A(n12620), .ZN(n12622) );
  XNOR2_X1 U15123 ( .A(n12624), .B(n12752), .ZN(n12625) );
  OAI21_X1 U15124 ( .B1(n11276), .B2(n12626), .A(n12625), .ZN(n12633) );
  NAND2_X1 U15125 ( .A1(n15502), .A2(n12627), .ZN(n12629) );
  NAND3_X1 U15126 ( .A1(n12629), .A2(n12742), .A3(n12628), .ZN(n12632) );
  NAND3_X1 U15127 ( .A1(n12974), .A2(n15513), .A3(n12742), .ZN(n12630) );
  NAND2_X1 U15128 ( .A1(n15489), .A2(n12630), .ZN(n12631) );
  AOI21_X1 U15129 ( .B1(n12633), .B2(n12632), .A(n12631), .ZN(n12636) );
  AOI21_X1 U15130 ( .B1(n11644), .B2(n8548), .A(n12752), .ZN(n12635) );
  OAI21_X1 U15131 ( .B1(n12636), .B2(n12635), .A(n12634), .ZN(n12640) );
  INV_X1 U15132 ( .A(n12637), .ZN(n12638) );
  NAND2_X1 U15133 ( .A1(n12638), .A2(n12752), .ZN(n12639) );
  NAND2_X1 U15134 ( .A1(n12640), .A2(n12639), .ZN(n12642) );
  OAI211_X1 U15135 ( .C1(n12742), .C2(n8548), .A(n12642), .B(n12641), .ZN(
        n12650) );
  NOR2_X1 U15136 ( .A1(n12973), .A2(n12752), .ZN(n12644) );
  AND2_X1 U15137 ( .A1(n12973), .A2(n12752), .ZN(n12643) );
  MUX2_X1 U15138 ( .A(n12644), .B(n12643), .S(n15472), .Z(n12646) );
  NOR2_X1 U15139 ( .A1(n12646), .A2(n12645), .ZN(n12649) );
  AOI21_X1 U15140 ( .B1(n12658), .B2(n12647), .A(n12742), .ZN(n12648) );
  AOI21_X1 U15141 ( .B1(n12650), .B2(n12649), .A(n12648), .ZN(n12655) );
  INV_X1 U15142 ( .A(n12651), .ZN(n12654) );
  INV_X1 U15143 ( .A(n12652), .ZN(n12653) );
  OAI22_X1 U15144 ( .A1(n12655), .A2(n12654), .B1(n12752), .B2(n12653), .ZN(
        n12657) );
  OAI211_X1 U15145 ( .C1(n12752), .C2(n12658), .A(n12657), .B(n12656), .ZN(
        n12664) );
  INV_X1 U15146 ( .A(n12659), .ZN(n12661) );
  MUX2_X1 U15147 ( .A(n12661), .B(n12660), .S(n12752), .Z(n12663) );
  INV_X1 U15148 ( .A(n12665), .ZN(n12668) );
  INV_X1 U15149 ( .A(n12666), .ZN(n12667) );
  MUX2_X1 U15150 ( .A(n12668), .B(n12667), .S(n12742), .Z(n12669) );
  NOR2_X1 U15151 ( .A1(n12670), .A2(n12669), .ZN(n12683) );
  MUX2_X1 U15152 ( .A(n12672), .B(n12671), .S(n12742), .Z(n12681) );
  INV_X1 U15153 ( .A(n12673), .ZN(n12676) );
  INV_X1 U15154 ( .A(n12674), .ZN(n12675) );
  MUX2_X1 U15155 ( .A(n12676), .B(n12675), .S(n12742), .Z(n12677) );
  INV_X1 U15156 ( .A(n12677), .ZN(n12678) );
  OAI211_X1 U15157 ( .C1(n12681), .C2(n12680), .A(n12679), .B(n12678), .ZN(
        n12682) );
  NAND2_X1 U15158 ( .A1(n12689), .A2(n12684), .ZN(n12687) );
  NAND2_X1 U15159 ( .A1(n12688), .A2(n12685), .ZN(n12686) );
  MUX2_X1 U15160 ( .A(n12687), .B(n12686), .S(n12752), .Z(n12692) );
  MUX2_X1 U15161 ( .A(n12689), .B(n12688), .S(n12742), .Z(n12690) );
  MUX2_X1 U15162 ( .A(n12694), .B(n12693), .S(n12742), .Z(n12696) );
  INV_X1 U15163 ( .A(n12697), .ZN(n12699) );
  MUX2_X1 U15164 ( .A(n12699), .B(n12698), .S(n12752), .Z(n12700) );
  OAI21_X1 U15165 ( .B1(n13373), .B2(n12955), .A(n12701), .ZN(n12702) );
  NAND2_X1 U15166 ( .A1(n12702), .A2(n12742), .ZN(n12704) );
  INV_X1 U15167 ( .A(n12706), .ZN(n12703) );
  AOI21_X1 U15168 ( .B1(n12706), .B2(n12705), .A(n12742), .ZN(n12708) );
  NAND2_X1 U15169 ( .A1(n13283), .A2(n12752), .ZN(n12707) );
  OAI22_X1 U15170 ( .A1(n12709), .A2(n12708), .B1(n13373), .B2(n12707), .ZN(
        n12710) );
  AND3_X1 U15171 ( .A1(n12710), .A2(n13259), .A3(n7348), .ZN(n12721) );
  INV_X1 U15172 ( .A(n12711), .ZN(n12712) );
  NAND2_X1 U15173 ( .A1(n12714), .A2(n12712), .ZN(n12713) );
  NAND3_X1 U15174 ( .A1(n6591), .A2(n13228), .A3(n12713), .ZN(n12717) );
  OAI211_X1 U15175 ( .C1(n13254), .C2(n12715), .A(n12714), .B(n12718), .ZN(
        n12716) );
  MUX2_X1 U15176 ( .A(n12717), .B(n12716), .S(n12742), .Z(n12720) );
  INV_X1 U15177 ( .A(n13218), .ZN(n13220) );
  MUX2_X1 U15178 ( .A(n6591), .B(n12718), .S(n12752), .Z(n12719) );
  OAI211_X1 U15179 ( .C1(n12721), .C2(n12720), .A(n13220), .B(n12719), .ZN(
        n12725) );
  MUX2_X1 U15180 ( .A(n12723), .B(n12722), .S(n12752), .Z(n12724) );
  MUX2_X1 U15181 ( .A(n12726), .B(n6610), .S(n12742), .Z(n12727) );
  MUX2_X1 U15182 ( .A(n12729), .B(n12728), .S(n12752), .Z(n12730) );
  MUX2_X1 U15183 ( .A(n13168), .B(n12742), .S(n13339), .Z(n12733) );
  NAND2_X1 U15184 ( .A1(n13168), .A2(n12742), .ZN(n12732) );
  NAND2_X1 U15185 ( .A1(n12733), .A2(n12732), .ZN(n12734) );
  OAI211_X1 U15186 ( .C1(n12737), .C2(n12736), .A(n12735), .B(n12734), .ZN(
        n12741) );
  MUX2_X1 U15187 ( .A(n12739), .B(n12738), .S(n12742), .Z(n12740) );
  NAND2_X1 U15188 ( .A1(n12964), .A2(n12742), .ZN(n12743) );
  NOR2_X1 U15189 ( .A1(n13333), .A2(n12743), .ZN(n12744) );
  NAND3_X1 U15190 ( .A1(n12747), .A2(n12752), .A3(n12746), .ZN(n12749) );
  NAND2_X1 U15191 ( .A1(n12749), .A2(n12748), .ZN(n12750) );
  INV_X1 U15192 ( .A(n13108), .ZN(n12962) );
  NAND3_X1 U15193 ( .A1(n12764), .A2(n12763), .A3(n13489), .ZN(n12765) );
  OAI211_X1 U15194 ( .C1(n12766), .C2(n12768), .A(n12765), .B(P3_B_REG_SCAN_IN), .ZN(n12767) );
  INV_X1 U15195 ( .A(n12769), .ZN(n12771) );
  OAI222_X1 U15196 ( .A1(n13495), .A2(n12771), .B1(n12770), .B2(P3_U3151), 
        .C1(n15606), .C2(n13487), .ZN(P3_U3265) );
  AND2_X1 U15197 ( .A1(n12863), .A2(n12772), .ZN(n12930) );
  XOR2_X1 U15198 ( .A(n12773), .B(n12971), .Z(n12929) );
  NAND2_X1 U15199 ( .A1(n12930), .A2(n12929), .ZN(n12928) );
  NAND2_X1 U15200 ( .A1(n12928), .A2(n12774), .ZN(n12830) );
  XNOR2_X1 U15201 ( .A(n12830), .B(n12829), .ZN(n12775) );
  NAND2_X1 U15202 ( .A1(n12775), .A2(n7163), .ZN(n12783) );
  AOI21_X1 U15203 ( .B1(n12958), .B2(n12777), .A(n12776), .ZN(n12782) );
  AOI22_X1 U15204 ( .A1(n12951), .A2(n12971), .B1(n12933), .B2(n12969), .ZN(
        n12781) );
  INV_X1 U15205 ( .A(n12778), .ZN(n12779) );
  NAND2_X1 U15206 ( .A1(n12952), .A2(n12779), .ZN(n12780) );
  NAND4_X1 U15207 ( .A1(n12783), .A2(n12782), .A3(n12781), .A4(n12780), .ZN(
        P3_U3153) );
  XOR2_X1 U15208 ( .A(n12785), .B(n12784), .Z(n12790) );
  AOI22_X1 U15209 ( .A1(n12933), .A2(n13128), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12787) );
  NAND2_X1 U15210 ( .A1(n12951), .A2(n13129), .ZN(n12786) );
  OAI211_X1 U15211 ( .C1(n12944), .C2(n13132), .A(n12787), .B(n12786), .ZN(
        n12788) );
  AOI21_X1 U15212 ( .B1(n13333), .B2(n12958), .A(n12788), .ZN(n12789) );
  OAI21_X1 U15213 ( .B1(n12790), .B2(n12960), .A(n12789), .ZN(P3_U3154) );
  INV_X1 U15214 ( .A(n12791), .ZN(n12792) );
  XNOR2_X1 U15215 ( .A(n12885), .B(n12913), .ZN(n12798) );
  AOI22_X1 U15216 ( .A1(n12965), .A2(n12933), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12795) );
  NAND2_X1 U15217 ( .A1(n13190), .A2(n12952), .ZN(n12794) );
  OAI211_X1 U15218 ( .C1(n13180), .C2(n12922), .A(n12795), .B(n12794), .ZN(
        n12796) );
  AOI21_X1 U15219 ( .B1(n13189), .B2(n12958), .A(n12796), .ZN(n12797) );
  OAI21_X1 U15220 ( .B1(n12798), .B2(n12960), .A(n12797), .ZN(P3_U3156) );
  AND2_X1 U15221 ( .A1(n12799), .A2(n12800), .ZN(n12803) );
  OAI211_X1 U15222 ( .C1(n12803), .C2(n12802), .A(n7163), .B(n12801), .ZN(
        n12810) );
  AOI21_X1 U15223 ( .B1(n12958), .B2(n12805), .A(n12804), .ZN(n12809) );
  AOI22_X1 U15224 ( .A1(n12951), .A2(n12968), .B1(n12933), .B2(n13314), .ZN(
        n12808) );
  NAND2_X1 U15225 ( .A1(n12952), .A2(n12806), .ZN(n12807) );
  NAND4_X1 U15226 ( .A1(n12810), .A2(n12809), .A3(n12808), .A4(n12807), .ZN(
        P3_U3157) );
  AND2_X1 U15227 ( .A1(n12812), .A2(n12811), .ZN(n12815) );
  OAI211_X1 U15228 ( .C1(n12815), .C2(n12814), .A(n7163), .B(n12813), .ZN(
        n12820) );
  AOI21_X1 U15229 ( .B1(n12958), .B2(n7378), .A(n12816), .ZN(n12819) );
  AOI22_X1 U15230 ( .A1(n12951), .A2(n15506), .B1(n12933), .B2(n12973), .ZN(
        n12818) );
  NAND2_X1 U15231 ( .A1(n12952), .A2(n15768), .ZN(n12817) );
  NAND4_X1 U15232 ( .A1(n12820), .A2(n12819), .A3(n12818), .A4(n12817), .ZN(
        P3_U3158) );
  OAI211_X1 U15233 ( .C1(n12823), .C2(n12822), .A(n12821), .B(n7163), .ZN(
        n12828) );
  AOI21_X1 U15234 ( .B1(n12933), .B2(n13207), .A(n12824), .ZN(n12825) );
  OAI21_X1 U15235 ( .B1(n13232), .B2(n12922), .A(n12825), .ZN(n12826) );
  AOI21_X1 U15236 ( .B1(n13237), .B2(n12952), .A(n12826), .ZN(n12827) );
  OAI211_X1 U15237 ( .C1(n12926), .C2(n13432), .A(n12828), .B(n12827), .ZN(
        P3_U3159) );
  MUX2_X1 U15238 ( .A(n12830), .B(n12970), .S(n12829), .Z(n12832) );
  XNOR2_X1 U15239 ( .A(n12832), .B(n12831), .ZN(n12833) );
  NAND2_X1 U15240 ( .A1(n12833), .A2(n7163), .ZN(n12839) );
  AOI21_X1 U15241 ( .B1(n12958), .B2(n7141), .A(n12834), .ZN(n12838) );
  AOI22_X1 U15242 ( .A1(n12951), .A2(n12970), .B1(n12933), .B2(n12968), .ZN(
        n12837) );
  NAND2_X1 U15243 ( .A1(n12952), .A2(n12835), .ZN(n12836) );
  NAND4_X1 U15244 ( .A1(n12839), .A2(n12838), .A3(n12837), .A4(n12836), .ZN(
        P3_U3161) );
  XOR2_X1 U15245 ( .A(n12841), .B(n12840), .Z(n12846) );
  AOI22_X1 U15246 ( .A1(n12951), .A2(n13207), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12843) );
  NAND2_X1 U15247 ( .A1(n12952), .A2(n13211), .ZN(n12842) );
  OAI211_X1 U15248 ( .C1(n13180), .C2(n12956), .A(n12843), .B(n12842), .ZN(
        n12844) );
  AOI21_X1 U15249 ( .B1(n13417), .B2(n12958), .A(n12844), .ZN(n12845) );
  OAI21_X1 U15250 ( .B1(n12846), .B2(n12960), .A(n12845), .ZN(P3_U3163) );
  XOR2_X1 U15251 ( .A(n12848), .B(n12847), .Z(n12853) );
  NAND2_X1 U15252 ( .A1(n12965), .A2(n12951), .ZN(n12850) );
  AOI22_X1 U15253 ( .A1(n12933), .A2(n13129), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12849) );
  OAI211_X1 U15254 ( .C1(n12944), .C2(n13161), .A(n12850), .B(n12849), .ZN(
        n12851) );
  AOI21_X1 U15255 ( .B1(n13339), .B2(n12958), .A(n12851), .ZN(n12852) );
  OAI21_X1 U15256 ( .B1(n12853), .B2(n12960), .A(n12852), .ZN(P3_U3165) );
  XNOR2_X1 U15257 ( .A(n12854), .B(n12955), .ZN(n12855) );
  XNOR2_X1 U15258 ( .A(n12856), .B(n12855), .ZN(n12862) );
  AND2_X1 U15259 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13058) );
  AOI21_X1 U15260 ( .B1(n12933), .B2(n12857), .A(n13058), .ZN(n12859) );
  NAND2_X1 U15261 ( .A1(n12952), .A2(n13274), .ZN(n12858) );
  OAI211_X1 U15262 ( .C1(n13272), .C2(n12922), .A(n12859), .B(n12858), .ZN(
        n12860) );
  AOI21_X1 U15263 ( .B1(n13373), .B2(n12958), .A(n12860), .ZN(n12861) );
  OAI21_X1 U15264 ( .B1(n12862), .B2(n12960), .A(n12861), .ZN(P3_U3166) );
  OAI21_X1 U15265 ( .B1(n12865), .B2(n12864), .A(n12863), .ZN(n12866) );
  NAND2_X1 U15266 ( .A1(n12866), .A2(n7163), .ZN(n12873) );
  AOI21_X1 U15267 ( .B1(n12958), .B2(n12868), .A(n12867), .ZN(n12872) );
  AOI22_X1 U15268 ( .A1(n12951), .A2(n12973), .B1(n12933), .B2(n12971), .ZN(
        n12871) );
  NAND2_X1 U15269 ( .A1(n12952), .A2(n12869), .ZN(n12870) );
  NAND4_X1 U15270 ( .A1(n12873), .A2(n12872), .A3(n12871), .A4(n12870), .ZN(
        P3_U3167) );
  INV_X1 U15271 ( .A(n13436), .ZN(n12882) );
  AOI21_X1 U15272 ( .B1(n12875), .B2(n12874), .A(n12960), .ZN(n12877) );
  NAND2_X1 U15273 ( .A1(n12877), .A2(n12876), .ZN(n12881) );
  AND2_X1 U15274 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13070) );
  AOI21_X1 U15275 ( .B1(n12933), .B2(n13261), .A(n13070), .ZN(n12878) );
  OAI21_X1 U15276 ( .B1(n12955), .B2(n12922), .A(n12878), .ZN(n12879) );
  AOI21_X1 U15277 ( .B1(n13264), .B2(n12952), .A(n12879), .ZN(n12880) );
  OAI211_X1 U15278 ( .C1(n12882), .C2(n12926), .A(n12881), .B(n12880), .ZN(
        P3_U3168) );
  AOI22_X1 U15279 ( .A1(n12933), .A2(n13168), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12888) );
  NAND2_X1 U15280 ( .A1(n13173), .A2(n12952), .ZN(n12887) );
  OAI211_X1 U15281 ( .C1(n12913), .C2(n12922), .A(n12888), .B(n12887), .ZN(
        n12889) );
  AOI21_X1 U15282 ( .B1(n8571), .B2(n12958), .A(n12889), .ZN(n12890) );
  INV_X1 U15283 ( .A(n12799), .ZN(n12891) );
  AOI21_X1 U15284 ( .B1(n12893), .B2(n12892), .A(n12891), .ZN(n12894) );
  OR2_X1 U15285 ( .A1(n12894), .A2(n12960), .ZN(n12901) );
  AOI21_X1 U15286 ( .B1(n12958), .B2(n12896), .A(n12895), .ZN(n12900) );
  AOI22_X1 U15287 ( .A1(n12951), .A2(n12969), .B1(n12933), .B2(n12967), .ZN(
        n12899) );
  NAND2_X1 U15288 ( .A1(n12952), .A2(n12897), .ZN(n12898) );
  NAND4_X1 U15289 ( .A1(n12901), .A2(n12900), .A3(n12899), .A4(n12898), .ZN(
        P3_U3171) );
  AOI21_X1 U15290 ( .B1(n12903), .B2(n12902), .A(n6627), .ZN(n12909) );
  AOI22_X1 U15291 ( .A1(n13222), .A2(n12933), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12905) );
  NAND2_X1 U15292 ( .A1(n12952), .A2(n13225), .ZN(n12904) );
  OAI211_X1 U15293 ( .C1(n12906), .C2(n12922), .A(n12905), .B(n12904), .ZN(
        n12907) );
  AOI21_X1 U15294 ( .B1(n13423), .B2(n12958), .A(n12907), .ZN(n12908) );
  OAI21_X1 U15295 ( .B1(n12909), .B2(n12960), .A(n12908), .ZN(P3_U3173) );
  XNOR2_X1 U15296 ( .A(n12910), .B(n13208), .ZN(n12916) );
  AOI22_X1 U15297 ( .A1(n13222), .A2(n12951), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12912) );
  NAND2_X1 U15298 ( .A1(n12952), .A2(n13201), .ZN(n12911) );
  OAI211_X1 U15299 ( .C1(n12913), .C2(n12956), .A(n12912), .B(n12911), .ZN(
        n12914) );
  AOI21_X1 U15300 ( .B1(n13411), .B2(n12958), .A(n12914), .ZN(n12915) );
  OAI21_X1 U15301 ( .B1(n12916), .B2(n12960), .A(n12915), .ZN(P3_U3175) );
  INV_X1 U15302 ( .A(n13247), .ZN(n12927) );
  OAI211_X1 U15303 ( .C1(n12919), .C2(n12918), .A(n12917), .B(n7163), .ZN(
        n12925) );
  AND2_X1 U15304 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13085) );
  AOI21_X1 U15305 ( .B1(n12933), .B2(n13243), .A(n13085), .ZN(n12921) );
  OAI21_X1 U15306 ( .B1(n13273), .B2(n12922), .A(n12921), .ZN(n12923) );
  AOI21_X1 U15307 ( .B1(n13248), .B2(n12952), .A(n12923), .ZN(n12924) );
  OAI211_X1 U15308 ( .C1(n12927), .C2(n12926), .A(n12925), .B(n12924), .ZN(
        P3_U3178) );
  OAI211_X1 U15309 ( .C1(n12930), .C2(n12929), .A(n12928), .B(n7163), .ZN(
        n12938) );
  AOI21_X1 U15310 ( .B1(n12958), .B2(n12932), .A(n12931), .ZN(n12937) );
  AOI22_X1 U15311 ( .A1(n12951), .A2(n12972), .B1(n12933), .B2(n12970), .ZN(
        n12936) );
  NAND2_X1 U15312 ( .A1(n12952), .A2(n12934), .ZN(n12935) );
  NAND4_X1 U15313 ( .A1(n12938), .A2(n12937), .A3(n12936), .A4(n12935), .ZN(
        P3_U3179) );
  XOR2_X1 U15314 ( .A(n12940), .B(n12939), .Z(n12947) );
  OAI22_X1 U15315 ( .A1(n12956), .A2(n13143), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12941), .ZN(n12942) );
  AOI21_X1 U15316 ( .B1(n12951), .B2(n13168), .A(n12942), .ZN(n12943) );
  OAI21_X1 U15317 ( .B1(n12944), .B2(n13144), .A(n12943), .ZN(n12945) );
  AOI21_X1 U15318 ( .B1(n8574), .B2(n12958), .A(n12945), .ZN(n12946) );
  OAI21_X1 U15319 ( .B1(n12947), .B2(n12960), .A(n12946), .ZN(P3_U3180) );
  XNOR2_X1 U15320 ( .A(n12948), .B(n13272), .ZN(n12949) );
  XNOR2_X1 U15321 ( .A(n12950), .B(n12949), .ZN(n12961) );
  AND2_X1 U15322 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13033) );
  AOI21_X1 U15323 ( .B1(n12951), .B2(n13305), .A(n13033), .ZN(n12954) );
  NAND2_X1 U15324 ( .A1(n12952), .A2(n13286), .ZN(n12953) );
  OAI211_X1 U15325 ( .C1(n12956), .C2(n12955), .A(n12954), .B(n12953), .ZN(
        n12957) );
  AOI21_X1 U15326 ( .B1(n13446), .B2(n12958), .A(n12957), .ZN(n12959) );
  OAI21_X1 U15327 ( .B1(n12961), .B2(n12960), .A(n12959), .ZN(P3_U3181) );
  MUX2_X1 U15328 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12962), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15329 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12963), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15330 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13128), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15331 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12964), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15332 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13168), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15333 ( .A(n12965), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12966), .Z(
        P3_U3515) );
  MUX2_X1 U15334 ( .A(n13198), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12966), .Z(
        P3_U3514) );
  MUX2_X1 U15335 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13208), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15336 ( .A(n13222), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12966), .Z(
        P3_U3512) );
  MUX2_X1 U15337 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13207), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15338 ( .A(n13243), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12966), .Z(
        P3_U3510) );
  MUX2_X1 U15339 ( .A(n13261), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12966), .Z(
        P3_U3509) );
  MUX2_X1 U15340 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13283), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15341 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13295), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15342 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13306), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15343 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13314), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15344 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12967), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15345 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12968), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15346 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12969), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15347 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12970), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15348 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12971), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15349 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12972), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15350 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12973), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15351 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15506), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15352 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12974), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15353 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15505), .S(P3_U3897), .Z(
        P3_U3491) );
  XOR2_X1 U15354 ( .A(n12977), .B(n12976), .Z(n12990) );
  OAI21_X1 U15355 ( .B1(n6699), .B2(P3_REG2_REG_11__SCAN_IN), .A(n12978), .ZN(
        n12988) );
  INV_X1 U15356 ( .A(n12979), .ZN(n12980) );
  AOI21_X1 U15357 ( .B1(n15467), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12980), 
        .ZN(n12981) );
  OAI21_X1 U15358 ( .B1(n13088), .B2(n12982), .A(n12981), .ZN(n12987) );
  AOI21_X1 U15359 ( .B1(n15739), .B2(n12984), .A(n12983), .ZN(n12985) );
  NOR2_X1 U15360 ( .A1(n12985), .A2(n13046), .ZN(n12986) );
  AOI211_X1 U15361 ( .C1(n13090), .C2(n12988), .A(n12987), .B(n12986), .ZN(
        n12989) );
  OAI21_X1 U15362 ( .B1(n12990), .B2(n13030), .A(n12989), .ZN(P3_U3193) );
  AOI21_X1 U15363 ( .B1(n15767), .B2(n12992), .A(n12991), .ZN(n13005) );
  OAI21_X1 U15364 ( .B1(n12995), .B2(n12994), .A(n12993), .ZN(n13000) );
  NAND2_X1 U15365 ( .A1(n15467), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n12996) );
  OAI211_X1 U15366 ( .C1(n13088), .C2(n12998), .A(n12997), .B(n12996), .ZN(
        n12999) );
  AOI21_X1 U15367 ( .B1(n13000), .B2(n13095), .A(n12999), .ZN(n13004) );
  OAI21_X1 U15368 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n13001), .A(n13017), 
        .ZN(n13002) );
  NAND2_X1 U15369 ( .A1(n13002), .A2(n13090), .ZN(n13003) );
  OAI211_X1 U15370 ( .C1(n13005), .C2(n13046), .A(n13004), .B(n13003), .ZN(
        P3_U3195) );
  INV_X1 U15371 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15175) );
  OAI21_X1 U15372 ( .B1(n13007), .B2(n15175), .A(n13006), .ZN(n13012) );
  AOI211_X1 U15373 ( .C1(n13010), .C2(n13009), .A(n13030), .B(n13008), .ZN(
        n13011) );
  AOI211_X1 U15374 ( .C1(n13014), .C2(n13013), .A(n13012), .B(n13011), .ZN(
        n13027) );
  AND3_X1 U15375 ( .A1(n13017), .A2(n13016), .A3(n13015), .ZN(n13018) );
  OAI21_X1 U15376 ( .B1(n13019), .B2(n13018), .A(n13090), .ZN(n13026) );
  INV_X1 U15377 ( .A(n13020), .ZN(n13024) );
  NOR3_X1 U15378 ( .A1(n12991), .A2(n13022), .A3(n13021), .ZN(n13023) );
  OAI21_X1 U15379 ( .B1(n13024), .B2(n13023), .A(n13100), .ZN(n13025) );
  NAND3_X1 U15380 ( .A1(n13027), .A2(n13026), .A3(n13025), .ZN(P3_U3196) );
  INV_X1 U15381 ( .A(n13052), .ZN(n13028) );
  AOI21_X1 U15382 ( .B1(n13285), .B2(n13029), .A(n13028), .ZN(n13043) );
  AOI21_X1 U15383 ( .B1(n13032), .B2(n13031), .A(n13030), .ZN(n13038) );
  AOI21_X1 U15384 ( .B1(n15467), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13033), 
        .ZN(n13034) );
  OAI21_X1 U15385 ( .B1(n13088), .B2(n13035), .A(n13034), .ZN(n13036) );
  AOI21_X1 U15386 ( .B1(n13038), .B2(n13037), .A(n13036), .ZN(n13042) );
  OAI21_X1 U15387 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n13039), .A(n13045), 
        .ZN(n13040) );
  NAND2_X1 U15388 ( .A1(n13040), .A2(n13100), .ZN(n13041) );
  OAI211_X1 U15389 ( .C1(n13043), .C2(n13077), .A(n13042), .B(n13041), .ZN(
        P3_U3197) );
  NAND3_X1 U15390 ( .A1(n13045), .A2(n6717), .A3(n13044), .ZN(n13047) );
  AOI21_X1 U15391 ( .B1(n13048), .B2(n13047), .A(n13046), .ZN(n13064) );
  INV_X1 U15392 ( .A(n13049), .ZN(n13051) );
  NAND3_X1 U15393 ( .A1(n13052), .A2(n13051), .A3(n13050), .ZN(n13053) );
  AOI21_X1 U15394 ( .B1(n13054), .B2(n13053), .A(n13077), .ZN(n13063) );
  OAI211_X1 U15395 ( .C1(n13057), .C2(n13056), .A(n13055), .B(n13095), .ZN(
        n13060) );
  AOI21_X1 U15396 ( .B1(n15467), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n13058), 
        .ZN(n13059) );
  OAI211_X1 U15397 ( .C1(n13088), .C2(n13061), .A(n13060), .B(n13059), .ZN(
        n13062) );
  OR3_X1 U15398 ( .A1(n13064), .A2(n13063), .A3(n13062), .ZN(P3_U3198) );
  INV_X1 U15399 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13263) );
  INV_X1 U15400 ( .A(n13082), .ZN(n13065) );
  AOI21_X1 U15401 ( .B1(n13263), .B2(n13066), .A(n13065), .ZN(n13078) );
  OAI21_X1 U15402 ( .B1(n6551), .B2(P3_REG1_REG_17__SCAN_IN), .A(n13099), .ZN(
        n13075) );
  OAI211_X1 U15403 ( .C1(n13069), .C2(n13068), .A(n13067), .B(n13095), .ZN(
        n13072) );
  AOI21_X1 U15404 ( .B1(n15467), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13070), 
        .ZN(n13071) );
  OAI211_X1 U15405 ( .C1(n13088), .C2(n13073), .A(n13072), .B(n13071), .ZN(
        n13074) );
  AOI21_X1 U15406 ( .B1(n13075), .B2(n13100), .A(n13074), .ZN(n13076) );
  OAI21_X1 U15407 ( .B1(n13078), .B2(n13077), .A(n13076), .ZN(P3_U3199) );
  INV_X1 U15408 ( .A(n13079), .ZN(n13080) );
  NAND3_X1 U15409 ( .A1(n13082), .A2(n13081), .A3(n13080), .ZN(n13083) );
  NAND2_X1 U15410 ( .A1(n13084), .A2(n13083), .ZN(n13091) );
  AOI21_X1 U15411 ( .B1(n15467), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n13085), 
        .ZN(n13086) );
  OAI21_X1 U15412 ( .B1(n13088), .B2(n13087), .A(n13086), .ZN(n13089) );
  AOI21_X1 U15413 ( .B1(n13091), .B2(n13090), .A(n13089), .ZN(n13105) );
  OAI21_X1 U15414 ( .B1(n13094), .B2(n13093), .A(n13092), .ZN(n13096) );
  NAND2_X1 U15415 ( .A1(n13096), .A2(n13095), .ZN(n13104) );
  AND3_X1 U15416 ( .A1(n13099), .A2(n13098), .A3(n13097), .ZN(n13101) );
  OAI21_X1 U15417 ( .B1(n13102), .B2(n13101), .A(n13100), .ZN(n13103) );
  NAND3_X1 U15418 ( .A1(n13105), .A2(n13104), .A3(n13103), .ZN(P3_U3200) );
  NAND2_X1 U15419 ( .A1(n12587), .A2(n6529), .ZN(n13109) );
  NOR2_X1 U15420 ( .A1(n15486), .A2(n13106), .ZN(n13114) );
  NOR2_X1 U15421 ( .A1(n13108), .A2(n13107), .ZN(n13392) );
  OAI21_X1 U15422 ( .B1(n13114), .B2(n13392), .A(n15500), .ZN(n13111) );
  OAI211_X1 U15423 ( .C1(n15500), .C2(n13110), .A(n13109), .B(n13111), .ZN(
        P3_U3202) );
  NAND2_X1 U15424 ( .A1(n13395), .A2(n6529), .ZN(n13112) );
  OAI211_X1 U15425 ( .C1(n15500), .C2(n15807), .A(n13112), .B(n13111), .ZN(
        P3_U3203) );
  NOR2_X1 U15426 ( .A1(n15500), .A2(n15589), .ZN(n13113) );
  AOI211_X1 U15427 ( .C1(n13115), .C2(n13252), .A(n13114), .B(n13113), .ZN(
        n13118) );
  NAND2_X1 U15428 ( .A1(n13116), .A2(n15500), .ZN(n13117) );
  OAI211_X1 U15429 ( .C1(n13119), .C2(n13327), .A(n13118), .B(n13117), .ZN(
        P3_U3204) );
  AOI22_X1 U15430 ( .A1(n8579), .A2(n6529), .B1(n15516), .B2(n13121), .ZN(
        n13122) );
  OAI211_X1 U15431 ( .C1(n13124), .C2(n13327), .A(n13123), .B(n13122), .ZN(
        P3_U3205) );
  INV_X1 U15432 ( .A(n13335), .ZN(n13137) );
  XNOR2_X1 U15433 ( .A(n13127), .B(n13125), .ZN(n13131) );
  AOI22_X1 U15434 ( .A1(n15504), .A2(n13129), .B1(n13128), .B2(n13320), .ZN(
        n13130) );
  NAND2_X1 U15435 ( .A1(n13334), .A2(n15500), .ZN(n13136) );
  OAI22_X1 U15436 ( .A1(n15500), .A2(n13133), .B1(n13132), .B2(n15486), .ZN(
        n13134) );
  AOI21_X1 U15437 ( .B1(n13333), .B2(n6529), .A(n13134), .ZN(n13135) );
  OAI211_X1 U15438 ( .C1(n13137), .C2(n13188), .A(n13136), .B(n13135), .ZN(
        P3_U3206) );
  XNOR2_X1 U15439 ( .A(n13138), .B(n13140), .ZN(n13403) );
  XNOR2_X1 U15440 ( .A(n13141), .B(n13140), .ZN(n13142) );
  NAND2_X1 U15441 ( .A1(n13337), .A2(n15500), .ZN(n13148) );
  OAI22_X1 U15442 ( .A1(n15500), .A2(n13145), .B1(n13144), .B2(n15486), .ZN(
        n13146) );
  AOI21_X1 U15443 ( .B1(n8574), .B2(n6529), .A(n13146), .ZN(n13147) );
  OAI211_X1 U15444 ( .C1(n13403), .C2(n13327), .A(n13148), .B(n13147), .ZN(
        P3_U3207) );
  NAND2_X1 U15445 ( .A1(n13153), .A2(n13150), .ZN(n13151) );
  AOI21_X1 U15446 ( .B1(n13151), .B2(n13159), .A(n15508), .ZN(n13157) );
  NAND2_X1 U15447 ( .A1(n13153), .A2(n13152), .ZN(n13156) );
  OAI22_X1 U15448 ( .A1(n13181), .A2(n15492), .B1(n13154), .B2(n15491), .ZN(
        n13155) );
  AOI21_X1 U15449 ( .B1(n13157), .B2(n13156), .A(n13155), .ZN(n13341) );
  OAI21_X1 U15450 ( .B1(n13160), .B2(n13159), .A(n13158), .ZN(n13340) );
  INV_X1 U15451 ( .A(n13161), .ZN(n13162) );
  AOI22_X1 U15452 ( .A1(n15519), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15516), 
        .B2(n13162), .ZN(n13163) );
  OAI21_X1 U15453 ( .B1(n13164), .B2(n15483), .A(n13163), .ZN(n13165) );
  AOI21_X1 U15454 ( .B1(n13340), .B2(n13255), .A(n13165), .ZN(n13166) );
  OAI21_X1 U15455 ( .B1(n13341), .B2(n15519), .A(n13166), .ZN(P3_U3208) );
  XNOR2_X1 U15456 ( .A(n13171), .B(n13167), .ZN(n13169) );
  AOI222_X1 U15457 ( .A1(n13308), .A2(n13169), .B1(n13198), .B2(n15504), .C1(
        n13168), .C2(n13320), .ZN(n13345) );
  OAI21_X1 U15458 ( .B1(n13172), .B2(n13171), .A(n13170), .ZN(n13343) );
  INV_X1 U15459 ( .A(n8571), .ZN(n13175) );
  AOI22_X1 U15460 ( .A1(n13173), .A2(n15516), .B1(n15519), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13174) );
  OAI21_X1 U15461 ( .B1(n13175), .B2(n15483), .A(n13174), .ZN(n13176) );
  AOI21_X1 U15462 ( .B1(n13343), .B2(n13255), .A(n13176), .ZN(n13177) );
  OAI21_X1 U15463 ( .B1(n13345), .B2(n15519), .A(n13177), .ZN(P3_U3209) );
  XNOR2_X1 U15464 ( .A(n13179), .B(n13178), .ZN(n13183) );
  OAI22_X1 U15465 ( .A1(n13181), .A2(n15491), .B1(n13180), .B2(n15492), .ZN(
        n13182) );
  AOI21_X1 U15466 ( .B1(n13183), .B2(n13308), .A(n13182), .ZN(n13187) );
  XNOR2_X1 U15467 ( .A(n13184), .B(n13185), .ZN(n13346) );
  NAND2_X1 U15468 ( .A1(n13346), .A2(n15511), .ZN(n13186) );
  INV_X1 U15469 ( .A(n13188), .ZN(n13193) );
  INV_X1 U15470 ( .A(n13189), .ZN(n13408) );
  AOI22_X1 U15471 ( .A1(n13190), .A2(n15516), .B1(n15519), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13191) );
  OAI21_X1 U15472 ( .B1(n13408), .B2(n15483), .A(n13191), .ZN(n13192) );
  AOI21_X1 U15473 ( .B1(n13346), .B2(n13193), .A(n13192), .ZN(n13194) );
  OAI21_X1 U15474 ( .B1(n13348), .B2(n15519), .A(n13194), .ZN(P3_U3210) );
  XOR2_X1 U15475 ( .A(n13196), .B(n13195), .Z(n13414) );
  XOR2_X1 U15476 ( .A(n13197), .B(n13196), .Z(n13199) );
  AOI222_X1 U15477 ( .A1(n13308), .A2(n13199), .B1(n13198), .B2(n13320), .C1(
        n13222), .C2(n15504), .ZN(n13409) );
  MUX2_X1 U15478 ( .A(n13200), .B(n13409), .S(n15500), .Z(n13203) );
  AOI22_X1 U15479 ( .A1(n13411), .A2(n6529), .B1(n15516), .B2(n13201), .ZN(
        n13202) );
  OAI211_X1 U15480 ( .C1(n13414), .C2(n13327), .A(n13203), .B(n13202), .ZN(
        P3_U3211) );
  XNOR2_X1 U15481 ( .A(n13204), .B(n13205), .ZN(n13420) );
  XNOR2_X1 U15482 ( .A(n13206), .B(n13205), .ZN(n13209) );
  AOI222_X1 U15483 ( .A1(n13308), .A2(n13209), .B1(n13208), .B2(n13320), .C1(
        n13207), .C2(n15504), .ZN(n13415) );
  MUX2_X1 U15484 ( .A(n13210), .B(n13415), .S(n15500), .Z(n13213) );
  AOI22_X1 U15485 ( .A1(n13417), .A2(n6529), .B1(n15516), .B2(n13211), .ZN(
        n13212) );
  OAI211_X1 U15486 ( .C1(n13420), .C2(n13327), .A(n13213), .B(n13212), .ZN(
        P3_U3212) );
  OR2_X1 U15487 ( .A1(n13214), .A2(n13215), .ZN(n13217) );
  AND2_X1 U15488 ( .A1(n13217), .A2(n13216), .ZN(n13219) );
  XNOR2_X1 U15489 ( .A(n13219), .B(n13218), .ZN(n13426) );
  INV_X1 U15490 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13224) );
  XNOR2_X1 U15491 ( .A(n13221), .B(n13220), .ZN(n13223) );
  AOI222_X1 U15492 ( .A1(n13308), .A2(n13223), .B1(n13243), .B2(n15504), .C1(
        n13222), .C2(n13320), .ZN(n13421) );
  MUX2_X1 U15493 ( .A(n13224), .B(n13421), .S(n15500), .Z(n13227) );
  AOI22_X1 U15494 ( .A1(n13423), .A2(n6529), .B1(n15516), .B2(n13225), .ZN(
        n13226) );
  OAI211_X1 U15495 ( .C1(n13426), .C2(n13327), .A(n13227), .B(n13226), .ZN(
        P3_U3213) );
  NAND2_X1 U15496 ( .A1(n13365), .A2(n13228), .ZN(n13229) );
  XNOR2_X1 U15497 ( .A(n13229), .B(n13230), .ZN(n13429) );
  INV_X1 U15498 ( .A(n13429), .ZN(n13363) );
  XNOR2_X1 U15499 ( .A(n13231), .B(n13230), .ZN(n13235) );
  OAI22_X1 U15500 ( .A1(n13233), .A2(n15491), .B1(n13232), .B2(n15492), .ZN(
        n13234) );
  AOI21_X1 U15501 ( .B1(n13235), .B2(n13308), .A(n13234), .ZN(n13428) );
  MUX2_X1 U15502 ( .A(n13428), .B(n13236), .S(n15519), .Z(n13239) );
  INV_X1 U15503 ( .A(n13432), .ZN(n13360) );
  AOI22_X1 U15504 ( .A1(n13360), .A2(n6529), .B1(n15516), .B2(n13237), .ZN(
        n13238) );
  OAI211_X1 U15505 ( .C1(n13363), .C2(n13327), .A(n13239), .B(n13238), .ZN(
        P3_U3214) );
  NAND2_X1 U15506 ( .A1(n13240), .A2(n7348), .ZN(n13241) );
  NAND2_X1 U15507 ( .A1(n13242), .A2(n13241), .ZN(n13246) );
  NAND2_X1 U15508 ( .A1(n13243), .A2(n13320), .ZN(n13244) );
  OAI21_X1 U15509 ( .B1(n13273), .B2(n15492), .A(n13244), .ZN(n13245) );
  AOI21_X1 U15510 ( .B1(n13246), .B2(n13308), .A(n13245), .ZN(n13369) );
  NAND2_X1 U15511 ( .A1(n13247), .A2(n13374), .ZN(n13366) );
  INV_X1 U15512 ( .A(n13366), .ZN(n13253) );
  INV_X1 U15513 ( .A(n13248), .ZN(n13249) );
  OAI22_X1 U15514 ( .A1(n15500), .A2(n13250), .B1(n13249), .B2(n15486), .ZN(
        n13251) );
  AOI21_X1 U15515 ( .B1(n13253), .B2(n13252), .A(n13251), .ZN(n13257) );
  NAND2_X1 U15516 ( .A1(n13214), .A2(n13254), .ZN(n13364) );
  NAND3_X1 U15517 ( .A1(n13365), .A2(n13364), .A3(n13255), .ZN(n13256) );
  OAI211_X1 U15518 ( .C1(n13369), .C2(n15519), .A(n13257), .B(n13256), .ZN(
        P3_U3215) );
  XOR2_X1 U15519 ( .A(n13258), .B(n13259), .Z(n13439) );
  XOR2_X1 U15520 ( .A(n13260), .B(n13259), .Z(n13262) );
  AOI222_X1 U15521 ( .A1(n13308), .A2(n13262), .B1(n13261), .B2(n13320), .C1(
        n13283), .C2(n15504), .ZN(n13434) );
  MUX2_X1 U15522 ( .A(n13263), .B(n13434), .S(n15500), .Z(n13266) );
  AOI22_X1 U15523 ( .A1(n13436), .A2(n6529), .B1(n15516), .B2(n13264), .ZN(
        n13265) );
  OAI211_X1 U15524 ( .C1(n13439), .C2(n13327), .A(n13266), .B(n13265), .ZN(
        P3_U3216) );
  OAI21_X1 U15525 ( .B1(n13268), .B2(n13270), .A(n13267), .ZN(n13269) );
  INV_X1 U15526 ( .A(n13269), .ZN(n13443) );
  OAI222_X1 U15527 ( .A1(n15491), .A2(n13273), .B1(n15492), .B2(n13272), .C1(
        n15508), .C2(n13271), .ZN(n13372) );
  NAND2_X1 U15528 ( .A1(n13372), .A2(n15500), .ZN(n13279) );
  INV_X1 U15529 ( .A(n13274), .ZN(n13275) );
  OAI22_X1 U15530 ( .A1(n15500), .A2(n13276), .B1(n13275), .B2(n15486), .ZN(
        n13277) );
  AOI21_X1 U15531 ( .B1(n13373), .B2(n6529), .A(n13277), .ZN(n13278) );
  OAI211_X1 U15532 ( .C1(n13443), .C2(n13327), .A(n13279), .B(n13278), .ZN(
        P3_U3217) );
  XNOR2_X1 U15533 ( .A(n13280), .B(n7409), .ZN(n13449) );
  XNOR2_X1 U15534 ( .A(n13282), .B(n13281), .ZN(n13284) );
  AOI222_X1 U15535 ( .A1(n13308), .A2(n13284), .B1(n13283), .B2(n13320), .C1(
        n13305), .C2(n15504), .ZN(n13444) );
  MUX2_X1 U15536 ( .A(n13285), .B(n13444), .S(n15500), .Z(n13288) );
  AOI22_X1 U15537 ( .A1(n13446), .A2(n6529), .B1(n15516), .B2(n13286), .ZN(
        n13287) );
  OAI211_X1 U15538 ( .C1(n13449), .C2(n13327), .A(n13288), .B(n13287), .ZN(
        P3_U3218) );
  XNOR2_X1 U15539 ( .A(n13289), .B(n7305), .ZN(n13455) );
  INV_X1 U15540 ( .A(n13291), .ZN(n13292) );
  OAI21_X1 U15541 ( .B1(n13290), .B2(n13293), .A(n13292), .ZN(n13294) );
  XNOR2_X1 U15542 ( .A(n13294), .B(n7305), .ZN(n13296) );
  AOI222_X1 U15543 ( .A1(n13308), .A2(n13296), .B1(n13295), .B2(n13320), .C1(
        n13319), .C2(n15504), .ZN(n13450) );
  MUX2_X1 U15544 ( .A(n13297), .B(n13450), .S(n15500), .Z(n13300) );
  AOI22_X1 U15545 ( .A1(n13452), .A2(n6529), .B1(n15516), .B2(n13298), .ZN(
        n13299) );
  OAI211_X1 U15546 ( .C1(n13455), .C2(n13327), .A(n13300), .B(n13299), .ZN(
        P3_U3219) );
  XNOR2_X1 U15547 ( .A(n13301), .B(n13303), .ZN(n13462) );
  NOR2_X1 U15548 ( .A1(n13290), .A2(n13316), .ZN(n13315) );
  NOR2_X1 U15549 ( .A1(n13315), .A2(n13302), .ZN(n13304) );
  XNOR2_X1 U15550 ( .A(n13304), .B(n13303), .ZN(n13307) );
  AOI222_X1 U15551 ( .A1(n13308), .A2(n13307), .B1(n13306), .B2(n15504), .C1(
        n13305), .C2(n13320), .ZN(n13456) );
  MUX2_X1 U15552 ( .A(n13309), .B(n13456), .S(n15500), .Z(n13312) );
  AOI22_X1 U15553 ( .A1(n6529), .A2(n13457), .B1(n15516), .B2(n13310), .ZN(
        n13311) );
  OAI211_X1 U15554 ( .C1(n13462), .C2(n13327), .A(n13312), .B(n13311), .ZN(
        P3_U3220) );
  XNOR2_X1 U15555 ( .A(n13313), .B(n13316), .ZN(n13466) );
  INV_X1 U15556 ( .A(n13466), .ZN(n13328) );
  AND2_X1 U15557 ( .A1(n13314), .A2(n15504), .ZN(n13318) );
  AOI211_X1 U15558 ( .C1(n13316), .C2(n13290), .A(n15508), .B(n13315), .ZN(
        n13317) );
  AOI211_X1 U15559 ( .C1(n13320), .C2(n13319), .A(n13318), .B(n13317), .ZN(
        n13463) );
  MUX2_X1 U15560 ( .A(n13321), .B(n13463), .S(n15500), .Z(n13326) );
  INV_X1 U15561 ( .A(n13469), .ZN(n13323) );
  AOI22_X1 U15562 ( .A1(n6529), .A2(n13323), .B1(n15516), .B2(n13322), .ZN(
        n13325) );
  OAI211_X1 U15563 ( .C1(n13328), .C2(n13327), .A(n13326), .B(n13325), .ZN(
        P3_U3221) );
  NAND2_X1 U15564 ( .A1(n12587), .A2(n13383), .ZN(n13329) );
  NAND2_X1 U15565 ( .A1(n15549), .A2(n13392), .ZN(n13331) );
  OAI211_X1 U15566 ( .C1(n15549), .C2(n13330), .A(n13329), .B(n13331), .ZN(
        P3_U3490) );
  NAND2_X1 U15567 ( .A1(n13395), .A2(n13383), .ZN(n13332) );
  OAI211_X1 U15568 ( .C1(n15549), .C2(n10384), .A(n13332), .B(n13331), .ZN(
        P3_U3489) );
  INV_X1 U15569 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13336) );
  INV_X1 U15570 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U15571 ( .A1(n13340), .A2(n15537), .B1(n13374), .B2(n13339), .ZN(
        n13342) );
  NAND2_X1 U15572 ( .A1(n13342), .A2(n13341), .ZN(n13404) );
  MUX2_X1 U15573 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13404), .S(n15549), .Z(
        P3_U3484) );
  AOI22_X1 U15574 ( .A1(n13343), .A2(n15537), .B1(n13374), .B2(n8571), .ZN(
        n13344) );
  NAND2_X1 U15575 ( .A1(n13345), .A2(n13344), .ZN(n13405) );
  MUX2_X1 U15576 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13405), .S(n15549), .Z(
        P3_U3483) );
  NAND2_X1 U15577 ( .A1(n13346), .A2(n6716), .ZN(n13347) );
  MUX2_X1 U15578 ( .A(n15797), .B(n13406), .S(n15549), .Z(n13349) );
  OAI21_X1 U15579 ( .B1(n13408), .B2(n13391), .A(n13349), .ZN(P3_U3482) );
  INV_X1 U15580 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13350) );
  MUX2_X1 U15581 ( .A(n13350), .B(n13409), .S(n15549), .Z(n13352) );
  NAND2_X1 U15582 ( .A1(n13411), .A2(n13383), .ZN(n13351) );
  OAI211_X1 U15583 ( .C1(n13386), .C2(n13414), .A(n13352), .B(n13351), .ZN(
        P3_U3481) );
  INV_X1 U15584 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13353) );
  MUX2_X1 U15585 ( .A(n13353), .B(n13415), .S(n15549), .Z(n13355) );
  NAND2_X1 U15586 ( .A1(n13417), .A2(n13383), .ZN(n13354) );
  OAI211_X1 U15587 ( .C1(n13386), .C2(n13420), .A(n13355), .B(n13354), .ZN(
        P3_U3480) );
  INV_X1 U15588 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13356) );
  MUX2_X1 U15589 ( .A(n13356), .B(n13421), .S(n15549), .Z(n13358) );
  NAND2_X1 U15590 ( .A1(n13423), .A2(n13383), .ZN(n13357) );
  OAI211_X1 U15591 ( .C1(n13386), .C2(n13426), .A(n13358), .B(n13357), .ZN(
        P3_U3479) );
  INV_X1 U15592 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13359) );
  MUX2_X1 U15593 ( .A(n13359), .B(n13428), .S(n15549), .Z(n13362) );
  NAND2_X1 U15594 ( .A1(n13360), .A2(n13383), .ZN(n13361) );
  OAI211_X1 U15595 ( .C1(n13363), .C2(n13386), .A(n13362), .B(n13361), .ZN(
        P3_U3478) );
  NAND3_X1 U15596 ( .A1(n13365), .A2(n13364), .A3(n15537), .ZN(n13367) );
  AND2_X1 U15597 ( .A1(n13367), .A2(n13366), .ZN(n13368) );
  NAND2_X1 U15598 ( .A1(n13369), .A2(n13368), .ZN(n13433) );
  MUX2_X1 U15599 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13433), .S(n15549), .Z(
        P3_U3477) );
  MUX2_X1 U15600 ( .A(n6930), .B(n13434), .S(n15549), .Z(n13371) );
  NAND2_X1 U15601 ( .A1(n13436), .A2(n13383), .ZN(n13370) );
  OAI211_X1 U15602 ( .C1(n13386), .C2(n13439), .A(n13371), .B(n13370), .ZN(
        P3_U3476) );
  INV_X1 U15603 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13375) );
  AOI21_X1 U15604 ( .B1(n13374), .B2(n13373), .A(n13372), .ZN(n13440) );
  MUX2_X1 U15605 ( .A(n13375), .B(n13440), .S(n15549), .Z(n13376) );
  OAI21_X1 U15606 ( .B1(n13443), .B2(n13386), .A(n13376), .ZN(P3_U3475) );
  MUX2_X1 U15607 ( .A(n13377), .B(n13444), .S(n15549), .Z(n13379) );
  NAND2_X1 U15608 ( .A1(n13446), .A2(n13383), .ZN(n13378) );
  OAI211_X1 U15609 ( .C1(n13386), .C2(n13449), .A(n13379), .B(n13378), .ZN(
        P3_U3474) );
  MUX2_X1 U15610 ( .A(n13380), .B(n13450), .S(n15549), .Z(n13382) );
  NAND2_X1 U15611 ( .A1(n13452), .A2(n13383), .ZN(n13381) );
  OAI211_X1 U15612 ( .C1(n13455), .C2(n13386), .A(n13382), .B(n13381), .ZN(
        P3_U3473) );
  MUX2_X1 U15613 ( .A(n15767), .B(n13456), .S(n15549), .Z(n13385) );
  NAND2_X1 U15614 ( .A1(n13457), .A2(n13383), .ZN(n13384) );
  OAI211_X1 U15615 ( .C1(n13386), .C2(n13462), .A(n13385), .B(n13384), .ZN(
        P3_U3472) );
  MUX2_X1 U15616 ( .A(n13387), .B(n13463), .S(n15549), .Z(n13390) );
  NAND2_X1 U15617 ( .A1(n13466), .A2(n13388), .ZN(n13389) );
  OAI211_X1 U15618 ( .C1(n13391), .C2(n13469), .A(n13390), .B(n13389), .ZN(
        P3_U3471) );
  NAND2_X1 U15619 ( .A1(n12587), .A2(n13458), .ZN(n13393) );
  NAND2_X1 U15620 ( .A1(n15540), .A2(n13392), .ZN(n13396) );
  OAI211_X1 U15621 ( .C1(n15540), .C2(n13394), .A(n13393), .B(n13396), .ZN(
        P3_U3458) );
  NAND2_X1 U15622 ( .A1(n13395), .A2(n13458), .ZN(n13397) );
  OAI211_X1 U15623 ( .C1(n10385), .C2(n15540), .A(n13397), .B(n13396), .ZN(
        P3_U3457) );
  OAI21_X1 U15624 ( .B1(n13403), .B2(n13461), .A(n13402), .ZN(P3_U3453) );
  MUX2_X1 U15625 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13404), .S(n15540), .Z(
        P3_U3452) );
  MUX2_X1 U15626 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13405), .S(n15540), .Z(
        P3_U3451) );
  MUX2_X1 U15627 ( .A(n13406), .B(n15708), .S(n15539), .Z(n13407) );
  OAI21_X1 U15628 ( .B1(n13408), .B2(n13470), .A(n13407), .ZN(P3_U3450) );
  INV_X1 U15629 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13410) );
  MUX2_X1 U15630 ( .A(n13410), .B(n13409), .S(n15540), .Z(n13413) );
  NAND2_X1 U15631 ( .A1(n13411), .A2(n13458), .ZN(n13412) );
  OAI211_X1 U15632 ( .C1(n13414), .C2(n13461), .A(n13413), .B(n13412), .ZN(
        P3_U3449) );
  INV_X1 U15633 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13416) );
  MUX2_X1 U15634 ( .A(n13416), .B(n13415), .S(n15540), .Z(n13419) );
  NAND2_X1 U15635 ( .A1(n13417), .A2(n13458), .ZN(n13418) );
  OAI211_X1 U15636 ( .C1(n13420), .C2(n13461), .A(n13419), .B(n13418), .ZN(
        P3_U3448) );
  MUX2_X1 U15637 ( .A(n13422), .B(n13421), .S(n15540), .Z(n13425) );
  NAND2_X1 U15638 ( .A1(n13423), .A2(n13458), .ZN(n13424) );
  OAI211_X1 U15639 ( .C1(n13426), .C2(n13461), .A(n13425), .B(n13424), .ZN(
        P3_U3447) );
  INV_X1 U15640 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13427) );
  MUX2_X1 U15641 ( .A(n13428), .B(n13427), .S(n15539), .Z(n13431) );
  NAND2_X1 U15642 ( .A1(n13429), .A2(n13465), .ZN(n13430) );
  OAI211_X1 U15643 ( .C1(n13470), .C2(n13432), .A(n13431), .B(n13430), .ZN(
        P3_U3446) );
  MUX2_X1 U15644 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13433), .S(n15540), .Z(
        P3_U3444) );
  INV_X1 U15645 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13435) );
  MUX2_X1 U15646 ( .A(n13435), .B(n13434), .S(n15540), .Z(n13438) );
  NAND2_X1 U15647 ( .A1(n13436), .A2(n13458), .ZN(n13437) );
  OAI211_X1 U15648 ( .C1(n13439), .C2(n13461), .A(n13438), .B(n13437), .ZN(
        P3_U3441) );
  MUX2_X1 U15649 ( .A(n13441), .B(n13440), .S(n15540), .Z(n13442) );
  OAI21_X1 U15650 ( .B1(n13443), .B2(n13461), .A(n13442), .ZN(P3_U3438) );
  INV_X1 U15651 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13445) );
  MUX2_X1 U15652 ( .A(n13445), .B(n13444), .S(n15540), .Z(n13448) );
  NAND2_X1 U15653 ( .A1(n13446), .A2(n13458), .ZN(n13447) );
  OAI211_X1 U15654 ( .C1(n13449), .C2(n13461), .A(n13448), .B(n13447), .ZN(
        P3_U3435) );
  MUX2_X1 U15655 ( .A(n13451), .B(n13450), .S(n15540), .Z(n13454) );
  NAND2_X1 U15656 ( .A1(n13458), .A2(n13452), .ZN(n13453) );
  OAI211_X1 U15657 ( .C1(n13455), .C2(n13461), .A(n13454), .B(n13453), .ZN(
        P3_U3432) );
  MUX2_X1 U15658 ( .A(n15737), .B(n13456), .S(n15540), .Z(n13460) );
  NAND2_X1 U15659 ( .A1(n13458), .A2(n13457), .ZN(n13459) );
  OAI211_X1 U15660 ( .C1(n13462), .C2(n13461), .A(n13460), .B(n13459), .ZN(
        P3_U3429) );
  MUX2_X1 U15661 ( .A(n13464), .B(n13463), .S(n15540), .Z(n13468) );
  NAND2_X1 U15662 ( .A1(n13466), .A2(n13465), .ZN(n13467) );
  OAI211_X1 U15663 ( .C1(n13470), .C2(n13469), .A(n13468), .B(n13467), .ZN(
        P3_U3426) );
  MUX2_X1 U15664 ( .A(n13471), .B(P3_D_REG_1__SCAN_IN), .S(n13472), .Z(
        P3_U3377) );
  MUX2_X1 U15665 ( .A(n13473), .B(P3_D_REG_0__SCAN_IN), .S(n13472), .Z(
        P3_U3376) );
  NAND4_X1 U15666 ( .A1(n13475), .A2(n13474), .A3(P3_STATE_REG_SCAN_IN), .A4(
        P3_IR_REG_31__SCAN_IN), .ZN(n13477) );
  OAI22_X1 U15667 ( .A1(n13478), .A2(n13477), .B1(n13476), .B2(n13487), .ZN(
        n13479) );
  AOI21_X1 U15668 ( .B1(n13481), .B2(n13480), .A(n13479), .ZN(n13482) );
  INV_X1 U15669 ( .A(n13482), .ZN(P3_U3264) );
  INV_X1 U15670 ( .A(n13483), .ZN(n13485) );
  OAI222_X1 U15671 ( .A1(n13487), .A2(n15777), .B1(n13495), .B2(n13485), .C1(
        P3_U3151), .C2(n13484), .ZN(P3_U3266) );
  INV_X1 U15672 ( .A(n13486), .ZN(n13490) );
  OAI222_X1 U15673 ( .A1(n13495), .A2(n13490), .B1(n13489), .B2(P3_U3151), 
        .C1(n13488), .C2(n13487), .ZN(P3_U3268) );
  INV_X1 U15674 ( .A(n13491), .ZN(n13494) );
  OAI222_X1 U15675 ( .A1(n13495), .A2(n13494), .B1(P3_U3151), .B2(n13493), 
        .C1(n13492), .C2(n13487), .ZN(P3_U3269) );
  XNOR2_X1 U15676 ( .A(n6680), .B(n13496), .ZN(n13502) );
  OAI22_X1 U15677 ( .A1(n13782), .A2(n13618), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13497), .ZN(n13498) );
  AOI21_X1 U15678 ( .B1(n13966), .B2(n13634), .A(n13498), .ZN(n13499) );
  OAI21_X1 U15679 ( .B1(n13793), .B2(n13621), .A(n13499), .ZN(n13500) );
  AOI21_X1 U15680 ( .B1(n14211), .B2(n13623), .A(n13500), .ZN(n13501) );
  OAI21_X1 U15681 ( .B1(n13502), .B2(n13625), .A(n13501), .ZN(P2_U3186) );
  INV_X1 U15682 ( .A(n13503), .ZN(n13504) );
  AOI21_X1 U15683 ( .B1(n13506), .B2(n13505), .A(n13504), .ZN(n13512) );
  AOI22_X1 U15684 ( .A1(n13605), .A2(n13896), .B1(n13634), .B2(n13507), .ZN(
        n13509) );
  OAI211_X1 U15685 ( .C1(n13733), .C2(n13621), .A(n13509), .B(n13508), .ZN(
        n13510) );
  AOI21_X1 U15686 ( .B1(n13724), .B2(n13623), .A(n13510), .ZN(n13511) );
  OAI21_X1 U15687 ( .B1(n13512), .B2(n13625), .A(n13511), .ZN(P2_U3187) );
  XNOR2_X1 U15688 ( .A(n13568), .B(n13513), .ZN(n13572) );
  XNOR2_X1 U15689 ( .A(n13572), .B(n13571), .ZN(n13518) );
  OAI22_X1 U15690 ( .A1(n14025), .A2(n13621), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13514), .ZN(n13516) );
  OAI22_X1 U15691 ( .A1(n14024), .A2(n13618), .B1(n14031), .B2(n13599), .ZN(
        n13515) );
  AOI211_X1 U15692 ( .C1(n14034), .C2(n13623), .A(n13516), .B(n13515), .ZN(
        n13517) );
  OAI21_X1 U15693 ( .B1(n13518), .B2(n13625), .A(n13517), .ZN(P2_U3188) );
  NAND2_X1 U15694 ( .A1(n13520), .A2(n13519), .ZN(n13522) );
  XOR2_X1 U15695 ( .A(n13522), .B(n13521), .Z(n13527) );
  OAI21_X1 U15696 ( .B1(n13618), .B2(n14091), .A(n13523), .ZN(n13525) );
  INV_X1 U15697 ( .A(n14057), .ZN(n14093) );
  OAI22_X1 U15698 ( .A1(n13621), .A2(n14093), .B1(n13599), .B2(n14099), .ZN(
        n13524) );
  AOI211_X1 U15699 ( .C1(n14257), .C2(n13623), .A(n13525), .B(n13524), .ZN(
        n13526) );
  OAI21_X1 U15700 ( .B1(n13527), .B2(n13625), .A(n13526), .ZN(P2_U3191) );
  XNOR2_X1 U15701 ( .A(n13529), .B(n13528), .ZN(n13534) );
  OAI22_X1 U15702 ( .A1(n14024), .A2(n13621), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13530), .ZN(n13532) );
  OAI22_X1 U15703 ( .A1(n13618), .A2(n14093), .B1(n13599), .B2(n14061), .ZN(
        n13531) );
  AOI211_X1 U15704 ( .C1(n14246), .C2(n13623), .A(n13532), .B(n13531), .ZN(
        n13533) );
  OAI21_X1 U15705 ( .B1(n13534), .B2(n13625), .A(n13533), .ZN(P2_U3195) );
  XNOR2_X1 U15706 ( .A(n13536), .B(n13535), .ZN(n13542) );
  NAND2_X1 U15707 ( .A1(n13999), .A2(n13537), .ZN(n13539) );
  AOI22_X1 U15708 ( .A1(n13998), .A2(n13605), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13538) );
  OAI211_X1 U15709 ( .C1(n13599), .C2(n13989), .A(n13539), .B(n13538), .ZN(
        n13540) );
  AOI21_X1 U15710 ( .B1(n14225), .B2(n13623), .A(n13540), .ZN(n13541) );
  OAI21_X1 U15711 ( .B1(n13542), .B2(n13625), .A(n13541), .ZN(P2_U3197) );
  XNOR2_X1 U15712 ( .A(n13544), .B(n13543), .ZN(n13549) );
  INV_X1 U15713 ( .A(n13545), .ZN(n13547) );
  XNOR2_X1 U15714 ( .A(n13546), .B(n13545), .ZN(n13630) );
  NAND2_X1 U15715 ( .A1(n13630), .A2(n13629), .ZN(n13628) );
  OAI21_X1 U15716 ( .B1(n13547), .B2(n13546), .A(n13628), .ZN(n13548) );
  NOR2_X1 U15717 ( .A1(n13548), .A2(n13549), .ZN(n13559) );
  AOI21_X1 U15718 ( .B1(n13549), .B2(n13548), .A(n13559), .ZN(n13555) );
  OAI22_X1 U15719 ( .A1(n13743), .A2(n14094), .B1(n13733), .B2(n14092), .ZN(
        n14273) );
  NAND2_X1 U15720 ( .A1(n13550), .A2(n14273), .ZN(n13551) );
  OAI211_X1 U15721 ( .C1(n13599), .C2(n14147), .A(n13552), .B(n13551), .ZN(
        n13553) );
  AOI21_X1 U15722 ( .B1(n14274), .B2(n13623), .A(n13553), .ZN(n13554) );
  OAI21_X1 U15723 ( .B1(n13555), .B2(n13625), .A(n13554), .ZN(P2_U3198) );
  INV_X1 U15724 ( .A(n13556), .ZN(n13558) );
  NOR3_X1 U15725 ( .A1(n13559), .A2(n13558), .A3(n13557), .ZN(n13562) );
  INV_X1 U15726 ( .A(n13560), .ZN(n13561) );
  OAI21_X1 U15727 ( .B1(n13562), .B2(n13561), .A(n13627), .ZN(n13567) );
  AND2_X1 U15728 ( .A1(n13893), .A2(n14106), .ZN(n13563) );
  AOI21_X1 U15729 ( .B1(n13892), .B2(n14108), .A(n13563), .ZN(n14126) );
  OAI21_X1 U15730 ( .B1(n13632), .B2(n14126), .A(n13564), .ZN(n13565) );
  AOI21_X1 U15731 ( .B1(n13634), .B2(n14132), .A(n13565), .ZN(n13566) );
  OAI211_X1 U15732 ( .C1(n13742), .C2(n13637), .A(n13567), .B(n13566), .ZN(
        P2_U3200) );
  INV_X1 U15733 ( .A(n13568), .ZN(n13570) );
  OAI22_X1 U15734 ( .A1(n13572), .A2(n13571), .B1(n13570), .B2(n13569), .ZN(
        n13576) );
  XNOR2_X1 U15735 ( .A(n13574), .B(n13573), .ZN(n13575) );
  XNOR2_X1 U15736 ( .A(n13576), .B(n13575), .ZN(n13582) );
  OAI22_X1 U15737 ( .A1(n13977), .A2(n13621), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13577), .ZN(n13580) );
  INV_X1 U15738 ( .A(n14015), .ZN(n13578) );
  OAI22_X1 U15739 ( .A1(n13578), .A2(n13599), .B1(n13597), .B2(n13618), .ZN(
        n13579) );
  AOI211_X1 U15740 ( .C1(n14230), .C2(n13623), .A(n13580), .B(n13579), .ZN(
        n13581) );
  OAI21_X1 U15741 ( .B1(n13582), .B2(n13625), .A(n13581), .ZN(P2_U3201) );
  INV_X1 U15742 ( .A(n13583), .ZN(n13584) );
  AOI21_X1 U15743 ( .B1(n13586), .B2(n13585), .A(n13584), .ZN(n13591) );
  OAI22_X1 U15744 ( .A1(n13621), .A2(n13600), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13587), .ZN(n13589) );
  OAI22_X1 U15745 ( .A1(n13618), .A2(n13607), .B1(n13599), .B2(n14072), .ZN(
        n13588) );
  AOI211_X1 U15746 ( .C1(n14252), .C2(n13623), .A(n13589), .B(n13588), .ZN(
        n13590) );
  OAI21_X1 U15747 ( .B1(n13591), .B2(n13625), .A(n13590), .ZN(P2_U3205) );
  XOR2_X1 U15748 ( .A(n13593), .B(n13592), .Z(n13594) );
  XNOR2_X1 U15749 ( .A(n13595), .B(n13594), .ZN(n13604) );
  OAI22_X1 U15750 ( .A1(n13597), .A2(n13621), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13596), .ZN(n13602) );
  INV_X1 U15751 ( .A(n14048), .ZN(n13598) );
  OAI22_X1 U15752 ( .A1(n13600), .A2(n13618), .B1(n13599), .B2(n13598), .ZN(
        n13601) );
  AOI211_X1 U15753 ( .C1(n14049), .C2(n13623), .A(n13602), .B(n13601), .ZN(
        n13603) );
  OAI21_X1 U15754 ( .B1(n13604), .B2(n13625), .A(n13603), .ZN(P2_U3207) );
  AOI22_X1 U15755 ( .A1(n13605), .A2(n14107), .B1(n13634), .B2(n14113), .ZN(
        n13606) );
  NAND2_X1 U15756 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13926)
         );
  OAI211_X1 U15757 ( .C1(n13607), .C2(n13621), .A(n13606), .B(n13926), .ZN(
        n13613) );
  INV_X1 U15758 ( .A(n13608), .ZN(n13609) );
  AOI211_X1 U15759 ( .C1(n13611), .C2(n13610), .A(n13625), .B(n13609), .ZN(
        n13612) );
  AOI211_X1 U15760 ( .C1(n14262), .C2(n13623), .A(n13613), .B(n13612), .ZN(
        n13614) );
  INV_X1 U15761 ( .A(n13614), .ZN(P2_U3210) );
  AOI21_X1 U15762 ( .B1(n13617), .B2(n13616), .A(n13615), .ZN(n13626) );
  OAI22_X1 U15763 ( .A1(n13977), .A2(n13618), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15702), .ZN(n13619) );
  AOI21_X1 U15764 ( .B1(n13979), .B2(n13634), .A(n13619), .ZN(n13620) );
  OAI21_X1 U15765 ( .B1(n13978), .B2(n13621), .A(n13620), .ZN(n13622) );
  AOI21_X1 U15766 ( .B1(n14220), .B2(n13623), .A(n13622), .ZN(n13624) );
  OAI21_X1 U15767 ( .B1(n13626), .B2(n13625), .A(n13624), .ZN(P2_U3212) );
  OAI211_X1 U15768 ( .C1(n13630), .C2(n13629), .A(n13628), .B(n13627), .ZN(
        n13636) );
  AOI22_X1 U15769 ( .A1(n13893), .A2(n14108), .B1(n14106), .B2(n13895), .ZN(
        n14161) );
  OAI21_X1 U15770 ( .B1(n13632), .B2(n14161), .A(n13631), .ZN(n13633) );
  AOI21_X1 U15771 ( .B1(n13634), .B2(n14168), .A(n13633), .ZN(n13635) );
  OAI211_X1 U15772 ( .C1(n14280), .C2(n13637), .A(n13636), .B(n13635), .ZN(
        P2_U3213) );
  MUX2_X1 U15773 ( .A(n11068), .B(n13639), .S(n6533), .Z(n13649) );
  NAND2_X1 U15774 ( .A1(n10686), .A2(n13640), .ZN(n13646) );
  NAND2_X1 U15775 ( .A1(n13641), .A2(n13792), .ZN(n13645) );
  NAND3_X1 U15776 ( .A1(n13646), .A2(n13643), .A3(n13642), .ZN(n13644) );
  OAI211_X1 U15777 ( .C1(n13792), .C2(n13646), .A(n13645), .B(n13644), .ZN(
        n13647) );
  NAND2_X1 U15778 ( .A1(n13649), .A2(n13648), .ZN(n13651) );
  NAND3_X1 U15779 ( .A1(n13652), .A2(n13651), .A3(n13650), .ZN(n13658) );
  AOI21_X1 U15780 ( .B1(n13906), .B2(n13792), .A(n10867), .ZN(n13655) );
  OAI21_X1 U15781 ( .B1(n13792), .B2(n13906), .A(n10867), .ZN(n13653) );
  INV_X1 U15782 ( .A(n13653), .ZN(n13654) );
  OAI21_X1 U15783 ( .B1(n13655), .B2(n13654), .A(n13845), .ZN(n13656) );
  INV_X1 U15784 ( .A(n13656), .ZN(n13657) );
  NAND2_X1 U15785 ( .A1(n13658), .A2(n13657), .ZN(n13668) );
  AOI21_X1 U15786 ( .B1(n13660), .B2(n13792), .A(n13659), .ZN(n13661) );
  INV_X1 U15787 ( .A(n13661), .ZN(n13665) );
  AOI21_X1 U15788 ( .B1(n13808), .B2(n13905), .A(n13662), .ZN(n13663) );
  INV_X1 U15789 ( .A(n13663), .ZN(n13664) );
  NAND2_X1 U15790 ( .A1(n13668), .A2(n13667), .ZN(n13673) );
  AND2_X1 U15791 ( .A1(n13792), .A2(n13904), .ZN(n13671) );
  OAI21_X1 U15792 ( .B1(n13792), .B2(n13904), .A(n13670), .ZN(n13669) );
  OAI21_X1 U15793 ( .B1(n13671), .B2(n13670), .A(n13669), .ZN(n13672) );
  NAND3_X1 U15794 ( .A1(n13673), .A2(n13672), .A3(n13852), .ZN(n13682) );
  OAI21_X1 U15795 ( .B1(n13675), .B2(n6533), .A(n13674), .ZN(n13679) );
  NAND2_X1 U15796 ( .A1(n13675), .A2(n13792), .ZN(n13677) );
  NAND2_X1 U15797 ( .A1(n13677), .A2(n13676), .ZN(n13678) );
  NAND2_X1 U15798 ( .A1(n13679), .A2(n13678), .ZN(n13681) );
  NAND3_X1 U15799 ( .A1(n13682), .A2(n13681), .A3(n13680), .ZN(n13686) );
  AND2_X1 U15800 ( .A1(n6532), .A2(n13902), .ZN(n13684) );
  OAI21_X1 U15801 ( .B1(n13902), .B2(n13792), .A(n15438), .ZN(n13683) );
  OAI21_X1 U15802 ( .B1(n13684), .B2(n15438), .A(n13683), .ZN(n13685) );
  NAND2_X1 U15803 ( .A1(n13686), .A2(n13685), .ZN(n13689) );
  MUX2_X1 U15804 ( .A(n13687), .B(n13901), .S(n13792), .Z(n13690) );
  MUX2_X1 U15805 ( .A(n13687), .B(n13901), .S(n13810), .Z(n13688) );
  XNOR2_X1 U15806 ( .A(n14314), .B(n6832), .ZN(n13691) );
  NOR2_X1 U15807 ( .A1(n13810), .A2(n13692), .ZN(n13694) );
  OAI21_X1 U15808 ( .B1(n6832), .B2(n13792), .A(n14314), .ZN(n13693) );
  OAI21_X1 U15809 ( .B1(n13694), .B2(n14314), .A(n13693), .ZN(n13695) );
  MUX2_X1 U15810 ( .A(n14307), .B(n13900), .S(n6533), .Z(n13698) );
  MUX2_X1 U15811 ( .A(n13900), .B(n14307), .S(n6532), .Z(n13696) );
  INV_X1 U15812 ( .A(n13698), .ZN(n13699) );
  MUX2_X1 U15813 ( .A(n13899), .B(n14302), .S(n6532), .Z(n13703) );
  MUX2_X1 U15814 ( .A(n14302), .B(n13899), .S(n6533), .Z(n13700) );
  NAND2_X1 U15815 ( .A1(n13701), .A2(n13700), .ZN(n13708) );
  INV_X1 U15816 ( .A(n13702), .ZN(n13705) );
  INV_X1 U15817 ( .A(n13703), .ZN(n13704) );
  NAND2_X1 U15818 ( .A1(n13705), .A2(n13704), .ZN(n13707) );
  NAND3_X1 U15819 ( .A1(n13708), .A2(n13707), .A3(n13706), .ZN(n13714) );
  NOR2_X1 U15820 ( .A1(n13709), .A2(n6533), .ZN(n13712) );
  OAI21_X1 U15821 ( .B1(n13810), .B2(n13898), .A(n13711), .ZN(n13710) );
  OAI21_X1 U15822 ( .B1(n13712), .B2(n13711), .A(n13710), .ZN(n13713) );
  MUX2_X1 U15823 ( .A(n13897), .B(n14297), .S(n6532), .Z(n13719) );
  XNOR2_X1 U15824 ( .A(n14292), .B(n13896), .ZN(n13715) );
  NOR2_X1 U15825 ( .A1(n13720), .A2(n13792), .ZN(n13722) );
  OAI21_X1 U15826 ( .B1(n13810), .B2(n13896), .A(n14292), .ZN(n13721) );
  OAI21_X1 U15827 ( .B1(n13722), .B2(n14292), .A(n13721), .ZN(n13723) );
  MUX2_X1 U15828 ( .A(n13895), .B(n13724), .S(n13792), .Z(n13728) );
  NAND2_X1 U15829 ( .A1(n13727), .A2(n13728), .ZN(n13726) );
  MUX2_X1 U15830 ( .A(n13895), .B(n13724), .S(n13810), .Z(n13725) );
  NAND2_X1 U15831 ( .A1(n13726), .A2(n13725), .ZN(n13732) );
  INV_X1 U15832 ( .A(n13727), .ZN(n13730) );
  INV_X1 U15833 ( .A(n13728), .ZN(n13729) );
  NAND2_X1 U15834 ( .A1(n13730), .A2(n13729), .ZN(n13731) );
  NAND2_X1 U15835 ( .A1(n13732), .A2(n13731), .ZN(n13736) );
  MUX2_X1 U15836 ( .A(n13894), .B(n14170), .S(n13810), .Z(n13735) );
  OAI21_X1 U15837 ( .B1(n13736), .B2(n13735), .A(n13864), .ZN(n13741) );
  MUX2_X1 U15838 ( .A(n13733), .B(n14280), .S(n6533), .Z(n13734) );
  AOI21_X1 U15839 ( .B1(n13736), .B2(n13735), .A(n13734), .ZN(n13740) );
  AND2_X1 U15840 ( .A1(n13893), .A2(n6532), .ZN(n13738) );
  OAI21_X1 U15841 ( .B1(n13893), .B2(n13792), .A(n14274), .ZN(n13737) );
  OAI21_X1 U15842 ( .B1(n13738), .B2(n14274), .A(n13737), .ZN(n13739) );
  MUX2_X1 U15843 ( .A(n14107), .B(n14268), .S(n13810), .Z(n13747) );
  MUX2_X1 U15844 ( .A(n13743), .B(n13742), .S(n13792), .Z(n13744) );
  INV_X1 U15845 ( .A(n13744), .ZN(n13745) );
  INV_X1 U15846 ( .A(n13747), .ZN(n13748) );
  MUX2_X1 U15847 ( .A(n13892), .B(n14262), .S(n6532), .Z(n13750) );
  MUX2_X1 U15848 ( .A(n14091), .B(n14115), .S(n13810), .Z(n13749) );
  MUX2_X1 U15849 ( .A(n14109), .B(n14257), .S(n13810), .Z(n13753) );
  MUX2_X1 U15850 ( .A(n14109), .B(n14257), .S(n6533), .Z(n13752) );
  INV_X1 U15851 ( .A(n13753), .ZN(n13754) );
  MUX2_X1 U15852 ( .A(n14057), .B(n14252), .S(n6533), .Z(n13758) );
  NAND2_X1 U15853 ( .A1(n13757), .A2(n13758), .ZN(n13756) );
  MUX2_X1 U15854 ( .A(n14057), .B(n14252), .S(n13810), .Z(n13755) );
  INV_X1 U15855 ( .A(n13757), .ZN(n13760) );
  INV_X1 U15856 ( .A(n13758), .ZN(n13759) );
  MUX2_X1 U15857 ( .A(n14081), .B(n14246), .S(n13810), .Z(n13762) );
  MUX2_X1 U15858 ( .A(n14081), .B(n14246), .S(n13792), .Z(n13761) );
  INV_X1 U15859 ( .A(n13762), .ZN(n13763) );
  MUX2_X1 U15860 ( .A(n14058), .B(n14049), .S(n6533), .Z(n13766) );
  MUX2_X1 U15861 ( .A(n14058), .B(n14049), .S(n13810), .Z(n13764) );
  MUX2_X1 U15862 ( .A(n14041), .B(n14034), .S(n13810), .Z(n13768) );
  MUX2_X1 U15863 ( .A(n14041), .B(n14034), .S(n6532), .Z(n13767) );
  INV_X1 U15864 ( .A(n13768), .ZN(n13769) );
  MUX2_X1 U15865 ( .A(n13998), .B(n14230), .S(n6532), .Z(n13773) );
  NAND2_X1 U15866 ( .A1(n13772), .A2(n13773), .ZN(n13771) );
  MUX2_X1 U15867 ( .A(n13998), .B(n14230), .S(n13808), .Z(n13770) );
  NAND2_X1 U15868 ( .A1(n13771), .A2(n13770), .ZN(n13777) );
  INV_X1 U15869 ( .A(n13772), .ZN(n13775) );
  INV_X1 U15870 ( .A(n13773), .ZN(n13774) );
  NAND2_X1 U15871 ( .A1(n13775), .A2(n13774), .ZN(n13776) );
  NAND2_X1 U15872 ( .A1(n13777), .A2(n13776), .ZN(n13778) );
  MUX2_X1 U15873 ( .A(n14007), .B(n14225), .S(n13810), .Z(n13779) );
  MUX2_X1 U15874 ( .A(n14007), .B(n14225), .S(n6532), .Z(n13780) );
  MUX2_X1 U15875 ( .A(n13782), .B(n13781), .S(n6533), .Z(n13784) );
  MUX2_X1 U15876 ( .A(n14220), .B(n13999), .S(n13792), .Z(n13783) );
  MUX2_X1 U15877 ( .A(n13978), .B(n13968), .S(n6533), .Z(n13795) );
  MUX2_X1 U15878 ( .A(n13891), .B(n14211), .S(n13810), .Z(n13794) );
  NAND2_X1 U15879 ( .A1(n15156), .A2(n13785), .ZN(n13787) );
  NAND2_X1 U15880 ( .A1(n9913), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13786) );
  NAND2_X2 U15881 ( .A1(n13787), .A2(n13786), .ZN(n14196) );
  NAND2_X1 U15882 ( .A1(n9653), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n13791) );
  NAND2_X1 U15883 ( .A1(n9974), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n13790) );
  NAND2_X1 U15884 ( .A1(n13788), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n13789) );
  NAND3_X1 U15885 ( .A1(n13791), .A2(n13790), .A3(n13789), .ZN(n13933) );
  XNOR2_X1 U15886 ( .A(n14196), .B(n13933), .ZN(n13841) );
  MUX2_X1 U15887 ( .A(n13961), .B(n14207), .S(n6532), .Z(n13819) );
  MUX2_X1 U15888 ( .A(n13793), .B(n13953), .S(n13808), .Z(n13820) );
  INV_X1 U15889 ( .A(n13794), .ZN(n13797) );
  INV_X1 U15890 ( .A(n13795), .ZN(n13796) );
  AOI22_X1 U15891 ( .A1(n13819), .A2(n13820), .B1(n13797), .B2(n13796), .ZN(
        n13809) );
  MUX2_X1 U15892 ( .A(n13799), .B(n13798), .S(n13810), .Z(n13814) );
  INV_X1 U15893 ( .A(n13799), .ZN(n13890) );
  MUX2_X1 U15894 ( .A(n13890), .B(n14203), .S(n6532), .Z(n13813) );
  NAND2_X1 U15895 ( .A1(n13814), .A2(n13813), .ZN(n13822) );
  NAND2_X1 U15896 ( .A1(n9913), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13801) );
  MUX2_X1 U15897 ( .A(n13889), .B(n13942), .S(n13792), .Z(n13816) );
  NAND2_X1 U15898 ( .A1(n13792), .A2(n13933), .ZN(n13830) );
  OAI211_X1 U15899 ( .C1(n13803), .C2(n10080), .A(n13877), .B(n13835), .ZN(
        n13804) );
  INV_X1 U15900 ( .A(n13804), .ZN(n13806) );
  INV_X1 U15901 ( .A(n13889), .ZN(n13805) );
  AOI21_X1 U15902 ( .B1(n13830), .B2(n13806), .A(n13805), .ZN(n13807) );
  AOI21_X1 U15903 ( .B1(n13942), .B2(n13810), .A(n13807), .ZN(n13815) );
  NAND2_X1 U15904 ( .A1(n13816), .A2(n13815), .ZN(n13824) );
  INV_X1 U15905 ( .A(n13933), .ZN(n13812) );
  MUX2_X1 U15906 ( .A(n13933), .B(n13808), .S(n14196), .Z(n13811) );
  OAI21_X1 U15907 ( .B1(n13812), .B2(n6533), .A(n13811), .ZN(n13818) );
  OAI22_X1 U15908 ( .A1(n13816), .A2(n13815), .B1(n13814), .B2(n13813), .ZN(
        n13817) );
  NAND2_X1 U15909 ( .A1(n13818), .A2(n13817), .ZN(n13827) );
  INV_X1 U15910 ( .A(n13819), .ZN(n13823) );
  INV_X1 U15911 ( .A(n13820), .ZN(n13821) );
  NAND4_X1 U15912 ( .A1(n13841), .A2(n13823), .A3(n13822), .A4(n13821), .ZN(
        n13826) );
  INV_X1 U15913 ( .A(n13824), .ZN(n13825) );
  AOI21_X1 U15914 ( .B1(n13827), .B2(n13826), .A(n13825), .ZN(n13828) );
  MUX2_X1 U15915 ( .A(n13933), .B(n13792), .S(n14196), .Z(n13829) );
  INV_X1 U15916 ( .A(n13829), .ZN(n13832) );
  INV_X1 U15917 ( .A(n13830), .ZN(n13831) );
  MUX2_X1 U15918 ( .A(n13877), .B(n13884), .S(n13833), .Z(n13834) );
  INV_X1 U15919 ( .A(n13835), .ZN(n13837) );
  AOI211_X1 U15920 ( .C1(n13877), .C2(n14152), .A(n13837), .B(n13638), .ZN(
        n13838) );
  INV_X1 U15921 ( .A(n13841), .ZN(n13875) );
  INV_X1 U15922 ( .A(n13955), .ZN(n13871) );
  NAND2_X1 U15923 ( .A1(n13843), .A2(n13842), .ZN(n13982) );
  INV_X1 U15924 ( .A(n13844), .ZN(n14065) );
  NAND4_X1 U15925 ( .A1(n13847), .A2(n10080), .A3(n13846), .A4(n13845), .ZN(
        n13849) );
  NOR4_X1 U15926 ( .A1(n13851), .A2(n13850), .A3(n13849), .A4(n13848), .ZN(
        n13855) );
  NAND4_X1 U15927 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        n13857) );
  NOR2_X1 U15928 ( .A1(n13857), .A2(n13856), .ZN(n13859) );
  NAND3_X1 U15929 ( .A1(n13860), .A2(n13859), .A3(n13858), .ZN(n13863) );
  NOR3_X1 U15930 ( .A1(n13863), .A2(n13862), .A3(n14189), .ZN(n13865) );
  INV_X1 U15931 ( .A(n14130), .ZN(n14124) );
  NAND4_X1 U15932 ( .A1(n13866), .A2(n13865), .A3(n14124), .A4(n13864), .ZN(
        n13867) );
  NOR4_X1 U15933 ( .A1(n12504), .A2(n14165), .A3(n13867), .A4(n14089), .ZN(
        n13868) );
  NAND4_X1 U15934 ( .A1(n14044), .A2(n14065), .A3(n13868), .A4(n14076), .ZN(
        n13869) );
  NOR4_X1 U15935 ( .A1(n13982), .A2(n14012), .A3(n14029), .A4(n13869), .ZN(
        n13870) );
  NAND4_X1 U15936 ( .A1(n13871), .A2(n13870), .A3(n13959), .A4(n13994), .ZN(
        n13874) );
  XOR2_X1 U15937 ( .A(n13889), .B(n13942), .Z(n13873) );
  NOR4_X1 U15938 ( .A1(n13875), .A2(n13874), .A3(n13873), .A4(n13872), .ZN(
        n13876) );
  XNOR2_X1 U15939 ( .A(n13876), .B(n9912), .ZN(n13878) );
  NOR3_X1 U15940 ( .A1(n13878), .A2(n13877), .A3(n13887), .ZN(n13879) );
  OAI21_X1 U15941 ( .B1(n13880), .B2(n10080), .A(n13879), .ZN(n13886) );
  NAND3_X1 U15942 ( .A1(n13882), .A2(n13881), .A3(n14106), .ZN(n13883) );
  OAI211_X1 U15943 ( .C1(n13884), .C2(n13887), .A(n13883), .B(P2_B_REG_SCAN_IN), .ZN(n13885) );
  OAI211_X1 U15944 ( .C1(n13888), .C2(n13887), .A(n13886), .B(n13885), .ZN(
        P2_U3328) );
  MUX2_X1 U15945 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13933), .S(n13907), .Z(
        P2_U3562) );
  MUX2_X1 U15946 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13889), .S(n13907), .Z(
        P2_U3561) );
  MUX2_X1 U15947 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13890), .S(n13907), .Z(
        P2_U3560) );
  MUX2_X1 U15948 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13961), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15949 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13891), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15950 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13999), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15951 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n14007), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15952 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13998), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15953 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n14041), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15954 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14058), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15955 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n14081), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15956 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n14057), .S(n13907), .Z(
        P2_U3551) );
  CLKBUF_X2 U15957 ( .A(P2_U3947), .Z(n13907) );
  MUX2_X1 U15958 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n14109), .S(n13907), .Z(
        P2_U3550) );
  MUX2_X1 U15959 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13892), .S(n13907), .Z(
        P2_U3549) );
  MUX2_X1 U15960 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n14107), .S(n13907), .Z(
        P2_U3548) );
  MUX2_X1 U15961 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13893), .S(n13907), .Z(
        P2_U3547) );
  MUX2_X1 U15962 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13894), .S(n13907), .Z(
        P2_U3546) );
  MUX2_X1 U15963 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13895), .S(n13907), .Z(
        P2_U3545) );
  MUX2_X1 U15964 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13896), .S(n13907), .Z(
        P2_U3544) );
  MUX2_X1 U15965 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13897), .S(n13907), .Z(
        P2_U3543) );
  MUX2_X1 U15966 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13898), .S(n13907), .Z(
        P2_U3542) );
  MUX2_X1 U15967 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13899), .S(n13907), .Z(
        P2_U3541) );
  MUX2_X1 U15968 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13900), .S(n13907), .Z(
        P2_U3540) );
  MUX2_X1 U15969 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n6832), .S(n13907), .Z(
        P2_U3539) );
  MUX2_X1 U15970 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13901), .S(n13907), .Z(
        P2_U3538) );
  MUX2_X1 U15971 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13902), .S(n13907), .Z(
        P2_U3537) );
  MUX2_X1 U15972 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13903), .S(n13907), .Z(
        P2_U3536) );
  MUX2_X1 U15973 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13904), .S(n13907), .Z(
        P2_U3535) );
  MUX2_X1 U15974 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13905), .S(n13907), .Z(
        P2_U3534) );
  MUX2_X1 U15975 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13906), .S(n13907), .Z(
        P2_U3533) );
  MUX2_X1 U15976 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6543), .S(n13907), .Z(
        P2_U3532) );
  MUX2_X1 U15977 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n10686), .S(n13907), .Z(
        P2_U3531) );
  AOI22_X1 U15978 ( .A1(n15408), .A2(P2_ADDR_REG_7__SCAN_IN), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(P2_U3088), .ZN(n13921) );
  NAND2_X1 U15979 ( .A1(n13908), .A2(n13913), .ZN(n13920) );
  MUX2_X1 U15980 ( .A(n11729), .B(P2_REG2_REG_7__SCAN_IN), .S(n13913), .Z(
        n13909) );
  NAND3_X1 U15981 ( .A1(n15381), .A2(n13910), .A3(n13909), .ZN(n13911) );
  NAND3_X1 U15982 ( .A1(n15394), .A2(n13912), .A3(n13911), .ZN(n13919) );
  MUX2_X1 U15983 ( .A(n10610), .B(P2_REG1_REG_7__SCAN_IN), .S(n13913), .Z(
        n13914) );
  NAND3_X1 U15984 ( .A1(n15378), .A2(n13915), .A3(n13914), .ZN(n13916) );
  NAND3_X1 U15985 ( .A1(n15398), .A2(n13917), .A3(n13916), .ZN(n13918) );
  NAND4_X1 U15986 ( .A1(n13921), .A2(n13920), .A3(n13919), .A4(n13918), .ZN(
        P2_U3221) );
  INV_X1 U15987 ( .A(n13922), .ZN(n13923) );
  AOI21_X1 U15988 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13924), .A(n13923), 
        .ZN(n13932) );
  XOR2_X1 U15989 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13925), .Z(n13930) );
  NAND2_X1 U15990 ( .A1(n15408), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n13927) );
  OAI211_X1 U15991 ( .C1(n15412), .C2(n13928), .A(n13927), .B(n13926), .ZN(
        n13929) );
  AOI21_X1 U15992 ( .B1(n13930), .B2(n15398), .A(n13929), .ZN(n13931) );
  OAI21_X1 U15993 ( .B1(n13932), .B2(n15414), .A(n13931), .ZN(P2_U3232) );
  NAND2_X1 U15994 ( .A1(n14201), .A2(n13938), .ZN(n13937) );
  XNOR2_X1 U15995 ( .A(n14196), .B(n13937), .ZN(n14198) );
  NAND2_X1 U15996 ( .A1(n13934), .A2(n13933), .ZN(n14199) );
  NOR2_X1 U15997 ( .A1(n14186), .A2(n14199), .ZN(n13940) );
  AOI21_X1 U15998 ( .B1(n14186), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13940), 
        .ZN(n13936) );
  NAND2_X1 U15999 ( .A1(n14196), .A2(n14169), .ZN(n13935) );
  OAI211_X1 U16000 ( .C1(n14198), .C2(n14052), .A(n13936), .B(n13935), .ZN(
        P2_U3234) );
  OAI211_X1 U16001 ( .C1(n14201), .C2(n13938), .A(n14308), .B(n13937), .ZN(
        n14200) );
  NOR2_X1 U16002 ( .A1(n14135), .A2(n13939), .ZN(n13941) );
  AOI211_X1 U16003 ( .C1(n13942), .C2(n14169), .A(n13941), .B(n13940), .ZN(
        n13943) );
  OAI21_X1 U16004 ( .B1(n14200), .B2(n14173), .A(n13943), .ZN(P2_U3235) );
  AOI21_X1 U16005 ( .B1(n13944), .B2(n13955), .A(n14162), .ZN(n13947) );
  NAND2_X1 U16006 ( .A1(n14207), .A2(n13963), .ZN(n13948) );
  OAI22_X1 U16007 ( .A1(n13950), .A2(n14146), .B1(n13949), .B2(n14135), .ZN(
        n13951) );
  INV_X1 U16008 ( .A(n13951), .ZN(n13952) );
  OAI21_X1 U16009 ( .B1(n13953), .B2(n14188), .A(n13952), .ZN(n13957) );
  NOR2_X1 U16010 ( .A1(n14210), .A2(n14191), .ZN(n13956) );
  OAI21_X1 U16011 ( .B1(n14209), .B2(n14186), .A(n13958), .ZN(P2_U3237) );
  XNOR2_X1 U16012 ( .A(n13960), .B(n13959), .ZN(n13962) );
  INV_X1 U16013 ( .A(n13973), .ZN(n13965) );
  INV_X1 U16014 ( .A(n13963), .ZN(n13964) );
  AOI21_X1 U16015 ( .B1(n14211), .B2(n13965), .A(n13964), .ZN(n14212) );
  AOI22_X1 U16016 ( .A1(n13966), .A2(n14184), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14186), .ZN(n13967) );
  OAI21_X1 U16017 ( .B1(n13968), .B2(n14188), .A(n13967), .ZN(n13969) );
  AOI21_X1 U16018 ( .B1(n14212), .B2(n14122), .A(n13969), .ZN(n13972) );
  NAND3_X1 U16019 ( .A1(n14214), .A2(n14213), .A3(n14019), .ZN(n13971) );
  OAI211_X1 U16020 ( .C1(n14217), .C2(n14186), .A(n13972), .B(n13971), .ZN(
        P2_U3238) );
  INV_X1 U16021 ( .A(n13988), .ZN(n13974) );
  AOI211_X1 U16022 ( .C1(n14220), .C2(n13974), .A(n15453), .B(n13973), .ZN(
        n14219) );
  XNOR2_X1 U16023 ( .A(n13975), .B(n13982), .ZN(n13976) );
  OAI222_X1 U16024 ( .A1(n14094), .A2(n13978), .B1(n14092), .B2(n13977), .C1(
        n13976), .C2(n14162), .ZN(n14218) );
  AOI21_X1 U16025 ( .B1(n14219), .B2(n14152), .A(n14218), .ZN(n13986) );
  INV_X1 U16026 ( .A(n13979), .ZN(n13980) );
  OAI22_X1 U16027 ( .A1(n13980), .A2(n14146), .B1(n15583), .B2(n14135), .ZN(
        n13984) );
  XOR2_X1 U16028 ( .A(n13982), .B(n13981), .Z(n14223) );
  NOR2_X1 U16029 ( .A1(n14223), .A2(n14191), .ZN(n13983) );
  AOI211_X1 U16030 ( .C1(n14169), .C2(n14220), .A(n13984), .B(n13983), .ZN(
        n13985) );
  OAI21_X1 U16031 ( .B1(n13986), .B2(n14186), .A(n13985), .ZN(P2_U3239) );
  XOR2_X1 U16032 ( .A(n13987), .B(n13994), .Z(n14228) );
  AOI211_X1 U16033 ( .C1(n14225), .C2(n14013), .A(n15453), .B(n13988), .ZN(
        n14224) );
  INV_X1 U16034 ( .A(n14225), .ZN(n13992) );
  INV_X1 U16035 ( .A(n13989), .ZN(n13990) );
  AOI22_X1 U16036 ( .A1(n13990), .A2(n14184), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14186), .ZN(n13991) );
  OAI21_X1 U16037 ( .B1(n13992), .B2(n14188), .A(n13991), .ZN(n14002) );
  INV_X1 U16038 ( .A(n13994), .ZN(n13996) );
  NAND3_X1 U16039 ( .A1(n14004), .A2(n13996), .A3(n13995), .ZN(n13997) );
  NAND2_X1 U16040 ( .A1(n13993), .A2(n13997), .ZN(n14000) );
  AOI222_X1 U16041 ( .A1(n14180), .A2(n14000), .B1(n13999), .B2(n14108), .C1(
        n13998), .C2(n14106), .ZN(n14227) );
  NOR2_X1 U16042 ( .A1(n14227), .A2(n14186), .ZN(n14001) );
  OAI21_X1 U16043 ( .B1(n14228), .B2(n14191), .A(n14003), .ZN(P2_U3240) );
  OAI21_X1 U16044 ( .B1(n14006), .B2(n14005), .A(n14004), .ZN(n14008) );
  AOI222_X1 U16045 ( .A1(n14180), .A2(n14008), .B1(n14041), .B2(n14106), .C1(
        n14007), .C2(n14108), .ZN(n14232) );
  AND2_X1 U16046 ( .A1(n14028), .A2(n14009), .ZN(n14011) );
  OAI21_X1 U16047 ( .B1(n14012), .B2(n14011), .A(n14010), .ZN(n14233) );
  INV_X1 U16048 ( .A(n14233), .ZN(n14020) );
  AOI21_X1 U16049 ( .B1(n6616), .B2(n14230), .A(n15453), .ZN(n14014) );
  AND2_X1 U16050 ( .A1(n14014), .A2(n14013), .ZN(n14229) );
  NAND2_X1 U16051 ( .A1(n14229), .A2(n14194), .ZN(n14017) );
  AOI22_X1 U16052 ( .A1(n14015), .A2(n14184), .B1(n14186), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n14016) );
  OAI211_X1 U16053 ( .C1(n7588), .C2(n14188), .A(n14017), .B(n14016), .ZN(
        n14018) );
  AOI21_X1 U16054 ( .B1(n14020), .B2(n14019), .A(n14018), .ZN(n14021) );
  OAI21_X1 U16055 ( .B1(n14232), .B2(n14186), .A(n14021), .ZN(P2_U3241) );
  XOR2_X1 U16056 ( .A(n14029), .B(n14022), .Z(n14023) );
  OAI222_X1 U16057 ( .A1(n14094), .A2(n14025), .B1(n14092), .B2(n14024), .C1(
        n14023), .C2(n14162), .ZN(n14236) );
  INV_X1 U16058 ( .A(n14236), .ZN(n14038) );
  AND2_X1 U16059 ( .A1(n14026), .A2(n14027), .ZN(n14030) );
  OAI21_X1 U16060 ( .B1(n14030), .B2(n14029), .A(n14028), .ZN(n14238) );
  OAI211_X1 U16061 ( .C1(n14047), .C2(n14235), .A(n14308), .B(n6616), .ZN(
        n14234) );
  OAI22_X1 U16062 ( .A1(n14032), .A2(n14135), .B1(n14031), .B2(n14146), .ZN(
        n14033) );
  AOI21_X1 U16063 ( .B1(n14034), .B2(n14169), .A(n14033), .ZN(n14035) );
  OAI21_X1 U16064 ( .B1(n14234), .B2(n14173), .A(n14035), .ZN(n14036) );
  AOI21_X1 U16065 ( .B1(n14238), .B2(n14019), .A(n14036), .ZN(n14037) );
  OAI21_X1 U16066 ( .B1(n14038), .B2(n14186), .A(n14037), .ZN(P2_U3242) );
  OAI211_X1 U16067 ( .C1(n14040), .C2(n14044), .A(n14039), .B(n14180), .ZN(
        n14043) );
  AOI22_X1 U16068 ( .A1(n14041), .A2(n14108), .B1(n14106), .B2(n14081), .ZN(
        n14042) );
  NAND2_X1 U16069 ( .A1(n14043), .A2(n14042), .ZN(n14245) );
  NAND2_X1 U16070 ( .A1(n14045), .A2(n14044), .ZN(n14240) );
  AND3_X1 U16071 ( .A1(n14026), .A2(n14019), .A3(n14240), .ZN(n14054) );
  NOR2_X1 U16072 ( .A1(n14060), .A2(n14241), .ZN(n14046) );
  OR2_X1 U16073 ( .A1(n14047), .A2(n14046), .ZN(n14242) );
  AOI22_X1 U16074 ( .A1(n14186), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14048), 
        .B2(n14184), .ZN(n14051) );
  NAND2_X1 U16075 ( .A1(n14049), .A2(n14169), .ZN(n14050) );
  OAI211_X1 U16076 ( .C1(n14242), .C2(n14052), .A(n14051), .B(n14050), .ZN(
        n14053) );
  AOI211_X1 U16077 ( .C1(n14245), .C2(n14135), .A(n14054), .B(n14053), .ZN(
        n14055) );
  INV_X1 U16078 ( .A(n14055), .ZN(P2_U3243) );
  XNOR2_X1 U16079 ( .A(n14056), .B(n14065), .ZN(n14059) );
  AOI222_X1 U16080 ( .A1(n14180), .A2(n14059), .B1(n14058), .B2(n14108), .C1(
        n14057), .C2(n14106), .ZN(n14249) );
  AOI21_X1 U16081 ( .B1(n14246), .B2(n14071), .A(n14060), .ZN(n14247) );
  INV_X1 U16082 ( .A(n14061), .ZN(n14062) );
  AOI22_X1 U16083 ( .A1(n14186), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14062), 
        .B2(n14184), .ZN(n14063) );
  OAI21_X1 U16084 ( .B1(n14064), .B2(n14188), .A(n14063), .ZN(n14068) );
  XNOR2_X1 U16085 ( .A(n14066), .B(n14065), .ZN(n14250) );
  NOR2_X1 U16086 ( .A1(n14250), .A2(n14191), .ZN(n14067) );
  AOI211_X1 U16087 ( .C1(n14247), .C2(n14122), .A(n14068), .B(n14067), .ZN(
        n14069) );
  OAI21_X1 U16088 ( .B1(n14249), .B2(n14186), .A(n14069), .ZN(P2_U3244) );
  XOR2_X1 U16089 ( .A(n14070), .B(n14076), .Z(n14255) );
  AOI211_X1 U16090 ( .C1(n14252), .C2(n14095), .A(n15453), .B(n12543), .ZN(
        n14251) );
  INV_X1 U16091 ( .A(n14072), .ZN(n14073) );
  AOI22_X1 U16092 ( .A1(n14186), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14073), 
        .B2(n14184), .ZN(n14074) );
  OAI21_X1 U16093 ( .B1(n14075), .B2(n14188), .A(n14074), .ZN(n14084) );
  INV_X1 U16094 ( .A(n14076), .ZN(n14078) );
  NAND2_X1 U16095 ( .A1(n14078), .A2(n14077), .ZN(n14080) );
  OAI21_X1 U16096 ( .B1(n14087), .B2(n14080), .A(n14079), .ZN(n14082) );
  AOI222_X1 U16097 ( .A1(n14180), .A2(n14082), .B1(n14081), .B2(n14108), .C1(
        n14109), .C2(n14106), .ZN(n14254) );
  NOR2_X1 U16098 ( .A1(n14254), .A2(n14186), .ZN(n14083) );
  AOI211_X1 U16099 ( .C1(n14251), .C2(n14194), .A(n14084), .B(n14083), .ZN(
        n14085) );
  OAI21_X1 U16100 ( .B1(n14255), .B2(n14191), .A(n14085), .ZN(P2_U3245) );
  XOR2_X1 U16101 ( .A(n14086), .B(n14089), .Z(n14261) );
  AOI21_X1 U16102 ( .B1(n14089), .B2(n14088), .A(n14087), .ZN(n14090) );
  OAI222_X1 U16103 ( .A1(n14094), .A2(n14093), .B1(n14092), .B2(n14091), .C1(
        n14162), .C2(n14090), .ZN(n14256) );
  NAND2_X1 U16104 ( .A1(n14256), .A2(n14135), .ZN(n14104) );
  INV_X1 U16105 ( .A(n14112), .ZN(n14097) );
  INV_X1 U16106 ( .A(n14095), .ZN(n14096) );
  AOI21_X1 U16107 ( .B1(n14257), .B2(n14097), .A(n14096), .ZN(n14258) );
  NOR2_X1 U16108 ( .A1(n14098), .A2(n14188), .ZN(n14102) );
  OAI22_X1 U16109 ( .A1(n14135), .A2(n14100), .B1(n14099), .B2(n14146), .ZN(
        n14101) );
  AOI211_X1 U16110 ( .C1(n14258), .C2(n14122), .A(n14102), .B(n14101), .ZN(
        n14103) );
  OAI211_X1 U16111 ( .C1(n14261), .C2(n14191), .A(n14104), .B(n14103), .ZN(
        P2_U3246) );
  XNOR2_X1 U16112 ( .A(n14105), .B(n12504), .ZN(n14110) );
  AOI222_X1 U16113 ( .A1(n14180), .A2(n14110), .B1(n14109), .B2(n14108), .C1(
        n14107), .C2(n14106), .ZN(n14265) );
  AND2_X1 U16114 ( .A1(n14139), .A2(n14262), .ZN(n14111) );
  NOR2_X1 U16115 ( .A1(n14112), .A2(n14111), .ZN(n14263) );
  AOI22_X1 U16116 ( .A1(n14186), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14113), 
        .B2(n14184), .ZN(n14114) );
  OAI21_X1 U16117 ( .B1(n14115), .B2(n14188), .A(n14114), .ZN(n14121) );
  INV_X1 U16118 ( .A(n14116), .ZN(n14117) );
  AOI21_X1 U16119 ( .B1(n14119), .B2(n14118), .A(n14117), .ZN(n14266) );
  NOR2_X1 U16120 ( .A1(n14266), .A2(n14191), .ZN(n14120) );
  AOI211_X1 U16121 ( .C1(n14263), .C2(n14122), .A(n14121), .B(n14120), .ZN(
        n14123) );
  OAI21_X1 U16122 ( .B1(n14265), .B2(n14186), .A(n14123), .ZN(P2_U3247) );
  XNOR2_X1 U16123 ( .A(n14125), .B(n14124), .ZN(n14128) );
  INV_X1 U16124 ( .A(n14126), .ZN(n14127) );
  AOI21_X1 U16125 ( .B1(n14128), .B2(n14180), .A(n14127), .ZN(n14270) );
  OAI21_X1 U16126 ( .B1(n14131), .B2(n14130), .A(n14129), .ZN(n14271) );
  INV_X1 U16127 ( .A(n14132), .ZN(n14133) );
  OAI22_X1 U16128 ( .A1(n14135), .A2(n14134), .B1(n14133), .B2(n14146), .ZN(
        n14136) );
  AOI21_X1 U16129 ( .B1(n14268), .B2(n14169), .A(n14136), .ZN(n14141) );
  AOI21_X1 U16130 ( .B1(n14144), .B2(n14268), .A(n15453), .ZN(n14138) );
  AND2_X1 U16131 ( .A1(n14139), .A2(n14138), .ZN(n14267) );
  NAND2_X1 U16132 ( .A1(n14267), .A2(n14194), .ZN(n14140) );
  OAI211_X1 U16133 ( .C1(n14271), .C2(n14191), .A(n14141), .B(n14140), .ZN(
        n14142) );
  INV_X1 U16134 ( .A(n14142), .ZN(n14143) );
  OAI21_X1 U16135 ( .B1(n14270), .B2(n14186), .A(n14143), .ZN(P2_U3248) );
  AOI211_X1 U16136 ( .C1(n14274), .C2(n6565), .A(n15453), .B(n14137), .ZN(
        n14272) );
  INV_X1 U16137 ( .A(n14273), .ZN(n14145) );
  OAI21_X1 U16138 ( .B1(n14147), .B2(n14146), .A(n14145), .ZN(n14151) );
  XNOR2_X1 U16139 ( .A(n14148), .B(n14153), .ZN(n14149) );
  NAND2_X1 U16140 ( .A1(n14149), .A2(n14180), .ZN(n14278) );
  INV_X1 U16141 ( .A(n14278), .ZN(n14150) );
  AOI211_X1 U16142 ( .C1(n14272), .C2(n14152), .A(n14151), .B(n14150), .ZN(
        n14158) );
  AOI22_X1 U16143 ( .A1(n14274), .A2(n14169), .B1(P2_REG2_REG_16__SCAN_IN), 
        .B2(n14186), .ZN(n14157) );
  OR2_X1 U16144 ( .A1(n14154), .A2(n14153), .ZN(n14275) );
  NAND3_X1 U16145 ( .A1(n14275), .A2(n14019), .A3(n14155), .ZN(n14156) );
  OAI211_X1 U16146 ( .C1(n14158), .C2(n14186), .A(n14157), .B(n14156), .ZN(
        P2_U3249) );
  XOR2_X1 U16147 ( .A(n14160), .B(n14165), .Z(n14163) );
  OAI21_X1 U16148 ( .B1(n14163), .B2(n14162), .A(n14161), .ZN(n14281) );
  INV_X1 U16149 ( .A(n14281), .ZN(n14176) );
  OAI21_X1 U16150 ( .B1(n14166), .B2(n14165), .A(n14164), .ZN(n14283) );
  OAI211_X1 U16151 ( .C1(n14167), .C2(n14280), .A(n14308), .B(n6565), .ZN(
        n14279) );
  AOI22_X1 U16152 ( .A1(n14186), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n14168), 
        .B2(n14184), .ZN(n14172) );
  NAND2_X1 U16153 ( .A1(n14170), .A2(n14169), .ZN(n14171) );
  OAI211_X1 U16154 ( .C1(n14279), .C2(n14173), .A(n14172), .B(n14171), .ZN(
        n14174) );
  AOI21_X1 U16155 ( .B1(n14283), .B2(n14019), .A(n14174), .ZN(n14175) );
  OAI21_X1 U16156 ( .B1(n14176), .B2(n14186), .A(n14175), .ZN(P2_U3250) );
  XNOR2_X1 U16157 ( .A(n14177), .B(n14189), .ZN(n14181) );
  INV_X1 U16158 ( .A(n14178), .ZN(n14179) );
  AOI21_X1 U16159 ( .B1(n14181), .B2(n14180), .A(n14179), .ZN(n14294) );
  AOI211_X1 U16160 ( .C1(n14292), .C2(n14183), .A(n15453), .B(n14182), .ZN(
        n14291) );
  AOI22_X1 U16161 ( .A1(n14186), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n14185), 
        .B2(n14184), .ZN(n14187) );
  OAI21_X1 U16162 ( .B1(n7578), .B2(n14188), .A(n14187), .ZN(n14193) );
  XNOR2_X1 U16163 ( .A(n14190), .B(n14189), .ZN(n14295) );
  NOR2_X1 U16164 ( .A1(n14295), .A2(n14191), .ZN(n14192) );
  AOI211_X1 U16165 ( .C1(n14291), .C2(n14194), .A(n14193), .B(n14192), .ZN(
        n14195) );
  OAI21_X1 U16166 ( .B1(n14294), .B2(n14186), .A(n14195), .ZN(P2_U3252) );
  NAND2_X1 U16167 ( .A1(n14196), .A2(n14315), .ZN(n14197) );
  OAI211_X1 U16168 ( .C1(n14198), .C2(n15453), .A(n14199), .B(n14197), .ZN(
        n14321) );
  MUX2_X1 U16169 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14321), .S(n15466), .Z(
        P2_U3530) );
  OAI211_X1 U16170 ( .C1(n14201), .C2(n15451), .A(n14200), .B(n14199), .ZN(
        n14322) );
  MUX2_X1 U16171 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14322), .S(n15466), .Z(
        P2_U3529) );
  AOI21_X1 U16172 ( .B1(n14315), .B2(n14203), .A(n14202), .ZN(n14204) );
  AOI21_X1 U16173 ( .B1(n14315), .B2(n14207), .A(n14206), .ZN(n14208) );
  AOI22_X1 U16174 ( .A1(n14212), .A2(n14308), .B1(n14315), .B2(n14211), .ZN(
        n14216) );
  NAND3_X1 U16175 ( .A1(n14214), .A2(n14213), .A3(n15458), .ZN(n14215) );
  MUX2_X1 U16176 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14324), .S(n15466), .Z(
        P2_U3526) );
  INV_X1 U16177 ( .A(n14218), .ZN(n14222) );
  AOI21_X1 U16178 ( .B1(n14315), .B2(n14220), .A(n14219), .ZN(n14221) );
  OAI211_X1 U16179 ( .C1(n14319), .C2(n14223), .A(n14222), .B(n14221), .ZN(
        n14325) );
  MUX2_X1 U16180 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14325), .S(n15466), .Z(
        P2_U3525) );
  AOI21_X1 U16181 ( .B1(n14315), .B2(n14225), .A(n14224), .ZN(n14226) );
  OAI211_X1 U16182 ( .C1(n14319), .C2(n14228), .A(n14227), .B(n14226), .ZN(
        n14326) );
  MUX2_X1 U16183 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14326), .S(n15466), .Z(
        P2_U3524) );
  AOI21_X1 U16184 ( .B1(n14315), .B2(n14230), .A(n14229), .ZN(n14231) );
  OAI211_X1 U16185 ( .C1(n14319), .C2(n14233), .A(n14232), .B(n14231), .ZN(
        n14327) );
  MUX2_X1 U16186 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14327), .S(n15466), .Z(
        P2_U3523) );
  OAI21_X1 U16187 ( .B1(n14235), .B2(n15451), .A(n14234), .ZN(n14237) );
  AOI211_X1 U16188 ( .C1(n15458), .C2(n14238), .A(n14237), .B(n14236), .ZN(
        n14239) );
  INV_X1 U16189 ( .A(n14239), .ZN(n14328) );
  MUX2_X1 U16190 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14328), .S(n15466), .Z(
        P2_U3522) );
  AND3_X1 U16191 ( .A1(n14026), .A2(n15458), .A3(n14240), .ZN(n14244) );
  OAI22_X1 U16192 ( .A1(n14242), .A2(n15453), .B1(n14241), .B2(n15451), .ZN(
        n14243) );
  MUX2_X1 U16193 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n14329), .S(n15466), .Z(
        P2_U3521) );
  AOI22_X1 U16194 ( .A1(n14247), .A2(n14308), .B1(n14315), .B2(n14246), .ZN(
        n14248) );
  OAI211_X1 U16195 ( .C1(n14319), .C2(n14250), .A(n14249), .B(n14248), .ZN(
        n14330) );
  MUX2_X1 U16196 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14330), .S(n15466), .Z(
        P2_U3520) );
  AOI21_X1 U16197 ( .B1(n14315), .B2(n14252), .A(n14251), .ZN(n14253) );
  OAI211_X1 U16198 ( .C1(n14319), .C2(n14255), .A(n14254), .B(n14253), .ZN(
        n14331) );
  MUX2_X1 U16199 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14331), .S(n15466), .Z(
        P2_U3519) );
  INV_X1 U16200 ( .A(n14256), .ZN(n14260) );
  AOI22_X1 U16201 ( .A1(n14258), .A2(n14308), .B1(n14315), .B2(n14257), .ZN(
        n14259) );
  OAI211_X1 U16202 ( .C1(n14319), .C2(n14261), .A(n14260), .B(n14259), .ZN(
        n14332) );
  MUX2_X1 U16203 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14332), .S(n15466), .Z(
        P2_U3518) );
  AOI22_X1 U16204 ( .A1(n14263), .A2(n14308), .B1(n14315), .B2(n14262), .ZN(
        n14264) );
  OAI211_X1 U16205 ( .C1(n14319), .C2(n14266), .A(n14265), .B(n14264), .ZN(
        n14333) );
  MUX2_X1 U16206 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14333), .S(n15466), .Z(
        P2_U3517) );
  AOI21_X1 U16207 ( .B1(n14315), .B2(n14268), .A(n14267), .ZN(n14269) );
  OAI211_X1 U16208 ( .C1(n14319), .C2(n14271), .A(n14270), .B(n14269), .ZN(
        n14334) );
  MUX2_X1 U16209 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14334), .S(n15466), .Z(
        P2_U3516) );
  AOI211_X1 U16210 ( .C1(n14315), .C2(n14274), .A(n14273), .B(n14272), .ZN(
        n14277) );
  NAND3_X1 U16211 ( .A1(n14275), .A2(n15458), .A3(n14155), .ZN(n14276) );
  NAND3_X1 U16212 ( .A1(n14278), .A2(n14277), .A3(n14276), .ZN(n14335) );
  MUX2_X1 U16213 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14335), .S(n15466), .Z(
        P2_U3515) );
  OAI21_X1 U16214 ( .B1(n14280), .B2(n15451), .A(n14279), .ZN(n14282) );
  AOI211_X1 U16215 ( .C1(n15458), .C2(n14283), .A(n14282), .B(n14281), .ZN(
        n14284) );
  INV_X1 U16216 ( .A(n14284), .ZN(n14336) );
  MUX2_X1 U16217 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14336), .S(n15466), .Z(
        P2_U3514) );
  OAI22_X1 U16218 ( .A1(n14286), .A2(n15453), .B1(n14285), .B2(n15451), .ZN(
        n14287) );
  INV_X1 U16219 ( .A(n14287), .ZN(n14288) );
  OAI211_X1 U16220 ( .C1(n14319), .C2(n14290), .A(n14289), .B(n14288), .ZN(
        n14337) );
  MUX2_X1 U16221 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14337), .S(n15466), .Z(
        P2_U3513) );
  AOI21_X1 U16222 ( .B1(n14315), .B2(n14292), .A(n14291), .ZN(n14293) );
  OAI211_X1 U16223 ( .C1(n14319), .C2(n14295), .A(n14294), .B(n14293), .ZN(
        n14338) );
  MUX2_X1 U16224 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14338), .S(n15466), .Z(
        P2_U3512) );
  AOI21_X1 U16225 ( .B1(n14315), .B2(n14297), .A(n14296), .ZN(n14298) );
  OAI211_X1 U16226 ( .C1(n14301), .C2(n14300), .A(n14299), .B(n14298), .ZN(
        n14339) );
  MUX2_X1 U16227 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14339), .S(n15466), .Z(
        P2_U3511) );
  AOI22_X1 U16228 ( .A1(n14303), .A2(n14308), .B1(n14315), .B2(n14302), .ZN(
        n14304) );
  OAI211_X1 U16229 ( .C1(n14319), .C2(n14306), .A(n14305), .B(n14304), .ZN(
        n14340) );
  MUX2_X1 U16230 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n14340), .S(n15466), .Z(
        P2_U3509) );
  AOI22_X1 U16231 ( .A1(n14309), .A2(n14308), .B1(n14315), .B2(n14307), .ZN(
        n14310) );
  OAI211_X1 U16232 ( .C1(n14319), .C2(n14312), .A(n14311), .B(n14310), .ZN(
        n14341) );
  MUX2_X1 U16233 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14341), .S(n15466), .Z(
        P2_U3508) );
  AOI21_X1 U16234 ( .B1(n14315), .B2(n14314), .A(n14313), .ZN(n14316) );
  OAI211_X1 U16235 ( .C1(n14319), .C2(n14318), .A(n14317), .B(n14316), .ZN(
        n14342) );
  MUX2_X1 U16236 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n14342), .S(n15466), .Z(
        P2_U3507) );
  MUX2_X1 U16237 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n14320), .S(n15466), .Z(
        P2_U3503) );
  MUX2_X1 U16238 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14321), .S(n15462), .Z(
        P2_U3498) );
  MUX2_X1 U16239 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14322), .S(n15462), .Z(
        P2_U3497) );
  MUX2_X1 U16240 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14324), .S(n15462), .Z(
        P2_U3494) );
  MUX2_X1 U16241 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14325), .S(n15462), .Z(
        P2_U3493) );
  MUX2_X1 U16242 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14326), .S(n15462), .Z(
        P2_U3492) );
  MUX2_X1 U16243 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14327), .S(n15462), .Z(
        P2_U3491) );
  MUX2_X1 U16244 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14328), .S(n15462), .Z(
        P2_U3490) );
  MUX2_X1 U16245 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14329), .S(n15462), .Z(
        P2_U3489) );
  MUX2_X1 U16246 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14330), .S(n15462), .Z(
        P2_U3488) );
  MUX2_X1 U16247 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14331), .S(n15462), .Z(
        P2_U3487) );
  MUX2_X1 U16248 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14332), .S(n15462), .Z(
        P2_U3486) );
  MUX2_X1 U16249 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14333), .S(n15462), .Z(
        P2_U3484) );
  MUX2_X1 U16250 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14334), .S(n15462), .Z(
        P2_U3481) );
  MUX2_X1 U16251 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14335), .S(n15462), .Z(
        P2_U3478) );
  MUX2_X1 U16252 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14336), .S(n15462), .Z(
        P2_U3475) );
  MUX2_X1 U16253 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14337), .S(n15462), .Z(
        P2_U3472) );
  MUX2_X1 U16254 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n14338), .S(n15462), .Z(
        P2_U3469) );
  MUX2_X1 U16255 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n14339), .S(n15462), .Z(
        P2_U3466) );
  MUX2_X1 U16256 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n14340), .S(n15462), .Z(
        P2_U3460) );
  MUX2_X1 U16257 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n14341), .S(n15462), .Z(
        P2_U3457) );
  MUX2_X1 U16258 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n14342), .S(n15462), .Z(
        P2_U3454) );
  INV_X1 U16259 ( .A(n15156), .ZN(n14351) );
  NAND4_X1 U16260 ( .A1(n14345), .A2(n14344), .A3(n14343), .A4(
        P2_IR_REG_31__SCAN_IN), .ZN(n14346) );
  NOR4_X1 U16261 ( .A1(n14348), .A2(n14347), .A3(P2_U3088), .A4(n14346), .ZN(
        n14349) );
  AOI21_X1 U16262 ( .B1(n14356), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14349), 
        .ZN(n14350) );
  OAI21_X1 U16263 ( .B1(n14351), .B2(n14360), .A(n14350), .ZN(P2_U3296) );
  INV_X1 U16264 ( .A(n14352), .ZN(n15159) );
  OAI222_X1 U16265 ( .A1(n15159), .A2(n14360), .B1(P2_U3088), .B2(n14354), 
        .C1(n14353), .C2(n14362), .ZN(P2_U3298) );
  INV_X1 U16266 ( .A(n14355), .ZN(n15162) );
  NAND2_X1 U16267 ( .A1(n14356), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14358) );
  OAI211_X1 U16268 ( .C1(n15162), .C2(n14360), .A(n14358), .B(n14357), .ZN(
        P2_U3299) );
  OAI222_X1 U16269 ( .A1(P2_U3088), .A2(n14363), .B1(n14362), .B2(n14361), 
        .C1(n14360), .C2(n14359), .ZN(P2_U3300) );
  MUX2_X1 U16270 ( .A(n7845), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XNOR2_X1 U16271 ( .A(n14365), .B(n14364), .ZN(n14372) );
  INV_X1 U16272 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14366) );
  OAI22_X1 U16273 ( .A1(n14367), .A2(n14528), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14366), .ZN(n14369) );
  NOR2_X1 U16274 ( .A1(n15110), .A2(n14524), .ZN(n14368) );
  AOI211_X1 U16275 ( .C1(n14497), .C2(n14370), .A(n14369), .B(n14368), .ZN(
        n14371) );
  OAI21_X1 U16276 ( .B1(n14372), .B2(n14546), .A(n14371), .ZN(P1_U3214) );
  NOR2_X1 U16277 ( .A1(n14426), .A2(n14373), .ZN(n14374) );
  NOR2_X1 U16278 ( .A1(n14375), .A2(n14374), .ZN(n14376) );
  AND2_X1 U16279 ( .A1(n14375), .A2(n14374), .ZN(n14427) );
  OAI21_X1 U16280 ( .B1(n14376), .B2(n14427), .A(n14515), .ZN(n14381) );
  OAI22_X1 U16281 ( .A1(n14435), .A2(n14909), .B1(n14377), .B2(n14907), .ZN(
        n14963) );
  NOR2_X1 U16282 ( .A1(n14528), .A2(n14968), .ZN(n14378) );
  AOI211_X1 U16283 ( .C1(n14497), .C2(n14963), .A(n14379), .B(n14378), .ZN(
        n14380) );
  OAI211_X1 U16284 ( .C1(n7500), .C2(n14524), .A(n14381), .B(n14380), .ZN(
        P1_U3215) );
  XOR2_X1 U16285 ( .A(n14383), .B(n14382), .Z(n14388) );
  AOI22_X1 U16286 ( .A1(n14552), .A2(n14940), .B1(n14939), .B2(n14554), .ZN(
        n14794) );
  NOR2_X1 U16287 ( .A1(n14794), .A2(n14458), .ZN(n14386) );
  OAI22_X1 U16288 ( .A1(n14791), .A2(n14528), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14384), .ZN(n14385) );
  AOI211_X1 U16289 ( .C1(n14800), .C2(n14544), .A(n14386), .B(n14385), .ZN(
        n14387) );
  OAI21_X1 U16290 ( .B1(n14388), .B2(n14546), .A(n14387), .ZN(P1_U3216) );
  AOI22_X1 U16291 ( .A1(n14556), .A2(n14940), .B1(n14939), .B2(n14558), .ZN(
        n14872) );
  NAND2_X1 U16292 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14696)
         );
  INV_X1 U16293 ( .A(n14876), .ZN(n14389) );
  NAND2_X1 U16294 ( .A1(n14539), .A2(n14389), .ZN(n14390) );
  OAI211_X1 U16295 ( .C1(n14872), .C2(n14458), .A(n14696), .B(n14390), .ZN(
        n14395) );
  AOI211_X1 U16296 ( .C1(n14393), .C2(n7102), .A(n14546), .B(n14391), .ZN(
        n14394) );
  AOI211_X1 U16297 ( .C1(n14875), .C2(n14544), .A(n14395), .B(n14394), .ZN(
        n14396) );
  INV_X1 U16298 ( .A(n14396), .ZN(P1_U3219) );
  OAI21_X1 U16299 ( .B1(n14399), .B2(n14398), .A(n14397), .ZN(n14400) );
  NAND2_X1 U16300 ( .A1(n14400), .A2(n14515), .ZN(n14408) );
  NAND2_X1 U16301 ( .A1(n14554), .A2(n14940), .ZN(n14403) );
  OR2_X1 U16302 ( .A1(n14401), .A2(n14907), .ZN(n14402) );
  NAND2_X1 U16303 ( .A1(n14403), .A2(n14402), .ZN(n14831) );
  INV_X1 U16304 ( .A(n14836), .ZN(n14405) );
  INV_X1 U16305 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14404) );
  OAI22_X1 U16306 ( .A1(n14405), .A2(n14528), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14404), .ZN(n14406) );
  AOI21_X1 U16307 ( .B1(n14831), .B2(n14497), .A(n14406), .ZN(n14407) );
  OAI211_X1 U16308 ( .C1(n15127), .C2(n14524), .A(n14408), .B(n14407), .ZN(
        P1_U3223) );
  AND2_X1 U16309 ( .A1(n14500), .A2(n14410), .ZN(n14413) );
  OAI211_X1 U16310 ( .C1(n14413), .C2(n14412), .A(n14515), .B(n14411), .ZN(
        n14419) );
  AOI21_X1 U16311 ( .B1(n14521), .B2(n14559), .A(n14414), .ZN(n14418) );
  AOI22_X1 U16312 ( .A1(n14539), .A2(n14415), .B1(n14538), .B2(n14561), .ZN(
        n14417) );
  NAND2_X1 U16313 ( .A1(n14974), .A2(n14544), .ZN(n14416) );
  NAND4_X1 U16314 ( .A1(n14419), .A2(n14418), .A3(n14417), .A4(n14416), .ZN(
        P1_U3224) );
  AOI22_X1 U16315 ( .A1(n14551), .A2(n14940), .B1(n14939), .B2(n14552), .ZN(
        n14762) );
  NOR2_X1 U16316 ( .A1(n14762), .A2(n14458), .ZN(n14423) );
  OAI22_X1 U16317 ( .A1(n14767), .A2(n14528), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14421), .ZN(n14422) );
  AOI211_X1 U16318 ( .C1(n14765), .C2(n14544), .A(n14423), .B(n14422), .ZN(
        n14424) );
  OAI21_X1 U16319 ( .B1(n14425), .B2(n14546), .A(n14424), .ZN(P1_U3225) );
  NOR2_X1 U16320 ( .A1(n14427), .A2(n14426), .ZN(n14429) );
  XOR2_X1 U16321 ( .A(n14428), .B(n14429), .Z(n14537) );
  AOI22_X1 U16322 ( .A1(n14537), .A2(n14536), .B1(n14429), .B2(n14428), .ZN(
        n14433) );
  NAND2_X1 U16323 ( .A1(n14431), .A2(n14430), .ZN(n14432) );
  XNOR2_X1 U16324 ( .A(n14433), .B(n14432), .ZN(n14439) );
  OAI21_X1 U16325 ( .B1(n14542), .B2(n14884), .A(n14434), .ZN(n14437) );
  INV_X1 U16326 ( .A(n14538), .ZN(n14518) );
  OAI22_X1 U16327 ( .A1(n14518), .A2(n14435), .B1(n14927), .B2(n14528), .ZN(
        n14436) );
  AOI211_X1 U16328 ( .C1(n15060), .C2(n14544), .A(n14437), .B(n14436), .ZN(
        n14438) );
  OAI21_X1 U16329 ( .B1(n14439), .B2(n14546), .A(n14438), .ZN(P1_U3226) );
  INV_X1 U16330 ( .A(n14443), .ZN(n14440) );
  NOR2_X1 U16331 ( .A1(n14441), .A2(n14440), .ZN(n14446) );
  AOI21_X1 U16332 ( .B1(n14444), .B2(n14443), .A(n14442), .ZN(n14445) );
  OAI21_X1 U16333 ( .B1(n14446), .B2(n14445), .A(n14515), .ZN(n14452) );
  INV_X1 U16334 ( .A(n14447), .ZN(n14448) );
  AOI21_X1 U16335 ( .B1(n14521), .B2(n14558), .A(n14448), .ZN(n14451) );
  AOI22_X1 U16336 ( .A1(n14539), .A2(n14911), .B1(n14538), .B2(n14941), .ZN(
        n14450) );
  NAND2_X1 U16337 ( .A1(n15055), .A2(n14544), .ZN(n14449) );
  NAND4_X1 U16338 ( .A1(n14452), .A2(n14451), .A3(n14450), .A4(n14449), .ZN(
        P1_U3228) );
  AND2_X1 U16339 ( .A1(n14553), .A2(n14939), .ZN(n14455) );
  AOI21_X1 U16340 ( .B1(n14747), .B2(n14940), .A(n14455), .ZN(n14776) );
  INV_X1 U16341 ( .A(n14456), .ZN(n14784) );
  AOI22_X1 U16342 ( .A1(n14784), .A2(n14539), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14457) );
  OAI21_X1 U16343 ( .B1(n14776), .B2(n14458), .A(n14457), .ZN(n14459) );
  AOI21_X1 U16344 ( .B1(n15117), .B2(n14544), .A(n14459), .ZN(n14460) );
  OAI211_X1 U16345 ( .C1(n14463), .C2(n14462), .A(n14461), .B(n14515), .ZN(
        n14470) );
  AOI22_X1 U16346 ( .A1(n14544), .A2(n14464), .B1(n14538), .B2(n14569), .ZN(
        n14469) );
  AOI22_X1 U16347 ( .A1(n14521), .A2(n14567), .B1(P1_REG3_REG_4__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14468) );
  INV_X1 U16348 ( .A(n14465), .ZN(n14466) );
  NAND2_X1 U16349 ( .A1(n14539), .A2(n14466), .ZN(n14467) );
  NAND4_X1 U16350 ( .A1(n14470), .A2(n14469), .A3(n14468), .A4(n14467), .ZN(
        P1_U3230) );
  AOI22_X1 U16351 ( .A1(n14555), .A2(n14940), .B1(n14939), .B2(n14557), .ZN(
        n15035) );
  INV_X1 U16352 ( .A(n15035), .ZN(n14859) );
  AOI22_X1 U16353 ( .A1(n14859), .A2(n14497), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14471) );
  OAI21_X1 U16354 ( .B1(n14472), .B2(n14528), .A(n14471), .ZN(n14476) );
  AOI211_X1 U16355 ( .C1(n14474), .C2(n14473), .A(n14546), .B(n6623), .ZN(
        n14475) );
  AOI211_X1 U16356 ( .C1(n14858), .C2(n14544), .A(n14476), .B(n14475), .ZN(
        n14477) );
  INV_X1 U16357 ( .A(n14477), .ZN(P1_U3233) );
  XNOR2_X1 U16358 ( .A(n14479), .B(n14478), .ZN(n14487) );
  NAND2_X1 U16359 ( .A1(n14939), .A2(n14560), .ZN(n14482) );
  OR2_X1 U16360 ( .A1(n14480), .A2(n14909), .ZN(n14481) );
  NAND2_X1 U16361 ( .A1(n14482), .A2(n14481), .ZN(n15073) );
  NAND2_X1 U16362 ( .A1(n14497), .A2(n15073), .ZN(n14483) );
  OAI211_X1 U16363 ( .C1(n14528), .C2(n14985), .A(n14484), .B(n14483), .ZN(
        n14485) );
  AOI21_X1 U16364 ( .B1(n14984), .B2(n14544), .A(n14485), .ZN(n14486) );
  OAI21_X1 U16365 ( .B1(n14487), .B2(n14546), .A(n14486), .ZN(P1_U3234) );
  OAI21_X1 U16366 ( .B1(n14490), .B2(n14489), .A(n14488), .ZN(n14491) );
  NAND2_X1 U16367 ( .A1(n14491), .A2(n14515), .ZN(n14499) );
  NAND2_X1 U16368 ( .A1(n14553), .A2(n14940), .ZN(n14493) );
  NAND2_X1 U16369 ( .A1(n14555), .A2(n14939), .ZN(n14492) );
  NAND2_X1 U16370 ( .A1(n14493), .A2(n14492), .ZN(n15025) );
  INV_X1 U16371 ( .A(n14814), .ZN(n14495) );
  OAI22_X1 U16372 ( .A1(n14495), .A2(n14528), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14494), .ZN(n14496) );
  AOI21_X1 U16373 ( .B1(n15025), .B2(n14497), .A(n14496), .ZN(n14498) );
  OAI211_X1 U16374 ( .C1(n14524), .C2(n14817), .A(n14499), .B(n14498), .ZN(
        P1_U3235) );
  OAI21_X1 U16375 ( .B1(n14502), .B2(n14501), .A(n14500), .ZN(n14503) );
  NAND2_X1 U16376 ( .A1(n14503), .A2(n14515), .ZN(n14511) );
  AOI21_X1 U16377 ( .B1(n14521), .B2(n14560), .A(n14504), .ZN(n14510) );
  INV_X1 U16378 ( .A(n14505), .ZN(n14506) );
  AOI22_X1 U16379 ( .A1(n14539), .A2(n14506), .B1(n14538), .B2(n14562), .ZN(
        n14509) );
  NAND2_X1 U16380 ( .A1(n14544), .A2(n14507), .ZN(n14508) );
  NAND4_X1 U16381 ( .A1(n14511), .A2(n14510), .A3(n14509), .A4(n14508), .ZN(
        P1_U3236) );
  OAI21_X1 U16382 ( .B1(n14514), .B2(n14513), .A(n14512), .ZN(n14516) );
  NAND2_X1 U16383 ( .A1(n14516), .A2(n14515), .ZN(n14523) );
  NAND2_X1 U16384 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14690)
         );
  INV_X1 U16385 ( .A(n14690), .ZN(n14520) );
  INV_X1 U16386 ( .A(n14892), .ZN(n14517) );
  OAI22_X1 U16387 ( .A1(n14518), .A2(n14884), .B1(n14517), .B2(n14528), .ZN(
        n14519) );
  AOI211_X1 U16388 ( .C1(n14521), .C2(n14557), .A(n14520), .B(n14519), .ZN(
        n14522) );
  OAI211_X1 U16389 ( .C1(n14894), .C2(n14524), .A(n14523), .B(n14522), .ZN(
        P1_U3238) );
  XOR2_X1 U16390 ( .A(n14526), .B(n14525), .Z(n14535) );
  OAI22_X1 U16391 ( .A1(n14529), .A2(n14528), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14527), .ZN(n14530) );
  AOI21_X1 U16392 ( .B1(n14538), .B2(n14747), .A(n14530), .ZN(n14531) );
  OAI21_X1 U16393 ( .B1(n14532), .B2(n14542), .A(n14531), .ZN(n14533) );
  AOI21_X1 U16394 ( .B1(n14753), .B2(n14544), .A(n14533), .ZN(n14534) );
  OAI21_X1 U16395 ( .B1(n14535), .B2(n14546), .A(n14534), .ZN(P1_U3240) );
  XNOR2_X1 U16396 ( .A(n14537), .B(n14536), .ZN(n14547) );
  AOI22_X1 U16397 ( .A1(n14539), .A2(n14946), .B1(n14538), .B2(n14938), .ZN(
        n14541) );
  OAI211_X1 U16398 ( .C1(n14908), .C2(n14542), .A(n14541), .B(n14540), .ZN(
        n14543) );
  AOI21_X1 U16399 ( .B1(n9456), .B2(n14544), .A(n14543), .ZN(n14545) );
  OAI21_X1 U16400 ( .B1(n14547), .B2(n14546), .A(n14545), .ZN(P1_U3241) );
  MUX2_X1 U16401 ( .A(n14719), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14570), .Z(
        P1_U3591) );
  MUX2_X1 U16402 ( .A(n14548), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14570), .Z(
        P1_U3590) );
  MUX2_X1 U16403 ( .A(n14549), .B(P1_DATAO_REG_29__SCAN_IN), .S(n14570), .Z(
        P1_U3589) );
  MUX2_X1 U16404 ( .A(n14550), .B(P1_DATAO_REG_28__SCAN_IN), .S(n14570), .Z(
        P1_U3588) );
  MUX2_X1 U16405 ( .A(n14748), .B(P1_DATAO_REG_27__SCAN_IN), .S(n14570), .Z(
        P1_U3587) );
  MUX2_X1 U16406 ( .A(n14551), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14570), .Z(
        P1_U3586) );
  MUX2_X1 U16407 ( .A(n14747), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14570), .Z(
        P1_U3585) );
  MUX2_X1 U16408 ( .A(n14552), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14570), .Z(
        P1_U3584) );
  MUX2_X1 U16409 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14553), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16410 ( .A(n14554), .B(P1_DATAO_REG_22__SCAN_IN), .S(n14570), .Z(
        P1_U3582) );
  MUX2_X1 U16411 ( .A(n14555), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14570), .Z(
        P1_U3581) );
  MUX2_X1 U16412 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14556), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16413 ( .A(n14557), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14570), .Z(
        P1_U3579) );
  MUX2_X1 U16414 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14558), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16415 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14925), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16416 ( .A(n14941), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14570), .Z(
        P1_U3576) );
  MUX2_X1 U16417 ( .A(n14924), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14570), .Z(
        P1_U3575) );
  MUX2_X1 U16418 ( .A(n14938), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14570), .Z(
        P1_U3574) );
  MUX2_X1 U16419 ( .A(n14559), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14570), .Z(
        P1_U3573) );
  MUX2_X1 U16420 ( .A(n14560), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14570), .Z(
        P1_U3572) );
  MUX2_X1 U16421 ( .A(n14561), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14570), .Z(
        P1_U3571) );
  MUX2_X1 U16422 ( .A(n14562), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14570), .Z(
        P1_U3570) );
  MUX2_X1 U16423 ( .A(n14563), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14570), .Z(
        P1_U3569) );
  MUX2_X1 U16424 ( .A(n14564), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14570), .Z(
        P1_U3568) );
  MUX2_X1 U16425 ( .A(n14565), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14570), .Z(
        P1_U3567) );
  MUX2_X1 U16426 ( .A(n14566), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14570), .Z(
        P1_U3566) );
  MUX2_X1 U16427 ( .A(n14567), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14570), .Z(
        P1_U3565) );
  MUX2_X1 U16428 ( .A(n14568), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14570), .Z(
        P1_U3564) );
  MUX2_X1 U16429 ( .A(n14569), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14570), .Z(
        P1_U3563) );
  MUX2_X1 U16430 ( .A(n9433), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14570), .Z(
        P1_U3562) );
  MUX2_X1 U16431 ( .A(n8757), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14570), .Z(
        P1_U3561) );
  OAI22_X1 U16432 ( .A1(n14650), .A2(n14572), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14571), .ZN(n14573) );
  AOI21_X1 U16433 ( .B1(n14574), .B2(n14653), .A(n14573), .ZN(n14581) );
  OAI211_X1 U16434 ( .C1(n14576), .C2(n14575), .A(n14708), .B(n14598), .ZN(
        n14580) );
  NAND2_X1 U16435 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14583) );
  INV_X1 U16436 ( .A(n14583), .ZN(n14578) );
  OAI211_X1 U16437 ( .C1(n14578), .C2(n14577), .A(n14677), .B(n14593), .ZN(
        n14579) );
  NAND3_X1 U16438 ( .A1(n14581), .A2(n14580), .A3(n14579), .ZN(P1_U3244) );
  INV_X1 U16439 ( .A(n14582), .ZN(n14585) );
  AOI21_X1 U16440 ( .B1(n15236), .B2(n14583), .A(n15163), .ZN(n14584) );
  OAI21_X1 U16441 ( .B1(n14585), .B2(n15236), .A(n14584), .ZN(n14589) );
  OR2_X1 U16442 ( .A1(n14586), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14588) );
  NAND2_X1 U16443 ( .A1(n14588), .A2(n14587), .ZN(n15237) );
  NAND2_X1 U16444 ( .A1(n15237), .A2(n15239), .ZN(n15242) );
  NAND3_X1 U16445 ( .A1(n14589), .A2(P1_U4016), .A3(n15242), .ZN(n14632) );
  INV_X1 U16446 ( .A(n14596), .ZN(n14591) );
  OAI22_X1 U16447 ( .A1(n14650), .A2(n15554), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11356), .ZN(n14590) );
  AOI21_X1 U16448 ( .B1(n14591), .B2(n14653), .A(n14590), .ZN(n14603) );
  MUX2_X1 U16449 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10749), .S(n14596), .Z(
        n14594) );
  NAND3_X1 U16450 ( .A1(n14594), .A2(n14593), .A3(n14592), .ZN(n14595) );
  NAND3_X1 U16451 ( .A1(n14677), .A2(n14610), .A3(n14595), .ZN(n14602) );
  MUX2_X1 U16452 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10720), .S(n14596), .Z(
        n14599) );
  NAND3_X1 U16453 ( .A1(n14599), .A2(n14598), .A3(n14597), .ZN(n14600) );
  NAND3_X1 U16454 ( .A1(n14708), .A2(n14606), .A3(n14600), .ZN(n14601) );
  NAND4_X1 U16455 ( .A1(n14632), .A2(n14603), .A3(n14602), .A4(n14601), .ZN(
        P1_U3245) );
  MUX2_X1 U16456 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10723), .S(n14612), .Z(
        n14604) );
  NAND3_X1 U16457 ( .A1(n14606), .A2(n14605), .A3(n14604), .ZN(n14607) );
  NAND3_X1 U16458 ( .A1(n14708), .A2(n14622), .A3(n14607), .ZN(n14617) );
  MUX2_X1 U16459 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10752), .S(n14612), .Z(
        n14608) );
  NAND3_X1 U16460 ( .A1(n14610), .A2(n14609), .A3(n14608), .ZN(n14611) );
  NAND3_X1 U16461 ( .A1(n14677), .A2(n14628), .A3(n14611), .ZN(n14616) );
  AOI22_X1 U16462 ( .A1(n15244), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n14615) );
  INV_X1 U16463 ( .A(n14612), .ZN(n14613) );
  NAND2_X1 U16464 ( .A1(n14653), .A2(n14613), .ZN(n14614) );
  NAND4_X1 U16465 ( .A1(n14617), .A2(n14616), .A3(n14615), .A4(n14614), .ZN(
        P1_U3246) );
  AND2_X1 U16466 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14619) );
  NOR2_X1 U16467 ( .A1(n14650), .A2(n15556), .ZN(n14618) );
  AOI211_X1 U16468 ( .C1(n14653), .C2(n14625), .A(n14619), .B(n14618), .ZN(
        n14633) );
  MUX2_X1 U16469 ( .A(n10726), .B(P1_REG1_REG_4__SCAN_IN), .S(n14625), .Z(
        n14621) );
  NAND3_X1 U16470 ( .A1(n14622), .A2(n14621), .A3(n14620), .ZN(n14623) );
  NAND3_X1 U16471 ( .A1(n14708), .A2(n14624), .A3(n14623), .ZN(n14631) );
  MUX2_X1 U16472 ( .A(n11305), .B(P1_REG2_REG_4__SCAN_IN), .S(n14625), .Z(
        n14627) );
  NAND3_X1 U16473 ( .A1(n14628), .A2(n14627), .A3(n14626), .ZN(n14629) );
  NAND3_X1 U16474 ( .A1(n14677), .A2(n14640), .A3(n14629), .ZN(n14630) );
  NAND4_X1 U16475 ( .A1(n14633), .A2(n14632), .A3(n14631), .A4(n14630), .ZN(
        P1_U3247) );
  OAI21_X1 U16476 ( .B1(n14650), .B2(n14635), .A(n14634), .ZN(n14636) );
  AOI21_X1 U16477 ( .B1(n14637), .B2(n14653), .A(n14636), .ZN(n14648) );
  MUX2_X1 U16478 ( .A(n10757), .B(P1_REG2_REG_5__SCAN_IN), .S(n14637), .Z(
        n14638) );
  NAND3_X1 U16479 ( .A1(n14640), .A2(n14639), .A3(n14638), .ZN(n14641) );
  NAND3_X1 U16480 ( .A1(n14677), .A2(n14659), .A3(n14641), .ZN(n14647) );
  OAI21_X1 U16481 ( .B1(n14644), .B2(n14643), .A(n14642), .ZN(n14645) );
  NAND2_X1 U16482 ( .A1(n14708), .A2(n14645), .ZN(n14646) );
  NAND3_X1 U16483 ( .A1(n14648), .A2(n14647), .A3(n14646), .ZN(P1_U3248) );
  NOR2_X1 U16484 ( .A1(n14650), .A2(n14649), .ZN(n14651) );
  AOI211_X1 U16485 ( .C1(n14653), .C2(n14656), .A(n14652), .B(n14651), .ZN(
        n14663) );
  OAI211_X1 U16486 ( .C1(n14655), .C2(n14654), .A(n14708), .B(n14668), .ZN(
        n14662) );
  MUX2_X1 U16487 ( .A(n11456), .B(P1_REG2_REG_6__SCAN_IN), .S(n14656), .Z(
        n14657) );
  NAND3_X1 U16488 ( .A1(n14659), .A2(n14658), .A3(n14657), .ZN(n14660) );
  NAND3_X1 U16489 ( .A1(n14677), .A2(n14674), .A3(n14660), .ZN(n14661) );
  NAND3_X1 U16490 ( .A1(n14663), .A2(n14662), .A3(n14661), .ZN(P1_U3249) );
  NOR2_X1 U16491 ( .A1(n14709), .A2(n14671), .ZN(n14664) );
  AOI211_X1 U16492 ( .C1(n15244), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n14665), .B(
        n14664), .ZN(n14680) );
  MUX2_X1 U16493 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10732), .S(n14671), .Z(
        n14666) );
  NAND3_X1 U16494 ( .A1(n14668), .A2(n14667), .A3(n14666), .ZN(n14669) );
  NAND3_X1 U16495 ( .A1(n14708), .A2(n14670), .A3(n14669), .ZN(n14679) );
  MUX2_X1 U16496 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10761), .S(n14671), .Z(
        n14672) );
  NAND3_X1 U16497 ( .A1(n14674), .A2(n14673), .A3(n14672), .ZN(n14675) );
  NAND3_X1 U16498 ( .A1(n14677), .A2(n14676), .A3(n14675), .ZN(n14678) );
  NAND3_X1 U16499 ( .A1(n14680), .A2(n14679), .A3(n14678), .ZN(P1_U3250) );
  NAND2_X1 U16500 ( .A1(n14685), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14681) );
  XNOR2_X1 U16501 ( .A(n14698), .B(n14691), .ZN(n14697) );
  XNOR2_X1 U16502 ( .A(n14697), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n14695) );
  NAND2_X1 U16503 ( .A1(n14684), .A2(n14683), .ZN(n14687) );
  NAND2_X1 U16504 ( .A1(n14685), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n14686) );
  NAND2_X1 U16505 ( .A1(n14687), .A2(n14686), .ZN(n14704) );
  XNOR2_X1 U16506 ( .A(n14704), .B(n14691), .ZN(n14702) );
  XOR2_X1 U16507 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14702), .Z(n14688) );
  NAND2_X1 U16508 ( .A1(n14708), .A2(n14688), .ZN(n14689) );
  NAND2_X1 U16509 ( .A1(n14690), .A2(n14689), .ZN(n14693) );
  NOR2_X1 U16510 ( .A1(n14709), .A2(n14691), .ZN(n14692) );
  AOI211_X1 U16511 ( .C1(n15244), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n14693), 
        .B(n14692), .ZN(n14694) );
  OAI21_X1 U16512 ( .B1(n14695), .B2(n14712), .A(n14694), .ZN(P1_U3261) );
  INV_X1 U16513 ( .A(n14696), .ZN(n14716) );
  NAND2_X1 U16514 ( .A1(n14697), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n14700) );
  NAND2_X1 U16515 ( .A1(n14698), .A2(n14703), .ZN(n14699) );
  NAND2_X1 U16516 ( .A1(n14700), .A2(n14699), .ZN(n14701) );
  XNOR2_X1 U16517 ( .A(n14701), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n14713) );
  INV_X1 U16518 ( .A(n14713), .ZN(n14711) );
  NAND2_X1 U16519 ( .A1(n14702), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14706) );
  NAND2_X1 U16520 ( .A1(n14704), .A2(n14703), .ZN(n14705) );
  NAND2_X1 U16521 ( .A1(n14706), .A2(n14705), .ZN(n14707) );
  XNOR2_X1 U16522 ( .A(n14707), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n14715) );
  NAND2_X1 U16523 ( .A1(n14715), .A2(n14708), .ZN(n14710) );
  NOR2_X1 U16524 ( .A1(n14718), .A2(n15323), .ZN(n14993) );
  NAND2_X1 U16525 ( .A1(n14993), .A2(n15289), .ZN(n14723) );
  AND2_X1 U16526 ( .A1(n14720), .A2(n14719), .ZN(n14996) );
  INV_X1 U16527 ( .A(n14996), .ZN(n14721) );
  NOR2_X1 U16528 ( .A1(n6538), .A2(n14721), .ZN(n14728) );
  AOI21_X1 U16529 ( .B1(n6538), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14728), .ZN(
        n14722) );
  OAI211_X1 U16530 ( .C1(n7494), .C2(n15283), .A(n14723), .B(n14722), .ZN(
        P1_U3263) );
  INV_X1 U16531 ( .A(n14724), .ZN(n14726) );
  XNOR2_X1 U16532 ( .A(n14726), .B(n14725), .ZN(n14997) );
  NAND2_X1 U16533 ( .A1(n14997), .A2(n14727), .ZN(n14730) );
  AOI21_X1 U16534 ( .B1(n6538), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14728), .ZN(
        n14729) );
  OAI211_X1 U16535 ( .C1(n15107), .C2(n15283), .A(n14730), .B(n14729), .ZN(
        P1_U3264) );
  NOR2_X1 U16536 ( .A1(n14732), .A2(n14731), .ZN(n14733) );
  OAI21_X1 U16537 ( .B1(n14734), .B2(n14733), .A(n14987), .ZN(n14740) );
  OAI22_X1 U16538 ( .A1(n14987), .A2(n14736), .B1(n14735), .B2(n15280), .ZN(
        n14737) );
  AOI21_X1 U16539 ( .B1(n14738), .B2(n14752), .A(n14737), .ZN(n14739) );
  OAI211_X1 U16540 ( .C1(n14953), .C2(n14741), .A(n14740), .B(n14739), .ZN(
        P1_U3265) );
  XNOR2_X1 U16541 ( .A(n14742), .B(n14744), .ZN(n15006) );
  XOR2_X1 U16542 ( .A(n14744), .B(n14743), .Z(n15004) );
  OAI211_X1 U16543 ( .C1(n15002), .C2(n14746), .A(n14745), .B(n10110), .ZN(
        n15001) );
  AOI22_X1 U16544 ( .A1(n14748), .A2(n14940), .B1(n14939), .B2(n14747), .ZN(
        n15000) );
  AOI22_X1 U16545 ( .A1(n14749), .A2(n14945), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n6538), .ZN(n14750) );
  OAI21_X1 U16546 ( .B1(n15000), .B2(n6538), .A(n14750), .ZN(n14751) );
  AOI21_X1 U16547 ( .B1(n14753), .B2(n14752), .A(n14751), .ZN(n14754) );
  OAI21_X1 U16548 ( .B1(n15001), .B2(n15265), .A(n14754), .ZN(n14755) );
  AOI21_X1 U16549 ( .B1(n15004), .B2(n14905), .A(n14755), .ZN(n14756) );
  OAI21_X1 U16550 ( .B1(n15006), .B2(n14953), .A(n14756), .ZN(P1_U3267) );
  OAI21_X1 U16551 ( .B1(n14758), .B2(n14761), .A(n14757), .ZN(n15007) );
  OAI21_X1 U16552 ( .B1(n14763), .B2(n15276), .A(n14762), .ZN(n15008) );
  NAND2_X1 U16553 ( .A1(n15008), .A2(n14987), .ZN(n14771) );
  XNOR2_X1 U16554 ( .A(n14783), .B(n14765), .ZN(n14764) );
  NOR2_X1 U16555 ( .A1(n14764), .A2(n15323), .ZN(n15009) );
  NOR2_X1 U16556 ( .A1(n7507), .A2(n15283), .ZN(n14769) );
  OAI22_X1 U16557 ( .A1(n14767), .A2(n15280), .B1(n14766), .B2(n14987), .ZN(
        n14768) );
  AOI211_X1 U16558 ( .C1(n15009), .C2(n15289), .A(n14769), .B(n14768), .ZN(
        n14770) );
  OAI211_X1 U16559 ( .C1(n15007), .C2(n14953), .A(n14771), .B(n14770), .ZN(
        P1_U3268) );
  NAND2_X1 U16560 ( .A1(n14772), .A2(n14773), .ZN(n14774) );
  NAND3_X1 U16561 ( .A1(n14775), .A2(n15331), .A3(n14774), .ZN(n14777) );
  NAND2_X1 U16562 ( .A1(n14779), .A2(n14778), .ZN(n14780) );
  NAND2_X1 U16563 ( .A1(n14781), .A2(n14780), .ZN(n15013) );
  INV_X1 U16564 ( .A(n15117), .ZN(n14787) );
  AOI21_X1 U16565 ( .B1(n14797), .B2(n15117), .A(n15323), .ZN(n14782) );
  AND2_X1 U16566 ( .A1(n14783), .A2(n14782), .ZN(n15012) );
  NAND2_X1 U16567 ( .A1(n15012), .A2(n15289), .ZN(n14786) );
  AOI22_X1 U16568 ( .A1(n14784), .A2(n14945), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n6538), .ZN(n14785) );
  OAI211_X1 U16569 ( .C1(n14787), .C2(n15283), .A(n14786), .B(n14785), .ZN(
        n14788) );
  AOI21_X1 U16570 ( .B1(n15013), .B2(n14789), .A(n14788), .ZN(n14790) );
  OAI21_X1 U16571 ( .B1(n15015), .B2(n6538), .A(n14790), .ZN(P1_U3269) );
  INV_X1 U16572 ( .A(n14791), .ZN(n14796) );
  XNOR2_X1 U16573 ( .A(n14792), .B(n14793), .ZN(n14795) );
  OAI21_X1 U16574 ( .B1(n14795), .B2(n15276), .A(n14794), .ZN(n15019) );
  AOI21_X1 U16575 ( .B1(n14796), .B2(n14945), .A(n15019), .ZN(n14809) );
  INV_X1 U16576 ( .A(n14797), .ZN(n14798) );
  AOI211_X1 U16577 ( .C1(n14800), .C2(n14799), .A(n15323), .B(n14798), .ZN(
        n15020) );
  INV_X1 U16578 ( .A(n14800), .ZN(n15122) );
  OAI22_X1 U16579 ( .A1(n15122), .A2(n15283), .B1(n14801), .B2(n14987), .ZN(
        n14802) );
  AOI21_X1 U16580 ( .B1(n15020), .B2(n15289), .A(n14802), .ZN(n14808) );
  INV_X1 U16581 ( .A(n14803), .ZN(n14804) );
  AOI21_X1 U16582 ( .B1(n14806), .B2(n14805), .A(n14804), .ZN(n15021) );
  NAND2_X1 U16583 ( .A1(n15021), .A2(n14990), .ZN(n14807) );
  OAI211_X1 U16584 ( .C1(n14809), .C2(n6538), .A(n14808), .B(n14807), .ZN(
        P1_U3270) );
  INV_X1 U16585 ( .A(n14810), .ZN(n14811) );
  AOI21_X1 U16586 ( .B1(n14820), .B2(n14812), .A(n14811), .ZN(n15029) );
  INV_X1 U16587 ( .A(n14905), .ZN(n14867) );
  XNOR2_X1 U16588 ( .A(n14834), .B(n7511), .ZN(n14813) );
  AOI22_X1 U16589 ( .A1(n14814), .A2(n14945), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n6538), .ZN(n14816) );
  NAND2_X1 U16590 ( .A1(n15025), .A2(n14987), .ZN(n14815) );
  OAI211_X1 U16591 ( .C1(n14817), .C2(n15283), .A(n14816), .B(n14815), .ZN(
        n14818) );
  AOI21_X1 U16592 ( .B1(n15024), .B2(n15289), .A(n14818), .ZN(n14823) );
  OAI21_X1 U16593 ( .B1(n14821), .B2(n14820), .A(n14819), .ZN(n15026) );
  NAND2_X1 U16594 ( .A1(n15026), .A2(n14990), .ZN(n14822) );
  OAI211_X1 U16595 ( .C1(n15029), .C2(n14867), .A(n14823), .B(n14822), .ZN(
        P1_U3271) );
  XNOR2_X1 U16596 ( .A(n14824), .B(n14827), .ZN(n15032) );
  INV_X1 U16597 ( .A(n15032), .ZN(n14841) );
  INV_X1 U16598 ( .A(n14827), .ZN(n14829) );
  NAND3_X1 U16599 ( .A1(n14826), .A2(n14829), .A3(n14828), .ZN(n14830) );
  NAND3_X1 U16600 ( .A1(n14825), .A2(n15331), .A3(n14830), .ZN(n14833) );
  INV_X1 U16601 ( .A(n14831), .ZN(n14832) );
  NAND2_X1 U16602 ( .A1(n14833), .A2(n14832), .ZN(n15030) );
  OAI21_X1 U16603 ( .B1(n14856), .B2(n15127), .A(n10110), .ZN(n14835) );
  NOR2_X1 U16604 ( .A1(n14835), .A2(n14834), .ZN(n15031) );
  NAND2_X1 U16605 ( .A1(n15031), .A2(n15289), .ZN(n14838) );
  AOI22_X1 U16606 ( .A1(n14836), .A2(n14945), .B1(n6538), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n14837) );
  OAI211_X1 U16607 ( .C1(n15127), .C2(n15283), .A(n14838), .B(n14837), .ZN(
        n14839) );
  AOI21_X1 U16608 ( .B1(n15030), .B2(n14987), .A(n14839), .ZN(n14840) );
  OAI21_X1 U16609 ( .B1(n14841), .B2(n14953), .A(n14840), .ZN(P1_U3272) );
  INV_X1 U16610 ( .A(n14842), .ZN(n14845) );
  AOI21_X1 U16611 ( .B1(n14845), .B2(n14844), .A(n14843), .ZN(n14848) );
  INV_X1 U16612 ( .A(n14846), .ZN(n14847) );
  NOR2_X1 U16613 ( .A1(n14848), .A2(n14847), .ZN(n14849) );
  OAI21_X1 U16614 ( .B1(n14849), .B2(n14855), .A(n14826), .ZN(n15041) );
  NAND2_X1 U16615 ( .A1(n14850), .A2(n14851), .ZN(n14854) );
  INV_X1 U16616 ( .A(n14852), .ZN(n14853) );
  AOI21_X1 U16617 ( .B1(n14855), .B2(n14854), .A(n14853), .ZN(n15039) );
  AOI211_X1 U16618 ( .C1(n14858), .C2(n14857), .A(n15323), .B(n14856), .ZN(
        n15038) );
  NAND2_X1 U16619 ( .A1(n15038), .A2(n15289), .ZN(n14864) );
  AOI21_X1 U16620 ( .B1(n14860), .B2(n14945), .A(n14859), .ZN(n14861) );
  MUX2_X1 U16621 ( .A(n14862), .B(n14861), .S(n14987), .Z(n14863) );
  OAI211_X1 U16622 ( .C1(n15036), .C2(n15283), .A(n14864), .B(n14863), .ZN(
        n14865) );
  AOI21_X1 U16623 ( .B1(n15039), .B2(n14990), .A(n14865), .ZN(n14866) );
  OAI21_X1 U16624 ( .B1(n15041), .B2(n14867), .A(n14866), .ZN(P1_U3273) );
  XNOR2_X1 U16625 ( .A(n14868), .B(n9368), .ZN(n15044) );
  INV_X1 U16626 ( .A(n15044), .ZN(n14882) );
  INV_X1 U16627 ( .A(n14901), .ZN(n14904) );
  NOR2_X1 U16628 ( .A1(n14842), .A2(n14904), .ZN(n14903) );
  NOR2_X1 U16629 ( .A1(n14903), .A2(n14869), .ZN(n14883) );
  OR2_X1 U16630 ( .A1(n14883), .A2(n14895), .ZN(n14887) );
  NAND2_X1 U16631 ( .A1(n14887), .A2(n14870), .ZN(n14871) );
  XNOR2_X1 U16632 ( .A(n14871), .B(n9368), .ZN(n14873) );
  OAI21_X1 U16633 ( .B1(n14873), .B2(n15276), .A(n14872), .ZN(n15042) );
  NAND2_X1 U16634 ( .A1(n15042), .A2(n14987), .ZN(n14881) );
  XNOR2_X1 U16635 ( .A(n14889), .B(n14875), .ZN(n14874) );
  NOR2_X1 U16636 ( .A1(n14874), .A2(n15323), .ZN(n15043) );
  INV_X1 U16637 ( .A(n14875), .ZN(n15132) );
  NOR2_X1 U16638 ( .A1(n15132), .A2(n15283), .ZN(n14879) );
  OAI22_X1 U16639 ( .A1(n14987), .A2(n14877), .B1(n14876), .B2(n15280), .ZN(
        n14878) );
  AOI211_X1 U16640 ( .C1(n15043), .C2(n15289), .A(n14879), .B(n14878), .ZN(
        n14880) );
  OAI211_X1 U16641 ( .C1(n14882), .C2(n14953), .A(n14881), .B(n14880), .ZN(
        P1_U3274) );
  AOI21_X1 U16642 ( .B1(n14883), .B2(n14895), .A(n15276), .ZN(n14888) );
  OAI22_X1 U16643 ( .A1(n14885), .A2(n14909), .B1(n14884), .B2(n14907), .ZN(
        n14886) );
  AOI21_X1 U16644 ( .B1(n14888), .B2(n14887), .A(n14886), .ZN(n15050) );
  INV_X1 U16645 ( .A(n14906), .ZN(n14891) );
  INV_X1 U16646 ( .A(n14889), .ZN(n14890) );
  AOI211_X1 U16647 ( .C1(n15048), .C2(n14891), .A(n15323), .B(n14890), .ZN(
        n15047) );
  AOI22_X1 U16648 ( .A1(n6538), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14892), 
        .B2(n14945), .ZN(n14893) );
  OAI21_X1 U16649 ( .B1(n14894), .B2(n15283), .A(n14893), .ZN(n14899) );
  XNOR2_X1 U16650 ( .A(n14896), .B(n14895), .ZN(n15051) );
  NOR2_X1 U16651 ( .A1(n15051), .A2(n14897), .ZN(n14898) );
  AOI211_X1 U16652 ( .C1(n15047), .C2(n15289), .A(n14899), .B(n14898), .ZN(
        n14900) );
  OAI21_X1 U16653 ( .B1(n15050), .B2(n6538), .A(n14900), .ZN(P1_U3275) );
  XNOR2_X1 U16654 ( .A(n14902), .B(n14901), .ZN(n15058) );
  AOI21_X1 U16655 ( .B1(n14904), .B2(n14842), .A(n14903), .ZN(n15052) );
  NAND2_X1 U16656 ( .A1(n15052), .A2(n14905), .ZN(n14916) );
  AOI211_X1 U16657 ( .C1(n15055), .C2(n14929), .A(n15323), .B(n14906), .ZN(
        n15053) );
  OAI22_X1 U16658 ( .A1(n14910), .A2(n14909), .B1(n14908), .B2(n14907), .ZN(
        n15054) );
  AOI22_X1 U16659 ( .A1(n14987), .A2(n15054), .B1(n14911), .B2(n14945), .ZN(
        n14913) );
  NAND2_X1 U16660 ( .A1(n6538), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14912) );
  OAI211_X1 U16661 ( .C1(n7090), .C2(n15283), .A(n14913), .B(n14912), .ZN(
        n14914) );
  AOI21_X1 U16662 ( .B1(n15053), .B2(n15289), .A(n14914), .ZN(n14915) );
  OAI211_X1 U16663 ( .C1(n15058), .C2(n14953), .A(n14916), .B(n14915), .ZN(
        P1_U3276) );
  OAI21_X1 U16664 ( .B1(n14919), .B2(n14918), .A(n14917), .ZN(n14920) );
  INV_X1 U16665 ( .A(n14920), .ZN(n15063) );
  OAI21_X1 U16666 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n14926) );
  AOI222_X1 U16667 ( .A1(n15331), .A2(n14926), .B1(n14925), .B2(n14940), .C1(
        n14924), .C2(n14939), .ZN(n15062) );
  OAI21_X1 U16668 ( .B1(n14927), .B2(n15280), .A(n15062), .ZN(n14928) );
  NAND2_X1 U16669 ( .A1(n14928), .A2(n14987), .ZN(n14935) );
  INV_X1 U16670 ( .A(n14929), .ZN(n14930) );
  AOI211_X1 U16671 ( .C1(n15060), .C2(n14931), .A(n15323), .B(n14930), .ZN(
        n15059) );
  OAI22_X1 U16672 ( .A1(n7498), .A2(n15283), .B1(n14932), .B2(n14987), .ZN(
        n14933) );
  AOI21_X1 U16673 ( .B1(n15059), .B2(n15289), .A(n14933), .ZN(n14934) );
  OAI211_X1 U16674 ( .C1(n15063), .C2(n14953), .A(n14935), .B(n14934), .ZN(
        P1_U3277) );
  OAI211_X1 U16675 ( .C1(n14937), .C2(n14952), .A(n14936), .B(n15331), .ZN(
        n14943) );
  AOI22_X1 U16676 ( .A1(n14941), .A2(n14940), .B1(n14939), .B2(n14938), .ZN(
        n14942) );
  XNOR2_X1 U16677 ( .A(n6558), .B(n14948), .ZN(n14944) );
  NOR2_X1 U16678 ( .A1(n14944), .A2(n15323), .ZN(n15064) );
  AOI22_X1 U16679 ( .A1(n6538), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14946), 
        .B2(n14945), .ZN(n14947) );
  OAI21_X1 U16680 ( .B1(n14948), .B2(n15283), .A(n14947), .ZN(n14955) );
  NOR2_X1 U16681 ( .A1(n14949), .A2(n14967), .ZN(n14966) );
  NOR2_X1 U16682 ( .A1(n14966), .A2(n14950), .ZN(n14951) );
  XNOR2_X1 U16683 ( .A(n14952), .B(n14951), .ZN(n15067) );
  NOR2_X1 U16684 ( .A1(n15067), .A2(n14953), .ZN(n14954) );
  AOI211_X1 U16685 ( .C1(n15064), .C2(n15289), .A(n14955), .B(n14954), .ZN(
        n14956) );
  OAI21_X1 U16686 ( .B1(n6538), .B2(n15066), .A(n14956), .ZN(P1_U3278) );
  AOI211_X1 U16687 ( .C1(n14957), .C2(n14977), .A(n15323), .B(n6558), .ZN(
        n15069) );
  NAND3_X1 U16688 ( .A1(n14959), .A2(n14961), .A3(n14960), .ZN(n14962) );
  NAND3_X1 U16689 ( .A1(n14958), .A2(n15331), .A3(n14962), .ZN(n14965) );
  INV_X1 U16690 ( .A(n14963), .ZN(n14964) );
  NAND2_X1 U16691 ( .A1(n14965), .A2(n14964), .ZN(n15068) );
  AOI21_X1 U16692 ( .B1(n15069), .B2(n8984), .A(n15068), .ZN(n14973) );
  AOI21_X1 U16693 ( .B1(n14967), .B2(n14949), .A(n14966), .ZN(n15070) );
  NOR2_X1 U16694 ( .A1(n7500), .A2(n15283), .ZN(n14971) );
  OAI22_X1 U16695 ( .A1(n14987), .A2(n14969), .B1(n14968), .B2(n15280), .ZN(
        n14970) );
  AOI211_X1 U16696 ( .C1(n15070), .C2(n14990), .A(n14971), .B(n14970), .ZN(
        n14972) );
  OAI21_X1 U16697 ( .B1(n14973), .B2(n6538), .A(n14972), .ZN(P1_U3279) );
  OAI21_X1 U16698 ( .B1(n14975), .B2(n14974), .A(n14984), .ZN(n14976) );
  NAND3_X1 U16699 ( .A1(n14977), .A2(n14976), .A3(n10110), .ZN(n15075) );
  INV_X1 U16700 ( .A(n15075), .ZN(n14980) );
  NAND3_X1 U16701 ( .A1(n12051), .A2(n14982), .A3(n14978), .ZN(n14979) );
  AOI211_X1 U16702 ( .C1(n14980), .C2(n8984), .A(n15073), .B(n15076), .ZN(
        n14992) );
  OAI21_X1 U16703 ( .B1(n14983), .B2(n14982), .A(n14981), .ZN(n15078) );
  INV_X1 U16704 ( .A(n14984), .ZN(n15143) );
  NOR2_X1 U16705 ( .A1(n15143), .A2(n15283), .ZN(n14989) );
  OAI22_X1 U16706 ( .A1(n14987), .A2(n14986), .B1(n14985), .B2(n15280), .ZN(
        n14988) );
  AOI211_X1 U16707 ( .C1(n15078), .C2(n14990), .A(n14989), .B(n14988), .ZN(
        n14991) );
  OAI21_X1 U16708 ( .B1(n14992), .B2(n6538), .A(n14991), .ZN(P1_U3280) );
  INV_X1 U16709 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14994) );
  NOR2_X1 U16710 ( .A1(n14993), .A2(n14996), .ZN(n15102) );
  MUX2_X1 U16711 ( .A(n14994), .B(n15102), .S(n15348), .Z(n14995) );
  OAI21_X1 U16712 ( .B1(n7494), .B2(n15086), .A(n14995), .ZN(P1_U3559) );
  INV_X1 U16713 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14998) );
  AOI21_X1 U16714 ( .B1(n14997), .B2(n10110), .A(n14996), .ZN(n15104) );
  MUX2_X1 U16715 ( .A(n14998), .B(n15104), .S(n15348), .Z(n14999) );
  OAI21_X1 U16716 ( .B1(n15107), .B2(n15086), .A(n14999), .ZN(P1_U3558) );
  OAI211_X1 U16717 ( .C1(n15002), .C2(n15335), .A(n15001), .B(n15000), .ZN(
        n15003) );
  AOI21_X1 U16718 ( .B1(n15004), .B2(n15331), .A(n15003), .ZN(n15005) );
  OAI21_X1 U16719 ( .B1(n15100), .B2(n15006), .A(n15005), .ZN(n15111) );
  MUX2_X1 U16720 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15111), .S(n15348), .Z(
        P1_U3554) );
  INV_X1 U16721 ( .A(n15007), .ZN(n15010) );
  OAI21_X1 U16722 ( .B1(n7507), .B2(n15086), .A(n15011), .ZN(P1_U3553) );
  INV_X1 U16723 ( .A(n15086), .ZN(n15017) );
  AOI21_X1 U16724 ( .B1(n15013), .B2(n15339), .A(n15012), .ZN(n15014) );
  NAND2_X1 U16725 ( .A1(n15015), .A2(n15014), .ZN(n15115) );
  MUX2_X1 U16726 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15115), .S(n15348), .Z(
        n15016) );
  AOI21_X1 U16727 ( .B1(n15017), .B2(n15117), .A(n15016), .ZN(n15018) );
  INV_X1 U16728 ( .A(n15018), .ZN(P1_U3552) );
  INV_X1 U16729 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n15022) );
  AOI211_X1 U16730 ( .C1(n15021), .C2(n15339), .A(n15020), .B(n15019), .ZN(
        n15119) );
  MUX2_X1 U16731 ( .A(n15022), .B(n15119), .S(n15348), .Z(n15023) );
  OAI21_X1 U16732 ( .B1(n15122), .B2(n15086), .A(n15023), .ZN(P1_U3551) );
  AOI211_X1 U16733 ( .C1(n15295), .C2(n7511), .A(n15025), .B(n15024), .ZN(
        n15028) );
  NAND2_X1 U16734 ( .A1(n15026), .A2(n15339), .ZN(n15027) );
  OAI211_X1 U16735 ( .C1(n15029), .C2(n15276), .A(n15028), .B(n15027), .ZN(
        n15123) );
  MUX2_X1 U16736 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15123), .S(n15348), .Z(
        P1_U3550) );
  INV_X1 U16737 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n15033) );
  AOI211_X1 U16738 ( .C1(n15339), .C2(n15032), .A(n15031), .B(n15030), .ZN(
        n15124) );
  MUX2_X1 U16739 ( .A(n15033), .B(n15124), .S(n15348), .Z(n15034) );
  OAI21_X1 U16740 ( .B1(n15127), .B2(n15086), .A(n15034), .ZN(P1_U3549) );
  OAI21_X1 U16741 ( .B1(n15036), .B2(n15335), .A(n15035), .ZN(n15037) );
  AOI211_X1 U16742 ( .C1(n15039), .C2(n15339), .A(n15038), .B(n15037), .ZN(
        n15040) );
  OAI21_X1 U16743 ( .B1(n15041), .B2(n15276), .A(n15040), .ZN(n15128) );
  MUX2_X1 U16744 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15128), .S(n15348), .Z(
        P1_U3548) );
  INV_X1 U16745 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n15045) );
  AOI211_X1 U16746 ( .C1(n15339), .C2(n15044), .A(n15043), .B(n15042), .ZN(
        n15129) );
  MUX2_X1 U16747 ( .A(n15045), .B(n15129), .S(n15348), .Z(n15046) );
  OAI21_X1 U16748 ( .B1(n15132), .B2(n15086), .A(n15046), .ZN(P1_U3547) );
  AOI21_X1 U16749 ( .B1(n15295), .B2(n15048), .A(n15047), .ZN(n15049) );
  OAI211_X1 U16750 ( .C1(n15100), .C2(n15051), .A(n15050), .B(n15049), .ZN(
        n15133) );
  MUX2_X1 U16751 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15133), .S(n15348), .Z(
        P1_U3546) );
  NAND2_X1 U16752 ( .A1(n15052), .A2(n15331), .ZN(n15057) );
  AOI211_X1 U16753 ( .C1(n15295), .C2(n15055), .A(n15054), .B(n15053), .ZN(
        n15056) );
  OAI211_X1 U16754 ( .C1(n15100), .C2(n15058), .A(n15057), .B(n15056), .ZN(
        n15134) );
  MUX2_X1 U16755 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15134), .S(n15348), .Z(
        P1_U3545) );
  AOI21_X1 U16756 ( .B1(n15295), .B2(n15060), .A(n15059), .ZN(n15061) );
  OAI211_X1 U16757 ( .C1(n15100), .C2(n15063), .A(n15062), .B(n15061), .ZN(
        n15135) );
  MUX2_X1 U16758 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15135), .S(n15348), .Z(
        P1_U3544) );
  AOI21_X1 U16759 ( .B1(n15295), .B2(n9456), .A(n15064), .ZN(n15065) );
  OAI211_X1 U16760 ( .C1(n15100), .C2(n15067), .A(n15066), .B(n15065), .ZN(
        n15136) );
  MUX2_X1 U16761 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15136), .S(n15348), .Z(
        P1_U3543) );
  AOI211_X1 U16762 ( .C1(n15070), .C2(n15339), .A(n15069), .B(n15068), .ZN(
        n15137) );
  MUX2_X1 U16763 ( .A(n15071), .B(n15137), .S(n15348), .Z(n15072) );
  OAI21_X1 U16764 ( .B1(n7500), .B2(n15086), .A(n15072), .ZN(P1_U3542) );
  INV_X1 U16765 ( .A(n15073), .ZN(n15074) );
  NAND2_X1 U16766 ( .A1(n15075), .A2(n15074), .ZN(n15077) );
  AOI211_X1 U16767 ( .C1(n15339), .C2(n15078), .A(n15077), .B(n15076), .ZN(
        n15140) );
  MUX2_X1 U16768 ( .A(n15079), .B(n15140), .S(n15348), .Z(n15080) );
  OAI21_X1 U16769 ( .B1(n15143), .B2(n15086), .A(n15080), .ZN(P1_U3541) );
  AOI211_X1 U16770 ( .C1(n15339), .C2(n15083), .A(n15082), .B(n15081), .ZN(
        n15144) );
  MUX2_X1 U16771 ( .A(n15084), .B(n15144), .S(n15348), .Z(n15085) );
  OAI21_X1 U16772 ( .B1(n15148), .B2(n15086), .A(n15085), .ZN(P1_U3540) );
  OAI22_X1 U16773 ( .A1(n15088), .A2(n15323), .B1(n15087), .B2(n15335), .ZN(
        n15090) );
  AOI211_X1 U16774 ( .C1(n15339), .C2(n15091), .A(n15090), .B(n15089), .ZN(
        n15092) );
  INV_X1 U16775 ( .A(n15092), .ZN(n15149) );
  MUX2_X1 U16776 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15149), .S(n15348), .Z(
        P1_U3539) );
  NAND3_X1 U16777 ( .A1(n11516), .A2(n15093), .A3(n15331), .ZN(n15098) );
  AOI211_X1 U16778 ( .C1(n15295), .C2(n15096), .A(n15095), .B(n15094), .ZN(
        n15097) );
  OAI211_X1 U16779 ( .C1(n15100), .C2(n15099), .A(n15098), .B(n15097), .ZN(
        n15150) );
  MUX2_X1 U16780 ( .A(n15150), .B(P1_REG1_REG_10__SCAN_IN), .S(n9548), .Z(
        P1_U3538) );
  MUX2_X1 U16781 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n15101), .S(n15348), .Z(
        P1_U3528) );
  MUX2_X1 U16782 ( .A(n15782), .B(n15102), .S(n15342), .Z(n15103) );
  OAI21_X1 U16783 ( .B1(n7494), .B2(n15147), .A(n15103), .ZN(P1_U3527) );
  INV_X1 U16784 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15105) );
  MUX2_X1 U16785 ( .A(n15105), .B(n15104), .S(n15342), .Z(n15106) );
  OAI21_X1 U16786 ( .B1(n15107), .B2(n15147), .A(n15106), .ZN(P1_U3526) );
  INV_X1 U16787 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n15109) );
  MUX2_X1 U16788 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15111), .S(n15342), .Z(
        P1_U3522) );
  INV_X1 U16789 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n15113) );
  MUX2_X1 U16790 ( .A(n15113), .B(n15112), .S(n15342), .Z(n15114) );
  OAI21_X1 U16791 ( .B1(n7507), .B2(n15147), .A(n15114), .ZN(P1_U3521) );
  MUX2_X1 U16792 ( .A(n15115), .B(P1_REG0_REG_24__SCAN_IN), .S(n9554), .Z(
        n15116) );
  AOI21_X1 U16793 ( .B1(n7110), .B2(n15117), .A(n15116), .ZN(n15118) );
  INV_X1 U16794 ( .A(n15118), .ZN(P1_U3520) );
  INV_X1 U16795 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n15120) );
  MUX2_X1 U16796 ( .A(n15120), .B(n15119), .S(n15342), .Z(n15121) );
  OAI21_X1 U16797 ( .B1(n15122), .B2(n15147), .A(n15121), .ZN(P1_U3519) );
  MUX2_X1 U16798 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15123), .S(n15342), .Z(
        P1_U3518) );
  INV_X1 U16799 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n15125) );
  MUX2_X1 U16800 ( .A(n15125), .B(n15124), .S(n15342), .Z(n15126) );
  OAI21_X1 U16801 ( .B1(n15127), .B2(n15147), .A(n15126), .ZN(P1_U3517) );
  MUX2_X1 U16802 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15128), .S(n15342), .Z(
        P1_U3516) );
  INV_X1 U16803 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n15130) );
  MUX2_X1 U16804 ( .A(n15130), .B(n15129), .S(n15342), .Z(n15131) );
  OAI21_X1 U16805 ( .B1(n15132), .B2(n15147), .A(n15131), .ZN(P1_U3515) );
  MUX2_X1 U16806 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15133), .S(n15342), .Z(
        P1_U3513) );
  MUX2_X1 U16807 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15134), .S(n15342), .Z(
        P1_U3510) );
  MUX2_X1 U16808 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15135), .S(n15342), .Z(
        P1_U3507) );
  MUX2_X1 U16809 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15136), .S(n15342), .Z(
        P1_U3504) );
  MUX2_X1 U16810 ( .A(n15138), .B(n15137), .S(n15342), .Z(n15139) );
  OAI21_X1 U16811 ( .B1(n7500), .B2(n15147), .A(n15139), .ZN(P1_U3501) );
  INV_X1 U16812 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n15141) );
  MUX2_X1 U16813 ( .A(n15141), .B(n15140), .S(n15342), .Z(n15142) );
  OAI21_X1 U16814 ( .B1(n15143), .B2(n15147), .A(n15142), .ZN(P1_U3498) );
  INV_X1 U16815 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n15145) );
  MUX2_X1 U16816 ( .A(n15145), .B(n15144), .S(n15342), .Z(n15146) );
  OAI21_X1 U16817 ( .B1(n15148), .B2(n15147), .A(n15146), .ZN(P1_U3495) );
  MUX2_X1 U16818 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15149), .S(n15342), .Z(
        P1_U3492) );
  MUX2_X1 U16819 ( .A(n15150), .B(P1_REG0_REG_10__SCAN_IN), .S(n9554), .Z(
        P1_U3489) );
  NAND3_X1 U16820 ( .A1(n15152), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n15153) );
  OAI22_X1 U16821 ( .A1(n15151), .A2(n15153), .B1(n15682), .B2(n15161), .ZN(
        n15154) );
  AOI21_X1 U16822 ( .B1(n15156), .B2(n15155), .A(n15154), .ZN(n15157) );
  INV_X1 U16823 ( .A(n15157), .ZN(P1_U3324) );
  OAI222_X1 U16824 ( .A1(P1_U3086), .A2(n15160), .B1(n12474), .B2(n15159), 
        .C1(n15158), .C2(n15161), .ZN(P1_U3326) );
  OAI222_X1 U16825 ( .A1(n15163), .A2(P1_U3086), .B1(n12474), .B2(n15162), 
        .C1(n15840), .C2(n15161), .ZN(P1_U3327) );
  MUX2_X1 U16826 ( .A(n15165), .B(n15164), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16827 ( .A(n15166), .ZN(n15167) );
  MUX2_X1 U16828 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15167), .S(P1_U3086), .Z(
        P1_U3355) );
  XOR2_X1 U16829 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15168), .Z(SUB_1596_U53) );
  INV_X1 U16830 ( .A(n15170), .ZN(n15172) );
  INV_X1 U16831 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15171) );
  NAND2_X1 U16832 ( .A1(n15175), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n15176) );
  NAND2_X1 U16833 ( .A1(n15177), .A2(n15176), .ZN(n15187) );
  XNOR2_X1 U16834 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n15178) );
  XNOR2_X1 U16835 ( .A(n15187), .B(n15178), .ZN(n15179) );
  INV_X1 U16836 ( .A(n15194), .ZN(n15184) );
  INV_X1 U16837 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15180) );
  INV_X1 U16838 ( .A(n15181), .ZN(n15182) );
  OAI21_X1 U16839 ( .B1(n15182), .B2(n15184), .A(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n15183) );
  OAI21_X1 U16840 ( .B1(n15184), .B2(n15195), .A(n15183), .ZN(SUB_1596_U65) );
  NAND2_X1 U16841 ( .A1(n15195), .A2(n15194), .ZN(n15192) );
  NOR2_X1 U16842 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15185), .ZN(n15186) );
  NAND2_X1 U16843 ( .A1(n15185), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n15188) );
  NAND2_X1 U16844 ( .A1(n15189), .A2(n15188), .ZN(n15205) );
  INV_X1 U16845 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15202) );
  NOR2_X1 U16846 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15202), .ZN(n15204) );
  AOI21_X1 U16847 ( .B1(n15202), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n15204), 
        .ZN(n15190) );
  XNOR2_X1 U16848 ( .A(n15205), .B(n15190), .ZN(n15193) );
  INV_X1 U16849 ( .A(n15193), .ZN(n15191) );
  NAND2_X1 U16850 ( .A1(n15192), .A2(n15191), .ZN(n15200) );
  NAND2_X1 U16851 ( .A1(n15196), .A2(n15195), .ZN(n15199) );
  NAND2_X1 U16852 ( .A1(n15200), .A2(n15199), .ZN(n15197) );
  XNOR2_X1 U16853 ( .A(n15197), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  INV_X1 U16854 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15198) );
  NAND2_X1 U16855 ( .A1(n15199), .A2(n15198), .ZN(n15201) );
  NAND2_X1 U16856 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15202), .ZN(n15203) );
  OAI21_X1 U16857 ( .B1(n15205), .B2(n15204), .A(n15203), .ZN(n15214) );
  XNOR2_X1 U16858 ( .A(n15214), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n15213) );
  XNOR2_X1 U16859 ( .A(n15213), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15206) );
  INV_X1 U16860 ( .A(n15209), .ZN(n15207) );
  NAND2_X1 U16861 ( .A1(n15207), .A2(n15210), .ZN(n15208) );
  XNOR2_X1 U16862 ( .A(n15208), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  AOI21_X1 U16863 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n15210), .A(n15209), 
        .ZN(n15222) );
  INV_X1 U16864 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15211) );
  NOR2_X1 U16865 ( .A1(n15211), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n15224) );
  INV_X1 U16866 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15223) );
  NOR2_X1 U16867 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15223), .ZN(n15212) );
  NOR2_X1 U16868 ( .A1(n15224), .A2(n15212), .ZN(n15217) );
  INV_X1 U16869 ( .A(n15213), .ZN(n15216) );
  NOR2_X1 U16870 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15214), .ZN(n15215) );
  AOI21_X1 U16871 ( .B1(n15216), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n15215), 
        .ZN(n15225) );
  XOR2_X1 U16872 ( .A(n15217), .B(n15225), .Z(n15219) );
  INV_X1 U16873 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15220) );
  XNOR2_X1 U16874 ( .A(n15219), .B(n15220), .ZN(n15218) );
  XNOR2_X1 U16875 ( .A(n15222), .B(n15218), .ZN(SUB_1596_U62) );
  NAND2_X1 U16876 ( .A1(n15219), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n15221) );
  OAI22_X1 U16877 ( .A1(n15225), .A2(n15224), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n15223), .ZN(n15228) );
  XNOR2_X1 U16878 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n15226) );
  XNOR2_X1 U16879 ( .A(n15226), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n15227) );
  XNOR2_X1 U16880 ( .A(n15228), .B(n15227), .ZN(n15229) );
  XNOR2_X1 U16881 ( .A(n15230), .B(n15229), .ZN(SUB_1596_U4) );
  AOI21_X1 U16882 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15231) );
  OAI21_X1 U16883 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15231), 
        .ZN(U28) );
  AOI21_X1 U16884 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15232) );
  OAI21_X1 U16885 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15232), 
        .ZN(U29) );
  XOR2_X1 U16886 ( .A(n15234), .B(n15233), .Z(n15235) );
  XNOR2_X1 U16887 ( .A(n15235), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  NOR2_X1 U16888 ( .A1(n15236), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n15238) );
  OR2_X1 U16889 ( .A1(n15237), .A2(n15238), .ZN(n15241) );
  INV_X1 U16890 ( .A(n15238), .ZN(n15240) );
  MUX2_X1 U16891 ( .A(n15241), .B(n15240), .S(n15239), .Z(n15243) );
  NAND2_X1 U16892 ( .A1(n15243), .A2(n15242), .ZN(n15246) );
  AOI22_X1 U16893 ( .A1(n15244), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15245) );
  OAI21_X1 U16894 ( .B1(n15247), .B2(n15246), .A(n15245), .ZN(P1_U3243) );
  NOR2_X1 U16895 ( .A1(n15280), .A2(n15248), .ZN(n15249) );
  AOI21_X1 U16896 ( .B1(n6538), .B2(P1_REG2_REG_7__SCAN_IN), .A(n15249), .ZN(
        n15250) );
  OAI21_X1 U16897 ( .B1(n15283), .B2(n15251), .A(n15250), .ZN(n15252) );
  INV_X1 U16898 ( .A(n15252), .ZN(n15257) );
  OAI22_X1 U16899 ( .A1(n15254), .A2(n15285), .B1(n15265), .B2(n15253), .ZN(
        n15255) );
  INV_X1 U16900 ( .A(n15255), .ZN(n15256) );
  OAI211_X1 U16901 ( .C1(n6538), .C2(n15258), .A(n15257), .B(n15256), .ZN(
        P1_U3286) );
  NOR2_X1 U16902 ( .A1(n15280), .A2(n15259), .ZN(n15260) );
  AOI21_X1 U16903 ( .B1(n6538), .B2(P1_REG2_REG_5__SCAN_IN), .A(n15260), .ZN(
        n15261) );
  OAI21_X1 U16904 ( .B1(n15283), .B2(n15262), .A(n15261), .ZN(n15263) );
  INV_X1 U16905 ( .A(n15263), .ZN(n15269) );
  OAI22_X1 U16906 ( .A1(n15266), .A2(n15285), .B1(n15265), .B2(n15264), .ZN(
        n15267) );
  INV_X1 U16907 ( .A(n15267), .ZN(n15268) );
  OAI211_X1 U16908 ( .C1(n6538), .C2(n15270), .A(n15269), .B(n15268), .ZN(
        P1_U3288) );
  XNOR2_X1 U16909 ( .A(n15271), .B(n15275), .ZN(n15319) );
  INV_X1 U16910 ( .A(n15272), .ZN(n15279) );
  NAND3_X1 U16911 ( .A1(n11359), .A2(n15275), .A3(n15274), .ZN(n15277) );
  AOI21_X1 U16912 ( .B1(n15273), .B2(n15277), .A(n15276), .ZN(n15278) );
  AOI211_X1 U16913 ( .C1(n10368), .C2(n15319), .A(n15279), .B(n15278), .ZN(
        n15316) );
  NOR2_X1 U16914 ( .A1(n15280), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n15281) );
  AOI21_X1 U16915 ( .B1(n6538), .B2(P1_REG2_REG_3__SCAN_IN), .A(n15281), .ZN(
        n15282) );
  OAI21_X1 U16916 ( .B1(n15283), .B2(n15315), .A(n15282), .ZN(n15284) );
  INV_X1 U16917 ( .A(n15284), .ZN(n15292) );
  INV_X1 U16918 ( .A(n15285), .ZN(n15290) );
  OAI211_X1 U16919 ( .C1(n15287), .C2(n15315), .A(n15286), .B(n10110), .ZN(
        n15314) );
  INV_X1 U16920 ( .A(n15314), .ZN(n15288) );
  AOI22_X1 U16921 ( .A1(n15290), .A2(n15319), .B1(n15289), .B2(n15288), .ZN(
        n15291) );
  OAI211_X1 U16922 ( .C1(n6538), .C2(n15316), .A(n15292), .B(n15291), .ZN(
        P1_U3290) );
  INV_X1 U16923 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15776) );
  NOR2_X1 U16924 ( .A1(n15293), .A2(n15776), .ZN(P1_U3294) );
  AND2_X1 U16925 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15859), .ZN(P1_U3295) );
  INV_X1 U16926 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15836) );
  NOR2_X1 U16927 ( .A1(n15293), .A2(n15836), .ZN(P1_U3296) );
  INV_X1 U16928 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15841) );
  NOR2_X1 U16929 ( .A1(n15293), .A2(n15841), .ZN(P1_U3297) );
  AND2_X1 U16930 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15859), .ZN(P1_U3298) );
  AND2_X1 U16931 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15859), .ZN(P1_U3300) );
  AND2_X1 U16932 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15859), .ZN(P1_U3301) );
  AND2_X1 U16933 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15859), .ZN(P1_U3302) );
  AND2_X1 U16934 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15859), .ZN(P1_U3303) );
  AND2_X1 U16935 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15859), .ZN(P1_U3304) );
  AND2_X1 U16936 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15859), .ZN(P1_U3305) );
  AND2_X1 U16937 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15859), .ZN(P1_U3306) );
  AND2_X1 U16938 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15859), .ZN(P1_U3307) );
  AND2_X1 U16939 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15859), .ZN(P1_U3308) );
  AND2_X1 U16940 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15859), .ZN(P1_U3309) );
  AND2_X1 U16941 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15859), .ZN(P1_U3310) );
  AND2_X1 U16942 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15859), .ZN(P1_U3311) );
  AND2_X1 U16943 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15859), .ZN(P1_U3312) );
  AND2_X1 U16944 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15859), .ZN(P1_U3313) );
  AND2_X1 U16945 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15859), .ZN(P1_U3314) );
  AND2_X1 U16946 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15859), .ZN(P1_U3315) );
  AND2_X1 U16947 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15859), .ZN(P1_U3316) );
  INV_X1 U16948 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15626) );
  NOR2_X1 U16949 ( .A1(n15293), .A2(n15626), .ZN(P1_U3317) );
  AND2_X1 U16950 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15859), .ZN(P1_U3318) );
  AND2_X1 U16951 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15859), .ZN(P1_U3319) );
  AND2_X1 U16952 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15859), .ZN(P1_U3320) );
  AND2_X1 U16953 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15859), .ZN(P1_U3321) );
  AND2_X1 U16954 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15859), .ZN(P1_U3322) );
  INV_X1 U16955 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15780) );
  NOR2_X1 U16956 ( .A1(n15293), .A2(n15780), .ZN(P1_U3323) );
  NAND2_X1 U16957 ( .A1(n15295), .A2(n15294), .ZN(n15297) );
  OAI211_X1 U16958 ( .C1(n15298), .C2(n15323), .A(n15297), .B(n15296), .ZN(
        n15301) );
  INV_X1 U16959 ( .A(n15299), .ZN(n15300) );
  AOI211_X1 U16960 ( .C1(n15339), .C2(n15302), .A(n15301), .B(n15300), .ZN(
        n15343) );
  AOI22_X1 U16961 ( .A1(n15342), .A2(n15343), .B1(n8743), .B2(n9554), .ZN(
        P1_U3462) );
  INV_X1 U16962 ( .A(n15311), .ZN(n15313) );
  INV_X1 U16963 ( .A(n15303), .ZN(n15304) );
  OAI211_X1 U16964 ( .C1(n15306), .C2(n15335), .A(n15305), .B(n15304), .ZN(
        n15307) );
  AOI21_X1 U16965 ( .B1(n15308), .B2(n15331), .A(n15307), .ZN(n15309) );
  OAI21_X1 U16966 ( .B1(n15311), .B2(n15310), .A(n15309), .ZN(n15312) );
  AOI21_X1 U16967 ( .B1(n10368), .B2(n15313), .A(n15312), .ZN(n15344) );
  AOI22_X1 U16968 ( .A1(n15342), .A2(n15344), .B1(n8761), .B2(n9554), .ZN(
        P1_U3465) );
  OAI21_X1 U16969 ( .B1(n15315), .B2(n15335), .A(n15314), .ZN(n15318) );
  INV_X1 U16970 ( .A(n15316), .ZN(n15317) );
  AOI211_X1 U16971 ( .C1(n15320), .C2(n15319), .A(n15318), .B(n15317), .ZN(
        n15345) );
  AOI22_X1 U16972 ( .A1(n15342), .A2(n15345), .B1(n8785), .B2(n9554), .ZN(
        P1_U3468) );
  INV_X1 U16973 ( .A(n15321), .ZN(n15328) );
  OAI22_X1 U16974 ( .A1(n15324), .A2(n15323), .B1(n15322), .B2(n15335), .ZN(
        n15327) );
  INV_X1 U16975 ( .A(n15325), .ZN(n15326) );
  AOI211_X1 U16976 ( .C1(n15328), .C2(n15339), .A(n15327), .B(n15326), .ZN(
        n15346) );
  INV_X1 U16977 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15329) );
  AOI22_X1 U16978 ( .A1(n15342), .A2(n15346), .B1(n15329), .B2(n9554), .ZN(
        P1_U3471) );
  AND3_X1 U16979 ( .A1(n11495), .A2(n15331), .A3(n15330), .ZN(n15338) );
  INV_X1 U16980 ( .A(n15332), .ZN(n15333) );
  OAI211_X1 U16981 ( .C1(n15336), .C2(n15335), .A(n15334), .B(n15333), .ZN(
        n15337) );
  AOI211_X1 U16982 ( .C1(n15340), .C2(n15339), .A(n15338), .B(n15337), .ZN(
        n15347) );
  INV_X1 U16983 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15341) );
  AOI22_X1 U16984 ( .A1(n15342), .A2(n15347), .B1(n15341), .B2(n9554), .ZN(
        P1_U3483) );
  AOI22_X1 U16985 ( .A1(n15348), .A2(n15343), .B1(n10719), .B2(n9548), .ZN(
        P1_U3529) );
  AOI22_X1 U16986 ( .A1(n15348), .A2(n15344), .B1(n10720), .B2(n9548), .ZN(
        P1_U3530) );
  AOI22_X1 U16987 ( .A1(n15348), .A2(n15345), .B1(n10723), .B2(n9548), .ZN(
        P1_U3531) );
  AOI22_X1 U16988 ( .A1(n15348), .A2(n15346), .B1(n10726), .B2(n9548), .ZN(
        P1_U3532) );
  AOI22_X1 U16989 ( .A1(n15348), .A2(n15347), .B1(n10736), .B2(n9548), .ZN(
        P1_U3536) );
  NOR2_X1 U16990 ( .A1(n15408), .A2(P2_U3947), .ZN(P2_U3087) );
  NAND2_X1 U16991 ( .A1(n15349), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15376) );
  NAND2_X1 U16992 ( .A1(n15350), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15351) );
  OAI211_X1 U16993 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(P2_STATE_REG_SCAN_IN), 
        .A(n15376), .B(n15351), .ZN(n15361) );
  OAI211_X1 U16994 ( .C1(n15354), .C2(n15353), .A(n15398), .B(n15352), .ZN(
        n15360) );
  OAI211_X1 U16995 ( .C1(n15357), .C2(n15356), .A(n15394), .B(n15355), .ZN(
        n15359) );
  NAND2_X1 U16996 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(n15408), .ZN(n15358) );
  NAND4_X1 U16997 ( .A1(n15361), .A2(n15360), .A3(n15359), .A4(n15358), .ZN(
        P2_U3216) );
  NAND2_X1 U16998 ( .A1(n15362), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15363) );
  OAI211_X1 U16999 ( .C1(P2_REG3_REG_4__SCAN_IN), .C2(P2_STATE_REG_SCAN_IN), 
        .A(n15376), .B(n15363), .ZN(n15373) );
  OAI211_X1 U17000 ( .C1(n15366), .C2(n15365), .A(n15398), .B(n15364), .ZN(
        n15372) );
  NAND2_X1 U17001 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15408), .ZN(n15371) );
  OAI211_X1 U17002 ( .C1(n15369), .C2(n15368), .A(n15394), .B(n15367), .ZN(
        n15370) );
  NAND4_X1 U17003 ( .A1(n15373), .A2(n15372), .A3(n15371), .A4(n15370), .ZN(
        P2_U3218) );
  NAND2_X1 U17004 ( .A1(P2_U3088), .A2(n15374), .ZN(n15375) );
  OAI211_X1 U17005 ( .C1(n15377), .C2(P2_U3088), .A(n15376), .B(n15375), .ZN(
        n15387) );
  OAI211_X1 U17006 ( .C1(n15380), .C2(n15379), .A(n15398), .B(n15378), .ZN(
        n15386) );
  NAND2_X1 U17007 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n15408), .ZN(n15385) );
  OAI211_X1 U17008 ( .C1(n15383), .C2(n15382), .A(n15394), .B(n15381), .ZN(
        n15384) );
  NAND4_X1 U17009 ( .A1(n15387), .A2(n15386), .A3(n15385), .A4(n15384), .ZN(
        P2_U3220) );
  INV_X1 U17010 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15407) );
  INV_X1 U17011 ( .A(n15388), .ZN(n15390) );
  NAND3_X1 U17012 ( .A1(n15391), .A2(n15390), .A3(n15389), .ZN(n15392) );
  NAND2_X1 U17013 ( .A1(n15393), .A2(n15392), .ZN(n15395) );
  NAND2_X1 U17014 ( .A1(n15395), .A2(n15394), .ZN(n15401) );
  XNOR2_X1 U17015 ( .A(n15397), .B(n15396), .ZN(n15399) );
  NAND2_X1 U17016 ( .A1(n15399), .A2(n15398), .ZN(n15400) );
  OAI211_X1 U17017 ( .C1(n15412), .C2(n15402), .A(n15401), .B(n15400), .ZN(
        n15403) );
  INV_X1 U17018 ( .A(n15403), .ZN(n15405) );
  OAI211_X1 U17019 ( .C1(n15407), .C2(n15406), .A(n15405), .B(n15404), .ZN(
        P2_U3226) );
  NAND2_X1 U17020 ( .A1(n15408), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n15409) );
  OAI211_X1 U17021 ( .C1(n15412), .C2(n15411), .A(n15410), .B(n15409), .ZN(
        n15413) );
  INV_X1 U17022 ( .A(n15413), .ZN(n15426) );
  AOI21_X1 U17023 ( .B1(n15416), .B2(n15415), .A(n15414), .ZN(n15418) );
  NAND2_X1 U17024 ( .A1(n15418), .A2(n15417), .ZN(n15425) );
  AOI211_X1 U17025 ( .C1(n15422), .C2(n15421), .A(n15420), .B(n15419), .ZN(
        n15423) );
  INV_X1 U17026 ( .A(n15423), .ZN(n15424) );
  NAND3_X1 U17027 ( .A1(n15426), .A2(n15425), .A3(n15424), .ZN(P2_U3227) );
  AND2_X1 U17028 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15429), .ZN(P2_U3266) );
  AND2_X1 U17029 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15429), .ZN(P2_U3267) );
  INV_X1 U17030 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15831) );
  NOR2_X1 U17031 ( .A1(n15428), .A2(n15831), .ZN(P2_U3268) );
  AND2_X1 U17032 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15429), .ZN(P2_U3269) );
  AND2_X1 U17033 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15429), .ZN(P2_U3270) );
  AND2_X1 U17034 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15429), .ZN(P2_U3271) );
  AND2_X1 U17035 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15429), .ZN(P2_U3272) );
  AND2_X1 U17036 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15429), .ZN(P2_U3273) );
  INV_X1 U17037 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15664) );
  NOR2_X1 U17038 ( .A1(n15428), .A2(n15664), .ZN(P2_U3274) );
  AND2_X1 U17039 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15429), .ZN(P2_U3275) );
  AND2_X1 U17040 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15429), .ZN(P2_U3276) );
  INV_X1 U17041 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15765) );
  NOR2_X1 U17042 ( .A1(n15428), .A2(n15765), .ZN(P2_U3277) );
  AND2_X1 U17043 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15429), .ZN(P2_U3278) );
  AND2_X1 U17044 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15429), .ZN(P2_U3279) );
  AND2_X1 U17045 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15429), .ZN(P2_U3280) );
  INV_X1 U17046 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15811) );
  NOR2_X1 U17047 ( .A1(n15428), .A2(n15811), .ZN(P2_U3281) );
  AND2_X1 U17048 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15429), .ZN(P2_U3282) );
  AND2_X1 U17049 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15429), .ZN(P2_U3283) );
  AND2_X1 U17050 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15429), .ZN(P2_U3284) );
  AND2_X1 U17051 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15429), .ZN(P2_U3285) );
  AND2_X1 U17052 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15429), .ZN(P2_U3286) );
  AND2_X1 U17053 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15429), .ZN(P2_U3287) );
  AND2_X1 U17054 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15429), .ZN(P2_U3288) );
  AND2_X1 U17055 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15429), .ZN(P2_U3289) );
  AND2_X1 U17056 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15429), .ZN(P2_U3290) );
  AND2_X1 U17057 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15429), .ZN(P2_U3291) );
  INV_X1 U17058 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15717) );
  NOR2_X1 U17059 ( .A1(n15428), .A2(n15717), .ZN(P2_U3292) );
  AND2_X1 U17060 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15429), .ZN(P2_U3293) );
  AND2_X1 U17061 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15429), .ZN(P2_U3294) );
  AND2_X1 U17062 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15429), .ZN(P2_U3295) );
  AOI22_X1 U17063 ( .A1(n15432), .A2(n15431), .B1(n15430), .B2(n15434), .ZN(
        P2_U3416) );
  AOI21_X1 U17064 ( .B1(n15435), .B2(n15434), .A(n15433), .ZN(P2_U3417) );
  INV_X1 U17065 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15436) );
  AOI22_X1 U17066 ( .A1(n15462), .A2(n15437), .B1(n15436), .B2(n15460), .ZN(
        P2_U3430) );
  INV_X1 U17067 ( .A(n15438), .ZN(n15440) );
  OAI21_X1 U17068 ( .B1(n15440), .B2(n15451), .A(n15439), .ZN(n15441) );
  NOR2_X1 U17069 ( .A1(n15442), .A2(n15441), .ZN(n15448) );
  NAND2_X1 U17070 ( .A1(n15445), .A2(n15443), .ZN(n15447) );
  NAND2_X1 U17071 ( .A1(n15445), .A2(n15444), .ZN(n15446) );
  INV_X1 U17072 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15449) );
  AOI22_X1 U17073 ( .A1(n15462), .A2(n15463), .B1(n15449), .B2(n15460), .ZN(
        P2_U3448) );
  INV_X1 U17074 ( .A(n15450), .ZN(n15459) );
  OAI22_X1 U17075 ( .A1(n15454), .A2(n15453), .B1(n15452), .B2(n15451), .ZN(
        n15457) );
  INV_X1 U17076 ( .A(n15455), .ZN(n15456) );
  AOI211_X1 U17077 ( .C1(n15459), .C2(n15458), .A(n15457), .B(n15456), .ZN(
        n15465) );
  INV_X1 U17078 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15461) );
  AOI22_X1 U17079 ( .A1(n15462), .A2(n15465), .B1(n15461), .B2(n15460), .ZN(
        P2_U3451) );
  AOI22_X1 U17080 ( .A1(n15466), .A2(n15463), .B1(n10609), .B2(n15464), .ZN(
        P2_U3505) );
  AOI22_X1 U17081 ( .A1(n15466), .A2(n15465), .B1(n10610), .B2(n15464), .ZN(
        P2_U3506) );
  NOR2_X1 U17082 ( .A1(P3_U3897), .A2(n15467), .ZN(P3_U3150) );
  AOI21_X1 U17083 ( .B1(n15477), .B2(n15469), .A(n15468), .ZN(n15471) );
  OAI222_X1 U17084 ( .A1(n15472), .A2(n15483), .B1(n15519), .B2(n15471), .C1(
        n15486), .C2(n15470), .ZN(n15473) );
  INV_X1 U17085 ( .A(n15473), .ZN(n15474) );
  OAI21_X1 U17086 ( .B1(n15500), .B2(n15475), .A(n15474), .ZN(P3_U3229) );
  AOI21_X1 U17087 ( .B1(n15478), .B2(n15477), .A(n15476), .ZN(n15479) );
  MUX2_X1 U17088 ( .A(n15480), .B(n15479), .S(n15500), .Z(n15481) );
  OAI21_X1 U17089 ( .B1(n15483), .B2(n15482), .A(n15481), .ZN(n15484) );
  INV_X1 U17090 ( .A(n15484), .ZN(n15485) );
  OAI21_X1 U17091 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(n15486), .A(n15485), .ZN(
        P3_U3230) );
  XNOR2_X1 U17092 ( .A(n15487), .B(n15489), .ZN(n15496) );
  OAI21_X1 U17093 ( .B1(n15490), .B2(n15489), .A(n15488), .ZN(n15526) );
  OAI22_X1 U17094 ( .A1(n15493), .A2(n15492), .B1(n7381), .B2(n15491), .ZN(
        n15494) );
  AOI21_X1 U17095 ( .B1(n15526), .B2(n15511), .A(n15494), .ZN(n15495) );
  OAI21_X1 U17096 ( .B1(n15508), .B2(n15496), .A(n15495), .ZN(n15524) );
  NOR2_X1 U17097 ( .A1(n15497), .A2(n15512), .ZN(n15525) );
  AOI22_X1 U17098 ( .A1(n15526), .A2(n15515), .B1(n15525), .B2(n15514), .ZN(
        n15498) );
  INV_X1 U17099 ( .A(n15498), .ZN(n15499) );
  AOI211_X1 U17100 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15516), .A(n15524), .B(
        n15499), .ZN(n15501) );
  AOI22_X1 U17101 ( .A1(n15519), .A2(n6899), .B1(n15501), .B2(n15500), .ZN(
        P3_U3231) );
  XNOR2_X1 U17102 ( .A(n15502), .B(n11276), .ZN(n15523) );
  XNOR2_X1 U17103 ( .A(n11276), .B(n15503), .ZN(n15509) );
  AOI22_X1 U17104 ( .A1(n13320), .A2(n15506), .B1(n15505), .B2(n15504), .ZN(
        n15507) );
  OAI21_X1 U17105 ( .B1(n15509), .B2(n15508), .A(n15507), .ZN(n15510) );
  AOI21_X1 U17106 ( .B1(n15511), .B2(n15523), .A(n15510), .ZN(n15520) );
  NOR2_X1 U17107 ( .A1(n15513), .A2(n15512), .ZN(n15522) );
  AOI22_X1 U17108 ( .A1(n15523), .A2(n15515), .B1(n15522), .B2(n15514), .ZN(
        n15518) );
  AOI22_X1 U17109 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(n15516), .B1(
        P3_REG2_REG_1__SCAN_IN), .B2(n15519), .ZN(n15517) );
  OAI221_X1 U17110 ( .B1(n15519), .B2(n15520), .C1(n15519), .C2(n15518), .A(
        n15517), .ZN(P3_U3232) );
  INV_X1 U17111 ( .A(n15520), .ZN(n15521) );
  AOI211_X1 U17112 ( .C1(n6716), .C2(n15523), .A(n15522), .B(n15521), .ZN(
        n15542) );
  AOI22_X1 U17113 ( .A1(n15540), .A2(n15542), .B1(n15598), .B2(n15539), .ZN(
        P3_U3393) );
  AOI211_X1 U17114 ( .C1(n6716), .C2(n15526), .A(n15525), .B(n15524), .ZN(
        n15543) );
  INV_X1 U17115 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15527) );
  AOI22_X1 U17116 ( .A1(n15540), .A2(n15543), .B1(n15527), .B2(n15539), .ZN(
        P3_U3396) );
  INV_X1 U17117 ( .A(n15528), .ZN(n15531) );
  AOI211_X1 U17118 ( .C1(n15531), .C2(n6716), .A(n15530), .B(n15529), .ZN(
        n15545) );
  INV_X1 U17119 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15532) );
  AOI22_X1 U17120 ( .A1(n15540), .A2(n15545), .B1(n15532), .B2(n15539), .ZN(
        P3_U3405) );
  INV_X1 U17121 ( .A(n15533), .ZN(n15538) );
  INV_X1 U17122 ( .A(n15534), .ZN(n15535) );
  AOI211_X1 U17123 ( .C1(n15538), .C2(n15537), .A(n15536), .B(n15535), .ZN(
        n15548) );
  AOI22_X1 U17124 ( .A1(n15540), .A2(n15548), .B1(n8121), .B2(n15539), .ZN(
        P3_U3408) );
  AOI22_X1 U17125 ( .A1(n15549), .A2(n15542), .B1(n15541), .B2(n15546), .ZN(
        P3_U3460) );
  AOI22_X1 U17126 ( .A1(n15549), .A2(n15543), .B1(n7477), .B2(n15546), .ZN(
        P3_U3461) );
  AOI22_X1 U17127 ( .A1(n15549), .A2(n15545), .B1(n15544), .B2(n15546), .ZN(
        P3_U3464) );
  AOI22_X1 U17128 ( .A1(n15549), .A2(n15548), .B1(n15547), .B2(n15546), .ZN(
        P3_U3465) );
  OR4_X1 U17129 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .A3(
        n8873), .A4(n15779), .ZN(n15568) );
  INV_X1 U17130 ( .A(n15550), .ZN(n15567) );
  NAND4_X1 U17131 ( .A1(n15747), .A2(n15551), .A3(n15807), .A4(
        P1_REG3_REG_11__SCAN_IN), .ZN(n15553) );
  NAND4_X1 U17132 ( .A1(n15797), .A2(P1_DATAO_REG_17__SCAN_IN), .A3(
        P3_REG2_REG_5__SCAN_IN), .A4(P3_REG0_REG_14__SCAN_IN), .ZN(n15552) );
  NOR2_X1 U17133 ( .A1(n15553), .A2(n15552), .ZN(n15562) );
  AND4_X1 U17134 ( .A1(n15556), .A2(n15555), .A3(n15554), .A4(n15716), .ZN(
        n15560) );
  INV_X1 U17135 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n15813) );
  INV_X1 U17136 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n15557) );
  NOR4_X1 U17137 ( .A1(P2_REG1_REG_23__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), 
        .A3(n15813), .A4(n15557), .ZN(n15558) );
  AND4_X1 U17138 ( .A1(n15816), .A2(n15783), .A3(P3_B_REG_SCAN_IN), .A4(n15558), .ZN(n15559) );
  NAND4_X1 U17139 ( .A1(n15562), .A2(n15561), .A3(n15560), .A4(n15559), .ZN(
        n15566) );
  NAND2_X1 U17140 ( .A1(n15564), .A2(n15563), .ZN(n15565) );
  NOR4_X1 U17141 ( .A1(n15568), .A2(n15567), .A3(n15566), .A4(n15565), .ZN(
        n15620) );
  NAND4_X1 U17142 ( .A1(P3_ADDR_REG_19__SCAN_IN), .A2(P1_REG2_REG_5__SCAN_IN), 
        .A3(n15569), .A4(n10720), .ZN(n15570) );
  NOR3_X1 U17143 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(n15571), .A3(n15570), .ZN(
        n15581) );
  INV_X1 U17144 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n15839) );
  NOR4_X1 U17145 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(P2_REG1_REG_9__SCAN_IN), 
        .A3(P3_IR_REG_22__SCAN_IN), .A4(n15839), .ZN(n15572) );
  NAND3_X1 U17146 ( .A1(SI_0_), .A2(P1_D_REG_28__SCAN_IN), .A3(n15572), .ZN(
        n15579) );
  NOR4_X1 U17147 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(P3_REG1_REG_11__SCAN_IN), 
        .A3(P3_DATAO_REG_13__SCAN_IN), .A4(n10086), .ZN(n15577) );
  NOR4_X1 U17148 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(SI_29_), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_REG0_REG_31__SCAN_IN), .ZN(n15576) );
  NOR4_X1 U17149 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P1_DATAO_REG_16__SCAN_IN), 
        .A3(P1_REG2_REG_4__SCAN_IN), .A4(n15755), .ZN(n15573) );
  NAND3_X1 U17150 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P2_REG0_REG_18__SCAN_IN), 
        .A3(n15573), .ZN(n15574) );
  NOR3_X1 U17151 ( .A1(n15574), .A2(n15737), .A3(P1_REG2_REG_18__SCAN_IN), 
        .ZN(n15575) );
  NAND3_X1 U17152 ( .A1(n15577), .A2(n15576), .A3(n15575), .ZN(n15578) );
  NOR4_X1 U17153 ( .A1(P2_REG0_REG_28__SCAN_IN), .A2(P3_REG2_REG_23__SCAN_IN), 
        .A3(n15579), .A4(n15578), .ZN(n15580) );
  NAND4_X1 U17154 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(n15581), .A3(n15580), .A4(
        n7477), .ZN(n15618) );
  INV_X1 U17155 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n15582) );
  INV_X1 U17156 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n15652) );
  NAND4_X1 U17157 ( .A1(n15583), .A2(n15582), .A3(n15652), .A4(n15703), .ZN(
        n15588) );
  INV_X1 U17158 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n15584) );
  NAND4_X1 U17159 ( .A1(n15586), .A2(n15585), .A3(n15584), .A4(
        P2_REG1_REG_13__SCAN_IN), .ZN(n15587) );
  NOR3_X1 U17160 ( .A1(n15639), .A2(n15588), .A3(n15587), .ZN(n15605) );
  NAND4_X1 U17161 ( .A1(n15589), .A2(P2_DATAO_REG_6__SCAN_IN), .A3(
        P1_DATAO_REG_5__SCAN_IN), .A4(P3_REG1_REG_21__SCAN_IN), .ZN(n15597) );
  NOR4_X1 U17162 ( .A1(P3_REG0_REG_0__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .A3(n11705), .A4(n15717), .ZN(n15593) );
  NOR4_X1 U17163 ( .A1(P2_REG0_REG_10__SCAN_IN), .A2(P3_REG1_REG_0__SCAN_IN), 
        .A3(n15708), .A4(n15705), .ZN(n15592) );
  NOR4_X1 U17164 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(P2_DATAO_REG_18__SCAN_IN), .A3(P3_REG3_REG_22__SCAN_IN), .A4(P2_DATAO_REG_31__SCAN_IN), .ZN(n15591) );
  NOR4_X1 U17165 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(SI_28_), .A3(n15702), 
        .A4(n11626), .ZN(n15590) );
  AND4_X1 U17166 ( .A1(n15593), .A2(n15592), .A3(n15591), .A4(n15590), .ZN(
        n15594) );
  NAND3_X1 U17167 ( .A1(n15650), .A2(n15595), .A3(n15594), .ZN(n15596) );
  NOR2_X1 U17168 ( .A1(n15597), .A2(n15596), .ZN(n15604) );
  NAND4_X1 U17169 ( .A1(n15598), .A2(n15767), .A3(SI_18_), .A4(SI_11_), .ZN(
        n15602) );
  INV_X1 U17170 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n15599) );
  NAND4_X1 U17171 ( .A1(n15600), .A2(n15599), .A3(P2_IR_REG_6__SCAN_IN), .A4(
        P2_IR_REG_20__SCAN_IN), .ZN(n15601) );
  NOR2_X1 U17172 ( .A1(n15602), .A2(n15601), .ZN(n15603) );
  NAND4_X1 U17173 ( .A1(n15605), .A2(n15604), .A3(n15603), .A4(
        P3_DATAO_REG_17__SCAN_IN), .ZN(n15609) );
  NOR4_X1 U17174 ( .A1(P3_REG2_REG_26__SCAN_IN), .A2(P3_REG2_REG_22__SCAN_IN), 
        .A3(P1_REG3_REG_19__SCAN_IN), .A4(n15606), .ZN(n15607) );
  NAND3_X1 U17175 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P1_REG3_REG_20__SCAN_IN), 
        .A3(n15607), .ZN(n15608) );
  NOR2_X1 U17176 ( .A1(n15609), .A2(n15608), .ZN(n15613) );
  NOR4_X1 U17177 ( .A1(P3_REG2_REG_21__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .A3(n15664), .A4(n12398), .ZN(n15612) );
  INV_X1 U17178 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15623) );
  NAND4_X1 U17179 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_REG0_REG_22__SCAN_IN), 
        .A3(n15623), .A4(n15625), .ZN(n15610) );
  NOR3_X1 U17180 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n15629), .A3(n15610), 
        .ZN(n15611) );
  NAND3_X1 U17181 ( .A1(n15613), .A2(n15612), .A3(n15611), .ZN(n15617) );
  NOR4_X1 U17182 ( .A1(P3_D_REG_8__SCAN_IN), .A2(P3_IR_REG_30__SCAN_IN), .A3(
        n15764), .A4(n15765), .ZN(n15615) );
  NOR4_X1 U17183 ( .A1(P1_REG0_REG_9__SCAN_IN), .A2(n15693), .A3(n13133), .A4(
        n15691), .ZN(n15614) );
  NAND2_X1 U17184 ( .A1(n15615), .A2(n15614), .ZN(n15616) );
  NOR3_X1 U17185 ( .A1(n15618), .A2(n15617), .A3(n15616), .ZN(n15619) );
  AOI21_X1 U17186 ( .B1(n15620), .B2(n15619), .A(P3_IR_REG_25__SCAN_IN), .ZN(
        n15858) );
  INV_X1 U17187 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n15622) );
  AOI22_X1 U17188 ( .A1(n15623), .A2(keyinput95), .B1(keyinput105), .B2(n15622), .ZN(n15621) );
  OAI221_X1 U17189 ( .B1(n15623), .B2(keyinput95), .C1(n15622), .C2(
        keyinput105), .A(n15621), .ZN(n15635) );
  AOI22_X1 U17190 ( .A1(n15626), .A2(keyinput82), .B1(keyinput114), .B2(n15625), .ZN(n15624) );
  OAI221_X1 U17191 ( .B1(n15626), .B2(keyinput82), .C1(n15625), .C2(
        keyinput114), .A(n15624), .ZN(n15634) );
  AOI22_X1 U17192 ( .A1(n15629), .A2(keyinput41), .B1(n15628), .B2(keyinput80), 
        .ZN(n15627) );
  OAI221_X1 U17193 ( .B1(n15629), .B2(keyinput41), .C1(n15628), .C2(keyinput80), .A(n15627), .ZN(n15633) );
  XNOR2_X1 U17194 ( .A(P3_REG1_REG_21__SCAN_IN), .B(keyinput64), .ZN(n15631)
         );
  XNOR2_X1 U17195 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput110), .ZN(n15630) );
  NAND2_X1 U17196 ( .A1(n15631), .A2(n15630), .ZN(n15632) );
  NOR4_X1 U17197 ( .A1(n15635), .A2(n15634), .A3(n15633), .A4(n15632), .ZN(
        n15677) );
  AOI22_X1 U17198 ( .A1(n15589), .A2(keyinput68), .B1(n15637), .B2(keyinput26), 
        .ZN(n15636) );
  OAI221_X1 U17199 ( .B1(n15589), .B2(keyinput68), .C1(n15637), .C2(keyinput26), .A(n15636), .ZN(n15647) );
  AOI22_X1 U17200 ( .A1(n15640), .A2(keyinput93), .B1(keyinput14), .B2(n15639), 
        .ZN(n15638) );
  OAI221_X1 U17201 ( .B1(n15640), .B2(keyinput93), .C1(n15639), .C2(keyinput14), .A(n15638), .ZN(n15646) );
  AOI22_X1 U17202 ( .A1(n13200), .A2(keyinput125), .B1(n13145), .B2(keyinput0), 
        .ZN(n15641) );
  OAI221_X1 U17203 ( .B1(n13200), .B2(keyinput125), .C1(n13145), .C2(keyinput0), .A(n15641), .ZN(n15645) );
  XNOR2_X1 U17204 ( .A(P1_REG3_REG_20__SCAN_IN), .B(keyinput59), .ZN(n15643)
         );
  XNOR2_X1 U17205 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput101), .ZN(n15642) );
  NAND2_X1 U17206 ( .A1(n15643), .A2(n15642), .ZN(n15644) );
  NOR4_X1 U17207 ( .A1(n15647), .A2(n15646), .A3(n15645), .A4(n15644), .ZN(
        n15676) );
  AOI22_X1 U17208 ( .A1(n15650), .A2(keyinput85), .B1(keyinput33), .B2(n15649), 
        .ZN(n15648) );
  OAI221_X1 U17209 ( .B1(n15650), .B2(keyinput85), .C1(n15649), .C2(keyinput33), .A(n15648), .ZN(n15660) );
  XNOR2_X1 U17210 ( .A(n15651), .B(keyinput5), .ZN(n15659) );
  XNOR2_X1 U17211 ( .A(n15652), .B(keyinput90), .ZN(n15658) );
  XNOR2_X1 U17212 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput77), .ZN(n15656) );
  XNOR2_X1 U17213 ( .A(P1_REG3_REG_19__SCAN_IN), .B(keyinput53), .ZN(n15655)
         );
  XNOR2_X1 U17214 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput70), .ZN(n15654)
         );
  XNOR2_X1 U17215 ( .A(SI_30_), .B(keyinput27), .ZN(n15653) );
  NAND4_X1 U17216 ( .A1(n15656), .A2(n15655), .A3(n15654), .A4(n15653), .ZN(
        n15657) );
  NOR4_X1 U17217 ( .A1(n15660), .A2(n15659), .A3(n15658), .A4(n15657), .ZN(
        n15675) );
  AOI22_X1 U17218 ( .A1(n13210), .A2(keyinput126), .B1(keyinput38), .B2(n12398), .ZN(n15661) );
  OAI221_X1 U17219 ( .B1(n13210), .B2(keyinput126), .C1(n12398), .C2(
        keyinput38), .A(n15661), .ZN(n15673) );
  INV_X1 U17220 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n15663) );
  AOI22_X1 U17221 ( .A1(n15664), .A2(keyinput3), .B1(keyinput22), .B2(n15663), 
        .ZN(n15662) );
  OAI221_X1 U17222 ( .B1(n15664), .B2(keyinput3), .C1(n15663), .C2(keyinput22), 
        .A(n15662), .ZN(n15672) );
  AOI22_X1 U17223 ( .A1(n15667), .A2(keyinput91), .B1(keyinput69), .B2(n15666), 
        .ZN(n15665) );
  OAI221_X1 U17224 ( .B1(n15667), .B2(keyinput91), .C1(n15666), .C2(keyinput69), .A(n15665), .ZN(n15671) );
  XOR2_X1 U17225 ( .A(n15598), .B(keyinput13), .Z(n15669) );
  XNOR2_X1 U17226 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput78), .ZN(n15668) );
  NAND2_X1 U17227 ( .A1(n15669), .A2(n15668), .ZN(n15670) );
  NOR4_X1 U17228 ( .A1(n15673), .A2(n15672), .A3(n15671), .A4(n15670), .ZN(
        n15674) );
  NAND4_X1 U17229 ( .A1(n15677), .A2(n15676), .A3(n15675), .A4(n15674), .ZN(
        n15856) );
  INV_X1 U17230 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15679) );
  AOI22_X1 U17231 ( .A1(n8873), .A2(keyinput48), .B1(n15679), .B2(keyinput32), 
        .ZN(n15678) );
  OAI221_X1 U17232 ( .B1(n8873), .B2(keyinput48), .C1(n15679), .C2(keyinput32), 
        .A(n15678), .ZN(n15689) );
  AOI22_X1 U17233 ( .A1(n15682), .A2(keyinput10), .B1(n15681), .B2(keyinput7), 
        .ZN(n15680) );
  OAI221_X1 U17234 ( .B1(n15682), .B2(keyinput10), .C1(n15681), .C2(keyinput7), 
        .A(n15680), .ZN(n15688) );
  XOR2_X1 U17235 ( .A(n15585), .B(keyinput46), .Z(n15686) );
  XNOR2_X1 U17236 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(keyinput87), .ZN(n15685) );
  XNOR2_X1 U17237 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput99), .ZN(n15684) );
  XNOR2_X1 U17238 ( .A(P3_IR_REG_13__SCAN_IN), .B(keyinput56), .ZN(n15683) );
  NAND4_X1 U17239 ( .A1(n15686), .A2(n15685), .A3(n15684), .A4(n15683), .ZN(
        n15687) );
  NOR3_X1 U17240 ( .A1(n15689), .A2(n15688), .A3(n15687), .ZN(n15732) );
  AOI22_X1 U17241 ( .A1(n15691), .A2(keyinput119), .B1(keyinput40), .B2(n8914), 
        .ZN(n15690) );
  OAI221_X1 U17242 ( .B1(n15691), .B2(keyinput119), .C1(n8914), .C2(keyinput40), .A(n15690), .ZN(n15700) );
  AOI22_X1 U17243 ( .A1(n13133), .A2(keyinput102), .B1(keyinput31), .B2(n15693), .ZN(n15692) );
  OAI221_X1 U17244 ( .B1(n13133), .B2(keyinput102), .C1(n15693), .C2(
        keyinput31), .A(n15692), .ZN(n15699) );
  XOR2_X1 U17245 ( .A(n15551), .B(keyinput79), .Z(n15697) );
  XNOR2_X1 U17246 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput34), .ZN(n15696) );
  XNOR2_X1 U17247 ( .A(P2_REG0_REG_10__SCAN_IN), .B(keyinput121), .ZN(n15695)
         );
  XNOR2_X1 U17248 ( .A(P3_REG1_REG_0__SCAN_IN), .B(keyinput71), .ZN(n15694) );
  NAND4_X1 U17249 ( .A1(n15697), .A2(n15696), .A3(n15695), .A4(n15694), .ZN(
        n15698) );
  NOR3_X1 U17250 ( .A1(n15700), .A2(n15699), .A3(n15698), .ZN(n15731) );
  AOI22_X1 U17251 ( .A1(n15703), .A2(keyinput4), .B1(keyinput39), .B2(n15702), 
        .ZN(n15701) );
  OAI221_X1 U17252 ( .B1(n15703), .B2(keyinput4), .C1(n15702), .C2(keyinput39), 
        .A(n15701), .ZN(n15714) );
  AOI22_X1 U17253 ( .A1(n15705), .A2(keyinput81), .B1(n15583), .B2(keyinput19), 
        .ZN(n15704) );
  OAI221_X1 U17254 ( .B1(n15705), .B2(keyinput81), .C1(n15583), .C2(keyinput19), .A(n15704), .ZN(n15713) );
  AOI22_X1 U17255 ( .A1(n15708), .A2(keyinput58), .B1(n15707), .B2(keyinput127), .ZN(n15706) );
  OAI221_X1 U17256 ( .B1(n15708), .B2(keyinput58), .C1(n15707), .C2(
        keyinput127), .A(n15706), .ZN(n15712) );
  XNOR2_X1 U17257 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput97), .ZN(n15710)
         );
  XNOR2_X1 U17258 ( .A(P2_REG1_REG_19__SCAN_IN), .B(keyinput117), .ZN(n15709)
         );
  NAND2_X1 U17259 ( .A1(n15710), .A2(n15709), .ZN(n15711) );
  NOR4_X1 U17260 ( .A1(n15714), .A2(n15713), .A3(n15712), .A4(n15711), .ZN(
        n15730) );
  AOI22_X1 U17261 ( .A1(n11705), .A2(keyinput50), .B1(keyinput11), .B2(n15716), 
        .ZN(n15715) );
  OAI221_X1 U17262 ( .B1(n11705), .B2(keyinput50), .C1(n15716), .C2(keyinput11), .A(n15715), .ZN(n15721) );
  XNOR2_X1 U17263 ( .A(n15717), .B(keyinput103), .ZN(n15720) );
  XNOR2_X1 U17264 ( .A(n15718), .B(keyinput9), .ZN(n15719) );
  OR3_X1 U17265 ( .A1(n15721), .A2(n15720), .A3(n15719), .ZN(n15728) );
  AOI22_X1 U17266 ( .A1(n15723), .A2(keyinput124), .B1(keyinput8), .B2(n8065), 
        .ZN(n15722) );
  OAI221_X1 U17267 ( .B1(n15723), .B2(keyinput124), .C1(n8065), .C2(keyinput8), 
        .A(n15722), .ZN(n15727) );
  AOI22_X1 U17268 ( .A1(n11626), .A2(keyinput25), .B1(n15725), .B2(keyinput111), .ZN(n15724) );
  OAI221_X1 U17269 ( .B1(n11626), .B2(keyinput25), .C1(n15725), .C2(
        keyinput111), .A(n15724), .ZN(n15726) );
  NOR3_X1 U17270 ( .A1(n15728), .A2(n15727), .A3(n15726), .ZN(n15729) );
  NAND4_X1 U17271 ( .A1(n15732), .A2(n15731), .A3(n15730), .A4(n15729), .ZN(
        n15855) );
  AOI22_X1 U17272 ( .A1(n15735), .A2(keyinput47), .B1(keyinput76), .B2(n15734), 
        .ZN(n15733) );
  OAI221_X1 U17273 ( .B1(n15735), .B2(keyinput47), .C1(n15734), .C2(keyinput76), .A(n15733), .ZN(n15745) );
  AOI22_X1 U17274 ( .A1(n15737), .A2(keyinput83), .B1(keyinput65), .B2(n9004), 
        .ZN(n15736) );
  OAI221_X1 U17275 ( .B1(n15737), .B2(keyinput83), .C1(n9004), .C2(keyinput65), 
        .A(n15736), .ZN(n15744) );
  AOI22_X1 U17276 ( .A1(n15739), .A2(keyinput12), .B1(n10086), .B2(keyinput6), 
        .ZN(n15738) );
  OAI221_X1 U17277 ( .B1(n15739), .B2(keyinput12), .C1(n10086), .C2(keyinput6), 
        .A(n15738), .ZN(n15743) );
  XNOR2_X1 U17278 ( .A(P3_IR_REG_7__SCAN_IN), .B(keyinput29), .ZN(n15741) );
  XNOR2_X1 U17279 ( .A(P2_REG0_REG_18__SCAN_IN), .B(keyinput116), .ZN(n15740)
         );
  NAND2_X1 U17280 ( .A1(n15741), .A2(n15740), .ZN(n15742) );
  NOR4_X1 U17281 ( .A1(n15745), .A2(n15744), .A3(n15743), .A4(n15742), .ZN(
        n15793) );
  INV_X1 U17282 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n15747) );
  AOI22_X1 U17283 ( .A1(n15748), .A2(keyinput43), .B1(keyinput20), .B2(n15747), 
        .ZN(n15746) );
  OAI221_X1 U17284 ( .B1(n15748), .B2(keyinput43), .C1(n15747), .C2(keyinput20), .A(n15746), .ZN(n15751) );
  XNOR2_X1 U17285 ( .A(n15749), .B(keyinput61), .ZN(n15750) );
  NOR2_X1 U17286 ( .A1(n15751), .A2(n15750), .ZN(n15760) );
  AOI22_X1 U17287 ( .A1(n10720), .A2(keyinput60), .B1(n9566), .B2(keyinput66), 
        .ZN(n15752) );
  OAI221_X1 U17288 ( .B1(n10720), .B2(keyinput60), .C1(n9566), .C2(keyinput66), 
        .A(n15752), .ZN(n15753) );
  INV_X1 U17289 ( .A(n15753), .ZN(n15759) );
  AOI22_X1 U17290 ( .A1(n15755), .A2(keyinput51), .B1(keyinput17), .B2(n11305), 
        .ZN(n15754) );
  OAI221_X1 U17291 ( .B1(n15755), .B2(keyinput51), .C1(n11305), .C2(keyinput17), .A(n15754), .ZN(n15756) );
  INV_X1 U17292 ( .A(n15756), .ZN(n15758) );
  XNOR2_X1 U17293 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(keyinput37), .ZN(n15757)
         );
  AND4_X1 U17294 ( .A1(n15760), .A2(n15759), .A3(n15758), .A4(n15757), .ZN(
        n15792) );
  AOI22_X1 U17295 ( .A1(n15762), .A2(keyinput44), .B1(keyinput42), .B2(n13475), 
        .ZN(n15761) );
  OAI221_X1 U17296 ( .B1(n15762), .B2(keyinput44), .C1(n13475), .C2(keyinput42), .A(n15761), .ZN(n15774) );
  AOI22_X1 U17297 ( .A1(n15765), .A2(keyinput106), .B1(keyinput74), .B2(n15764), .ZN(n15763) );
  OAI221_X1 U17298 ( .B1(n15765), .B2(keyinput106), .C1(n15764), .C2(
        keyinput74), .A(n15763), .ZN(n15773) );
  AOI22_X1 U17299 ( .A1(n15768), .A2(keyinput88), .B1(keyinput107), .B2(n15767), .ZN(n15766) );
  OAI221_X1 U17300 ( .B1(n15768), .B2(keyinput88), .C1(n15767), .C2(
        keyinput107), .A(n15766), .ZN(n15772) );
  XNOR2_X1 U17301 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput98), .ZN(n15770) );
  XNOR2_X1 U17302 ( .A(P2_REG1_REG_22__SCAN_IN), .B(keyinput36), .ZN(n15769)
         );
  NAND2_X1 U17303 ( .A1(n15770), .A2(n15769), .ZN(n15771) );
  NOR4_X1 U17304 ( .A1(n15774), .A2(n15773), .A3(n15772), .A4(n15771), .ZN(
        n15791) );
  AOI22_X1 U17305 ( .A1(n15777), .A2(keyinput49), .B1(keyinput113), .B2(n15776), .ZN(n15775) );
  OAI221_X1 U17306 ( .B1(n15777), .B2(keyinput49), .C1(n15776), .C2(
        keyinput113), .A(n15775), .ZN(n15789) );
  AOI22_X1 U17307 ( .A1(n15780), .A2(keyinput30), .B1(keyinput84), .B2(n15779), 
        .ZN(n15778) );
  OAI221_X1 U17308 ( .B1(n15780), .B2(keyinput30), .C1(n15779), .C2(keyinput84), .A(n15778), .ZN(n15788) );
  AOI22_X1 U17309 ( .A1(n15783), .A2(keyinput92), .B1(keyinput16), .B2(n15782), 
        .ZN(n15781) );
  OAI221_X1 U17310 ( .B1(n15783), .B2(keyinput92), .C1(n15782), .C2(keyinput16), .A(n15781), .ZN(n15787) );
  XOR2_X1 U17311 ( .A(n14344), .B(keyinput108), .Z(n15785) );
  XNOR2_X1 U17312 ( .A(SI_11_), .B(keyinput67), .ZN(n15784) );
  NAND2_X1 U17313 ( .A1(n15785), .A2(n15784), .ZN(n15786) );
  NOR4_X1 U17314 ( .A1(n15789), .A2(n15788), .A3(n15787), .A4(n15786), .ZN(
        n15790) );
  NAND4_X1 U17315 ( .A1(n15793), .A2(n15792), .A3(n15791), .A4(n15790), .ZN(
        n15854) );
  AOI22_X1 U17316 ( .A1(n15795), .A2(keyinput62), .B1(keyinput23), .B2(n15555), 
        .ZN(n15794) );
  OAI221_X1 U17317 ( .B1(n15795), .B2(keyinput62), .C1(n15555), .C2(keyinput23), .A(n15794), .ZN(n15806) );
  AOI22_X1 U17318 ( .A1(n15798), .A2(keyinput94), .B1(keyinput24), .B2(n15797), 
        .ZN(n15796) );
  OAI221_X1 U17319 ( .B1(n15798), .B2(keyinput94), .C1(n15797), .C2(keyinput24), .A(n15796), .ZN(n15805) );
  INV_X1 U17320 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n15800) );
  AOI22_X1 U17321 ( .A1(n8414), .A2(keyinput115), .B1(n15800), .B2(keyinput18), 
        .ZN(n15799) );
  OAI221_X1 U17322 ( .B1(n8414), .B2(keyinput115), .C1(n15800), .C2(keyinput18), .A(n15799), .ZN(n15804) );
  XNOR2_X1 U17323 ( .A(P3_REG0_REG_14__SCAN_IN), .B(keyinput52), .ZN(n15802)
         );
  XNOR2_X1 U17324 ( .A(P3_B_REG_SCAN_IN), .B(keyinput123), .ZN(n15801) );
  NAND2_X1 U17325 ( .A1(n15802), .A2(n15801), .ZN(n15803) );
  NOR4_X1 U17326 ( .A1(n15806), .A2(n15805), .A3(n15804), .A4(n15803), .ZN(
        n15852) );
  XNOR2_X1 U17327 ( .A(n15807), .B(keyinput54), .ZN(n15809) );
  XOR2_X1 U17328 ( .A(P2_REG1_REG_25__SCAN_IN), .B(keyinput73), .Z(n15808) );
  AOI211_X1 U17329 ( .C1(keyinput45), .C2(n15810), .A(n15809), .B(n15808), 
        .ZN(n15822) );
  XOR2_X1 U17330 ( .A(keyinput15), .B(n15811), .Z(n15821) );
  INV_X1 U17331 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n15814) );
  AOI22_X1 U17332 ( .A1(n15814), .A2(keyinput72), .B1(n15813), .B2(keyinput118), .ZN(n15812) );
  OAI221_X1 U17333 ( .B1(n15814), .B2(keyinput72), .C1(n15813), .C2(
        keyinput118), .A(n15812), .ZN(n15819) );
  XNOR2_X1 U17334 ( .A(n15815), .B(keyinput109), .ZN(n15818) );
  XNOR2_X1 U17335 ( .A(n15816), .B(keyinput63), .ZN(n15817) );
  NOR3_X1 U17336 ( .A1(n15819), .A2(n15818), .A3(n15817), .ZN(n15820) );
  AND3_X1 U17337 ( .A1(n15822), .A2(n15821), .A3(n15820), .ZN(n15851) );
  XOR2_X1 U17338 ( .A(P1_REG2_REG_26__SCAN_IN), .B(keyinput86), .Z(n15826) );
  XOR2_X1 U17339 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput1), .Z(n15825) );
  XNOR2_X1 U17340 ( .A(n15823), .B(keyinput112), .ZN(n15824) );
  NOR3_X1 U17341 ( .A1(n15826), .A2(n15825), .A3(n15824), .ZN(n15829) );
  XNOR2_X1 U17342 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput96), .ZN(n15828) );
  XNOR2_X1 U17343 ( .A(P3_REG1_REG_7__SCAN_IN), .B(keyinput89), .ZN(n15827) );
  NAND3_X1 U17344 ( .A1(n15829), .A2(n15828), .A3(n15827), .ZN(n15834) );
  AOI22_X1 U17345 ( .A1(n7477), .A2(keyinput21), .B1(keyinput28), .B2(n10757), 
        .ZN(n15830) );
  OAI221_X1 U17346 ( .B1(n7477), .B2(keyinput21), .C1(n10757), .C2(keyinput28), 
        .A(n15830), .ZN(n15833) );
  XNOR2_X1 U17347 ( .A(n15831), .B(keyinput75), .ZN(n15832) );
  NOR3_X1 U17348 ( .A1(n15834), .A2(n15833), .A3(n15832), .ZN(n15850) );
  INV_X1 U17349 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n15837) );
  AOI22_X1 U17350 ( .A1(n15837), .A2(keyinput100), .B1(keyinput120), .B2(
        n15836), .ZN(n15835) );
  OAI221_X1 U17351 ( .B1(n15837), .B2(keyinput100), .C1(n15836), .C2(
        keyinput120), .A(n15835), .ZN(n15848) );
  AOI22_X1 U17352 ( .A1(n15840), .A2(keyinput35), .B1(keyinput57), .B2(n15839), 
        .ZN(n15838) );
  OAI221_X1 U17353 ( .B1(n15840), .B2(keyinput35), .C1(n15839), .C2(keyinput57), .A(n15838), .ZN(n15847) );
  XNOR2_X1 U17354 ( .A(n15841), .B(keyinput2), .ZN(n15846) );
  XNOR2_X1 U17355 ( .A(P3_IR_REG_22__SCAN_IN), .B(keyinput104), .ZN(n15844) );
  XNOR2_X1 U17356 ( .A(SI_0_), .B(keyinput122), .ZN(n15843) );
  XNOR2_X1 U17357 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(keyinput55), .ZN(n15842) );
  NAND3_X1 U17358 ( .A1(n15844), .A2(n15843), .A3(n15842), .ZN(n15845) );
  NOR4_X1 U17359 ( .A1(n15848), .A2(n15847), .A3(n15846), .A4(n15845), .ZN(
        n15849) );
  NAND4_X1 U17360 ( .A1(n15852), .A2(n15851), .A3(n15850), .A4(n15849), .ZN(
        n15853) );
  NOR4_X1 U17361 ( .A1(n15856), .A2(n15855), .A3(n15854), .A4(n15853), .ZN(
        n15857) );
  OAI21_X1 U17362 ( .B1(keyinput45), .B2(n15858), .A(n15857), .ZN(n15861) );
  NAND2_X1 U17363 ( .A1(n15859), .A2(P1_D_REG_26__SCAN_IN), .ZN(n15860) );
  XOR2_X1 U17364 ( .A(n15861), .B(n15860), .Z(P1_U3299) );
  AND2_X1 U17365 ( .A1(n15863), .A2(n15862), .ZN(n15864) );
  XOR2_X1 U17366 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15864), .Z(SUB_1596_U60) );
  AOI21_X1 U17367 ( .B1(n15867), .B2(n15866), .A(n15865), .ZN(SUB_1596_U5) );
  NAND2_X2 U7338 ( .A1(n6589), .A2(n7593), .ZN(n13906) );
  INV_X1 U7281 ( .A(n9912), .ZN(n14152) );
  INV_X1 U12061 ( .A(n10190), .ZN(n10270) );
  INV_X2 U7343 ( .A(n9316), .ZN(n8803) );
  XOR2_X1 U7280 ( .A(n10270), .B(n10184), .Z(n12292) );
  CLKBUF_X1 U7283 ( .A(n9655), .Z(n13788) );
  INV_X1 U7305 ( .A(n9324), .ZN(n9088) );
  CLKBUF_X1 U7654 ( .A(n10109), .Z(n15323) );
  CLKBUF_X1 U7683 ( .A(n8508), .Z(n7080) );
  NAND2_X1 U9123 ( .A1(n8933), .A2(n8936), .ZN(n10570) );
endmodule

