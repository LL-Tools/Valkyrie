

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, 
        DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, 
        DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, 
        DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, 
        DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, 
        DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, 
        DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_,
         DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_,
         DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_,
         DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_,
         DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_,
         DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
         HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN,
         P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN,
         P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN,
         P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN,
         P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN,
         P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN,
         P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN,
         P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN,
         P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN,
         P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
         P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
         P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
         P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
         P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
         P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
         P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
         P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
         P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
         P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
         P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN,
         P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
         P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
         P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
         P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN,
         P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
         P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
         P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN,
         P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
         P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
         P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN,
         P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
         P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
         P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN,
         P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN,
         P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN,
         P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN,
         P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN,
         P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
         P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
         P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN,
         P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
         P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
         P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN,
         P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
         P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
         P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN,
         P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
         P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
         P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
         P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
         P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330;

  OR2_X2 U11068 ( .A1(n21232), .A2(n21256), .ZN(n21259) );
  AND2_X1 U11069 ( .A1(n16333), .A2(n11191), .ZN(n15972) );
  NOR2_X1 U11070 ( .A1(n15747), .A2(n19922), .ZN(n15605) );
  NAND2_X1 U11071 ( .A1(n14055), .A2(n14054), .ZN(n15066) );
  INV_X1 U11072 ( .A(n18190), .ZN(n18189) );
  NAND2_X1 U11073 ( .A1(n13672), .A2(n13644), .ZN(n21821) );
  NAND2_X2 U11074 ( .A1(n13864), .A2(n10981), .ZN(n13869) );
  AND2_X1 U11075 ( .A1(n14025), .A2(n13591), .ZN(n11129) );
  NAND2_X2 U11076 ( .A1(n20652), .A2(n11634), .ZN(n20788) );
  CLKBUF_X2 U11077 ( .A(n11899), .Z(n12622) );
  INV_X2 U11078 ( .A(n12535), .ZN(n12689) );
  OR2_X1 U11079 ( .A1(n11926), .A2(n11925), .ZN(n11927) );
  OAI21_X1 U11080 ( .B1(n13590), .B2(n13550), .A(n13575), .ZN(n13576) );
  AOI21_X1 U11081 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11931), .ZN(n12261) );
  INV_X1 U11082 ( .A(n19642), .ZN(n12651) );
  INV_X1 U11083 ( .A(n12282), .ZN(n10980) );
  OR2_X1 U11084 ( .A1(n11889), .A2(n12641), .ZN(n11392) );
  INV_X1 U11085 ( .A(n13026), .ZN(n13108) );
  AND2_X1 U11086 ( .A1(n11975), .A2(n11832), .ZN(n13117) );
  AND2_X1 U11087 ( .A1(n11975), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13022) );
  AND2_X1 U11088 ( .A1(n15777), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11991) );
  AND2_X1 U11089 ( .A1(n11008), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13101) );
  AND2_X1 U11090 ( .A1(n13083), .A2(n11970), .ZN(n13102) );
  AND2_X1 U11091 ( .A1(n13083), .A2(n14939), .ZN(n11996) );
  CLKBUF_X2 U11092 ( .A(n11561), .Z(n10972) );
  NAND2_X1 U11093 ( .A1(n11877), .A2(n11876), .ZN(n11881) );
  INV_X2 U11094 ( .A(n17731), .ZN(n17850) );
  OR3_X1 U11095 ( .A1(n11420), .A2(n11421), .A3(n15640), .ZN(n11506) );
  BUF_X1 U11096 ( .A(n14419), .Z(n13529) );
  CLKBUF_X2 U11098 ( .A(n13519), .Z(n10970) );
  CLKBUF_X2 U11099 ( .A(n13604), .Z(n14770) );
  CLKBUF_X2 U11100 ( .A(n13514), .Z(n14479) );
  CLKBUF_X2 U11101 ( .A(n11561), .Z(n10971) );
  CLKBUF_X2 U11102 ( .A(n13431), .Z(n13513) );
  CLKBUF_X2 U11103 ( .A(n11869), .Z(n19703) );
  NOR2_X1 U11104 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20822), .ZN(
        n11469) );
  NAND2_X1 U11105 ( .A1(n13488), .A2(n13487), .ZN(n13836) );
  INV_X1 U11106 ( .A(n13491), .ZN(n21935) );
  AND4_X1 U11107 ( .A1(n13423), .A2(n13422), .A3(n13421), .A4(n13420), .ZN(
        n13428) );
  AND4_X1 U11108 ( .A1(n13409), .A2(n13408), .A3(n13407), .A4(n13406), .ZN(
        n11039) );
  AND2_X2 U11109 ( .A1(n14941), .A2(n14972), .ZN(n15791) );
  AND4_X1 U11110 ( .A1(n13374), .A2(n13373), .A3(n13372), .A4(n13371), .ZN(
        n13380) );
  AND4_X1 U11111 ( .A1(n13389), .A2(n13388), .A3(n13387), .A4(n13386), .ZN(
        n13390) );
  AND2_X1 U11112 ( .A1(n14771), .A2(n14915), .ZN(n13432) );
  BUF_X2 U11113 ( .A(n13445), .Z(n10975) );
  AND2_X2 U11114 ( .A1(n13375), .A2(n14915), .ZN(n13451) );
  AND2_X2 U11115 ( .A1(n14915), .A2(n14763), .ZN(n13433) );
  AND2_X2 U11116 ( .A1(n13551), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13381) );
  INV_X4 U11117 ( .A(n11764), .ZN(n10979) );
  NOR2_X1 U11119 ( .A1(n13495), .A2(n13429), .ZN(n13430) );
  AND2_X1 U11120 ( .A1(n14771), .A2(n11176), .ZN(n13514) );
  AND2_X1 U11121 ( .A1(n11176), .A2(n14764), .ZN(n13450) );
  AND3_X1 U11122 ( .A1(n13378), .A2(n13377), .A3(n13376), .ZN(n11418) );
  AND2_X2 U11123 ( .A1(n14941), .A2(n14972), .ZN(n10965) );
  BUF_X1 U11124 ( .A(n13484), .Z(n13786) );
  AND4_X1 U11125 ( .A1(n13405), .A2(n13404), .A3(n13403), .A4(n13402), .ZN(
        n13410) );
  NOR2_X1 U11126 ( .A1(n13603), .A2(n17186), .ZN(n13814) );
  AND2_X1 U11127 ( .A1(n15792), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12012) );
  NAND3_X1 U11128 ( .A1(n11902), .A2(n11887), .A3(n11392), .ZN(n11915) );
  NAND2_X1 U11129 ( .A1(n13711), .A2(n13710), .ZN(n13737) );
  AND3_X1 U11130 ( .A1(n13481), .A2(n13479), .A3(n13480), .ZN(n13494) );
  INV_X1 U11131 ( .A(n12400), .ZN(n12634) );
  NAND2_X1 U11132 ( .A1(n11780), .A2(n11779), .ZN(n12400) );
  NOR2_X1 U11133 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11422), .ZN(
        n11437) );
  NAND2_X1 U11135 ( .A1(n15925), .A2(n11326), .ZN(n15844) );
  CLKBUF_X3 U11137 ( .A(n12634), .Z(n12539) );
  INV_X1 U11138 ( .A(n12539), .ZN(n12357) );
  NOR2_X1 U11139 ( .A1(n16596), .A2(n11148), .ZN(n16591) );
  INV_X2 U11140 ( .A(n11506), .ZN(n17832) );
  CLKBUF_X2 U11141 ( .A(n13865), .Z(n10981) );
  NAND2_X1 U11142 ( .A1(n16350), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16349) );
  NAND2_X1 U11143 ( .A1(n20009), .A2(n13734), .ZN(n15527) );
  AOI21_X1 U11144 ( .B1(n13300), .B2(n15704), .A(n12931), .ZN(n15713) );
  OR2_X1 U11145 ( .A1(n21207), .A2(n20113), .ZN(n20101) );
  NOR2_X1 U11146 ( .A1(n20474), .A2(n20473), .ZN(n20486) );
  NOR2_X1 U11147 ( .A1(n20450), .A2(n20462), .ZN(n20460) );
  INV_X1 U11148 ( .A(n20596), .ZN(n20106) );
  NOR2_X1 U11149 ( .A1(n20723), .A2(n20717), .ZN(n20716) );
  INV_X1 U11150 ( .A(n21521), .ZN(n21560) );
  AOI211_X1 U11151 ( .C1(n20038), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20020), .B(n20019), .ZN(n20021) );
  BUF_X1 U11152 ( .A(n18180), .Z(n10978) );
  OAI21_X1 U11153 ( .B1(n17890), .B2(P3_STATE2_REG_0__SCAN_IN), .A(n21259), 
        .ZN(n18280) );
  AND2_X1 U11154 ( .A1(n13381), .A2(n14771), .ZN(n13519) );
  AND4_X1 U11155 ( .A1(n12031), .A2(n12032), .A3(n12033), .A4(n12030), .ZN(
        n10961) );
  AND2_X2 U11156 ( .A1(n12440), .A2(n11028), .ZN(n12457) );
  NAND2_X1 U11157 ( .A1(n12056), .A2(n12057), .ZN(n12058) );
  NOR2_X4 U11158 ( .A1(n17935), .A2(n11543), .ZN(n21138) );
  CLKBUF_X3 U11159 ( .A(n11004), .Z(n10962) );
  BUF_X4 U11160 ( .A(n11004), .Z(n10963) );
  AND2_X2 U11161 ( .A1(n11969), .A2(n17066), .ZN(n11004) );
  NOR3_X2 U11162 ( .A1(n20775), .A2(n20657), .A3(n20656), .ZN(n20764) );
  NAND2_X1 U11163 ( .A1(n11842), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12046) );
  AND2_X1 U11164 ( .A1(n14941), .A2(n14972), .ZN(n10964) );
  NAND2_X1 U11165 ( .A1(n15000), .A2(n18656), .ZN(n13256) );
  AND2_X4 U11166 ( .A1(n11970), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15792) );
  AOI211_X1 U11167 ( .C1(n21063), .C2(n21025), .A(n21024), .B(n21023), .ZN(
        n21027) );
  AND3_X2 U11168 ( .A1(n11893), .A2(n11892), .A3(n11891), .ZN(n11000) );
  NAND2_X2 U11169 ( .A1(n14723), .A2(n13578), .ZN(n13623) );
  NOR2_X2 U11170 ( .A1(n21237), .A2(n14562), .ZN(n20445) );
  INV_X1 U11171 ( .A(n20445), .ZN(n20450) );
  AND2_X1 U11172 ( .A1(n14978), .A2(n17066), .ZN(n10966) );
  AND2_X1 U11173 ( .A1(n14978), .A2(n17066), .ZN(n10967) );
  AND2_X1 U11174 ( .A1(n14978), .A2(n17066), .ZN(n15776) );
  INV_X2 U11175 ( .A(n12274), .ZN(n11899) );
  NAND2_X2 U11176 ( .A1(n13543), .A2(n13542), .ZN(n13580) );
  INV_X1 U11177 ( .A(n15777), .ZN(n10968) );
  NAND2_X1 U11178 ( .A1(n11970), .A2(n17066), .ZN(n15785) );
  NAND2_X1 U11179 ( .A1(n11780), .A2(n11779), .ZN(n10969) );
  NOR2_X1 U11180 ( .A1(n11430), .A2(n11429), .ZN(n11561) );
  BUF_X8 U11181 ( .A(n13433), .Z(n10974) );
  BUF_X8 U11182 ( .A(n13445), .Z(n10976) );
  NAND2_X2 U11183 ( .A1(n16622), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16596) );
  NOR2_X1 U11184 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11422), .ZN(
        n10977) );
  OR2_X1 U11185 ( .A1(n15715), .A2(n17411), .ZN(n11142) );
  NOR2_X1 U11186 ( .A1(n11374), .A2(n11373), .ZN(n11372) );
  NAND2_X1 U11187 ( .A1(n13758), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16080) );
  NAND2_X1 U11188 ( .A1(n13760), .A2(n16337), .ZN(n16107) );
  CLKBUF_X1 U11189 ( .A(n16623), .Z(n11001) );
  XNOR2_X1 U11190 ( .A(n12409), .B(n12395), .ZN(n15565) );
  OR2_X1 U11191 ( .A1(n15827), .A2(n14519), .ZN(n14527) );
  INV_X4 U11192 ( .A(n16337), .ZN(n16336) );
  AND2_X2 U11193 ( .A1(n14514), .A2(n15251), .ZN(n21521) );
  OR2_X1 U11194 ( .A1(n10988), .A2(n13671), .ZN(n10987) );
  INV_X4 U11195 ( .A(n13755), .ZN(n16337) );
  XNOR2_X1 U11196 ( .A(n13670), .B(n21311), .ZN(n19990) );
  NOR2_X1 U11198 ( .A1(n15862), .A2(n13961), .ZN(n15836) );
  INV_X1 U11199 ( .A(n20532), .ZN(n20582) );
  OR2_X1 U11200 ( .A1(n20101), .A2(n19087), .ZN(n14562) );
  INV_X1 U11201 ( .A(n21146), .ZN(n21187) );
  NAND2_X1 U11202 ( .A1(n14722), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14723) );
  NOR2_X2 U11203 ( .A1(n16331), .A2(n16330), .ZN(n16333) );
  OR2_X1 U11204 ( .A1(n16353), .A2(n15512), .ZN(n16331) );
  OR2_X1 U11205 ( .A1(n15384), .A2(n16351), .ZN(n16353) );
  NAND2_X1 U11206 ( .A1(n11017), .A2(n17168), .ZN(n21574) );
  AOI21_X2 U11207 ( .B1(n11662), .B2(n17881), .A(n11659), .ZN(n17125) );
  AND2_X1 U11208 ( .A1(n12905), .A2(n11871), .ZN(n11904) );
  AOI21_X1 U11209 ( .B1(n14720), .B2(n13864), .A(n11177), .ZN(n14864) );
  INV_X2 U11210 ( .A(n20622), .ZN(n20768) );
  CLKBUF_X2 U11211 ( .A(n12638), .Z(n12875) );
  BUF_X1 U11212 ( .A(n11804), .Z(n19376) );
  INV_X2 U11213 ( .A(n12046), .ZN(n13116) );
  BUF_X2 U11214 ( .A(n13450), .Z(n14477) );
  BUF_X2 U11215 ( .A(n13451), .Z(n11006) );
  BUF_X2 U11216 ( .A(n13443), .Z(n14478) );
  BUF_X2 U11217 ( .A(n13432), .Z(n14484) );
  CLKBUF_X2 U11218 ( .A(n13458), .Z(n14461) );
  CLKBUF_X2 U11219 ( .A(n11566), .Z(n17851) );
  CLKBUF_X3 U11220 ( .A(n11517), .Z(n17858) );
  CLKBUF_X1 U11221 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10990) );
  NAND2_X1 U11222 ( .A1(n16080), .A2(n13762), .ZN(n16045) );
  NAND2_X1 U11223 ( .A1(n11115), .A2(n11375), .ZN(n11374) );
  XNOR2_X1 U11224 ( .A(n11324), .B(n14504), .ZN(n15654) );
  AND2_X1 U11225 ( .A1(n16591), .A2(n12923), .ZN(n12931) );
  CLKBUF_X1 U11226 ( .A(n16113), .Z(n16114) );
  AND2_X2 U11227 ( .A1(n15933), .A2(n15936), .ZN(n15925) );
  NAND2_X1 U11228 ( .A1(n16106), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13759) );
  NOR2_X1 U11229 ( .A1(n16487), .A2(n13189), .ZN(n13231) );
  NAND2_X1 U11230 ( .A1(n16128), .A2(n16127), .ZN(n16129) );
  OR2_X1 U11231 ( .A1(n15599), .A2(n15600), .ZN(n15970) );
  NOR2_X1 U11232 ( .A1(n16489), .A2(n16488), .ZN(n16487) );
  NOR2_X1 U11233 ( .A1(n16522), .A2(n16509), .ZN(n16432) );
  NAND2_X1 U11234 ( .A1(n12179), .A2(n12178), .ZN(n15566) );
  XNOR2_X1 U11235 ( .A(n13188), .B(n11393), .ZN(n16489) );
  NOR2_X1 U11236 ( .A1(n15505), .A2(n13294), .ZN(n16520) );
  NAND2_X1 U11237 ( .A1(n15508), .A2(n14143), .ZN(n15586) );
  NOR2_X1 U11238 ( .A1(n12172), .A2(n12170), .ZN(n12171) );
  NOR2_X2 U11239 ( .A1(n15381), .A2(n14127), .ZN(n15457) );
  NAND2_X1 U11240 ( .A1(n11264), .A2(n12320), .ZN(n15503) );
  NOR2_X2 U11241 ( .A1(n15517), .A2(n15518), .ZN(n15519) );
  NOR2_X1 U11242 ( .A1(n18100), .A2(n21075), .ZN(n21051) );
  AND2_X1 U11243 ( .A1(n13747), .A2(n13744), .ZN(n11127) );
  AND2_X1 U11244 ( .A1(n13732), .A2(n13722), .ZN(n11381) );
  NAND2_X1 U11245 ( .A1(n15210), .A2(n18678), .ZN(n11352) );
  OAI21_X1 U11246 ( .B1(n12377), .B2(n11111), .A(n12380), .ZN(n11110) );
  AOI211_X1 U11247 ( .C1(n21551), .C2(P1_EBX_REG_29__SCAN_IN), .A(n15826), .B(
        n15825), .ZN(n15830) );
  AND2_X1 U11248 ( .A1(n11219), .A2(n11218), .ZN(n11559) );
  AOI211_X1 U11249 ( .C1(n20562), .C2(n20561), .A(n20574), .B(n20560), .ZN(
        n20566) );
  NAND2_X1 U11250 ( .A1(n13053), .A2(n11412), .ZN(n15517) );
  AND2_X1 U11251 ( .A1(n15367), .A2(n15450), .ZN(n13053) );
  AND2_X1 U11252 ( .A1(n15194), .A2(n15369), .ZN(n15367) );
  OR2_X1 U11253 ( .A1(n12184), .A2(n12183), .ZN(n12209) );
  NOR2_X1 U11254 ( .A1(n20557), .A2(n20556), .ZN(n20572) );
  XNOR2_X1 U11255 ( .A(n12184), .B(n12173), .ZN(n12393) );
  OR3_X1 U11256 ( .A1(n16162), .A2(n16158), .A3(n16321), .ZN(n16147) );
  NAND2_X1 U11257 ( .A1(n20724), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n20723) );
  NOR2_X2 U11258 ( .A1(n15193), .A2(n15195), .ZN(n15194) );
  NAND2_X2 U11259 ( .A1(n13737), .A2(n13736), .ZN(n13755) );
  XNOR2_X1 U11260 ( .A(n13737), .B(n13725), .ZN(n14020) );
  OR2_X2 U11261 ( .A1(n15078), .A2(n10992), .ZN(n15193) );
  AND2_X1 U11262 ( .A1(n12169), .A2(n12168), .ZN(n12173) );
  AOI22_X1 U11263 ( .A1(n21138), .A2(n18141), .B1(n18225), .B2(n18149), .ZN(
        n18180) );
  AND2_X1 U11264 ( .A1(n12132), .A2(n12131), .ZN(n12135) );
  NOR2_X1 U11265 ( .A1(n19225), .A2(n17097), .ZN(n19728) );
  NAND2_X1 U11266 ( .A1(n11240), .A2(n12966), .ZN(n14822) );
  NOR2_X1 U11267 ( .A1(n15197), .A2(n15198), .ZN(n15402) );
  OR2_X1 U11268 ( .A1(n12147), .A2(n12146), .ZN(n12169) );
  NAND2_X1 U11269 ( .A1(n13696), .A2(n13695), .ZN(n13713) );
  XNOR2_X1 U11270 ( .A(n14818), .B(n14817), .ZN(n19431) );
  NAND2_X1 U11271 ( .A1(n21506), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n21518) );
  AND2_X1 U11272 ( .A1(n15929), .A2(n15922), .ZN(n15920) );
  NOR2_X2 U11273 ( .A1(n21488), .A2(n21487), .ZN(n21506) );
  AND2_X1 U11274 ( .A1(n12965), .A2(n11241), .ZN(n14817) );
  AND2_X1 U11275 ( .A1(n12106), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11949) );
  NAND2_X1 U11276 ( .A1(n15879), .A2(n11095), .ZN(n21488) );
  NAND2_X1 U11277 ( .A1(n14828), .A2(n12963), .ZN(n14818) );
  BUF_X2 U11278 ( .A(n11962), .Z(n11009) );
  AND2_X1 U11279 ( .A1(n11964), .A2(n11957), .ZN(n15140) );
  AND2_X1 U11280 ( .A1(n11964), .A2(n11956), .ZN(n19288) );
  AND2_X1 U11281 ( .A1(n11960), .A2(n11963), .ZN(n19226) );
  AND2_X1 U11282 ( .A1(n11964), .A2(n11950), .ZN(n19273) );
  AND2_X1 U11283 ( .A1(n11964), .A2(n11963), .ZN(n19259) );
  AND2_X1 U11284 ( .A1(n11960), .A2(n11957), .ZN(n15231) );
  INV_X2 U11285 ( .A(n21050), .ZN(n21203) );
  OAI21_X1 U11286 ( .B1(n14926), .B2(n13550), .A(n13622), .ZN(n14871) );
  NAND2_X1 U11287 ( .A1(n14034), .A2(n14033), .ZN(n14780) );
  NOR2_X2 U11288 ( .A1(n11181), .A2(n13931), .ZN(n15951) );
  NAND2_X1 U11289 ( .A1(n20106), .A2(n21162), .ZN(n21050) );
  NAND2_X1 U11290 ( .A1(n15872), .A2(n11071), .ZN(n11181) );
  AND2_X1 U11291 ( .A1(n14809), .A2(n12959), .ZN(n14829) );
  NAND2_X1 U11292 ( .A1(n12949), .A2(n12948), .ZN(n12962) );
  OAI21_X1 U11293 ( .B1(n18205), .B2(n18204), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11694) );
  INV_X1 U11294 ( .A(n21007), .ZN(n21192) );
  NOR2_X2 U11295 ( .A1(n21187), .A2(n21204), .ZN(n21162) );
  NAND2_X1 U11296 ( .A1(n13588), .A2(n13587), .ZN(n14025) );
  XNOR2_X1 U11297 ( .A(n14842), .B(n12957), .ZN(n14804) );
  OR2_X1 U11298 ( .A1(n14681), .A2(n18393), .ZN(n11961) );
  NAND2_X2 U11299 ( .A1(n16039), .A2(n14884), .ZN(n16033) );
  NAND2_X1 U11300 ( .A1(n13641), .A2(n13640), .ZN(n14927) );
  OAI21_X1 U11301 ( .B1(n20599), .B2(n20598), .A(n20597), .ZN(n20621) );
  AND2_X1 U11302 ( .A1(n13591), .A2(n13617), .ZN(n11128) );
  OAI21_X1 U11303 ( .B1(n12950), .B2(n15129), .A(n12952), .ZN(n14842) );
  NAND2_X1 U11304 ( .A1(n11945), .A2(n11942), .ZN(n12950) );
  CLKBUF_X1 U11305 ( .A(n21718), .Z(n21722) );
  AND2_X1 U11306 ( .A1(n11914), .A2(n11118), .ZN(n11937) );
  XNOR2_X1 U11307 ( .A(n12261), .B(n12260), .ZN(n12259) );
  NAND2_X1 U11308 ( .A1(n11941), .A2(n11940), .ZN(n11942) );
  NOR2_X2 U11309 ( .A1(n19374), .A2(n19700), .ZN(n19375) );
  NAND2_X1 U11310 ( .A1(n11923), .A2(n11922), .ZN(n11926) );
  NAND2_X1 U11311 ( .A1(n11317), .A2(n13602), .ZN(n14748) );
  OR2_X1 U11312 ( .A1(n11317), .A2(n13602), .ZN(n11316) );
  NAND2_X1 U11313 ( .A1(n11117), .A2(n11903), .ZN(n11941) );
  NAND2_X2 U11314 ( .A1(n19989), .A2(n14882), .ZN(n15965) );
  NOR2_X2 U11315 ( .A1(n19218), .A2(n19700), .ZN(n15143) );
  OR2_X1 U11316 ( .A1(n12402), .A2(n11158), .ZN(n12412) );
  NAND2_X1 U11317 ( .A1(n21665), .A2(n14627), .ZN(n21262) );
  AOI221_X1 U11318 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17136), .C1(n17135), .C2(
        n17136), .A(n19362), .ZN(n17435) );
  INV_X2 U11319 ( .A(n20115), .ZN(n20166) );
  NAND2_X1 U11320 ( .A1(n13885), .A2(n13884), .ZN(n19975) );
  NAND2_X1 U11321 ( .A1(n13843), .A2(n11068), .ZN(n21665) );
  NAND2_X1 U11322 ( .A1(n13629), .A2(n13628), .ZN(n21784) );
  CLKBUF_X1 U11323 ( .A(n14037), .Z(n21772) );
  NOR2_X1 U11324 ( .A1(n18109), .A2(n20549), .ZN(n18108) );
  AND2_X1 U11325 ( .A1(n11202), .A2(n11051), .ZN(n18235) );
  AND2_X1 U11326 ( .A1(n13556), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13593) );
  INV_X1 U11327 ( .A(n15068), .ZN(n11188) );
  NAND3_X1 U11328 ( .A1(n13498), .A2(n13555), .A3(n13497), .ZN(n11126) );
  NAND2_X1 U11329 ( .A1(n12629), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11902) );
  NAND2_X1 U11330 ( .A1(n12628), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11887) );
  NOR2_X1 U11331 ( .A1(n11715), .A2(n11664), .ZN(n11636) );
  NOR2_X1 U11332 ( .A1(n18264), .A2(n18263), .ZN(n18262) );
  NAND2_X1 U11333 ( .A1(n11868), .A2(n11395), .ZN(n18657) );
  NAND2_X1 U11334 ( .A1(n11402), .A2(n12606), .ZN(n12899) );
  NAND2_X1 U11335 ( .A1(n13866), .A2(n13867), .ZN(n11177) );
  NAND2_X1 U11336 ( .A1(n11874), .A2(n11825), .ZN(n12892) );
  INV_X1 U11337 ( .A(n11881), .ZN(n15031) );
  AND3_X1 U11338 ( .A1(n11175), .A2(n11174), .A3(n11173), .ZN(n13808) );
  AND2_X1 U11339 ( .A1(n20788), .A2(n11132), .ZN(n11715) );
  NOR2_X1 U11340 ( .A1(n20651), .A2(n11680), .ZN(n11676) );
  INV_X1 U11341 ( .A(n15000), .ZN(n15291) );
  AND2_X1 U11342 ( .A1(n11395), .A2(n12627), .ZN(n11343) );
  NAND2_X1 U11343 ( .A1(n13603), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13806) );
  INV_X1 U11344 ( .A(n11869), .ZN(n12627) );
  AND2_X1 U11345 ( .A1(n12023), .A2(n12022), .ZN(n12663) );
  INV_X1 U11346 ( .A(n11804), .ZN(n14840) );
  INV_X1 U11347 ( .A(n12894), .ZN(n11867) );
  NAND2_X1 U11348 ( .A1(n11792), .A2(n11791), .ZN(n11804) );
  NAND2_X2 U11349 ( .A1(n11246), .A2(n11244), .ZN(n12635) );
  INV_X1 U11350 ( .A(n12901), .ZN(n11880) );
  OAI21_X1 U11351 ( .B1(n11813), .B2(n11245), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11244) );
  OAI21_X1 U11352 ( .B1(n11248), .B2(n11247), .A(n11832), .ZN(n11246) );
  INV_X2 U11353 ( .A(U214), .ZN(n20090) );
  NAND2_X2 U11354 ( .A1(U214), .A2(n20049), .ZN(n20098) );
  AND4_X1 U11355 ( .A1(n11056), .A2(n11027), .A3(n11163), .A4(n13455), .ZN(
        n13500) );
  NAND2_X2 U11356 ( .A1(n13391), .A2(n13390), .ZN(n13484) );
  AND4_X1 U11357 ( .A1(n13395), .A2(n13394), .A3(n13393), .A4(n13392), .ZN(
        n13401) );
  AND4_X1 U11358 ( .A1(n13399), .A2(n13398), .A3(n13397), .A4(n13396), .ZN(
        n13400) );
  AND4_X1 U11359 ( .A1(n13385), .A2(n13384), .A3(n13383), .A4(n13382), .ZN(
        n13391) );
  NOR2_X1 U11360 ( .A1(n18181), .A2(n11289), .ZN(n17930) );
  CLKBUF_X1 U11361 ( .A(n18532), .Z(n18500) );
  INV_X2 U11362 ( .A(n18358), .ZN(n18365) );
  NOR2_X2 U11363 ( .A1(n18808), .A2(n18821), .ZN(n19168) );
  INV_X2 U11364 ( .A(n19080), .ZN(U215) );
  BUF_X2 U11366 ( .A(n11566), .Z(n17791) );
  NOR2_X1 U11367 ( .A1(n17394), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18532) );
  INV_X2 U11368 ( .A(n13238), .ZN(n15793) );
  OR2_X2 U11369 ( .A1(n22328), .A2(n17192), .ZN(n17151) );
  INV_X1 U11370 ( .A(n20810), .ZN(n11422) );
  INV_X2 U11371 ( .A(n19820), .ZN(n19878) );
  AND2_X1 U11373 ( .A1(n14771), .A2(n13381), .ZN(n11417) );
  AND2_X2 U11374 ( .A1(n14771), .A2(n14762), .ZN(n14419) );
  OR2_X2 U11375 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17884), .ZN(n11764) );
  NAND2_X1 U11376 ( .A1(n20813), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11429) );
  AND2_X1 U11377 ( .A1(n11768), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14978) );
  NOR2_X1 U11378 ( .A1(n11768), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11969) );
  CLKBUF_X1 U11379 ( .A(n21868), .Z(n21896) );
  AND2_X1 U11380 ( .A1(n14776), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13375) );
  AND2_X2 U11381 ( .A1(n13370), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14771) );
  NAND3_X1 U11382 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20822) );
  NAND2_X1 U11383 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15640) );
  AND2_X2 U11384 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14939) );
  NOR2_X1 U11385 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13083) );
  NAND2_X1 U11386 ( .A1(n19991), .A2(n13671), .ZN(n19996) );
  NAND2_X1 U11387 ( .A1(n15031), .A2(n14717), .ZN(n11889) );
  NAND2_X1 U11388 ( .A1(n19703), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18377) );
  NOR2_X2 U11389 ( .A1(n18034), .A2(n18026), .ZN(n18063) );
  AND4_X2 U11390 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n11046) );
  NAND2_X1 U11393 ( .A1(n15457), .A2(n15509), .ZN(n15508) );
  CLKBUF_X1 U11394 ( .A(n11333), .Z(n10985) );
  NAND2_X2 U11395 ( .A1(n14840), .A2(n10969), .ZN(n11886) );
  NAND2_X1 U11396 ( .A1(n19990), .A2(n10989), .ZN(n10986) );
  AND2_X2 U11397 ( .A1(n10986), .A2(n10987), .ZN(n19997) );
  INV_X1 U11398 ( .A(n19998), .ZN(n10988) );
  AND2_X1 U11399 ( .A1(n19992), .A2(n19998), .ZN(n10989) );
  NAND2_X1 U11400 ( .A1(n11352), .A2(n12095), .ZN(n10991) );
  NAND2_X1 U11401 ( .A1(n11352), .A2(n12095), .ZN(n12137) );
  OR2_X1 U11402 ( .A1(n16684), .A2(n11403), .ZN(n15716) );
  OR2_X1 U11403 ( .A1(n12974), .A2(n11030), .ZN(n10992) );
  NOR2_X1 U11404 ( .A1(n16489), .A2(n16488), .ZN(n10993) );
  NOR2_X1 U11405 ( .A1(n13231), .A2(n13230), .ZN(n10994) );
  NOR2_X1 U11406 ( .A1(n13231), .A2(n13230), .ZN(n16474) );
  INV_X2 U11407 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13551) );
  NOR2_X2 U11408 ( .A1(n13292), .A2(n16847), .ZN(n16622) );
  INV_X1 U11409 ( .A(n13494), .ZN(n13502) );
  NAND2_X2 U11410 ( .A1(n16774), .A2(n12211), .ZN(n16764) );
  AND4_X2 U11411 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n12026), .ZN(
        n11045) );
  OAI21_X1 U11412 ( .B1(n15519), .B2(n11257), .A(n11085), .ZN(n11260) );
  NAND3_X2 U11413 ( .A1(n13380), .A2(n11418), .A3(n13379), .ZN(n13476) );
  AND2_X2 U11415 ( .A1(n14708), .A2(n13500), .ZN(n13506) );
  NOR2_X2 U11416 ( .A1(n13473), .A2(n13504), .ZN(n14708) );
  AND2_X4 U11417 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14762) );
  NAND2_X2 U11418 ( .A1(n15161), .A2(n12068), .ZN(n12092) );
  XNOR2_X2 U11419 ( .A(n12092), .B(n12093), .ZN(n15210) );
  NAND2_X1 U11420 ( .A1(n11879), .A2(n14717), .ZN(n11908) );
  NAND2_X2 U11421 ( .A1(n11243), .A2(n11242), .ZN(n12894) );
  INV_X2 U11422 ( .A(n11635), .ZN(n20652) );
  OR2_X2 U11423 ( .A1(n11428), .A2(n15640), .ZN(n11093) );
  NAND2_X1 U11424 ( .A1(n11421), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11428) );
  NOR2_X2 U11425 ( .A1(n20763), .A2(n20749), .ZN(n20748) );
  NAND2_X1 U11426 ( .A1(n15527), .A2(n13743), .ZN(n10995) );
  INV_X1 U11427 ( .A(n14755), .ZN(n10996) );
  BUF_X1 U11428 ( .A(n13495), .Z(n10997) );
  AND2_X2 U11429 ( .A1(n12882), .A2(n12895), .ZN(n12629) );
  NOR2_X2 U11430 ( .A1(n16676), .A2(n16649), .ZN(n16665) );
  NAND2_X2 U11431 ( .A1(n14025), .A2(n11128), .ZN(n13643) );
  NAND2_X1 U11432 ( .A1(n10995), .A2(n11382), .ZN(n10998) );
  NAND2_X1 U11433 ( .A1(n19997), .A2(n11054), .ZN(n10999) );
  NAND2_X1 U11434 ( .A1(n11384), .A2(n11382), .ZN(n15552) );
  NAND2_X1 U11435 ( .A1(n19997), .A2(n11054), .ZN(n20002) );
  AND3_X1 U11437 ( .A1(n11346), .A2(n11143), .A3(n11344), .ZN(n11003) );
  INV_X1 U11438 ( .A(n10962), .ZN(n11793) );
  OAI21_X2 U11439 ( .B1(n15264), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13571), 
        .ZN(n13590) );
  NAND2_X1 U11440 ( .A1(n14732), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11005) );
  NAND2_X1 U11441 ( .A1(n11944), .A2(n11914), .ZN(n11936) );
  AND2_X1 U11442 ( .A1(n11381), .A2(n10999), .ZN(n11007) );
  NAND2_X1 U11443 ( .A1(n19990), .A2(n19992), .ZN(n19991) );
  NAND2_X2 U11444 ( .A1(n11343), .A2(n11868), .ZN(n12599) );
  XNOR2_X2 U11445 ( .A(n11924), .B(n11926), .ZN(n11935) );
  NAND2_X4 U11446 ( .A1(n13596), .A2(n21752), .ZN(n15264) );
  NAND2_X2 U11447 ( .A1(n13642), .A2(n14927), .ZN(n13672) );
  XNOR2_X1 U11448 ( .A(n13651), .B(n21317), .ZN(n15090) );
  AND2_X4 U11449 ( .A1(n14978), .A2(n17066), .ZN(n11008) );
  NAND2_X2 U11450 ( .A1(n15092), .A2(n13652), .ZN(n13670) );
  XNOR2_X1 U11451 ( .A(n14733), .B(n13576), .ZN(n14722) );
  OAI21_X2 U11452 ( .B1(n14035), .B2(n13550), .A(n13549), .ZN(n14732) );
  INV_X2 U11453 ( .A(n12641), .ZN(n12633) );
  AND2_X1 U11454 ( .A1(n16732), .A2(n16730), .ZN(n16715) );
  OR2_X1 U11455 ( .A1(n16732), .A2(n13277), .ZN(n11335) );
  NAND2_X1 U11456 ( .A1(n14732), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14733) );
  XNOR2_X1 U11458 ( .A(n13623), .B(n21301), .ZN(n14870) );
  XNOR2_X2 U11459 ( .A(n13353), .B(n13351), .ZN(n16578) );
  NAND2_X2 U11460 ( .A1(n16590), .A2(n13350), .ZN(n13353) );
  XOR2_X2 U11461 ( .A(n15730), .B(n15729), .Z(n16055) );
  OAI21_X2 U11462 ( .B1(n11129), .B2(n13617), .A(n13643), .ZN(n14926) );
  AND2_X1 U11463 ( .A1(n13375), .A2(n11176), .ZN(n13431) );
  AND2_X1 U11464 ( .A1(n13375), .A2(n13381), .ZN(n13458) );
  AND3_X2 U11465 ( .A1(n13854), .A2(n11378), .A3(n13856), .ZN(n13555) );
  OAI21_X2 U11466 ( .B1(n16623), .B2(n16625), .A(n16624), .ZN(n16611) );
  NOR2_X2 U11467 ( .A1(n11009), .A2(n11961), .ZN(n12097) );
  NOR2_X2 U11468 ( .A1(n15100), .A2(n15124), .ZN(n15123) );
  AND3_X2 U11469 ( .A1(n13415), .A2(n13416), .A3(n13417), .ZN(n11049) );
  NAND3_X4 U11470 ( .A1(n13419), .A2(n13418), .A3(n11049), .ZN(n13473) );
  NAND2_X2 U11471 ( .A1(n15552), .A2(n11127), .ZN(n16135) );
  XOR2_X2 U11472 ( .A(n16342), .B(n16341), .Z(n20018) );
  OAI21_X2 U11473 ( .B1(n16135), .B2(n11391), .A(n11021), .ZN(n16128) );
  INV_X1 U11474 ( .A(n13238), .ZN(n11010) );
  INV_X1 U11475 ( .A(n11842), .ZN(n11011) );
  OR2_X1 U11476 ( .A1(n13590), .A2(n13589), .ZN(n13591) );
  AND2_X1 U11477 ( .A1(n14819), .A2(n11943), .ZN(n11964) );
  AND2_X1 U11478 ( .A1(n15331), .A2(n14819), .ZN(n11960) );
  OR2_X1 U11479 ( .A1(n14819), .A2(n11943), .ZN(n11330) );
  OR2_X1 U11480 ( .A1(n15331), .A2(n14819), .ZN(n11962) );
  AND2_X2 U11481 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14764) );
  XOR2_X1 U11482 ( .A(n20583), .B(n14559), .Z(n11012) );
  XOR2_X1 U11483 ( .A(n20583), .B(n14559), .Z(n11013) );
  XOR2_X2 U11484 ( .A(n20583), .B(n14559), .Z(n20523) );
  AND2_X2 U11485 ( .A1(n15831), .A2(n11322), .ZN(n15729) );
  NOR2_X4 U11486 ( .A1(n15844), .A2(n15846), .ZN(n15831) );
  AND2_X2 U11487 ( .A1(n21935), .A2(n13860), .ZN(n13547) );
  INV_X4 U11488 ( .A(n13500), .ZN(n13860) );
  AND2_X2 U11489 ( .A1(n11969), .A2(n13083), .ZN(n12077) );
  AND2_X1 U11490 ( .A1(n11379), .A2(n13857), .ZN(n11378) );
  NAND2_X1 U11491 ( .A1(n13845), .A2(n11052), .ZN(n11379) );
  OAI21_X1 U11492 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14776), .A(
        n13779), .ZN(n13783) );
  OAI21_X1 U11493 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13778), .A(
        n13782), .ZN(n13779) );
  NAND2_X1 U11494 ( .A1(n11003), .A2(n12135), .ZN(n12184) );
  AND2_X1 U11495 ( .A1(n17985), .A2(n21105), .ZN(n11213) );
  OR2_X1 U11496 ( .A1(n12637), .A2(n12539), .ZN(n12826) );
  NAND2_X1 U11497 ( .A1(n18997), .A2(n19087), .ZN(n11132) );
  NAND2_X1 U11498 ( .A1(n11092), .A2(n11238), .ZN(n12878) );
  INV_X1 U11499 ( .A(n12637), .ZN(n11238) );
  XNOR2_X1 U11500 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12230) );
  NAND2_X1 U11501 ( .A1(n12227), .A2(n12226), .ZN(n12231) );
  AOI21_X1 U11502 ( .B1(n13492), .B2(n13547), .A(n11044), .ZN(n13508) );
  OAI22_X1 U11503 ( .A1(n14027), .A2(n13686), .B1(n13806), .B2(n13685), .ZN(
        n13695) );
  NAND2_X1 U11504 ( .A1(n13860), .A2(n13475), .ZN(n13603) );
  AND2_X1 U11505 ( .A1(n12251), .A2(n12600), .ZN(n11875) );
  AND2_X1 U11506 ( .A1(n14840), .A2(n12941), .ZN(n13208) );
  NAND2_X1 U11507 ( .A1(n13784), .A2(n11408), .ZN(n13823) );
  OAI21_X1 U11508 ( .B1(n16102), .B2(n16058), .A(n16337), .ZN(n13762) );
  OR2_X1 U11509 ( .A1(n13540), .A2(n13539), .ZN(n13572) );
  AOI21_X1 U11510 ( .B1(n13474), .B2(n13470), .A(n13429), .ZN(n13480) );
  INV_X1 U11511 ( .A(n13032), .ZN(n13113) );
  INV_X1 U11512 ( .A(n13033), .ZN(n13114) );
  INV_X1 U11513 ( .A(n13030), .ZN(n13115) );
  OR2_X1 U11514 ( .A1(n13082), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13026) );
  NAND2_X1 U11515 ( .A1(n16496), .A2(n11394), .ZN(n13188) );
  OR2_X1 U11516 ( .A1(n13170), .A2(n11260), .ZN(n11394) );
  NAND2_X1 U11517 ( .A1(n11890), .A2(n12641), .ZN(n12282) );
  AND2_X1 U11518 ( .A1(n18544), .A2(n12689), .ZN(n13286) );
  AND2_X1 U11519 ( .A1(n12849), .A2(n12848), .ZN(n15198) );
  INV_X1 U11520 ( .A(n12209), .ZN(n12208) );
  INV_X1 U11521 ( .A(n11916), .ZN(n12346) );
  AND2_X1 U11522 ( .A1(n12024), .A2(n12055), .ZN(n11345) );
  NOR2_X1 U11523 ( .A1(n13149), .A2(n13172), .ZN(n12942) );
  AND2_X1 U11524 ( .A1(n18711), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12956) );
  NOR3_X1 U11525 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n11430), .ZN(n11566) );
  INV_X1 U11526 ( .A(n11557), .ZN(n11214) );
  NAND2_X1 U11527 ( .A1(n11213), .A2(n11555), .ZN(n11216) );
  AOI21_X1 U11528 ( .B1(n17914), .B2(n11546), .A(n18189), .ZN(n11554) );
  NOR2_X1 U11529 ( .A1(n17949), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17914) );
  AND2_X1 U11530 ( .A1(n11131), .A2(n11130), .ZN(n21221) );
  NAND2_X1 U11531 ( .A1(n21234), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11130) );
  NAND2_X1 U11532 ( .A1(n21218), .A2(n21217), .ZN(n11131) );
  NAND2_X1 U11533 ( .A1(n14514), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15248) );
  INV_X1 U11534 ( .A(n21592), .ZN(n14880) );
  AND2_X1 U11535 ( .A1(n21917), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14501) );
  AND2_X1 U11536 ( .A1(n14272), .A2(n14271), .ZN(n15956) );
  INV_X1 U11537 ( .A(n15239), .ZN(n11220) );
  NOR2_X2 U11538 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12246), .ZN(
        n13118) );
  AND2_X1 U11539 ( .A1(n12853), .A2(n12852), .ZN(n15494) );
  AND2_X1 U11540 ( .A1(n15403), .A2(n11405), .ZN(n11228) );
  NOR2_X1 U11541 ( .A1(n11237), .A2(n15308), .ZN(n11236) );
  NAND2_X1 U11542 ( .A1(n16957), .A2(n15427), .ZN(n11237) );
  XNOR2_X1 U11543 ( .A(n15279), .B(n15278), .ZN(n15761) );
  OR2_X1 U11544 ( .A1(n15277), .A2(n15276), .ZN(n15279) );
  NAND2_X1 U11545 ( .A1(n12532), .A2(n12531), .ZN(n13310) );
  AND2_X1 U11546 ( .A1(n12530), .A2(n13350), .ZN(n12531) );
  NAND2_X1 U11547 ( .A1(n14804), .A2(n14805), .ZN(n14809) );
  NAND2_X1 U11548 ( .A1(n11666), .A2(n11661), .ZN(n20114) );
  NOR2_X1 U11549 ( .A1(n18269), .A2(n11521), .ZN(n18264) );
  INV_X1 U11550 ( .A(n20788), .ZN(n11708) );
  INV_X1 U11551 ( .A(n21519), .ZN(n21572) );
  OR2_X1 U11552 ( .A1(n15022), .A2(n18718), .ZN(n18721) );
  NAND2_X1 U11553 ( .A1(n12874), .A2(n12873), .ZN(n12881) );
  AOI22_X1 U11554 ( .A1(n13458), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13373) );
  AOI22_X1 U11555 ( .A1(n13431), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13604), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13371) );
  AOI22_X1 U11556 ( .A1(n13432), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13450), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13374) );
  AOI22_X1 U11557 ( .A1(n13443), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13378) );
  INV_X1 U11558 ( .A(n13118), .ZN(n12191) );
  AOI21_X1 U11559 ( .B1(n21763), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13777), .ZN(n13788) );
  AOI21_X1 U11560 ( .B1(n13502), .B2(n21737), .A(n10997), .ZN(n13497) );
  AOI22_X1 U11561 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13451), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13388) );
  AOI22_X1 U11562 ( .A1(n13443), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13387) );
  NAND2_X1 U11563 ( .A1(n12403), .A2(n11159), .ZN(n11158) );
  INV_X1 U11564 ( .A(n12406), .ZN(n11159) );
  INV_X1 U11565 ( .A(n12173), .ZN(n12183) );
  AND2_X1 U11566 ( .A1(n11345), .A2(n12233), .ZN(n11344) );
  NAND2_X1 U11567 ( .A1(n11873), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11140) );
  INV_X1 U11568 ( .A(n12895), .ZN(n11897) );
  NAND2_X1 U11569 ( .A1(n11937), .A2(n11942), .ZN(n11944) );
  INV_X1 U11570 ( .A(n11837), .ZN(n11838) );
  INV_X1 U11571 ( .A(n13490), .ZN(n14152) );
  NOR2_X1 U11572 ( .A1(n13484), .A2(n13475), .ZN(n14707) );
  AND2_X1 U11573 ( .A1(n11066), .A2(n15856), .ZN(n11326) );
  INV_X1 U11574 ( .A(n15204), .ZN(n14083) );
  INV_X1 U11575 ( .A(n17185), .ZN(n14497) );
  NAND2_X1 U11576 ( .A1(n13754), .A2(n11094), .ZN(n13760) );
  AND2_X1 U11577 ( .A1(n15873), .A2(n11180), .ZN(n11179) );
  INV_X1 U11578 ( .A(n15960), .ZN(n11180) );
  AND2_X1 U11579 ( .A1(n16293), .A2(n11390), .ZN(n11021) );
  NAND2_X1 U11580 ( .A1(n16337), .A2(n11097), .ZN(n11390) );
  NOR2_X1 U11581 ( .A1(n16337), .A2(n16287), .ZN(n11391) );
  INV_X1 U11582 ( .A(n13712), .ZN(n13710) );
  INV_X1 U11583 ( .A(n13713), .ZN(n13711) );
  AOI21_X1 U11584 ( .B1(n15530), .B2(n13743), .A(n11383), .ZN(n11382) );
  INV_X1 U11585 ( .A(n15553), .ZN(n11383) );
  XNOR2_X1 U11586 ( .A(n13672), .B(n13673), .ZN(n14065) );
  NOR2_X1 U11587 ( .A1(n15069), .A2(n17193), .ZN(n11187) );
  NOR2_X2 U11588 ( .A1(n10981), .A2(n14721), .ZN(n13957) );
  OR2_X1 U11589 ( .A1(n13528), .A2(n13527), .ZN(n13739) );
  INV_X1 U11590 ( .A(n13806), .ZN(n13794) );
  AND2_X1 U11591 ( .A1(n13968), .A2(n13475), .ZN(n13471) );
  INV_X1 U11592 ( .A(n21759), .ZN(n21751) );
  INV_X1 U11593 ( .A(n14926), .ZN(n21820) );
  OR2_X1 U11594 ( .A1(n21872), .A2(n21871), .ZN(n21915) );
  INV_X1 U11595 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21763) );
  NOR2_X1 U11596 ( .A1(n12506), .A2(n12505), .ZN(n11153) );
  NAND2_X1 U11597 ( .A1(n11162), .A2(n12445), .ZN(n11161) );
  INV_X1 U11598 ( .A(n12449), .ZN(n11162) );
  NAND2_X1 U11599 ( .A1(n12358), .A2(n12357), .ZN(n12652) );
  NAND2_X1 U11600 ( .A1(n11842), .A2(n11832), .ZN(n13033) );
  NAND2_X1 U11601 ( .A1(n11977), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13032) );
  NAND2_X1 U11602 ( .A1(n15791), .A2(n11832), .ZN(n13030) );
  NAND2_X1 U11603 ( .A1(n12633), .A2(n12654), .ZN(n12637) );
  OAI211_X1 U11604 ( .C1(n16474), .C2(n16484), .A(n13251), .B(n16481), .ZN(
        n13249) );
  AND2_X1 U11605 ( .A1(n13128), .A2(n13127), .ZN(n13146) );
  AND2_X1 U11606 ( .A1(n11258), .A2(n11255), .ZN(n11254) );
  NAND2_X1 U11607 ( .A1(n11256), .A2(n11261), .ZN(n11255) );
  INV_X1 U11608 ( .A(n16504), .ZN(n11258) );
  INV_X1 U11609 ( .A(n16508), .ZN(n11256) );
  INV_X1 U11610 ( .A(n13208), .ZN(n13149) );
  NOR2_X1 U11611 ( .A1(n16447), .A2(n11299), .ZN(n11298) );
  NOR2_X1 U11612 ( .A1(n16768), .A2(n11307), .ZN(n11306) );
  INV_X1 U11613 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11307) );
  INV_X1 U11614 ( .A(n15281), .ZN(n11305) );
  INV_X1 U11615 ( .A(n15209), .ZN(n11111) );
  OR2_X1 U11616 ( .A1(n18595), .A2(n12535), .ZN(n12526) );
  NAND2_X1 U11617 ( .A1(n12290), .A2(n11269), .ZN(n11268) );
  INV_X1 U11618 ( .A(n15059), .ZN(n11269) );
  INV_X2 U11619 ( .A(n10980), .ZN(n12349) );
  NAND2_X1 U11620 ( .A1(n11124), .A2(n15343), .ZN(n12376) );
  NAND2_X1 U11621 ( .A1(n11879), .A2(n11137), .ZN(n11138) );
  NAND2_X1 U11622 ( .A1(n11873), .A2(n11136), .ZN(n11135) );
  NAND2_X1 U11623 ( .A1(n10980), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U11624 ( .A1(n13208), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12957) );
  NAND2_X1 U11625 ( .A1(n13208), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12960) );
  NAND2_X1 U11626 ( .A1(n11798), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11243) );
  NAND2_X1 U11627 ( .A1(n11803), .A2(n11832), .ZN(n11242) );
  NAND2_X1 U11628 ( .A1(n12238), .A2(n12237), .ZN(n12594) );
  NOR2_X1 U11629 ( .A1(n20517), .A2(n11287), .ZN(n11286) );
  INV_X1 U11630 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11287) );
  NOR2_X1 U11631 ( .A1(n20768), .A2(n18957), .ZN(n11707) );
  AOI21_X1 U11632 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17124), .A(
        n11722), .ZN(n11728) );
  NOR2_X1 U11633 ( .A1(n11541), .A2(n11544), .ZN(n11205) );
  AND2_X1 U11634 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11536), .ZN(
        n11537) );
  NOR2_X1 U11635 ( .A1(n18233), .A2(n11530), .ZN(n11533) );
  NAND2_X1 U11636 ( .A1(n11676), .A2(n20780), .ZN(n11365) );
  AOI22_X1 U11637 ( .A1(n11638), .A2(n11637), .B1(n11636), .B2(n11706), .ZN(
        n11657) );
  NOR2_X1 U11638 ( .A1(n20595), .A2(n20768), .ZN(n11660) );
  AND2_X1 U11639 ( .A1(n14738), .A2(n13830), .ZN(n14659) );
  NAND2_X1 U11640 ( .A1(n14522), .A2(n13860), .ZN(n11168) );
  OR2_X1 U11641 ( .A1(n15248), .A2(n11168), .ZN(n21403) );
  AND2_X1 U11642 ( .A1(n14696), .A2(n14695), .ZN(n19882) );
  AND2_X1 U11643 ( .A1(n11065), .A2(n15956), .ZN(n11319) );
  AND2_X1 U11644 ( .A1(n11318), .A2(n11065), .ZN(n15957) );
  AND2_X1 U11645 ( .A1(n16157), .A2(n16159), .ZN(n16293) );
  AND2_X1 U11646 ( .A1(n14096), .A2(n14095), .ZN(n15348) );
  NAND2_X1 U11647 ( .A1(n14074), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14097) );
  NAND2_X1 U11648 ( .A1(n14068), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14075) );
  NAND2_X1 U11649 ( .A1(n14926), .A2(n14024), .ZN(n11311) );
  NAND2_X1 U11650 ( .A1(n11386), .A2(n11070), .ZN(n13767) );
  INV_X1 U11651 ( .A(n14006), .ZN(n11387) );
  NAND2_X1 U11652 ( .A1(n15929), .A2(n11084), .ZN(n15862) );
  INV_X1 U11653 ( .A(n15860), .ZN(n11189) );
  NAND2_X1 U11654 ( .A1(n15872), .A2(n11179), .ZN(n15963) );
  AND2_X1 U11655 ( .A1(n11193), .A2(n11192), .ZN(n11191) );
  INV_X1 U11656 ( .A(n15973), .ZN(n11192) );
  NOR2_X1 U11657 ( .A1(n11022), .A2(n11183), .ZN(n11182) );
  INV_X1 U11658 ( .A(n19975), .ZN(n11184) );
  INV_X1 U11659 ( .A(n15385), .ZN(n11183) );
  NOR2_X1 U11660 ( .A1(n19975), .A2(n11022), .ZN(n15386) );
  NOR2_X1 U11661 ( .A1(n19975), .A2(n15206), .ZN(n15376) );
  INV_X1 U11662 ( .A(n13864), .ZN(n14721) );
  INV_X1 U11663 ( .A(n13814), .ZN(n14027) );
  INV_X1 U11664 ( .A(n14028), .ZN(n13587) );
  OR2_X1 U11665 ( .A1(n13825), .A2(n13806), .ZN(n13820) );
  OAI21_X1 U11666 ( .B1(n13825), .B2(n13818), .A(n13817), .ZN(n13819) );
  NAND2_X1 U11667 ( .A1(n21821), .A2(n14926), .ZN(n21781) );
  NAND2_X1 U11668 ( .A1(n21820), .A2(n14928), .ZN(n21810) );
  AND2_X1 U11669 ( .A1(n21759), .A2(n21750), .ZN(n21852) );
  INV_X1 U11670 ( .A(n21859), .ZN(n21853) );
  NOR2_X1 U11671 ( .A1(n21843), .A2(n22212), .ZN(n21907) );
  NAND2_X1 U11672 ( .A1(n21759), .A2(n14035), .ZN(n21894) );
  NAND2_X1 U11673 ( .A1(n21820), .A2(n14927), .ZN(n21895) );
  NAND2_X1 U11674 ( .A1(n17186), .A2(n21735), .ZN(n22212) );
  AND2_X1 U11675 ( .A1(n15006), .A2(n15004), .ZN(n15017) );
  CLKBUF_X1 U11676 ( .A(n15429), .Z(n18606) );
  NOR2_X1 U11677 ( .A1(n15189), .A2(n11251), .ZN(n11250) );
  INV_X1 U11678 ( .A(n15148), .ZN(n11251) );
  NAND2_X1 U11679 ( .A1(n13360), .A2(n13260), .ZN(n15703) );
  INV_X1 U11680 ( .A(n13170), .ZN(n11259) );
  NAND2_X1 U11681 ( .A1(n16515), .A2(n16508), .ZN(n11253) );
  NAND2_X1 U11682 ( .A1(n14817), .A2(n14818), .ZN(n11240) );
  AND2_X1 U11683 ( .A1(n13256), .A2(n18716), .ZN(n15015) );
  AND2_X1 U11684 ( .A1(n15019), .A2(n12895), .ZN(n12889) );
  AND2_X1 U11685 ( .A1(n14569), .A2(n14568), .ZN(n15298) );
  AND2_X1 U11686 ( .A1(n11033), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11302) );
  NOR2_X1 U11687 ( .A1(n16410), .A2(n16605), .ZN(n16411) );
  OR2_X1 U11688 ( .A1(n16408), .A2(n16407), .ZN(n16410) );
  AND2_X1 U11689 ( .A1(n12256), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16403) );
  NOR2_X1 U11690 ( .A1(n15474), .A2(n15473), .ZN(n15475) );
  NOR2_X1 U11691 ( .A1(n15286), .A2(n17418), .ZN(n15287) );
  NAND2_X1 U11692 ( .A1(n11353), .A2(n11352), .ZN(n12180) );
  AND2_X1 U11693 ( .A1(n11354), .A2(n12095), .ZN(n11353) );
  NOR2_X1 U11694 ( .A1(n12350), .A2(n12351), .ZN(n12626) );
  AND2_X1 U11695 ( .A1(n11414), .A2(n11090), .ZN(n13304) );
  INV_X1 U11696 ( .A(n13359), .ZN(n11275) );
  XNOR2_X1 U11697 ( .A(n12526), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13354) );
  INV_X1 U11698 ( .A(n16436), .ZN(n11224) );
  NAND2_X1 U11699 ( .A1(n16570), .A2(n11222), .ZN(n16548) );
  NOR2_X1 U11700 ( .A1(n11077), .A2(n11223), .ZN(n11222) );
  INV_X1 U11701 ( .A(n16545), .ZN(n11223) );
  INV_X1 U11702 ( .A(n11336), .ZN(n11334) );
  OAI21_X1 U11703 ( .B1(n12494), .B2(n11337), .A(n11409), .ZN(n11336) );
  NAND2_X1 U11704 ( .A1(n11340), .A2(n13277), .ZN(n11337) );
  INV_X1 U11705 ( .A(n15494), .ZN(n11227) );
  INV_X1 U11706 ( .A(n11150), .ZN(n11149) );
  OAI21_X1 U11707 ( .B1(n16775), .B2(n11151), .A(n16833), .ZN(n11150) );
  INV_X1 U11708 ( .A(n12211), .ZN(n11151) );
  INV_X1 U11709 ( .A(n13285), .ZN(n11375) );
  NAND2_X1 U11710 ( .A1(n16660), .A2(n11113), .ZN(n11115) );
  NOR2_X1 U11711 ( .A1(n11376), .A2(n11114), .ZN(n11113) );
  NAND2_X1 U11712 ( .A1(n11263), .A2(n11262), .ZN(n15505) );
  INV_X1 U11713 ( .A(n15502), .ZN(n11262) );
  INV_X1 U11714 ( .A(n15503), .ZN(n11263) );
  AND2_X1 U11715 ( .A1(n15317), .A2(n15396), .ZN(n15398) );
  NOR2_X1 U11716 ( .A1(n15697), .A2(n12555), .ZN(n11377) );
  AND3_X1 U11717 ( .A1(n12745), .A2(n12744), .A3(n12743), .ZN(n15308) );
  NOR2_X1 U11718 ( .A1(n14834), .A2(n11273), .ZN(n11272) );
  INV_X1 U11719 ( .A(n12263), .ZN(n11273) );
  AND2_X1 U11720 ( .A1(n12620), .A2(n15440), .ZN(n12933) );
  AND3_X1 U11721 ( .A1(n12613), .A2(n14953), .A3(n12612), .ZN(n12618) );
  AOI21_X1 U11722 ( .B1(n14681), .B2(n12956), .A(n12955), .ZN(n14805) );
  AOI21_X1 U11723 ( .B1(n12953), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12951), .ZN(n12952) );
  XNOR2_X1 U11724 ( .A(n12962), .B(n12960), .ZN(n14830) );
  NAND2_X1 U11725 ( .A1(n19431), .A2(n19579), .ZN(n19342) );
  NAND2_X1 U11726 ( .A1(n19431), .A2(n17426), .ZN(n19314) );
  NAND2_X1 U11727 ( .A1(n19424), .A2(n19425), .ZN(n17097) );
  NOR2_X1 U11728 ( .A1(n19424), .A2(n19694), .ZN(n19324) );
  NOR2_X1 U11729 ( .A1(n19424), .A2(n19425), .ZN(n17096) );
  INV_X1 U11730 ( .A(n19362), .ZN(n19700) );
  NAND2_X1 U11731 ( .A1(n19293), .A2(n12654), .ZN(n19355) );
  INV_X1 U11732 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17057) );
  NOR2_X1 U11733 ( .A1(n11478), .A2(n11477), .ZN(n11479) );
  INV_X1 U11734 ( .A(n11471), .ZN(n11481) );
  NOR2_X1 U11735 ( .A1(n11429), .A2(n11428), .ZN(n11560) );
  NOR2_X1 U11736 ( .A1(n14558), .A2(n20824), .ZN(n11517) );
  OR3_X1 U11737 ( .A1(n20596), .A2(n20595), .A3(n20594), .ZN(n20597) );
  XNOR2_X1 U11738 ( .A(n20774), .B(n20864), .ZN(n18270) );
  NAND2_X1 U11739 ( .A1(n11212), .A2(n11067), .ZN(n11219) );
  INV_X1 U11740 ( .A(n20625), .ZN(n17893) );
  NAND2_X1 U11741 ( .A1(n11547), .A2(n11545), .ZN(n17949) );
  NOR2_X1 U11742 ( .A1(n11524), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11199) );
  NAND2_X1 U11743 ( .A1(n18262), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11195) );
  NAND2_X1 U11744 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20780), .ZN(
        n18278) );
  NAND2_X1 U11745 ( .A1(n20797), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n20823) );
  NAND2_X1 U11746 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11427), .ZN(
        n20824) );
  INV_X1 U11747 ( .A(n21172), .ZN(n21204) );
  AOI211_X1 U11748 ( .C1(n15645), .C2(n15644), .A(n15643), .B(n15642), .ZN(
        n21234) );
  INV_X1 U11749 ( .A(n21256), .ZN(n21235) );
  NAND2_X1 U11750 ( .A1(n15857), .A2(n11103), .ZN(n15827) );
  NOR2_X1 U11751 ( .A1(n21454), .A2(n21453), .ZN(n21460) );
  OR2_X1 U11752 ( .A1(n11170), .A2(n11169), .ZN(n21454) );
  NAND2_X1 U11753 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n11169) );
  NOR2_X1 U11754 ( .A1(n15250), .A2(n16379), .ZN(n14513) );
  NAND2_X1 U11755 ( .A1(n21403), .A2(n14514), .ZN(n21567) );
  AND2_X1 U11756 ( .A1(n14524), .A2(n14516), .ZN(n21519) );
  NAND2_X1 U11757 ( .A1(n16039), .A2(n14888), .ZN(n16027) );
  OR2_X1 U11758 ( .A1(n14533), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21288) );
  AND2_X1 U11759 ( .A1(n13986), .A2(n13967), .ZN(n21345) );
  NAND2_X1 U11760 ( .A1(n11316), .A2(n14748), .ZN(n21872) );
  AND2_X1 U11761 ( .A1(n15017), .A2(n15440), .ZN(n18371) );
  NAND2_X1 U11762 ( .A1(n18634), .A2(n15429), .ZN(n18648) );
  NAND2_X1 U11763 ( .A1(n18618), .A2(n18619), .ZN(n18634) );
  INV_X1 U11764 ( .A(n18640), .ZN(n18598) );
  AND2_X1 U11765 ( .A1(n12760), .A2(n12759), .ZN(n15112) );
  AND2_X1 U11766 ( .A1(n12725), .A2(n12724), .ZN(n15054) );
  INV_X1 U11767 ( .A(n19694), .ZN(n19425) );
  NAND2_X1 U11768 ( .A1(n18721), .A2(n12254), .ZN(n17417) );
  AND2_X1 U11769 ( .A1(n17417), .A2(n14678), .ZN(n17407) );
  INV_X1 U11770 ( .A(n17407), .ZN(n16782) );
  AOI21_X1 U11771 ( .B1(n11040), .B2(n12928), .A(n12927), .ZN(n12929) );
  XNOR2_X1 U11772 ( .A(n12931), .B(n15280), .ZN(n15765) );
  OR2_X1 U11773 ( .A1(n15803), .A2(n18662), .ZN(n11231) );
  AOI21_X1 U11774 ( .B1(n15709), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11230), .ZN(n11229) );
  NAND2_X1 U11775 ( .A1(n15708), .A2(n15707), .ZN(n11230) );
  XNOR2_X1 U11776 ( .A(n12544), .B(n12543), .ZN(n15715) );
  OAI211_X1 U11777 ( .C1(n13319), .C2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13318), .B(n11397), .ZN(n13320) );
  INV_X1 U11778 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19353) );
  INV_X1 U11779 ( .A(n19579), .ZN(n17426) );
  OR4_X1 U11780 ( .A1(n17057), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .A4(P2_STATEBS16_REG_SCAN_IN), .ZN(n18701)
         );
  NAND2_X1 U11781 ( .A1(n20580), .A2(n20579), .ZN(n11293) );
  NAND2_X1 U11782 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21202), .ZN(n21256) );
  NAND2_X1 U11783 ( .A1(n21245), .A2(n11134), .ZN(n21250) );
  NAND2_X1 U11784 ( .A1(n21607), .A2(n17117), .ZN(n11134) );
  INV_X1 U11785 ( .A(n13828), .ZN(n11380) );
  INV_X1 U11786 ( .A(n13666), .ZN(n13687) );
  XNOR2_X1 U11787 ( .A(n11804), .B(n12400), .ZN(n12604) );
  NAND2_X1 U11788 ( .A1(n11351), .A2(n11867), .ZN(n12606) );
  INV_X1 U11789 ( .A(n12604), .ZN(n11351) );
  INV_X1 U11790 ( .A(n12582), .ZN(n12588) );
  OAI22_X1 U11791 ( .A1(n13789), .A2(n13788), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13370), .ZN(n13782) );
  AND2_X1 U11792 ( .A1(n13709), .A2(n13708), .ZN(n13712) );
  OR2_X1 U11793 ( .A1(n13806), .A2(n13707), .ZN(n13708) );
  NAND2_X1 U11794 ( .A1(n13814), .A2(n13822), .ZN(n11175) );
  OR2_X1 U11795 ( .A1(n13806), .A2(n13822), .ZN(n11173) );
  NOR2_X1 U11796 ( .A1(n11053), .A2(n11164), .ZN(n11163) );
  AOI22_X1 U11797 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13451), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13407) );
  AOI22_X1 U11798 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13450), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13408) );
  AOI22_X1 U11799 ( .A1(n13432), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13431), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13409) );
  AOI22_X1 U11800 ( .A1(n13443), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U11801 ( .A1(n13458), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13396) );
  AOI22_X1 U11802 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13379) );
  OR2_X1 U11803 ( .A1(n12002), .A2(n12001), .ZN(n12358) );
  NOR2_X1 U11804 ( .A1(n11139), .A2(n18711), .ZN(n11136) );
  AND2_X1 U11805 ( .A1(n14717), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11137) );
  AND2_X1 U11806 ( .A1(n19353), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12242) );
  OR2_X1 U11807 ( .A1(n12588), .A2(n12586), .ZN(n12585) );
  OR2_X1 U11808 ( .A1(n11330), .A2(n11959), .ZN(n12025) );
  AOI21_X1 U11809 ( .B1(n12231), .B2(n12230), .A(n12229), .ZN(n12236) );
  OAI21_X1 U11810 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n11420), .A(
        n11716), .ZN(n11724) );
  NOR2_X1 U11811 ( .A1(n11430), .A2(n15640), .ZN(n11473) );
  NOR2_X1 U11812 ( .A1(n20633), .A2(n11531), .ZN(n11535) );
  OR2_X1 U11813 ( .A1(n11528), .A2(n20638), .ZN(n11531) );
  NAND2_X1 U11814 ( .A1(n11526), .A2(n11676), .ZN(n11528) );
  INV_X1 U11815 ( .A(n11366), .ZN(n11675) );
  OR2_X1 U11816 ( .A1(n11679), .A2(n11667), .ZN(n11366) );
  NOR2_X1 U11817 ( .A1(n15648), .A2(n11323), .ZN(n11322) );
  INV_X1 U11818 ( .A(n15833), .ZN(n11323) );
  INV_X1 U11819 ( .A(n15910), .ZN(n11327) );
  NOR2_X1 U11820 ( .A1(n15917), .A2(n11329), .ZN(n11328) );
  INV_X1 U11821 ( .A(n15926), .ZN(n11329) );
  NAND2_X1 U11822 ( .A1(n14152), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14472) );
  INV_X1 U11823 ( .A(n14472), .ZN(n14493) );
  NOR2_X1 U11824 ( .A1(n14235), .A2(n14234), .ZN(n14236) );
  OR2_X1 U11825 ( .A1(n14205), .A2(n15600), .ZN(n14235) );
  AND2_X1 U11826 ( .A1(n14229), .A2(n14142), .ZN(n15511) );
  NAND2_X1 U11827 ( .A1(n14067), .A2(n14066), .ZN(n15100) );
  INV_X1 U11828 ( .A(n15102), .ZN(n14066) );
  INV_X1 U11829 ( .A(n15103), .ZN(n14067) );
  AND2_X1 U11830 ( .A1(n15911), .A2(n15922), .ZN(n11190) );
  NAND2_X1 U11831 ( .A1(n16129), .A2(n13753), .ZN(n16113) );
  INV_X1 U11832 ( .A(n15953), .ZN(n11178) );
  AND2_X1 U11833 ( .A1(n15739), .A2(n11194), .ZN(n11193) );
  INV_X1 U11834 ( .A(n15601), .ZN(n11194) );
  OR2_X1 U11835 ( .A1(n13755), .A2(n13748), .ZN(n16157) );
  AND2_X1 U11836 ( .A1(n13845), .A2(n13860), .ZN(n14505) );
  INV_X1 U11837 ( .A(n13739), .ZN(n13723) );
  NOR2_X1 U11838 ( .A1(n13475), .A2(n17186), .ZN(n13583) );
  OR2_X1 U11839 ( .A1(n13614), .A2(n13613), .ZN(n13618) );
  NAND2_X1 U11840 ( .A1(n13814), .A2(n13792), .ZN(n13818) );
  NAND2_X1 U11841 ( .A1(n13502), .A2(n11315), .ZN(n11314) );
  NAND2_X1 U11842 ( .A1(n13596), .A2(n13595), .ZN(n11317) );
  NAND2_X1 U11843 ( .A1(n13601), .A2(n13600), .ZN(n13602) );
  AOI22_X1 U11844 ( .A1(n11417), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13458), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13384) );
  NAND2_X1 U11845 ( .A1(n21823), .A2(n17186), .ZN(n13641) );
  INV_X1 U11846 ( .A(n12533), .ZN(n12538) );
  NOR2_X1 U11847 ( .A1(n16413), .A2(n11304), .ZN(n11303) );
  INV_X1 U11848 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11304) );
  NOR3_X1 U11849 ( .A1(n12455), .A2(n11161), .A3(n11160), .ZN(n12503) );
  OR2_X1 U11850 ( .A1(n11080), .A2(n12496), .ZN(n11160) );
  INV_X1 U11851 ( .A(n12468), .ZN(n11154) );
  NOR2_X1 U11852 ( .A1(n11158), .A2(n11157), .ZN(n11156) );
  INV_X1 U11853 ( .A(n12413), .ZN(n11157) );
  CLKBUF_X1 U11854 ( .A(n10963), .Z(n15780) );
  AND2_X1 U11855 ( .A1(n12130), .A2(n12129), .ZN(n12682) );
  AND2_X1 U11856 ( .A1(n15477), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12561) );
  INV_X1 U11857 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15473) );
  AND2_X1 U11858 ( .A1(n11277), .A2(n16419), .ZN(n11276) );
  AND3_X1 U11859 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n16811), .ZN(n13323) );
  AND2_X1 U11860 ( .A1(n16491), .A2(n16498), .ZN(n11277) );
  NAND2_X1 U11861 ( .A1(n12215), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11148) );
  INV_X1 U11862 ( .A(n16586), .ZN(n11347) );
  NAND2_X1 U11863 ( .A1(n12859), .A2(n11226), .ZN(n11225) );
  INV_X1 U11864 ( .A(n16652), .ZN(n11376) );
  INV_X1 U11865 ( .A(n16661), .ZN(n11114) );
  INV_X1 U11866 ( .A(n15184), .ZN(n11280) );
  INV_X1 U11867 ( .A(n15071), .ZN(n11279) );
  AND2_X1 U11868 ( .A1(n11341), .A2(n16719), .ZN(n11340) );
  OR2_X1 U11869 ( .A1(n13277), .A2(n16730), .ZN(n11341) );
  AND2_X1 U11870 ( .A1(n17021), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11349) );
  NAND2_X1 U11871 ( .A1(n11002), .A2(n15565), .ZN(n16758) );
  AND2_X1 U11872 ( .A1(n12167), .A2(n12166), .ZN(n12684) );
  OAI21_X1 U11873 ( .B1(n12389), .B2(n12689), .A(n15424), .ZN(n12390) );
  NAND2_X1 U11874 ( .A1(n12134), .A2(n12091), .ZN(n12093) );
  INV_X1 U11875 ( .A(n12826), .ZN(n12846) );
  NAND2_X1 U11876 ( .A1(n11000), .A2(n11894), .ZN(n11914) );
  OAI22_X1 U11877 ( .A1(n11921), .A2(n11900), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11899), .ZN(n11117) );
  OAI211_X1 U11878 ( .C1(n11913), .C2(n18711), .A(n11116), .B(n11912), .ZN(
        n11940) );
  NOR2_X1 U11879 ( .A1(n11911), .A2(n11910), .ZN(n11116) );
  INV_X1 U11880 ( .A(n11853), .ZN(n11874) );
  AND2_X1 U11881 ( .A1(n12649), .A2(n12648), .ZN(n12659) );
  NAND2_X1 U11882 ( .A1(n11092), .A2(n11239), .ZN(n12649) );
  NOR2_X1 U11883 ( .A1(n12637), .A2(n12646), .ZN(n11239) );
  INV_X1 U11884 ( .A(n12878), .ZN(n12870) );
  NAND2_X1 U11885 ( .A1(n11123), .A2(n11880), .ZN(n11122) );
  NAND2_X1 U11886 ( .A1(n11886), .A2(n12901), .ZN(n11121) );
  OR2_X1 U11887 ( .A1(n12888), .A2(n12887), .ZN(n14962) );
  NAND2_X1 U11888 ( .A1(n11804), .A2(n11867), .ZN(n11853) );
  INV_X1 U11889 ( .A(n12025), .ZN(n12096) );
  INV_X1 U11890 ( .A(n11961), .ZN(n11956) );
  INV_X1 U11891 ( .A(n11808), .ZN(n11247) );
  OAI21_X1 U11892 ( .B1(n11839), .B2(n11838), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11840) );
  INV_X1 U11893 ( .A(n18657), .ZN(n15020) );
  AND3_X1 U11894 ( .A1(n14840), .A2(n11867), .A3(n12634), .ZN(n11876) );
  NAND2_X1 U11895 ( .A1(n11420), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11430) );
  INV_X1 U11896 ( .A(n11473), .ZN(n17747) );
  NOR2_X1 U11897 ( .A1(n11430), .A2(n20824), .ZN(n11508) );
  NOR2_X1 U11898 ( .A1(n11427), .A2(n11422), .ZN(n11458) );
  NAND2_X1 U11899 ( .A1(n11370), .A2(n11369), .ZN(n17731) );
  INV_X1 U11900 ( .A(n15640), .ZN(n11369) );
  INV_X1 U11901 ( .A(n14558), .ZN(n11370) );
  NAND2_X1 U11902 ( .A1(n17930), .A2(n20348), .ZN(n17912) );
  NOR2_X1 U11903 ( .A1(n11678), .A2(n11680), .ZN(n11679) );
  INV_X1 U11904 ( .A(n21093), .ZN(n11217) );
  NOR2_X1 U11905 ( .A1(n17889), .A2(n11752), .ZN(n17961) );
  OR2_X1 U11906 ( .A1(n21135), .A2(n17920), .ZN(n17901) );
  INV_X1 U11907 ( .A(n20653), .ZN(n11634) );
  AND2_X1 U11908 ( .A1(n18190), .A2(n18192), .ZN(n17935) );
  XNOR2_X1 U11909 ( .A(n11528), .B(n20638), .ZN(n11529) );
  INV_X1 U11910 ( .A(n11731), .ZN(n11666) );
  INV_X1 U11911 ( .A(n20799), .ZN(n11701) );
  AND2_X1 U11912 ( .A1(n20114), .A2(n20803), .ZN(n20598) );
  OAI21_X1 U11913 ( .B1(n11730), .B2(n11729), .A(n11728), .ZN(n21226) );
  INV_X1 U11914 ( .A(n11658), .ZN(n11661) );
  CLKBUF_X1 U11915 ( .A(n14505), .Z(n14658) );
  NOR2_X1 U11916 ( .A1(n13827), .A2(n13826), .ZN(n14738) );
  NAND2_X1 U11917 ( .A1(n15951), .A2(n15944), .ZN(n15943) );
  NOR2_X1 U11918 ( .A1(n19927), .A2(n11172), .ZN(n11171) );
  INV_X1 U11919 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n11172) );
  NOR2_X1 U11920 ( .A1(n15248), .A2(n21737), .ZN(n14524) );
  CLKBUF_X1 U11921 ( .A(n13968), .Z(n14882) );
  OR2_X1 U11922 ( .A1(n13856), .A2(n21616), .ZN(n21663) );
  NOR2_X1 U11923 ( .A1(n11325), .A2(n11321), .ZN(n11320) );
  INV_X1 U11924 ( .A(n11322), .ZN(n11321) );
  INV_X1 U11925 ( .A(n15730), .ZN(n11325) );
  NAND2_X1 U11926 ( .A1(n14416), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14417) );
  INV_X1 U11927 ( .A(n14415), .ZN(n14416) );
  OR2_X1 U11928 ( .A1(n14417), .A2(n15847), .ZN(n14453) );
  NAND2_X1 U11929 ( .A1(n14375), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14377) );
  INV_X1 U11930 ( .A(n14374), .ZN(n14375) );
  OR2_X1 U11931 ( .A1(n14377), .A2(n14376), .ZN(n14415) );
  AND2_X1 U11932 ( .A1(n15925), .A2(n11066), .ZN(n15909) );
  NAND2_X1 U11933 ( .A1(n15925), .A2(n11328), .ZN(n15919) );
  NAND2_X1 U11934 ( .A1(n14350), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14352) );
  OR2_X1 U11935 ( .A1(n14352), .A2(n14351), .ZN(n14374) );
  NAND2_X1 U11936 ( .A1(n14304), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14305) );
  NOR2_X1 U11937 ( .A1(n14305), .A2(n16117), .ZN(n14350) );
  INV_X1 U11938 ( .A(n15947), .ZN(n14289) );
  INV_X1 U11939 ( .A(n15946), .ZN(n14290) );
  AND2_X1 U11940 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n14266), .ZN(
        n14304) );
  OR2_X1 U11941 ( .A1(n14237), .A2(n15875), .ZN(n14265) );
  OR2_X1 U11942 ( .A1(n14158), .A2(n15886), .ZN(n14237) );
  NAND2_X1 U11943 ( .A1(n14175), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14158) );
  NOR2_X1 U11944 ( .A1(n14190), .A2(n15607), .ZN(n14175) );
  NAND2_X1 U11945 ( .A1(n14206), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14190) );
  INV_X1 U11946 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15607) );
  INV_X1 U11947 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14220) );
  NOR2_X1 U11948 ( .A1(n14128), .A2(n21436), .ZN(n14129) );
  NAND2_X1 U11949 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n14129), .ZN(
        n14219) );
  NAND2_X1 U11950 ( .A1(n14111), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14128) );
  INV_X1 U11951 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21436) );
  AOI21_X1 U11952 ( .B1(n14020), .B2(n14229), .A(n14019), .ZN(n15204) );
  AOI21_X1 U11953 ( .B1(n14072), .B2(n14229), .A(n14071), .ZN(n15124) );
  CLKBUF_X1 U11954 ( .A(n15100), .Z(n15101) );
  NOR2_X1 U11955 ( .A1(n14047), .A2(n14015), .ZN(n14060) );
  INV_X1 U11956 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14015) );
  AOI21_X1 U11957 ( .B1(n14024), .B2(n14045), .A(n11313), .ZN(n11312) );
  INV_X1 U11958 ( .A(n14044), .ZN(n11313) );
  NAND2_X1 U11959 ( .A1(n14780), .A2(n14779), .ZN(n14867) );
  INV_X1 U11960 ( .A(n13767), .ZN(n13769) );
  NAND2_X1 U11961 ( .A1(n11072), .A2(n11018), .ZN(n11385) );
  NAND3_X1 U11962 ( .A1(n16080), .A2(n13762), .A3(n11018), .ZN(n11386) );
  NAND2_X1 U11963 ( .A1(n15929), .A2(n11190), .ZN(n15913) );
  AND2_X1 U11964 ( .A1(n13943), .A2(n13942), .ZN(n15928) );
  NAND2_X1 U11965 ( .A1(n11389), .A2(n11388), .ZN(n13751) );
  AOI21_X1 U11966 ( .B1(n11021), .B2(n11391), .A(n11098), .ZN(n11388) );
  AND2_X1 U11967 ( .A1(n13914), .A2(n13913), .ZN(n15973) );
  NAND2_X1 U11968 ( .A1(n16333), .A2(n11193), .ZN(n15974) );
  NAND2_X1 U11969 ( .A1(n16333), .A2(n15739), .ZN(n15738) );
  AND2_X1 U11970 ( .A1(n13755), .A2(n16133), .ZN(n16321) );
  NAND2_X1 U11971 ( .A1(n16385), .A2(n17186), .ZN(n14533) );
  INV_X1 U11972 ( .A(n19972), .ZN(n13884) );
  NAND2_X1 U11973 ( .A1(n14864), .A2(n14863), .ZN(n15068) );
  NAND2_X1 U11974 ( .A1(n11188), .A2(n11186), .ZN(n17194) );
  INV_X1 U11975 ( .A(n15069), .ZN(n11186) );
  AND2_X1 U11976 ( .A1(n16365), .A2(n16312), .ZN(n21285) );
  AND2_X1 U11977 ( .A1(n13987), .A2(n16366), .ZN(n21284) );
  INV_X1 U11978 ( .A(n16286), .ZN(n16328) );
  NAND2_X1 U11979 ( .A1(n13986), .A2(n14664), .ZN(n21289) );
  OAI211_X1 U11980 ( .C1(n13546), .C2(n13860), .A(n13545), .B(n13544), .ZN(
        n13579) );
  AOI22_X1 U11981 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13451), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13466) );
  CLKBUF_X1 U11982 ( .A(n13854), .Z(n13855) );
  OR2_X1 U11983 ( .A1(n21821), .A2(n21820), .ZN(n21859) );
  NAND2_X1 U11984 ( .A1(n21751), .A2(n21750), .ZN(n21891) );
  INV_X1 U11985 ( .A(n13484), .ZN(n22117) );
  INV_X1 U11986 ( .A(n21852), .ZN(n21809) );
  AOI21_X1 U11987 ( .B1(n21885), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n22212), 
        .ZN(n21926) );
  NAND2_X1 U11988 ( .A1(n21732), .A2(n21731), .ZN(n22217) );
  AND2_X1 U11989 ( .A1(n16379), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13841) );
  INV_X1 U11990 ( .A(n13841), .ZN(n17179) );
  INV_X2 U11991 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21917) );
  OR2_X1 U11992 ( .A1(n12523), .A2(n12516), .ZN(n12533) );
  NOR2_X1 U11993 ( .A1(n12515), .A2(n12514), .ZN(n12518) );
  NAND2_X1 U11994 ( .A1(n12518), .A2(n12519), .ZN(n12523) );
  NAND2_X1 U11995 ( .A1(n16411), .A2(n11303), .ZN(n16416) );
  NAND2_X1 U11996 ( .A1(n16411), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16414) );
  NAND2_X1 U11997 ( .A1(n11153), .A2(n11091), .ZN(n12515) );
  INV_X1 U11998 ( .A(n11153), .ZN(n12511) );
  INV_X1 U11999 ( .A(n12503), .ZN(n12499) );
  NAND2_X1 U12000 ( .A1(n15402), .A2(n15403), .ZN(n15451) );
  AND2_X1 U12001 ( .A1(n12464), .A2(n12461), .ZN(n18482) );
  NAND2_X1 U12002 ( .A1(n12440), .A2(n12471), .ZN(n12475) );
  NAND2_X1 U12003 ( .A1(n12440), .A2(n11023), .ZN(n12470) );
  AND2_X1 U12004 ( .A1(n15004), .A2(n15440), .ZN(n14569) );
  AND2_X1 U12005 ( .A1(n12804), .A2(n12803), .ZN(n12974) );
  AND2_X1 U12006 ( .A1(n16422), .A2(n13362), .ZN(n13360) );
  NOR2_X1 U12007 ( .A1(n16538), .A2(n16421), .ZN(n16422) );
  NAND2_X1 U12008 ( .A1(n11261), .A2(n16517), .ZN(n11252) );
  AND2_X1 U12009 ( .A1(n15519), .A2(n13080), .ZN(n16515) );
  NOR2_X1 U12010 ( .A1(n17030), .A2(n17029), .ZN(n17007) );
  AND3_X1 U12011 ( .A1(n12667), .A2(n11233), .A3(n15215), .ZN(n11232) );
  AND2_X1 U12012 ( .A1(n14716), .A2(n21630), .ZN(n17448) );
  NAND2_X1 U12013 ( .A1(n16403), .A2(n11034), .ZN(n16406) );
  NAND2_X1 U12014 ( .A1(n11300), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16408) );
  INV_X1 U12015 ( .A(n16406), .ZN(n11300) );
  NAND2_X1 U12016 ( .A1(n16403), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16402) );
  AND2_X1 U12017 ( .A1(n15477), .A2(n11032), .ZN(n16399) );
  AND2_X1 U12018 ( .A1(n15477), .A2(n11064), .ZN(n16398) );
  NAND2_X1 U12019 ( .A1(n15477), .A2(n11029), .ZN(n16397) );
  AND2_X1 U12020 ( .A1(n15475), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15477) );
  NAND2_X1 U12021 ( .A1(n11305), .A2(n11031), .ZN(n15474) );
  NAND2_X1 U12022 ( .A1(n11305), .A2(n11306), .ZN(n15470) );
  NOR2_X1 U12023 ( .A1(n15281), .A2(n16768), .ZN(n15288) );
  NOR2_X1 U12024 ( .A1(n17406), .A2(n11309), .ZN(n11308) );
  NAND2_X1 U12025 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11309) );
  INV_X1 U12026 ( .A(n11110), .ZN(n11109) );
  NOR2_X1 U12027 ( .A1(n14834), .A2(n11270), .ZN(n11271) );
  NAND2_X1 U12028 ( .A1(n14824), .A2(n12263), .ZN(n11270) );
  NOR2_X1 U12029 ( .A1(n15285), .A2(n15339), .ZN(n15219) );
  NAND2_X1 U12030 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15285) );
  NAND2_X1 U12031 ( .A1(n11146), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11145) );
  INV_X1 U12032 ( .A(n11148), .ZN(n11146) );
  AND2_X1 U12033 ( .A1(n11414), .A2(n16498), .ZN(n16500) );
  INV_X1 U12034 ( .A(n12215), .ZN(n11147) );
  INV_X1 U12035 ( .A(n16637), .ZN(n11332) );
  NAND2_X1 U12036 ( .A1(n16732), .A2(n11338), .ZN(n11333) );
  NOR2_X1 U12037 ( .A1(n12494), .A2(n11339), .ZN(n11338) );
  INV_X1 U12038 ( .A(n11340), .ZN(n11339) );
  AND2_X1 U12039 ( .A1(n13291), .A2(n11102), .ZN(n11358) );
  OR2_X1 U12040 ( .A1(n12480), .A2(n12479), .ZN(n13287) );
  INV_X1 U12041 ( .A(n13286), .ZN(n11373) );
  INV_X1 U12042 ( .A(n15370), .ZN(n11264) );
  NAND2_X1 U12043 ( .A1(n16692), .A2(n11358), .ZN(n16650) );
  NAND2_X1 U12044 ( .A1(n13284), .A2(n16671), .ZN(n16660) );
  NAND2_X1 U12045 ( .A1(n11279), .A2(n11278), .ZN(n15316) );
  AND2_X1 U12046 ( .A1(n11024), .A2(n12309), .ZN(n11278) );
  INV_X1 U12047 ( .A(n12559), .ZN(n12309) );
  INV_X1 U12048 ( .A(n16684), .ZN(n16676) );
  NAND2_X1 U12049 ( .A1(n11279), .A2(n11024), .ZN(n15186) );
  NOR2_X1 U12050 ( .A1(n11267), .A2(n11268), .ZN(n11266) );
  INV_X1 U12051 ( .A(n15108), .ZN(n11267) );
  NAND2_X1 U12053 ( .A1(n15425), .A2(n15427), .ZN(n15426) );
  AND2_X1 U12054 ( .A1(n12211), .A2(n12210), .ZN(n16775) );
  NAND2_X1 U12055 ( .A1(n16776), .A2(n16775), .ZN(n16774) );
  NAND2_X1 U12056 ( .A1(n15567), .A2(n12182), .ZN(n17022) );
  AND2_X1 U12057 ( .A1(n15353), .A2(n15352), .ZN(n15355) );
  INV_X1 U12058 ( .A(n15165), .ZN(n11233) );
  OAI211_X1 U12059 ( .C1(n12826), .C2(n14675), .A(n12640), .B(n12661), .ZN(
        n18386) );
  NAND2_X1 U12060 ( .A1(n12933), .A2(n12907), .ZN(n17002) );
  NAND2_X1 U12061 ( .A1(n12657), .A2(n12656), .ZN(n16460) );
  NAND2_X1 U12062 ( .A1(n12655), .A2(n12654), .ZN(n12657) );
  INV_X1 U12063 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14972) );
  INV_X1 U12064 ( .A(n15429), .ZN(n18517) );
  OR2_X1 U12065 ( .A1(n12943), .A2(n12942), .ZN(n11241) );
  INV_X1 U12066 ( .A(n19341), .ZN(n15233) );
  INV_X1 U12067 ( .A(n19641), .ZN(n19702) );
  NAND3_X1 U12068 ( .A1(n15131), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19361), 
        .ZN(n19706) );
  NAND3_X1 U12069 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n15130), .A3(n19361), 
        .ZN(n19707) );
  INV_X1 U12070 ( .A(n19225), .ZN(n19223) );
  INV_X1 U12071 ( .A(n19706), .ZN(n19698) );
  INV_X1 U12072 ( .A(n19707), .ZN(n19699) );
  NOR2_X1 U12073 ( .A1(n18377), .A2(n12594), .ZN(n12595) );
  NOR2_X1 U12074 ( .A1(n20595), .A2(n20106), .ZN(n11662) );
  OAI21_X1 U12075 ( .B1(n18364), .B2(n21648), .A(n18363), .ZN(n20105) );
  INV_X1 U12076 ( .A(n21226), .ZN(n21208) );
  AND2_X1 U12077 ( .A1(n17125), .A2(n20598), .ZN(n21207) );
  AOI21_X1 U12078 ( .B1(n20508), .B2(n11284), .A(n11282), .ZN(n11281) );
  OAI21_X1 U12079 ( .B1(n11283), .B2(n20523), .A(n20523), .ZN(n11282) );
  INV_X1 U12080 ( .A(n11284), .ZN(n11283) );
  AOI21_X1 U12081 ( .B1(n20523), .B2(n11285), .A(n20521), .ZN(n11284) );
  NOR2_X1 U12082 ( .A1(n17977), .A2(n17997), .ZN(n17995) );
  NAND2_X1 U12083 ( .A1(n17907), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n20430) );
  NOR2_X1 U12084 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20367), .ZN(n20385) );
  INV_X1 U12085 ( .A(n20586), .ZN(n20461) );
  AOI211_X1 U12086 ( .C1(n17725), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n11647), .B(n11646), .ZN(n11648) );
  NOR3_X1 U12087 ( .A1(n17125), .A2(n20105), .A3(n20113), .ZN(n18337) );
  OR2_X1 U12088 ( .A1(n21607), .A2(n20113), .ZN(n20599) );
  NOR2_X1 U12089 ( .A1(n21236), .A2(n20113), .ZN(n20115) );
  NAND2_X1 U12090 ( .A1(n18063), .A2(n11035), .ZN(n18109) );
  NAND2_X1 U12091 ( .A1(n18063), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18062) );
  NAND2_X1 U12092 ( .A1(n17995), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18026) );
  NAND2_X1 U12093 ( .A1(n17978), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17977) );
  NOR2_X1 U12094 ( .A1(n20430), .A2(n20169), .ZN(n17978) );
  NAND2_X1 U12095 ( .A1(n18118), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17891) );
  NOR2_X1 U12096 ( .A1(n17912), .A2(n20378), .ZN(n18118) );
  NAND2_X1 U12097 ( .A1(n20298), .A2(n11290), .ZN(n11289) );
  INV_X1 U12098 ( .A(n20269), .ZN(n11290) );
  INV_X1 U12099 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18156) );
  NAND2_X1 U12100 ( .A1(n18193), .A2(n11696), .ZN(n18149) );
  INV_X1 U12101 ( .A(n11694), .ZN(n11692) );
  NAND2_X1 U12102 ( .A1(n18214), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18181) );
  NAND3_X1 U12103 ( .A1(n11582), .A2(n11581), .A3(n11580), .ZN(n20596) );
  AOI22_X1 U12104 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17725), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11581) );
  AOI211_X1 U12105 ( .C1(n17823), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n11579), .B(n11578), .ZN(n11580) );
  INV_X1 U12106 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20181) );
  XNOR2_X1 U12107 ( .A(n11523), .B(n11522), .ZN(n18263) );
  INV_X1 U12108 ( .A(n18100), .ZN(n21057) );
  NOR2_X1 U12109 ( .A1(n11745), .A2(n11744), .ZN(n18097) );
  NOR2_X1 U12110 ( .A1(n17955), .A2(n21093), .ZN(n11215) );
  NAND2_X1 U12111 ( .A1(n17961), .A2(n11753), .ZN(n18012) );
  NOR2_X1 U12112 ( .A1(n18007), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11550) );
  INV_X1 U12113 ( .A(n11216), .ZN(n18023) );
  NOR2_X1 U12114 ( .A1(n11752), .A2(n20984), .ZN(n20839) );
  NAND2_X1 U12115 ( .A1(n18122), .A2(n18190), .ZN(n17985) );
  NAND2_X1 U12116 ( .A1(n17985), .A2(n17901), .ZN(n17899) );
  NOR2_X1 U12117 ( .A1(n11554), .A2(n11553), .ZN(n18123) );
  NOR2_X1 U12118 ( .A1(n11554), .A2(n11552), .ZN(n17920) );
  NOR2_X1 U12119 ( .A1(n20652), .A2(n20653), .ZN(n11736) );
  INV_X1 U12120 ( .A(n11740), .ZN(n21205) );
  NAND2_X1 U12121 ( .A1(n18149), .A2(n20958), .ZN(n18138) );
  NAND2_X1 U12122 ( .A1(n11542), .A2(n11207), .ZN(n11203) );
  NAND2_X1 U12123 ( .A1(n11206), .A2(n11205), .ZN(n11204) );
  NOR2_X1 U12124 ( .A1(n18201), .A2(n11541), .ZN(n18192) );
  NAND2_X1 U12125 ( .A1(n18216), .A2(n11691), .ZN(n18205) );
  OAI21_X1 U12126 ( .B1(n18227), .B2(n11209), .A(n11208), .ZN(n18212) );
  NAND2_X1 U12127 ( .A1(n11210), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11209) );
  NAND2_X1 U12128 ( .A1(n11534), .A2(n11210), .ZN(n11208) );
  XNOR2_X1 U12129 ( .A(n11533), .B(n11532), .ZN(n18227) );
  NOR2_X1 U12130 ( .A1(n18227), .A2(n20891), .ZN(n18226) );
  OR2_X1 U12131 ( .A1(n18232), .A2(n20883), .ZN(n18237) );
  NOR2_X1 U12132 ( .A1(n18249), .A2(n11197), .ZN(n11196) );
  INV_X1 U12133 ( .A(n11201), .ZN(n11197) );
  NOR2_X1 U12134 ( .A1(n11633), .A2(n11632), .ZN(n19087) );
  NOR2_X2 U12135 ( .A1(n11572), .A2(n11571), .ZN(n18997) );
  NOR2_X1 U12136 ( .A1(n11592), .A2(n11591), .ZN(n18957) );
  NOR2_X1 U12137 ( .A1(n11612), .A2(n11611), .ZN(n18916) );
  OR2_X1 U12138 ( .A1(n21221), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21219) );
  AOI22_X1 U12139 ( .A1(n21205), .A2(n21203), .B1(n21209), .B2(n20856), .ZN(
        n21232) );
  NOR2_X1 U12140 ( .A1(n17883), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n21202) );
  NAND2_X1 U12141 ( .A1(n20106), .A2(n11661), .ZN(n21236) );
  AND2_X1 U12142 ( .A1(n15857), .A2(n11101), .ZN(n15839) );
  AND2_X1 U12143 ( .A1(n15857), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15855) );
  NAND2_X1 U12144 ( .A1(n21556), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n21565) );
  INV_X1 U12145 ( .A(n21517), .ZN(n21529) );
  INV_X1 U12146 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15875) );
  AND2_X1 U12147 ( .A1(n15879), .A2(n11171), .ZN(n21483) );
  NAND2_X1 U12148 ( .A1(n15879), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15880) );
  NAND2_X1 U12149 ( .A1(n11167), .A2(n11166), .ZN(n11165) );
  INV_X1 U12150 ( .A(n15742), .ZN(n11166) );
  INV_X1 U12151 ( .A(n11168), .ZN(n11167) );
  INV_X1 U12152 ( .A(n21564), .ZN(n21546) );
  AND2_X1 U12153 ( .A1(n14514), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21564) );
  INV_X1 U12154 ( .A(n21476), .ZN(n21492) );
  NAND2_X1 U12155 ( .A1(n15872), .A2(n15873), .ZN(n15961) );
  AND2_X2 U12156 ( .A1(n14709), .A2(n14880), .ZN(n19989) );
  INV_X1 U12157 ( .A(n15658), .ZN(n16029) );
  INV_X2 U12158 ( .A(n15655), .ZN(n16039) );
  NOR2_X2 U12159 ( .A1(n14890), .A2(n15616), .ZN(n16040) );
  NOR2_X1 U12160 ( .A1(n19882), .A2(n21264), .ZN(n19894) );
  NOR2_X1 U12161 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15035), .ZN(n19897) );
  BUF_X1 U12162 ( .A(n19894), .Z(n19905) );
  BUF_X1 U12163 ( .A(n19897), .Z(n21264) );
  NAND2_X1 U12164 ( .A1(n11017), .A2(n14693), .ZN(n21720) );
  INV_X1 U12165 ( .A(n21720), .ZN(n21721) );
  XNOR2_X1 U12166 ( .A(n14512), .B(n14511), .ZN(n15250) );
  OAI21_X1 U12167 ( .B1(n15831), .B2(n15833), .A(n15832), .ZN(n16066) );
  INV_X1 U12168 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16117) );
  AND2_X1 U12169 ( .A1(n15958), .A2(n15946), .ZN(n21499) );
  INV_X1 U12170 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n21478) );
  OR2_X1 U12171 ( .A1(n15457), .A2(n15459), .ZN(n21440) );
  CLKBUF_X1 U12172 ( .A(n15379), .Z(n15380) );
  INV_X1 U12173 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15532) );
  AND2_X1 U12174 ( .A1(n16164), .A2(n14536), .ZN(n20033) );
  CLKBUF_X1 U12175 ( .A(n14872), .Z(n14873) );
  INV_X1 U12176 ( .A(n21574), .ZN(n20039) );
  OAI211_X1 U12177 ( .C1(n16045), .C2(n16048), .A(n16047), .B(n16046), .ZN(
        n16050) );
  INV_X1 U12178 ( .A(n21319), .ZN(n16358) );
  CLKBUF_X1 U12179 ( .A(n15090), .Z(n15091) );
  NOR2_X1 U12180 ( .A1(n21285), .A2(n14725), .ZN(n21302) );
  INV_X1 U12181 ( .A(n21289), .ZN(n21305) );
  INV_X1 U12182 ( .A(n21339), .ZN(n21346) );
  INV_X1 U12183 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21885) );
  INV_X1 U12184 ( .A(n21868), .ZN(n21923) );
  NAND2_X2 U12185 ( .A1(n14025), .A2(n14030), .ZN(n21759) );
  INV_X1 U12186 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17191) );
  OAI21_X1 U12187 ( .B1(n14925), .B2(n21578), .A(n22212), .ZN(n17190) );
  NAND2_X1 U12188 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13843), .ZN(n16380) );
  NOR2_X1 U12189 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16385) );
  OAI21_X1 U12190 ( .B1(n22245), .B2(n21790), .A(n21907), .ZN(n22247) );
  NOR2_X2 U12191 ( .A1(n21810), .A2(n21891), .ZN(n22257) );
  OAI211_X1 U12192 ( .C1(n22269), .C2(n21881), .A(n21849), .B(n21830), .ZN(
        n22272) );
  AOI22_X1 U12193 ( .A1(n21879), .A2(n21876), .B1(n21874), .B2(n21873), .ZN(
        n22302) );
  OAI211_X1 U12194 ( .C1(n22310), .C2(n21908), .A(n21907), .B(n21906), .ZN(
        n22313) );
  NOR2_X1 U12195 ( .A1(n22212), .A2(n21729), .ZN(n21922) );
  NOR2_X1 U12196 ( .A1(n22212), .A2(n21976), .ZN(n22017) );
  NOR2_X1 U12197 ( .A1(n22212), .A2(n22022), .ZN(n22063) );
  NOR2_X1 U12198 ( .A1(n22212), .A2(n22068), .ZN(n22109) );
  NOR2_X1 U12199 ( .A1(n22212), .A2(n22114), .ZN(n22159) );
  NOR2_X1 U12200 ( .A1(n22212), .A2(n22164), .ZN(n22206) );
  NOR2_X2 U12201 ( .A1(n21895), .A2(n21809), .ZN(n22322) );
  NOR2_X1 U12202 ( .A1(n22212), .A2(n22211), .ZN(n22319) );
  NAND2_X1 U12203 ( .A1(n13841), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21592) );
  NAND2_X1 U12204 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21667) );
  INV_X1 U12205 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21611) );
  INV_X1 U12206 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n19909) );
  NAND2_X1 U12207 ( .A1(n18607), .A2(n18608), .ZN(n18616) );
  NAND2_X1 U12208 ( .A1(n16417), .A2(n16580), .ZN(n18605) );
  NAND2_X1 U12209 ( .A1(n11297), .A2(n11295), .ZN(n18588) );
  AOI21_X1 U12210 ( .B1(n18606), .B2(n16608), .A(n11296), .ZN(n11295) );
  INV_X1 U12211 ( .A(n18590), .ZN(n11296) );
  NAND2_X1 U12212 ( .A1(n11294), .A2(n15429), .ZN(n18589) );
  OR2_X1 U12213 ( .A1(n16430), .A2(n16608), .ZN(n11294) );
  NAND2_X1 U12214 ( .A1(n16430), .A2(n15429), .ZN(n18578) );
  NAND2_X1 U12215 ( .A1(n18578), .A2(n18579), .ZN(n18577) );
  NAND2_X1 U12216 ( .A1(n16431), .A2(n16619), .ZN(n16430) );
  OR2_X1 U12217 ( .A1(n12654), .A2(n18639), .ZN(n18596) );
  NAND2_X1 U12218 ( .A1(n18567), .A2(n18568), .ZN(n18566) );
  NAND2_X1 U12219 ( .A1(n16443), .A2(n18606), .ZN(n18558) );
  NAND2_X1 U12220 ( .A1(n18558), .A2(n18559), .ZN(n18557) );
  NAND2_X1 U12221 ( .A1(n16445), .A2(n16444), .ZN(n16443) );
  NAND2_X1 U12222 ( .A1(n18606), .A2(n11407), .ZN(n18547) );
  NAND2_X1 U12223 ( .A1(n18547), .A2(n18546), .ZN(n18545) );
  AND2_X1 U12224 ( .A1(n11038), .A2(n12447), .ZN(n18544) );
  AND2_X1 U12225 ( .A1(n15298), .A2(n15297), .ZN(n18640) );
  OR2_X1 U12226 ( .A1(n18371), .A2(n15292), .ZN(n18627) );
  AND2_X1 U12227 ( .A1(n18371), .A2(n15307), .ZN(n18644) );
  INV_X1 U12229 ( .A(n18701), .ZN(n18617) );
  OR2_X1 U12230 ( .A1(n15302), .A2(n15301), .ZN(n18529) );
  AND2_X1 U12231 ( .A1(n15299), .A2(n15293), .ZN(n18645) );
  AND2_X1 U12232 ( .A1(n12823), .A2(n12822), .ZN(n15189) );
  NOR2_X1 U12233 ( .A1(n15188), .A2(n15189), .ZN(n15187) );
  INV_X1 U12234 ( .A(n16524), .ZN(n15147) );
  INV_X1 U12235 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n14843) );
  OR2_X2 U12236 ( .A1(n16513), .A2(n14813), .ZN(n16524) );
  NAND2_X1 U12237 ( .A1(n15402), .A2(n11228), .ZN(n15495) );
  INV_X1 U12238 ( .A(n13053), .ZN(n15493) );
  AND2_X1 U12239 ( .A1(n19188), .A2(n14617), .ZN(n19185) );
  INV_X1 U12240 ( .A(n19189), .ZN(n16574) );
  NOR3_X1 U12241 ( .A1(n11235), .A2(n15308), .A3(n11234), .ZN(n16958) );
  INV_X1 U12242 ( .A(n15427), .ZN(n11234) );
  AND2_X1 U12243 ( .A1(n19636), .A2(n19688), .ZN(n19220) );
  INV_X1 U12244 ( .A(n19686), .ZN(n19631) );
  INV_X1 U12245 ( .A(n19688), .ZN(n19633) );
  NAND2_X1 U12246 ( .A1(n13255), .A2(n15440), .ZN(n13258) );
  NAND2_X1 U12247 ( .A1(n19686), .A2(n14813), .ZN(n19688) );
  OAI21_X2 U12249 ( .B1(n14574), .B2(n21624), .A(n14714), .ZN(n14630) );
  INV_X1 U12250 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16605) );
  INV_X1 U12251 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16768) );
  INV_X1 U12252 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17418) );
  AND2_X1 U12253 ( .A1(n11152), .A2(n12180), .ZN(n17401) );
  AOI22_X1 U12254 ( .A1(n16578), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n13353), .B2(n13352), .ZN(n13356) );
  NOR2_X1 U12255 ( .A1(n13334), .A2(n11077), .ZN(n16546) );
  AND2_X1 U12256 ( .A1(n16692), .A2(n11357), .ZN(n13293) );
  AND2_X1 U12257 ( .A1(n11358), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11357) );
  AND2_X1 U12258 ( .A1(n15370), .A2(n15372), .ZN(n18520) );
  NAND2_X1 U12259 ( .A1(n13282), .A2(n13281), .ZN(n15696) );
  NAND2_X1 U12260 ( .A1(n11274), .A2(n12263), .ZN(n14835) );
  NAND2_X1 U12261 ( .A1(n15323), .A2(n12667), .ZN(n15164) );
  NAND2_X1 U12262 ( .A1(n12090), .A2(n12058), .ZN(n11356) );
  NAND2_X1 U12263 ( .A1(n12933), .A2(n15010), .ZN(n17005) );
  AND2_X1 U12264 ( .A1(n14809), .A2(n14808), .ZN(n19424) );
  INV_X1 U12265 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19257) );
  OR2_X1 U12266 ( .A1(n19314), .A2(n19424), .ZN(n19298) );
  INV_X1 U12267 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17137) );
  NOR2_X1 U12268 ( .A1(n14842), .A2(n14841), .ZN(n19694) );
  NAND2_X1 U12269 ( .A1(n14828), .A2(n14831), .ZN(n19579) );
  INV_X1 U12270 ( .A(n19620), .ZN(n19788) );
  NAND2_X1 U12271 ( .A1(n19309), .A2(n19308), .ZN(n19769) );
  INV_X1 U12272 ( .A(n19613), .ZN(n19774) );
  OAI21_X1 U12273 ( .B1(n19276), .B2(n19275), .A(n19274), .ZN(n19740) );
  AOI22_X1 U12274 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19699), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19698), .ZN(n19624) );
  INV_X1 U12275 ( .A(n19744), .ZN(n19733) );
  NOR2_X1 U12276 ( .A1(n19248), .A2(n19247), .ZN(n19651) );
  INV_X1 U12277 ( .A(n19630), .ZN(n19621) );
  AOI22_X1 U12278 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19698), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19699), .ZN(n19677) );
  INV_X1 U12279 ( .A(n19684), .ZN(n19674) );
  NAND2_X1 U12280 ( .A1(n19223), .A2(n15233), .ZN(n19724) );
  OAI22_X1 U12281 ( .A1(n22119), .A2(n19707), .B1(n20660), .B2(n19706), .ZN(
        n19476) );
  AOI22_X1 U12282 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19699), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19698), .ZN(n19409) );
  OAI22_X1 U12283 ( .A1(n22166), .A2(n19707), .B1(n20706), .B2(n19706), .ZN(
        n19415) );
  INV_X1 U12284 ( .A(n19724), .ZN(n19590) );
  NAND2_X1 U12285 ( .A1(n19241), .A2(n19240), .ZN(n19715) );
  OAI22_X1 U12286 ( .A1(n21747), .A2(n19707), .B1(n20753), .B2(n19706), .ZN(
        n19810) );
  AOI22_X1 U12287 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19699), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19698), .ZN(n19818) );
  AOI22_X1 U12288 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19698), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19699), .ZN(n19630) );
  INV_X1 U12289 ( .A(n19624), .ZN(n19627) );
  INV_X1 U12290 ( .A(n19585), .ZN(n19625) );
  AOI22_X1 U12291 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19699), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19698), .ZN(n19571) );
  INV_X1 U12292 ( .A(n19568), .ZN(n19573) );
  AOI22_X1 U12293 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19699), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19698), .ZN(n19523) );
  INV_X1 U12294 ( .A(n19517), .ZN(n19527) );
  INV_X1 U12295 ( .A(n19462), .ZN(n19474) );
  INV_X1 U12296 ( .A(n19452), .ZN(n19473) );
  INV_X1 U12297 ( .A(n19476), .ZN(n19472) );
  INV_X1 U12298 ( .A(n19817), .ZN(n19709) );
  INV_X1 U12299 ( .A(n19409), .ZN(n19414) );
  AND2_X1 U12300 ( .A1(n19376), .A2(n19702), .ZN(n19413) );
  INV_X1 U12301 ( .A(n19415), .ZN(n19412) );
  INV_X1 U12302 ( .A(n19281), .ZN(n19357) );
  NAND2_X1 U12303 ( .A1(n19223), .A2(n17096), .ZN(n19817) );
  INV_X1 U12304 ( .A(n19712), .ZN(n19714) );
  OR2_X1 U12305 ( .A1(n15128), .A2(n12654), .ZN(n18706) );
  NAND3_X1 U12306 ( .A1(n17057), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18718) );
  INV_X1 U12307 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19293) );
  INV_X1 U12308 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n12654) );
  NOR2_X1 U12309 ( .A1(n11663), .A2(n11662), .ZN(n20108) );
  NAND2_X1 U12310 ( .A1(n21235), .A2(n21208), .ZN(n20113) );
  NAND2_X1 U12311 ( .A1(n20522), .A2(n20523), .ZN(n20524) );
  OAI21_X1 U12312 ( .B1(n20508), .B2(n20556), .A(n11284), .ZN(n20530) );
  NOR2_X1 U12313 ( .A1(n20515), .A2(n20514), .ZN(n20558) );
  NAND2_X1 U12314 ( .A1(n20508), .A2(n20509), .ZN(n20522) );
  NOR2_X1 U12315 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n20475), .ZN(n20489) );
  NAND2_X1 U12316 ( .A1(n20465), .A2(n20466), .ZN(n20480) );
  NAND2_X1 U12317 ( .A1(n20455), .A2(n20456), .ZN(n20464) );
  NOR2_X1 U12318 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n20426), .ZN(n20439) );
  NOR2_X1 U12319 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20285), .ZN(n20306) );
  INV_X1 U12320 ( .A(n21243), .ZN(n20561) );
  NOR2_X1 U12321 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20254), .ZN(n20275) );
  INV_X1 U12322 ( .A(n20587), .ZN(n20564) );
  NAND4_X1 U12323 ( .A1(n11764), .A2(n20101), .A3(n21243), .A4(n21253), .ZN(
        n20586) );
  NOR3_X1 U12324 ( .A1(n20491), .A2(n20476), .A3(n17784), .ZN(n17779) );
  NAND2_X1 U12325 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17803), .ZN(n17784) );
  AND2_X1 U12326 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17790), .ZN(n17803) );
  NOR3_X1 U12327 ( .A1(n20106), .A2(n19087), .A3(n20594), .ZN(n17874) );
  INV_X1 U12328 ( .A(n20701), .ZN(n20724) );
  NOR2_X1 U12329 ( .A1(n20731), .A2(n20691), .ZN(n20697) );
  OR2_X1 U12330 ( .A1(n20728), .A2(n20729), .ZN(n20731) );
  NOR2_X1 U12331 ( .A1(n20676), .A2(n20681), .ZN(n20675) );
  INV_X1 U12332 ( .A(n20686), .ZN(n20682) );
  INV_X1 U12333 ( .A(n20740), .ZN(n20747) );
  INV_X1 U12334 ( .A(n20627), .ZN(n20773) );
  INV_X1 U12335 ( .A(n20621), .ZN(n20775) );
  NOR2_X1 U12336 ( .A1(n20767), .A2(n20784), .ZN(n20627) );
  NOR2_X1 U12337 ( .A1(n11436), .A2(n11435), .ZN(n20625) );
  INV_X1 U12338 ( .A(n20782), .ZN(n20645) );
  AND3_X1 U12339 ( .A1(n11481), .A2(n11480), .A3(n11479), .ZN(n11484) );
  NAND3_X1 U12340 ( .A1(n11520), .A2(n11519), .A3(n11518), .ZN(n20780) );
  NOR2_X1 U12341 ( .A1(n20600), .A2(n20775), .ZN(n20782) );
  NOR2_X1 U12342 ( .A1(n20114), .A2(n20599), .ZN(n20149) );
  CLKBUF_X1 U12344 ( .A(n20130), .Z(n20163) );
  NAND2_X1 U12345 ( .A1(n11368), .A2(n11367), .ZN(n18100) );
  NOR2_X1 U12346 ( .A1(n21036), .A2(n18042), .ZN(n11367) );
  INV_X1 U12347 ( .A(n21040), .ZN(n11368) );
  NOR2_X1 U12348 ( .A1(n17891), .A2(n20401), .ZN(n17907) );
  NAND3_X1 U12349 ( .A1(n21602), .A2(n18280), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18116) );
  INV_X1 U12350 ( .A(n18144), .ZN(n18197) );
  NOR2_X1 U12351 ( .A1(n20196), .A2(n20225), .ZN(n18214) );
  INV_X1 U12352 ( .A(n18280), .ZN(n18251) );
  INV_X1 U12353 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20225) );
  NOR2_X1 U12354 ( .A1(n20596), .A2(n21259), .ZN(n18225) );
  AND2_X1 U12355 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18241) );
  INV_X1 U12356 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20180) );
  INV_X1 U12357 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20169) );
  INV_X1 U12358 ( .A(n18172), .ZN(n18275) );
  INV_X1 U12359 ( .A(n18253), .ZN(n18276) );
  INV_X1 U12360 ( .A(n18225), .ZN(n18285) );
  INV_X1 U12361 ( .A(n21137), .ZN(n21114) );
  NOR3_X1 U12362 ( .A1(n21066), .A2(n21061), .A3(n11362), .ZN(n11361) );
  NAND2_X1 U12363 ( .A1(n11363), .A2(n11083), .ZN(n11362) );
  OR2_X1 U12364 ( .A1(n21126), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11363) );
  OR2_X1 U12365 ( .A1(n18012), .A2(n11754), .ZN(n21040) );
  NOR2_X1 U12366 ( .A1(n18140), .A2(n18139), .ZN(n20976) );
  NOR2_X1 U12367 ( .A1(n18138), .A2(n18140), .ZN(n20974) );
  NAND2_X1 U12368 ( .A1(n17893), .A2(n20914), .ZN(n21168) );
  OAI21_X1 U12369 ( .B1(n20980), .B2(n20929), .A(n21171), .ZN(n21200) );
  INV_X1 U12370 ( .A(n21168), .ZN(n21196) );
  INV_X1 U12371 ( .A(n20992), .ZN(n21171) );
  CLKBUF_X1 U12372 ( .A(n20992), .Z(n21194) );
  INV_X1 U12373 ( .A(n21210), .ZN(n20856) );
  INV_X1 U12374 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18802) );
  INV_X1 U12375 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17124) );
  INV_X1 U12376 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20813) );
  OAI21_X1 U12377 ( .B1(n20823), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n20807), .ZN(n21218) );
  NOR2_X1 U12378 ( .A1(n14557), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n20810) );
  INV_X1 U12379 ( .A(n20803), .ZN(n15641) );
  AOI211_X2 U12380 ( .C1(n21235), .C2(n21217), .A(n18752), .B(n15646), .ZN(
        n20833) );
  INV_X1 U12381 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21246) );
  NAND2_X1 U12382 ( .A1(n21645), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n21651) );
  OR2_X1 U12383 ( .A1(n15131), .A2(n14556), .ZN(n20049) );
  INV_X1 U12385 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19821) );
  AOI21_X1 U12386 ( .B1(n15820), .B2(n21567), .A(n15819), .ZN(n15821) );
  OR2_X1 U12387 ( .A1(n21572), .A2(n16170), .ZN(n11185) );
  AND2_X1 U12388 ( .A1(n14013), .A2(n14012), .ZN(n14014) );
  AOI21_X1 U12389 ( .B1(n18648), .B2(n18649), .A(n18701), .ZN(n18635) );
  NAND2_X1 U12390 ( .A1(n12547), .A2(n11142), .ZN(P2_U2984) );
  NAND2_X1 U12391 ( .A1(n11043), .A2(n12546), .ZN(n13312) );
  NAND2_X1 U12392 ( .A1(n15765), .A2(n15725), .ZN(n12934) );
  AND2_X1 U12393 ( .A1(n11231), .A2(n11229), .ZN(n15710) );
  NAND2_X1 U12394 ( .A1(n11043), .A2(n13329), .ZN(n13330) );
  OAI21_X1 U12395 ( .B1(n20572), .B2(n11081), .A(n11291), .ZN(P3_U2640) );
  NOR2_X1 U12396 ( .A1(n20578), .A2(n11292), .ZN(n11291) );
  OAI21_X1 U12397 ( .B1(n21060), .B2(n21168), .A(n11359), .ZN(P3_U2833) );
  NOR2_X1 U12398 ( .A1(n11364), .A2(n11360), .ZN(n11359) );
  OR2_X1 U12399 ( .A1(n21059), .A2(n21058), .ZN(n11364) );
  NOR3_X1 U12400 ( .A1(n11361), .A2(n21075), .A3(n10979), .ZN(n11360) );
  OAI21_X1 U12401 ( .B1(n21250), .B2(n11096), .A(n11133), .ZN(n21254) );
  NAND2_X1 U12402 ( .A1(n21252), .A2(n17883), .ZN(n11133) );
  OR2_X1 U12403 ( .A1(n20049), .A2(n20090), .ZN(U212) );
  NAND2_X2 U12404 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11119), .ZN(
        n13238) );
  INV_X1 U12405 ( .A(n13238), .ZN(n11842) );
  AND2_X1 U12406 ( .A1(n17066), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11014) );
  INV_X1 U12407 ( .A(n15285), .ZN(n11310) );
  AND4_X1 U12408 ( .A1(n11310), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11015) );
  AND2_X1 U12409 ( .A1(n16411), .A2(n11033), .ZN(n11016) );
  AND2_X1 U12410 ( .A1(n13843), .A2(n14880), .ZN(n11017) );
  OR2_X1 U12411 ( .A1(n16336), .A2(n13763), .ZN(n11018) );
  OAI21_X1 U12412 ( .B1(n16776), .B2(n11151), .A(n11149), .ZN(n13292) );
  OR2_X1 U12413 ( .A1(n18023), .A2(n18189), .ZN(n11019) );
  AND3_X1 U12414 ( .A1(n13465), .A2(n13464), .A3(n13463), .ZN(n11020) );
  OR2_X1 U12415 ( .A1(n15206), .A2(n13892), .ZN(n11022) );
  AND2_X1 U12416 ( .A1(n12471), .A2(n11154), .ZN(n11023) );
  NOR2_X1 U12417 ( .A1(n15119), .A2(n11280), .ZN(n11024) );
  AND4_X1 U12418 ( .A1(n11968), .A2(n11967), .A3(n11966), .A4(n11965), .ZN(
        n11025) );
  OR3_X1 U12419 ( .A1(n12455), .A2(n11161), .A3(n11080), .ZN(n11026) );
  NAND2_X1 U12420 ( .A1(n10999), .A2(n13722), .ZN(n20008) );
  AND4_X1 U12421 ( .A1(n13442), .A2(n13441), .A3(n13440), .A4(n13439), .ZN(
        n11027) );
  AND2_X1 U12422 ( .A1(n15402), .A2(n11089), .ZN(n13335) );
  AND2_X1 U12423 ( .A1(n11023), .A2(n11078), .ZN(n11028) );
  NAND2_X1 U12424 ( .A1(n15325), .A2(n15324), .ZN(n15323) );
  OR2_X1 U12425 ( .A1(n16931), .A2(n11059), .ZN(n15464) );
  AND2_X1 U12426 ( .A1(n11064), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11029) );
  NAND2_X1 U12427 ( .A1(n11250), .A2(n11413), .ZN(n11030) );
  OR2_X1 U12428 ( .A1(n16931), .A2(n11073), .ZN(n15197) );
  AND2_X1 U12429 ( .A1(n17007), .A2(n17006), .ZN(n15425) );
  AND2_X1 U12430 ( .A1(n11306), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11031) );
  INV_X1 U12431 ( .A(n11120), .ZN(n12882) );
  INV_X1 U12432 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15339) );
  AND2_X1 U12433 ( .A1(n11029), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11032) );
  AND2_X1 U12434 ( .A1(n11303), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11033) );
  AND2_X1 U12435 ( .A1(n11088), .A2(n15323), .ZN(n15214) );
  AND2_X1 U12436 ( .A1(n11298), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11034) );
  AND2_X1 U12437 ( .A1(n11286), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11035) );
  INV_X1 U12438 ( .A(n11975), .ZN(n13081) );
  AND2_X2 U12439 ( .A1(n12641), .A2(n12654), .ZN(n12647) );
  INV_X1 U12440 ( .A(n10970), .ZN(n13520) );
  INV_X1 U12441 ( .A(n10976), .ZN(n13522) );
  INV_X1 U12442 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11427) );
  AND2_X1 U12443 ( .A1(n13491), .A2(n13860), .ZN(n13864) );
  AND2_X1 U12444 ( .A1(n12652), .A2(n12359), .ZN(n11036) );
  NAND2_X1 U12445 ( .A1(n10998), .A2(n13744), .ZN(n16146) );
  NAND2_X1 U12446 ( .A1(n13491), .A2(n13473), .ZN(n13865) );
  NOR3_X2 U12447 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n14558), .ZN(n11509) );
  NAND2_X1 U12448 ( .A1(n11335), .A2(n11340), .ZN(n12550) );
  AND2_X1 U12449 ( .A1(n11960), .A2(n11950), .ZN(n12099) );
  AND2_X1 U12450 ( .A1(n16692), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12549) );
  NAND2_X1 U12451 ( .A1(n11204), .A2(n11203), .ZN(n11547) );
  OR2_X1 U12452 ( .A1(n16596), .A2(n11147), .ZN(n11037) );
  NAND2_X1 U12453 ( .A1(n17022), .A2(n17021), .ZN(n17023) );
  AND2_X1 U12454 ( .A1(n11318), .A2(n14236), .ZN(n15612) );
  NAND2_X1 U12455 ( .A1(n11140), .A2(n11908), .ZN(n11921) );
  NAND2_X1 U12456 ( .A1(n15925), .A2(n15926), .ZN(n15916) );
  XNOR2_X1 U12457 ( .A(n15703), .B(n15702), .ZN(n15803) );
  OR2_X1 U12458 ( .A1(n12455), .A2(n11161), .ZN(n11038) );
  AND2_X1 U12459 ( .A1(n11216), .A2(n11215), .ZN(n18018) );
  XOR2_X1 U12460 ( .A(n12881), .B(n12880), .Z(n11040) );
  OR2_X1 U12461 ( .A1(n12455), .A2(n12449), .ZN(n11041) );
  AND4_X1 U12462 ( .A1(n13462), .A2(n13461), .A3(n13460), .A4(n13459), .ZN(
        n11042) );
  INV_X1 U12463 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14776) );
  NAND2_X1 U12464 ( .A1(n13616), .A2(n13615), .ZN(n13617) );
  XNOR2_X1 U12465 ( .A(n13311), .B(n13310), .ZN(n11043) );
  XNOR2_X1 U12466 ( .A(n11936), .B(n11935), .ZN(n12944) );
  NAND2_X1 U12467 ( .A1(n11155), .A2(n12403), .ZN(n12405) );
  NAND2_X1 U12468 ( .A1(n16764), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16726) );
  AND2_X1 U12469 ( .A1(n11960), .A2(n11956), .ZN(n12106) );
  NAND2_X1 U12470 ( .A1(n11334), .A2(n10985), .ZN(n16634) );
  NAND2_X1 U12471 ( .A1(n11386), .A2(n11385), .ZN(n14005) );
  AND2_X1 U12472 ( .A1(n13491), .A2(n13500), .ZN(n11044) );
  NAND2_X1 U12473 ( .A1(n11414), .A2(n11276), .ZN(n13358) );
  NAND2_X1 U12474 ( .A1(n14829), .A2(n14830), .ZN(n14828) );
  INV_X1 U12475 ( .A(n13476), .ZN(n13470) );
  NOR3_X1 U12476 ( .A1(n11765), .A2(n21168), .A3(n18046), .ZN(n11047) );
  OR2_X1 U12477 ( .A1(n15983), .A2(n21553), .ZN(n11048) );
  AND2_X1 U12478 ( .A1(n16660), .A2(n16661), .ZN(n11050) );
  OR2_X1 U12479 ( .A1(n11527), .A2(n11525), .ZN(n11051) );
  NAND2_X1 U12480 ( .A1(n13751), .A2(n16336), .ZN(n16106) );
  OAI21_X1 U12481 ( .B1(n16611), .B2(n16614), .A(n16612), .ZN(n16586) );
  INV_X1 U12482 ( .A(n11260), .ZN(n16503) );
  NAND2_X1 U12483 ( .A1(n14872), .A2(n13624), .ZN(n13651) );
  AND2_X1 U12484 ( .A1(n13860), .A2(n11380), .ZN(n11052) );
  AND2_X1 U12485 ( .A1(n13450), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11053) );
  AND2_X1 U12486 ( .A1(n13720), .A2(n13693), .ZN(n11054) );
  INV_X1 U12488 ( .A(n11144), .ZN(n13357) );
  NOR2_X1 U12489 ( .A1(n16596), .A2(n11145), .ZN(n11144) );
  AND2_X1 U12490 ( .A1(n11866), .A2(n12600), .ZN(n11055) );
  AND4_X1 U12491 ( .A1(n13437), .A2(n13436), .A3(n13435), .A4(n13434), .ZN(
        n11056) );
  NOR2_X1 U12492 ( .A1(n20309), .A2(n18156), .ZN(n20298) );
  INV_X1 U12493 ( .A(n11765), .ZN(n18081) );
  NAND2_X1 U12494 ( .A1(n14290), .A2(n14289), .ZN(n15941) );
  AND2_X1 U12495 ( .A1(n11414), .A2(n11277), .ZN(n16418) );
  NAND2_X1 U12496 ( .A1(n12184), .A2(n12136), .ZN(n12389) );
  INV_X1 U12497 ( .A(n12389), .ZN(n11354) );
  OR2_X1 U12498 ( .A1(n20582), .A2(n20583), .ZN(n11057) );
  AND2_X1 U12499 ( .A1(n16758), .A2(n12411), .ZN(n11058) );
  AND2_X1 U12500 ( .A1(n13375), .A2(n14762), .ZN(n13604) );
  OR2_X1 U12501 ( .A1(n21262), .A2(n14508), .ZN(n14514) );
  AND2_X1 U12502 ( .A1(n13494), .A2(n13483), .ZN(n13830) );
  AND2_X1 U12503 ( .A1(n13820), .A2(n13819), .ZN(n13843) );
  OR2_X1 U12504 ( .A1(n11221), .A2(n16932), .ZN(n11059) );
  AND2_X1 U12505 ( .A1(n15972), .A2(n15883), .ZN(n15872) );
  NOR3_X1 U12506 ( .A1(n16931), .A2(n11059), .A3(n15465), .ZN(n11060) );
  AND2_X1 U12507 ( .A1(n18063), .A2(n11286), .ZN(n11061) );
  INV_X1 U12508 ( .A(n20523), .ZN(n20556) );
  NOR2_X1 U12509 ( .A1(n15071), .A2(n15119), .ZN(n15118) );
  NOR2_X1 U12510 ( .A1(n16931), .A2(n16932), .ZN(n11062) );
  OR2_X1 U12511 ( .A1(n13334), .A2(n16569), .ZN(n11063) );
  NAND2_X1 U12512 ( .A1(n12392), .A2(n12391), .ZN(n15564) );
  NAND2_X1 U12513 ( .A1(n11112), .A2(n12377), .ZN(n15208) );
  AND2_X1 U12514 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11064) );
  AND2_X1 U12515 ( .A1(n12361), .A2(n12362), .ZN(n12382) );
  INV_X1 U12516 ( .A(n13807), .ZN(n11174) );
  AND2_X1 U12517 ( .A1(n14236), .A2(n15614), .ZN(n11065) );
  XNOR2_X1 U12518 ( .A(n11260), .B(n11259), .ZN(n16495) );
  AND2_X1 U12519 ( .A1(n11328), .A2(n11327), .ZN(n11066) );
  NAND3_X1 U12520 ( .A1(n11152), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n12180), .ZN(n17400) );
  OR2_X1 U12521 ( .A1(n15527), .A2(n15530), .ZN(n15528) );
  NAND2_X1 U12522 ( .A1(n15090), .A2(n15093), .ZN(n15092) );
  NAND2_X1 U12523 ( .A1(n11265), .A2(n12290), .ZN(n15039) );
  NAND2_X1 U12524 ( .A1(n15528), .A2(n13743), .ZN(n15551) );
  NOR2_X1 U12525 ( .A1(n13334), .A2(n11225), .ZN(n16435) );
  OR2_X1 U12526 ( .A1(n11557), .A2(n18190), .ZN(n11067) );
  NAND2_X1 U12527 ( .A1(n19997), .A2(n13693), .ZN(n20003) );
  NOR2_X1 U12528 ( .A1(n15316), .A2(n15315), .ZN(n15317) );
  AND2_X1 U12529 ( .A1(n14658), .A2(n14880), .ZN(n11068) );
  AND2_X1 U12530 ( .A1(n13766), .A2(n13765), .ZN(n11069) );
  AND2_X1 U12531 ( .A1(n11385), .A2(n11387), .ZN(n11070) );
  AND2_X1 U12532 ( .A1(n11179), .A2(n11178), .ZN(n11071) );
  AND2_X1 U12533 ( .A1(n16336), .A2(n16181), .ZN(n11072) );
  INV_X1 U12534 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16735) );
  INV_X1 U12535 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18711) );
  OR3_X1 U12536 ( .A1(n11059), .A2(n15465), .A3(n11220), .ZN(n11073) );
  NOR2_X1 U12537 ( .A1(n18192), .A2(n11542), .ZN(n11074) );
  AND2_X1 U12538 ( .A1(n11253), .A2(n11261), .ZN(n11075) );
  INV_X1 U12539 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17406) );
  INV_X1 U12540 ( .A(n11977), .ZN(n15787) );
  NAND3_X1 U12541 ( .A1(n11877), .A2(n11874), .A3(n12400), .ZN(n12251) );
  NOR2_X1 U12542 ( .A1(n15355), .A2(n15354), .ZN(n11076) );
  NOR2_X1 U12543 ( .A1(n15045), .A2(n15046), .ZN(n14896) );
  INV_X1 U12544 ( .A(n20509), .ZN(n11285) );
  NAND2_X1 U12545 ( .A1(n11249), .A2(n11250), .ZN(n15146) );
  NAND2_X1 U12546 ( .A1(n11184), .A2(n11182), .ZN(n15384) );
  OR2_X1 U12547 ( .A1(n11225), .A2(n11224), .ZN(n11077) );
  NOR2_X1 U12548 ( .A1(n15040), .A2(n11268), .ZN(n15058) );
  AND2_X1 U12549 ( .A1(n11274), .A2(n11272), .ZN(n14823) );
  NAND2_X1 U12550 ( .A1(n12300), .A2(n12299), .ZN(n15071) );
  OR2_X1 U12551 ( .A1(n12357), .A2(n12442), .ZN(n11078) );
  INV_X1 U12552 ( .A(n18666), .ZN(n18685) );
  NAND2_X1 U12553 ( .A1(n12933), .A2(n12632), .ZN(n18666) );
  NAND2_X1 U12554 ( .A1(n16411), .A2(n11302), .ZN(n15277) );
  AND2_X1 U12555 ( .A1(n16403), .A2(n11298), .ZN(n11079) );
  NAND2_X1 U12556 ( .A1(n21737), .A2(n21935), .ZN(n15814) );
  INV_X1 U12557 ( .A(n15814), .ZN(n11315) );
  AND2_X1 U12558 ( .A1(n12539), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11080) );
  NAND2_X1 U12559 ( .A1(n22167), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14045) );
  INV_X1 U12560 ( .A(n14045), .ZN(n14229) );
  OR2_X1 U12561 ( .A1(n20571), .A2(n20573), .ZN(n11081) );
  NAND2_X1 U12562 ( .A1(n11311), .A2(n11312), .ZN(n14866) );
  NOR2_X1 U12563 ( .A1(n18226), .A2(n11534), .ZN(n11082) );
  NOR2_X1 U12564 ( .A1(n21194), .A2(n21052), .ZN(n11083) );
  INV_X1 U12565 ( .A(n15425), .ZN(n11235) );
  BUF_X1 U12566 ( .A(n13500), .Z(n21737) );
  INV_X1 U12567 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n17186) );
  AND2_X1 U12568 ( .A1(n11190), .A2(n11189), .ZN(n11084) );
  INV_X1 U12569 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16679) );
  OR2_X1 U12570 ( .A1(n15248), .A2(n11165), .ZN(n11170) );
  AND2_X1 U12571 ( .A1(n11254), .A2(n11252), .ZN(n11085) );
  AND2_X1 U12572 ( .A1(n11187), .A2(n11188), .ZN(n11086) );
  INV_X1 U12573 ( .A(n11261), .ZN(n11257) );
  NAND2_X1 U12574 ( .A1(n13146), .A2(n19642), .ZN(n11261) );
  OR2_X1 U12575 ( .A1(n21236), .A2(n21237), .ZN(n11087) );
  AND2_X1 U12576 ( .A1(n12667), .A2(n11233), .ZN(n11088) );
  AND2_X1 U12577 ( .A1(n11228), .A2(n11227), .ZN(n11089) );
  AND2_X1 U12578 ( .A1(n11276), .A2(n11275), .ZN(n11090) );
  INV_X1 U12579 ( .A(n21732), .ZN(n20022) );
  AND2_X1 U12580 ( .A1(n14532), .A2(n21896), .ZN(n21732) );
  OR2_X1 U12581 ( .A1(n12357), .A2(n12509), .ZN(n11091) );
  NAND2_X1 U12582 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14557) );
  AND2_X1 U12583 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14941) );
  AND2_X1 U12584 ( .A1(n12539), .A2(n12635), .ZN(n11092) );
  AND2_X1 U12585 ( .A1(n13470), .A2(n14707), .ZN(n14661) );
  INV_X1 U12586 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11139) );
  AND2_X1 U12587 ( .A1(n12856), .A2(n12855), .ZN(n16569) );
  INV_X1 U12588 ( .A(n16569), .ZN(n11226) );
  INV_X1 U12589 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20918) );
  AND3_X1 U12590 ( .A1(n16276), .A2(n16122), .A3(n16253), .ZN(n11094) );
  NAND2_X1 U12591 ( .A1(n14553), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21731)
         );
  INV_X1 U12592 ( .A(n21731), .ZN(n21730) );
  AND2_X1 U12593 ( .A1(n11171), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n11095) );
  OR2_X1 U12594 ( .A1(n21251), .A2(n17883), .ZN(n11096) );
  OR2_X1 U12595 ( .A1(n16296), .A2(n13749), .ZN(n11097) );
  OR2_X1 U12596 ( .A1(n16242), .A2(n13750), .ZN(n11098) );
  AND2_X1 U12597 ( .A1(n16912), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11099) );
  AND2_X1 U12598 ( .A1(n11558), .A2(n11217), .ZN(n11100) );
  INV_X1 U12599 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11299) );
  INV_X1 U12600 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n17883) );
  AND2_X1 U12601 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n11101) );
  AND2_X1 U12602 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11102) );
  INV_X1 U12603 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11301) );
  AND2_X1 U12604 ( .A1(n11101), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n11103) );
  INV_X1 U12605 ( .A(n22064), .ZN(n11104) );
  INV_X1 U12606 ( .A(n11104), .ZN(n11105) );
  OAI22_X2 U12607 ( .A1(n22119), .A2(n22219), .B1(n22118), .B2(n22217), .ZN(
        n22160) );
  NOR3_X2 U12608 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21239), .A3(
        n18778), .ZN(n19119) );
  NOR3_X2 U12609 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21239), .A3(
        n18821), .ZN(n19165) );
  OAI22_X2 U12610 ( .A1(n21747), .A2(n22219), .B1(n21746), .B2(n22217), .ZN(
        n21929) );
  INV_X1 U12611 ( .A(n11106), .ZN(n21972) );
  NOR2_X1 U12612 ( .A1(n21936), .A2(n22217), .ZN(n11107) );
  NOR2_X1 U12613 ( .A1(n21937), .A2(n22219), .ZN(n11108) );
  NOR2_X1 U12614 ( .A1(n11107), .A2(n11108), .ZN(n11106) );
  NAND2_X1 U12615 ( .A1(n21732), .A2(n21730), .ZN(n22219) );
  NOR3_X2 U12616 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21239), .A3(
        n18803), .ZN(n19142) );
  OAI21_X2 U12617 ( .B1(n11112), .B2(n11111), .A(n11109), .ZN(n17398) );
  NAND2_X1 U12618 ( .A1(n15155), .A2(n15156), .ZN(n11112) );
  XNOR2_X2 U12619 ( .A(n11374), .B(n13286), .ZN(n16643) );
  NAND2_X1 U12620 ( .A1(n11895), .A2(n11896), .ZN(n11118) );
  NOR2_X1 U12621 ( .A1(n17066), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11119) );
  AND2_X1 U12622 ( .A1(n11014), .A2(n11969), .ZN(n12763) );
  NAND4_X1 U12623 ( .A1(n11885), .A2(n13256), .A3(n11121), .A4(n11122), .ZN(
        n11120) );
  NAND3_X1 U12624 ( .A1(n12634), .A2(n14840), .A3(n12627), .ZN(n11123) );
  XNOR2_X2 U12625 ( .A(n11141), .B(n12259), .ZN(n14819) );
  NAND2_X2 U12626 ( .A1(n11928), .A2(n11927), .ZN(n11141) );
  NAND3_X1 U12627 ( .A1(n12090), .A2(n12058), .A3(n12535), .ZN(n11124) );
  XNOR2_X2 U12628 ( .A(n11125), .B(n13593), .ZN(n21771) );
  OAI21_X2 U12629 ( .B1(n13554), .B2(n13551), .A(n13553), .ZN(n11125) );
  NAND2_X2 U12630 ( .A1(n11126), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13554) );
  NAND2_X1 U12631 ( .A1(n11381), .A2(n20002), .ZN(n20009) );
  NAND2_X1 U12632 ( .A1(n14871), .A2(n14870), .ZN(n14872) );
  NAND2_X2 U12633 ( .A1(n16107), .A2(n13759), .ZN(n16102) );
  NOR2_X2 U12634 ( .A1(n14558), .A2(n11429), .ZN(n17859) );
  NAND2_X2 U12635 ( .A1(n11421), .A2(n11420), .ZN(n14558) );
  INV_X2 U12636 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11420) );
  INV_X2 U12637 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11421) );
  OR2_X2 U12638 ( .A1(n20799), .A2(n11702), .ZN(n20803) );
  OR2_X2 U12639 ( .A1(n20802), .A2(n20820), .ZN(n20799) );
  NAND3_X1 U12640 ( .A1(n21255), .A2(n21235), .A3(n11087), .ZN(n21245) );
  NAND3_X1 U12641 ( .A1(n11135), .A2(n11883), .A3(n11138), .ZN(n11896) );
  NAND2_X1 U12642 ( .A1(n11141), .A2(n12259), .ZN(n11274) );
  NAND2_X1 U12643 ( .A1(n11143), .A2(n12024), .ZN(n12056) );
  NAND3_X1 U12644 ( .A1(n11346), .A2(n11143), .A3(n11345), .ZN(n12090) );
  NAND3_X1 U12645 ( .A1(n11346), .A2(n11143), .A3(n11344), .ZN(n12134) );
  NAND2_X2 U12646 ( .A1(n11046), .A2(n11025), .ZN(n11143) );
  OAI211_X2 U12647 ( .C1(n11350), .C2(n12182), .A(n11348), .B(n12206), .ZN(
        n16776) );
  NAND2_X1 U12648 ( .A1(n12137), .A2(n12389), .ZN(n11152) );
  NAND2_X1 U12649 ( .A1(n12171), .A2(n17400), .ZN(n12179) );
  NAND4_X1 U12650 ( .A1(n11347), .A2(n13354), .A3(n12512), .A4(n12525), .ZN(
        n12532) );
  INV_X1 U12651 ( .A(n12402), .ZN(n11155) );
  NAND2_X1 U12652 ( .A1(n11155), .A2(n11156), .ZN(n12423) );
  NAND3_X1 U12653 ( .A1(n13453), .A2(n13452), .A3(n13454), .ZN(n11164) );
  INV_X1 U12654 ( .A(n11170), .ZN(n21433) );
  AND2_X2 U12655 ( .A1(n11176), .A2(n14763), .ZN(n13443) );
  AND2_X2 U12656 ( .A1(n13797), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11176) );
  XNOR2_X1 U12657 ( .A(n11177), .B(n14705), .ZN(n14720) );
  INV_X1 U12658 ( .A(n11181), .ZN(n15954) );
  NAND3_X1 U12659 ( .A1(n11185), .A2(n15821), .A3(n11048), .ZN(P1_U2810) );
  XNOR2_X1 U12660 ( .A(n15736), .B(n15735), .ZN(n16170) );
  NAND3_X1 U12661 ( .A1(n11188), .A2(n11187), .A3(n15151), .ZN(n19973) );
  INV_X1 U12662 ( .A(n18262), .ZN(n11200) );
  NAND3_X1 U12663 ( .A1(n11198), .A2(n11201), .A3(n11195), .ZN(n18250) );
  NAND3_X1 U12664 ( .A1(n11198), .A2(n11196), .A3(n11195), .ZN(n11202) );
  NAND2_X1 U12665 ( .A1(n11200), .A2(n11199), .ZN(n11198) );
  NOR2_X1 U12666 ( .A1(n18262), .A2(n11524), .ZN(n11527) );
  NAND2_X1 U12667 ( .A1(n11524), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11201) );
  INV_X1 U12668 ( .A(n11202), .ZN(n18248) );
  INV_X1 U12669 ( .A(n18201), .ZN(n11206) );
  INV_X1 U12670 ( .A(n11544), .ZN(n11207) );
  INV_X1 U12671 ( .A(n18213), .ZN(n11210) );
  INV_X1 U12672 ( .A(n17955), .ZN(n11211) );
  NAND3_X1 U12673 ( .A1(n11211), .A2(n11216), .A3(n11100), .ZN(n11218) );
  NAND3_X1 U12674 ( .A1(n11555), .A2(n11214), .A3(n11213), .ZN(n11212) );
  NAND2_X1 U12675 ( .A1(n11555), .A2(n17985), .ZN(n18024) );
  INV_X1 U12676 ( .A(n16916), .ZN(n11221) );
  NAND2_X1 U12677 ( .A1(n15323), .A2(n11232), .ZN(n15412) );
  NAND2_X1 U12678 ( .A1(n15425), .A2(n11236), .ZN(n16945) );
  INV_X1 U12679 ( .A(n16945), .ZN(n12789) );
  INV_X1 U12680 ( .A(n11809), .ZN(n11245) );
  NAND2_X1 U12681 ( .A1(n12635), .A2(n12894), .ZN(n11884) );
  NAND3_X1 U12682 ( .A1(n11807), .A2(n11805), .A3(n11806), .ZN(n11248) );
  INV_X1 U12683 ( .A(n15188), .ZN(n11249) );
  INV_X1 U12684 ( .A(n15040), .ZN(n11265) );
  NAND2_X1 U12685 ( .A1(n11265), .A2(n11266), .ZN(n15072) );
  NAND2_X1 U12686 ( .A1(n11274), .A2(n11271), .ZN(n15045) );
  NAND2_X1 U12687 ( .A1(n20464), .A2(n20523), .ZN(n20465) );
  NAND2_X1 U12688 ( .A1(n20454), .A2(n20523), .ZN(n20455) );
  INV_X1 U12689 ( .A(n11281), .ZN(n20543) );
  INV_X1 U12690 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11288) );
  NAND3_X1 U12691 ( .A1(n20581), .A2(n11293), .A3(n11057), .ZN(n11292) );
  NAND2_X1 U12692 ( .A1(n16430), .A2(n15429), .ZN(n11297) );
  NAND3_X1 U12693 ( .A1(n11310), .A2(n11308), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15286) );
  NAND3_X1 U12694 ( .A1(n11310), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n15282) );
  NAND4_X1 U12695 ( .A1(n14780), .A2(n11311), .A3(n14779), .A4(n11312), .ZN(
        n14865) );
  NAND3_X1 U12696 ( .A1(n13975), .A2(n13976), .A3(n11314), .ZN(n14757) );
  NAND3_X1 U12697 ( .A1(n11316), .A2(n14748), .A3(n17186), .ZN(n13616) );
  NAND2_X1 U12698 ( .A1(n15586), .A2(n11319), .ZN(n15946) );
  CLKBUF_X1 U12699 ( .A(n15586), .Z(n11318) );
  NAND2_X1 U12700 ( .A1(n15831), .A2(n15833), .ZN(n15832) );
  NAND2_X1 U12701 ( .A1(n15831), .A2(n11320), .ZN(n11324) );
  XNOR2_X1 U12702 ( .A(n12390), .B(n18693), .ZN(n17397) );
  NOR2_X2 U12703 ( .A1(n11330), .A2(n11958), .ZN(n12098) );
  NOR2_X2 U12704 ( .A1(n11330), .A2(n11955), .ZN(n12104) );
  NOR2_X2 U12705 ( .A1(n11330), .A2(n11961), .ZN(n12105) );
  NAND2_X1 U12706 ( .A1(n11331), .A2(n16635), .ZN(n16623) );
  NAND3_X1 U12707 ( .A1(n11333), .A2(n11332), .A3(n11334), .ZN(n11331) );
  NAND2_X1 U12708 ( .A1(n12599), .A2(n11342), .ZN(n12628) );
  NAND4_X1 U12709 ( .A1(n13272), .A2(n15019), .A3(n12895), .A4(n12539), .ZN(
        n11342) );
  AND2_X2 U12710 ( .A1(n11880), .A2(n12600), .ZN(n12895) );
  NAND2_X2 U12711 ( .A1(n11045), .A2(n10961), .ZN(n11346) );
  NAND2_X1 U12712 ( .A1(n11346), .A2(n12055), .ZN(n12057) );
  NAND2_X1 U12713 ( .A1(n11347), .A2(n12512), .ZN(n16590) );
  NAND2_X1 U12714 ( .A1(n15566), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15567) );
  NAND2_X1 U12715 ( .A1(n15566), .A2(n11349), .ZN(n11348) );
  INV_X1 U12716 ( .A(n17021), .ZN(n11350) );
  NAND3_X1 U12717 ( .A1(n12090), .A2(n12058), .A3(n15160), .ZN(n15161) );
  NAND2_X1 U12718 ( .A1(n11356), .A2(n11355), .ZN(n15174) );
  INV_X1 U12719 ( .A(n15160), .ZN(n11355) );
  NAND2_X1 U12720 ( .A1(n16764), .A2(n11099), .ZN(n16705) );
  AND2_X2 U12721 ( .A1(n16692), .A2(n11102), .ZN(n16684) );
  NAND2_X1 U12722 ( .A1(n20974), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17889) );
  NAND2_X1 U12723 ( .A1(n11366), .A2(n11365), .ZN(n11677) );
  AOI22_X1 U12724 ( .A1(n19226), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12098), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U12725 ( .A1(n19226), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n19259), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12026) );
  NOR2_X4 U12726 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11970) );
  INV_X4 U12727 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n17066) );
  OAI21_X2 U12728 ( .B1(n12411), .B2(n12419), .A(n11371), .ZN(n16732) );
  NAND3_X1 U12729 ( .A1(n15564), .A2(n12420), .A3(n15565), .ZN(n11371) );
  NAND2_X1 U12730 ( .A1(n11055), .A2(n11868), .ZN(n11870) );
  AND2_X2 U12731 ( .A1(n11855), .A2(n11854), .ZN(n11868) );
  AOI21_X2 U12732 ( .B1(n16643), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11372), .ZN(n13290) );
  NAND2_X1 U12733 ( .A1(n13282), .A2(n11377), .ZN(n16673) );
  NAND2_X1 U12734 ( .A1(n16673), .A2(n13283), .ZN(n13284) );
  NOR2_X4 U12735 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14915) );
  NAND2_X1 U12736 ( .A1(n13469), .A2(n13468), .ZN(n13857) );
  NAND3_X1 U12737 ( .A1(n13494), .A2(n21935), .A3(n13483), .ZN(n13854) );
  NAND2_X1 U12738 ( .A1(n14505), .A2(n13491), .ZN(n13856) );
  INV_X1 U12739 ( .A(n13554), .ZN(n13597) );
  XNOR2_X1 U12740 ( .A(n13558), .B(n13512), .ZN(n14037) );
  OAI21_X2 U12741 ( .B1(n13554), .B2(n13797), .A(n13499), .ZN(n13558) );
  NAND2_X1 U12742 ( .A1(n15527), .A2(n13743), .ZN(n11384) );
  NAND2_X1 U12743 ( .A1(n16135), .A2(n11021), .ZN(n11389) );
  INV_X1 U12744 ( .A(n15179), .ZN(n14082) );
  NAND2_X1 U12745 ( .A1(n14865), .A2(n14044), .ZN(n15065) );
  CLKBUF_X1 U12746 ( .A(n15203), .Z(n15347) );
  AND3_X1 U12747 ( .A1(n11816), .A2(n11815), .A3(n11814), .ZN(n11817) );
  INV_X1 U12748 ( .A(n15792), .ZN(n13082) );
  NAND2_X1 U12749 ( .A1(n15123), .A2(n15178), .ZN(n15179) );
  NAND2_X1 U12750 ( .A1(n11936), .A2(n11935), .ZN(n11928) );
  AOI22_X1 U12751 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19333), .B1(
        n15140), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11967) );
  NAND2_X2 U12752 ( .A1(n12906), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12274) );
  AND2_X1 U12753 ( .A1(n13187), .A2(n13208), .ZN(n11393) );
  INV_X1 U12754 ( .A(n11509), .ZN(n11641) );
  CLKBUF_X3 U12755 ( .A(n11510), .Z(n17838) );
  AND4_X1 U12756 ( .A1(n11867), .A2(n12635), .A3(n17083), .A4(n12400), .ZN(
        n11395) );
  AND2_X1 U12757 ( .A1(n15722), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11396) );
  OR2_X1 U12758 ( .A1(n13317), .A2(n18662), .ZN(n11397) );
  NAND2_X1 U12759 ( .A1(n12933), .A2(n12886), .ZN(n18662) );
  INV_X1 U12760 ( .A(n18662), .ZN(n12928) );
  OR2_X1 U12761 ( .A1(n13332), .A2(n18688), .ZN(n11398) );
  AND2_X1 U12762 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11399) );
  OR2_X1 U12763 ( .A1(n13332), .A2(n17408), .ZN(n11400) );
  AND2_X1 U12764 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11401) );
  AND2_X1 U12765 ( .A1(n12601), .A2(n12635), .ZN(n11402) );
  INV_X1 U12766 ( .A(n14038), .ZN(n14081) );
  INV_X1 U12767 ( .A(n17411), .ZN(n12546) );
  NOR2_X1 U12768 ( .A1(n12549), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11403) );
  NAND2_X1 U12769 ( .A1(n18076), .A2(n18280), .ZN(n18117) );
  INV_X1 U12770 ( .A(n12586), .ZN(n12223) );
  INV_X2 U12771 ( .A(n19083), .ZN(n19082) );
  AND2_X1 U12772 ( .A1(n13117), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11404) );
  INV_X2 U12773 ( .A(n17878), .ZN(n17872) );
  NAND2_X1 U12774 ( .A1(n17893), .A2(n11538), .ZN(n18190) );
  INV_X2 U12775 ( .A(n16473), .ZN(n16513) );
  NAND2_X1 U12776 ( .A1(n12851), .A2(n12850), .ZN(n11405) );
  INV_X1 U12777 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11525) );
  OAI21_X1 U12778 ( .B1(n13269), .B2(n13268), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14617) );
  OR2_X1 U12779 ( .A1(n14006), .A2(n16042), .ZN(n11406) );
  OR2_X1 U12780 ( .A1(n18525), .A2(n18527), .ZN(n11407) );
  INV_X1 U12781 ( .A(n12647), .ZN(n12679) );
  INV_X1 U12782 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12524) );
  OR3_X1 U12783 ( .A1(n17191), .A2(n13783), .A3(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11408) );
  INV_X1 U12784 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13778) );
  INV_X2 U12785 ( .A(n17499), .ZN(n17495) );
  INV_X1 U12786 ( .A(n19979), .ZN(n19985) );
  NAND2_X1 U12787 ( .A1(n19989), .A2(n13429), .ZN(n19979) );
  AND2_X1 U12788 ( .A1(n13287), .A2(n12493), .ZN(n11409) );
  NAND2_X1 U12789 ( .A1(n21917), .A2(n21900), .ZN(n17185) );
  INV_X1 U12790 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11522) );
  AND2_X1 U12791 ( .A1(n12568), .A2(n13309), .ZN(n11410) );
  NAND3_X1 U12792 ( .A1(n12788), .A2(n12787), .A3(n12786), .ZN(n11411) );
  OR2_X1 U12793 ( .A1(n13052), .A2(n13051), .ZN(n11412) );
  INV_X1 U12794 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14986) );
  OR2_X1 U12795 ( .A1(n12987), .A2(n12986), .ZN(n11413) );
  AND2_X1 U12796 ( .A1(n16432), .A2(n12336), .ZN(n11414) );
  AND4_X1 U12797 ( .A1(n12110), .A2(n12109), .A3(n12108), .A4(n12107), .ZN(
        n11415) );
  AND4_X1 U12798 ( .A1(n12103), .A2(n12102), .A3(n12101), .A4(n12100), .ZN(
        n11416) );
  INV_X1 U12799 ( .A(n12393), .ZN(n12170) );
  AND4_X1 U12800 ( .A1(n13427), .A2(n13426), .A3(n13425), .A4(n13424), .ZN(
        n11419) );
  INV_X1 U12801 ( .A(n13475), .ZN(n13486) );
  INV_X1 U12802 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11768) );
  INV_X1 U12803 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13370) );
  INV_X1 U12804 ( .A(n13968), .ZN(n13429) );
  OR2_X1 U12805 ( .A1(n15871), .A2(n15869), .ZN(n14205) );
  INV_X1 U12806 ( .A(n13444), .ZN(n14396) );
  OR2_X1 U12807 ( .A1(n13684), .A2(n13683), .ZN(n13715) );
  NAND2_X1 U12808 ( .A1(n22117), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13800) );
  OR2_X1 U12809 ( .A1(n13706), .A2(n13705), .ZN(n13727) );
  OR2_X1 U12810 ( .A1(n13662), .A2(n13661), .ZN(n13666) );
  AOI22_X1 U12811 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13604), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13392) );
  OR2_X1 U12812 ( .A1(n13570), .A2(n13569), .ZN(n13584) );
  AND2_X1 U12813 ( .A1(n12241), .A2(n12240), .ZN(n12582) );
  NAND2_X1 U12814 ( .A1(n15291), .A2(n12663), .ZN(n12222) );
  INV_X1 U12815 ( .A(n12233), .ZN(n12675) );
  OAI21_X1 U12816 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20813), .A(
        n11717), .ZN(n11718) );
  AOI22_X1 U12817 ( .A1(n13514), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13443), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13426) );
  AND4_X1 U12818 ( .A1(n13449), .A2(n13448), .A3(n13447), .A4(n13446), .ZN(
        n13455) );
  INV_X1 U12819 ( .A(n15585), .ZN(n14234) );
  NOR2_X1 U12820 ( .A1(n16147), .A2(n13746), .ZN(n13747) );
  OAI22_X1 U12821 ( .A1(n14027), .A2(n13663), .B1(n13806), .B2(n13687), .ZN(
        n13673) );
  AND2_X1 U12822 ( .A1(n13800), .A2(n13491), .ZN(n13792) );
  OR2_X1 U12823 ( .A1(n13755), .A2(n13923), .ZN(n13753) );
  AOI22_X1 U12824 ( .A1(n13514), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13382) );
  INV_X1 U12825 ( .A(n16433), .ZN(n12336) );
  AND2_X1 U12826 ( .A1(n12651), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12941) );
  NAND2_X1 U12827 ( .A1(n17400), .A2(n12180), .ZN(n12181) );
  NAND2_X1 U12828 ( .A1(n11934), .A2(n11933), .ZN(n12260) );
  AND2_X1 U12829 ( .A1(n12218), .A2(n12217), .ZN(n12579) );
  INV_X1 U12830 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11832) );
  NAND2_X1 U12831 ( .A1(n11458), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11474) );
  INV_X1 U12832 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11543) );
  AND2_X1 U12833 ( .A1(n18189), .A2(n11543), .ZN(n11542) );
  AOI22_X1 U12834 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13423) );
  INV_X1 U12835 ( .A(n15458), .ZN(n14127) );
  NOR2_X1 U12836 ( .A1(n14453), .A2(n16065), .ZN(n14454) );
  OR2_X1 U12837 ( .A1(n21491), .A2(n17185), .ZN(n14271) );
  AND2_X1 U12838 ( .A1(n13786), .A2(n13491), .ZN(n13821) );
  OAI221_X1 U12839 ( .B1(n13783), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .C1(n13783), .C2(n17191), .A(n13780), .ZN(n13825) );
  OR2_X1 U12840 ( .A1(n13639), .A2(n13638), .ZN(n13664) );
  NAND2_X1 U12841 ( .A1(n11773), .A2(n11832), .ZN(n11780) );
  INV_X1 U12842 ( .A(n12585), .ZN(n12244) );
  AND2_X1 U12843 ( .A1(n13188), .A2(n11393), .ZN(n13189) );
  INV_X1 U12844 ( .A(n13022), .ZN(n13112) );
  INV_X1 U12845 ( .A(n12892), .ZN(n12890) );
  INV_X1 U12846 ( .A(n11915), .ZN(n11916) );
  AND2_X1 U12847 ( .A1(n11902), .A2(n11901), .ZN(n11903) );
  INV_X1 U12848 ( .A(n15488), .ZN(n12320) );
  AND3_X1 U12849 ( .A1(n12807), .A2(n12806), .A3(n12805), .ZN(n16932) );
  OAI21_X1 U12850 ( .B1(n10991), .B2(n12176), .A(n12175), .ZN(n12177) );
  NAND2_X1 U12851 ( .A1(n14986), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12656) );
  NAND2_X1 U12852 ( .A1(n12936), .A2(n12654), .ZN(n12953) );
  INV_X1 U12853 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17695) );
  INV_X1 U12854 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17730) );
  AND2_X1 U12855 ( .A1(n17936), .A2(n20952), .ZN(n11545) );
  NOR2_X1 U12856 ( .A1(n18189), .A2(n11543), .ZN(n11544) );
  INV_X1 U12857 ( .A(n20774), .ZN(n11680) );
  INV_X1 U12858 ( .A(n14081), .ZN(n14502) );
  NAND2_X1 U12859 ( .A1(n14454), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14509) );
  OR2_X1 U12860 ( .A1(n21543), .A2(n17185), .ZN(n14354) );
  NOR2_X1 U12861 ( .A1(n14265), .A2(n21478), .ZN(n14266) );
  INV_X1 U12862 ( .A(n21915), .ZN(n21904) );
  INV_X1 U12863 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21900) );
  AND2_X1 U12864 ( .A1(n12858), .A2(n12857), .ZN(n16562) );
  INV_X1 U12865 ( .A(n15041), .ZN(n12290) );
  INV_X1 U12866 ( .A(n15073), .ZN(n12299) );
  OR2_X1 U12867 ( .A1(n11881), .A2(n12627), .ZN(n12884) );
  NAND2_X1 U12868 ( .A1(n15287), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15281) );
  INV_X1 U12869 ( .A(n12926), .ZN(n12927) );
  NAND2_X1 U12870 ( .A1(n15398), .A2(n15371), .ZN(n15370) );
  AND2_X1 U12871 ( .A1(n12203), .A2(n12202), .ZN(n12535) );
  INV_X1 U12872 ( .A(n12358), .ZN(n12060) );
  AND3_X1 U12873 ( .A1(n12674), .A2(n12673), .A3(n12672), .ZN(n15165) );
  INV_X1 U12874 ( .A(n21236), .ZN(n11659) );
  AOI22_X1 U12875 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11582) );
  AND2_X1 U12876 ( .A1(n17960), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11556) );
  AND2_X1 U12877 ( .A1(n11535), .A2(n20629), .ZN(n11538) );
  INV_X1 U12878 ( .A(n20962), .ZN(n20958) );
  INV_X1 U12879 ( .A(n20943), .ZN(n21188) );
  NOR3_X1 U12880 ( .A1(n11665), .A2(n11732), .A3(n20801), .ZN(n15623) );
  INV_X1 U12881 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15886) );
  AND2_X1 U12882 ( .A1(n15250), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15251) );
  AND2_X1 U12883 ( .A1(n13929), .A2(n13928), .ZN(n15953) );
  OR2_X1 U12884 ( .A1(n14879), .A2(n14878), .ZN(n14881) );
  AND2_X1 U12885 ( .A1(n14355), .A2(n14354), .ZN(n15926) );
  OR2_X1 U12886 ( .A1(n15970), .A2(n15971), .ZN(n15968) );
  NOR2_X1 U12887 ( .A1(n14219), .A2(n14220), .ZN(n14206) );
  NOR2_X1 U12888 ( .A1(n14097), .A2(n15532), .ZN(n14111) );
  INV_X1 U12889 ( .A(n14075), .ZN(n14016) );
  NAND2_X1 U12890 ( .A1(n21574), .A2(n14534), .ZN(n16164) );
  OR2_X1 U12891 ( .A1(n21289), .A2(n15556), .ZN(n15536) );
  NAND2_X1 U12892 ( .A1(n13986), .A2(n17152), .ZN(n16365) );
  OAI21_X1 U12893 ( .B1(n21586), .B2(n14924), .A(n16380), .ZN(n21735) );
  AND2_X1 U12894 ( .A1(n14746), .A2(n14745), .ZN(n17161) );
  NOR2_X1 U12895 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21868) );
  AND2_X1 U12896 ( .A1(n13599), .A2(n13625), .ZN(n21738) );
  INV_X1 U12897 ( .A(n14035), .ZN(n21750) );
  INV_X1 U12898 ( .A(n15264), .ZN(n21903) );
  NAND2_X1 U12899 ( .A1(n21736), .A2(n21735), .ZN(n22215) );
  INV_X1 U12900 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16379) );
  INV_X1 U12901 ( .A(n14962), .ZN(n15010) );
  INV_X1 U12902 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16447) );
  AND2_X1 U12903 ( .A1(n12243), .A2(n12594), .ZN(n15004) );
  AND2_X1 U12904 ( .A1(n18371), .A2(n15291), .ZN(n15299) );
  AND2_X1 U12905 ( .A1(n19686), .A2(n13272), .ZN(n19188) );
  INV_X1 U12906 ( .A(n13352), .ZN(n13351) );
  NOR2_X1 U12907 ( .A1(n16587), .A2(n16601), .ZN(n12512) );
  NAND2_X1 U12908 ( .A1(n12208), .A2(n12207), .ZN(n12211) );
  NAND2_X1 U12909 ( .A1(n17419), .A2(n18705), .ZN(n15132) );
  AND2_X1 U12910 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19327) );
  AND2_X1 U12911 ( .A1(n19362), .A2(n19346), .ZN(n19361) );
  OR2_X1 U12912 ( .A1(n19431), .A2(n17426), .ZN(n19248) );
  OR2_X1 U12913 ( .A1(n19431), .A2(n19579), .ZN(n19225) );
  INV_X1 U12914 ( .A(n12956), .ZN(n15129) );
  NOR2_X1 U12915 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n20451), .ZN(n20468) );
  INV_X1 U12916 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20401) );
  INV_X1 U12917 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20274) );
  NOR2_X1 U12918 ( .A1(n20737), .A2(n20736), .ZN(n20735) );
  NAND3_X1 U12919 ( .A1(n11650), .A2(n11649), .A3(n11648), .ZN(n20622) );
  INV_X1 U12920 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18135) );
  NOR2_X1 U12921 ( .A1(n18081), .A2(n11743), .ZN(n18053) );
  NAND2_X1 U12922 ( .A1(n17899), .A2(n11556), .ZN(n17955) );
  NOR2_X2 U12923 ( .A1(n20819), .A2(n11749), .ZN(n21146) );
  NAND2_X1 U12924 ( .A1(n20856), .A2(n20625), .ZN(n21137) );
  NOR2_X1 U12925 ( .A1(n18202), .A2(n20918), .ZN(n18201) );
  NAND2_X1 U12926 ( .A1(n20108), .A2(n15623), .ZN(n21172) );
  OAI21_X1 U12927 ( .B1(n21248), .B2(n17885), .A(n20787), .ZN(n18751) );
  INV_X1 U12928 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18796) );
  AND2_X1 U12929 ( .A1(n21205), .A2(n15623), .ZN(n15643) );
  NOR2_X1 U12930 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21586) );
  INV_X1 U12931 ( .A(n21553), .ZN(n21568) );
  INV_X1 U12932 ( .A(n19989), .ZN(n17196) );
  AND2_X1 U12933 ( .A1(n15616), .A2(n21730), .ZN(n16030) );
  NAND2_X1 U12934 ( .A1(n14881), .A2(n14880), .ZN(n15655) );
  AND2_X1 U12935 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n14016), .ZN(
        n14074) );
  INV_X1 U12936 ( .A(n16164), .ZN(n20038) );
  OR2_X1 U12937 ( .A1(n13772), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13773) );
  AND2_X1 U12938 ( .A1(n13948), .A2(n13947), .ZN(n15922) );
  AND2_X1 U12939 ( .A1(n16280), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16277) );
  NAND2_X1 U12940 ( .A1(n13850), .A2(n13849), .ZN(n13986) );
  NAND2_X1 U12941 ( .A1(n15537), .A2(n15536), .ZN(n21319) );
  AND2_X1 U12942 ( .A1(n13830), .A2(n13491), .ZN(n17152) );
  NOR2_X2 U12943 ( .A1(n21781), .A2(n21867), .ZN(n22227) );
  INV_X1 U12944 ( .A(n22231), .ZN(n22233) );
  NOR2_X2 U12945 ( .A1(n21781), .A2(n21894), .ZN(n22239) );
  NOR2_X2 U12946 ( .A1(n21781), .A2(n21809), .ZN(n22246) );
  OAI211_X1 U12947 ( .C1(n22256), .C2(n21881), .A(n21907), .B(n21806), .ZN(
        n22258) );
  NOR2_X2 U12948 ( .A1(n21810), .A2(n21894), .ZN(n22264) );
  INV_X1 U12949 ( .A(n22268), .ZN(n22271) );
  NOR2_X2 U12950 ( .A1(n21859), .A2(n21891), .ZN(n22282) );
  NOR2_X2 U12951 ( .A1(n21859), .A2(n21894), .ZN(n22289) );
  INV_X1 U12952 ( .A(n22293), .ZN(n22297) );
  NAND2_X1 U12953 ( .A1(n21751), .A2(n14035), .ZN(n21867) );
  NOR2_X2 U12954 ( .A1(n21895), .A2(n21891), .ZN(n22312) );
  NOR2_X1 U12955 ( .A1(n22212), .A2(n21933), .ZN(n21971) );
  AND2_X1 U12956 ( .A1(n21619), .A2(n13457), .ZN(n13828) );
  INV_X1 U12957 ( .A(n22328), .ZN(n19938) );
  INV_X1 U12958 ( .A(n19946), .ZN(n19940) );
  NOR2_X1 U12959 ( .A1(n12614), .A2(n12595), .ZN(n15128) );
  NAND2_X1 U12960 ( .A1(n18616), .A2(n15429), .ZN(n18618) );
  INV_X1 U12961 ( .A(n18627), .ZN(n18639) );
  INV_X1 U12962 ( .A(n18529), .ZN(n18642) );
  INV_X1 U12963 ( .A(n18596), .ZN(n18641) );
  AND2_X1 U12964 ( .A1(n15316), .A2(n12560), .ZN(n15717) );
  INV_X1 U12965 ( .A(n18718), .ZN(n15440) );
  OR2_X1 U12966 ( .A1(n15049), .A2(n14895), .ZN(n15050) );
  OR2_X1 U12967 ( .A1(n14830), .A2(n14829), .ZN(n14831) );
  NOR2_X1 U12968 ( .A1(n12651), .A2(n13211), .ZN(n16484) );
  AND2_X1 U12969 ( .A1(n19188), .A2(n15130), .ZN(n19184) );
  INV_X1 U12970 ( .A(n19220), .ZN(n19419) );
  NAND2_X1 U12971 ( .A1(n19686), .A2(n11092), .ZN(n19189) );
  INV_X1 U12972 ( .A(n14630), .ZN(n14655) );
  INV_X1 U12973 ( .A(n14714), .ZN(n14622) );
  INV_X1 U12974 ( .A(n14617), .ZN(n15130) );
  AND2_X1 U12975 ( .A1(n16396), .A2(n16395), .ZN(n18497) );
  INV_X1 U12976 ( .A(n17417), .ZN(n16750) );
  INV_X1 U12977 ( .A(n18664), .ZN(n13329) );
  INV_X1 U12978 ( .A(n18688), .ZN(n15725) );
  OR2_X1 U12979 ( .A1(n12910), .A2(n12909), .ZN(n16990) );
  INV_X1 U12980 ( .A(n19355), .ZN(n19346) );
  OAI21_X2 U12981 ( .B1(n18706), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15132), 
        .ZN(n19362) );
  OAI21_X1 U12982 ( .B1(n17087), .B2(n17086), .A(n17085), .ZN(n19813) );
  INV_X1 U12983 ( .A(n19807), .ZN(n19811) );
  NOR2_X1 U12984 ( .A1(n19342), .A2(n19325), .ZN(n19617) );
  OAI21_X1 U12985 ( .B1(n17103), .B2(n17107), .A(n17102), .ZN(n19782) );
  INV_X1 U12986 ( .A(n19779), .ZN(n19781) );
  NOR2_X1 U12987 ( .A1(n19298), .A2(n19694), .ZN(n19608) );
  INV_X1 U12988 ( .A(n19760), .ZN(n19763) );
  INV_X1 U12989 ( .A(n19746), .ZN(n19739) );
  INV_X1 U12990 ( .A(n19248), .ZN(n19264) );
  OAI21_X1 U12991 ( .B1(n19254), .B2(n19253), .A(n19252), .ZN(n19727) );
  INV_X1 U12992 ( .A(n19571), .ZN(n19575) );
  INV_X1 U12993 ( .A(n19523), .ZN(n19525) );
  INV_X1 U12994 ( .A(n19677), .ZN(n19679) );
  NAND2_X1 U12995 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n17419) );
  NAND2_X1 U12996 ( .A1(n17496), .A2(n17477), .ZN(n21630) );
  INV_X1 U12997 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n17478) );
  NAND2_X1 U12998 ( .A1(n11666), .A2(n21162), .ZN(n21210) );
  NOR2_X1 U12999 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n20503), .ZN(n20520) );
  NOR2_X1 U13000 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20399), .ZN(n20418) );
  NOR2_X1 U13001 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20316), .ZN(n20332) );
  INV_X1 U13002 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20305) );
  NOR2_X1 U13003 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20226), .ZN(n20248) );
  INV_X1 U13004 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20189) );
  NOR2_X2 U13005 ( .A1(n21246), .A2(n20461), .ZN(n20532) );
  NOR2_X1 U13006 ( .A1(n20448), .A2(n17759), .ZN(n17790) );
  OAI21_X1 U13007 ( .B1(n15643), .B2(n15625), .A(n21235), .ZN(n20594) );
  NOR2_X1 U13008 ( .A1(n11602), .A2(n11601), .ZN(n20653) );
  NOR2_X1 U13009 ( .A1(n20772), .A2(n20773), .ZN(n20616) );
  NAND2_X1 U13010 ( .A1(n20622), .A2(n20621), .ZN(n20777) );
  INV_X1 U13011 ( .A(n19087), .ZN(n20595) );
  NOR2_X1 U13012 ( .A1(n20164), .A2(n20115), .ZN(n20130) );
  INV_X1 U13013 ( .A(n18116), .ZN(n18110) );
  OAI21_X1 U13014 ( .B1(n20169), .B2(n18117), .A(n19083), .ZN(n18074) );
  NAND2_X1 U13015 ( .A1(n18117), .A2(n18116), .ZN(n18253) );
  INV_X1 U13016 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21177) );
  NOR2_X1 U13017 ( .A1(n20928), .A2(n20927), .ZN(n20980) );
  NOR2_X1 U13018 ( .A1(n21194), .A2(n21210), .ZN(n20914) );
  NAND2_X1 U13019 ( .A1(n17883), .A2(n18751), .ZN(n18956) );
  INV_X1 U13020 ( .A(n19067), .ZN(n19178) );
  INV_X1 U13021 ( .A(n19152), .ZN(n19160) );
  INV_X1 U13022 ( .A(n19141), .ZN(n19148) );
  INV_X1 U13023 ( .A(n19112), .ZN(n19126) );
  INV_X1 U13024 ( .A(n19008), .ZN(n19120) );
  INV_X1 U13025 ( .A(n19106), .ZN(n19114) );
  INV_X1 U13026 ( .A(n19183), .ZN(n19092) );
  AND2_X1 U13027 ( .A1(n19084), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19074) );
  INV_X1 U13028 ( .A(n21652), .ZN(n21607) );
  INV_X1 U13029 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21654) );
  INV_X1 U13030 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n21645) );
  INV_X1 U13031 ( .A(n15130), .ZN(n15131) );
  NOR2_X1 U13032 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14556), .ZN(n18745)
         );
  INV_X1 U13033 ( .A(U212), .ZN(n20095) );
  INV_X1 U13034 ( .A(U212), .ZN(n20086) );
  NAND2_X1 U13035 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21614), .ZN(n22329) );
  NOR2_X1 U13036 ( .A1(n14529), .A2(n14528), .ZN(n14530) );
  NAND2_X1 U13037 ( .A1(n14514), .A2(n14513), .ZN(n21553) );
  INV_X1 U13038 ( .A(n21499), .ZN(n16022) );
  OR2_X1 U13039 ( .A1(n15594), .A2(n15593), .ZN(n21464) );
  AND2_X1 U13041 ( .A1(n14887), .A2(n14886), .ZN(n21729) );
  NAND2_X1 U13042 ( .A1(n21664), .A2(n11017), .ZN(n21724) );
  INV_X1 U13043 ( .A(n20033), .ZN(n20043) );
  NAND2_X1 U13044 ( .A1(n13986), .A2(n13859), .ZN(n21339) );
  INV_X1 U13045 ( .A(n21345), .ZN(n21338) );
  INV_X1 U13046 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21875) );
  INV_X1 U13047 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14922) );
  AOI22_X1 U13048 ( .A1(n21743), .A2(n21740), .B1(n21843), .B2(n21745), .ZN(
        n22224) );
  OR2_X1 U13049 ( .A1(n21781), .A2(n21891), .ZN(n22231) );
  AOI22_X1 U13050 ( .A1(n21764), .A2(n21766), .B1(n21801), .B2(n21843), .ZN(
        n22237) );
  INV_X1 U13051 ( .A(n21775), .ZN(n22243) );
  OR2_X1 U13052 ( .A1(n21810), .A2(n21867), .ZN(n22255) );
  AOI22_X1 U13053 ( .A1(n21805), .A2(n21802), .B1(n21801), .B2(n21874), .ZN(
        n22261) );
  OR2_X1 U13054 ( .A1(n21810), .A2(n21809), .ZN(n22268) );
  NAND2_X1 U13055 ( .A1(n21853), .A2(n21822), .ZN(n22280) );
  AOI22_X1 U13056 ( .A1(n21847), .A2(n21844), .B1(n21843), .B2(n21842), .ZN(
        n22286) );
  NAND2_X1 U13057 ( .A1(n21853), .A2(n21852), .ZN(n22293) );
  INV_X1 U13058 ( .A(n21971), .ZN(n21964) );
  INV_X1 U13059 ( .A(n22206), .ZN(n22198) );
  OR2_X1 U13060 ( .A1(n21895), .A2(n21867), .ZN(n22308) );
  OR2_X1 U13061 ( .A1(n21895), .A2(n21894), .ZN(n22326) );
  OR2_X1 U13062 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n13828), .ZN(n21617) );
  OR2_X1 U13063 ( .A1(n22329), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n19946) );
  INV_X1 U13064 ( .A(n15298), .ZN(n14574) );
  INV_X1 U13065 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n21597) );
  INV_X1 U13066 ( .A(n18645), .ZN(n18601) );
  INV_X1 U13067 ( .A(n18644), .ZN(n18638) );
  AND2_X1 U13068 ( .A1(n14812), .A2(n15440), .ZN(n16473) );
  AND2_X1 U13069 ( .A1(n13274), .A2(n13273), .ZN(n13275) );
  NAND2_X1 U13070 ( .A1(n19686), .A2(n13259), .ZN(n19636) );
  NAND2_X2 U13071 ( .A1(n13258), .A2(n13257), .ZN(n19686) );
  AND2_X1 U13072 ( .A1(n19190), .A2(n19189), .ZN(n19697) );
  NAND2_X1 U13073 ( .A1(n17448), .A2(n14717), .ZN(n14862) );
  INV_X1 U13074 ( .A(n17448), .ZN(n17475) );
  NAND2_X1 U13075 ( .A1(n15298), .A2(n19642), .ZN(n14714) );
  AOI21_X1 U13076 ( .B1(n16451), .B2(n16711), .A(n13298), .ZN(n13299) );
  OAI21_X1 U13077 ( .B1(n15728), .B2(n17411), .A(n12565), .ZN(n12566) );
  INV_X1 U13078 ( .A(n16766), .ZN(n17408) );
  NAND2_X1 U13079 ( .A1(n12545), .A2(n12651), .ZN(n17411) );
  XNOR2_X1 U13080 ( .A(n13356), .B(n13355), .ZN(n15758) );
  NOR2_X1 U13081 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  NAND2_X1 U13082 ( .A1(n12933), .A2(n12621), .ZN(n18664) );
  NAND2_X1 U13083 ( .A1(n12933), .A2(n12932), .ZN(n18688) );
  INV_X1 U13084 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18660) );
  AOI21_X1 U13085 ( .B1(n17082), .B2(n17091), .A(n19700), .ZN(n19680) );
  OR2_X1 U13086 ( .A1(n19342), .A2(n17097), .ZN(n19807) );
  INV_X1 U13087 ( .A(n19617), .ZN(n19799) );
  OR2_X1 U13088 ( .A1(n19342), .A2(n19247), .ZN(n19620) );
  AOI21_X1 U13089 ( .B1(n17108), .B2(n17107), .A(n17106), .ZN(n19786) );
  OR2_X1 U13090 ( .A1(n19314), .A2(n17097), .ZN(n19779) );
  OR2_X1 U13091 ( .A1(n19314), .A2(n19341), .ZN(n19613) );
  INV_X1 U13092 ( .A(n19608), .ZN(n19772) );
  NAND2_X1 U13093 ( .A1(n19279), .A2(n19694), .ZN(n19760) );
  NAND2_X1 U13094 ( .A1(n19264), .A2(n15127), .ZN(n19754) );
  NAND2_X1 U13095 ( .A1(n19264), .A2(n15233), .ZN(n19746) );
  NAND2_X1 U13096 ( .A1(n19264), .A2(n19324), .ZN(n19744) );
  INV_X1 U13097 ( .A(n19651), .ZN(n19737) );
  INV_X1 U13098 ( .A(n19810), .ZN(n19800) );
  INV_X1 U13099 ( .A(n19728), .ZN(n19495) );
  AOI22_X1 U13100 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19699), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19698), .ZN(n19517) );
  AOI22_X1 U13101 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19699), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19698), .ZN(n19684) );
  NAND2_X1 U13102 ( .A1(n19223), .A2(n19324), .ZN(n19712) );
  INV_X1 U13103 ( .A(n21600), .ZN(n17132) );
  INV_X1 U13104 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21640) );
  NAND2_X1 U13105 ( .A1(n17478), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n17499) );
  INV_X1 U13106 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21602) );
  OR3_X1 U13107 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n20370), .A3(n20372), .ZN(
        n20364) );
  INV_X1 U13108 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n20309) );
  INV_X1 U13109 ( .A(n20588), .ZN(n20516) );
  AND2_X1 U13110 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17779), .ZN(n17775) );
  NOR2_X1 U13111 ( .A1(n20400), .A2(n17817), .ZN(n17846) );
  INV_X1 U13112 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20251) );
  NOR2_X2 U13113 ( .A1(n17877), .A2(n20768), .ZN(n17878) );
  INV_X1 U13114 ( .A(n20744), .ZN(n20754) );
  INV_X1 U13115 ( .A(n20777), .ZN(n20757) );
  AND2_X1 U13116 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n20616), .ZN(n20619) );
  NOR2_X1 U13117 ( .A1(n11447), .A2(n11446), .ZN(n20633) );
  INV_X1 U13118 ( .A(n20781), .ZN(n20739) );
  NAND2_X1 U13119 ( .A1(n18337), .A2(n20595), .ZN(n18355) );
  INV_X1 U13120 ( .A(n18337), .ZN(n18336) );
  NAND2_X1 U13121 ( .A1(n17893), .A2(n18279), .ZN(n18144) );
  OR2_X1 U13122 ( .A1(n18956), .A2(n18798), .ZN(n19083) );
  NOR2_X1 U13123 ( .A1(n18037), .A2(n11047), .ZN(n11766) );
  OAI21_X1 U13124 ( .B1(n15642), .B2(n11741), .A(n21235), .ZN(n20992) );
  INV_X1 U13125 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21199) );
  INV_X1 U13126 ( .A(n19143), .ZN(n19130) );
  INV_X1 U13127 ( .A(n18791), .ZN(n18836) );
  INV_X1 U13128 ( .A(n18910), .ZN(n18908) );
  INV_X1 U13129 ( .A(n21605), .ZN(n17121) );
  OR2_X1 U13130 ( .A1(n12567), .A2(n12566), .ZN(P2_U2999) );
  NOR3_X2 U13131 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n11428), .ZN(n11510) );
  AOI22_X1 U13132 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17838), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11426) );
  INV_X4 U13133 ( .A(n11641), .ZN(n17824) );
  AOI22_X1 U13134 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U13135 ( .A1(n17832), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11424) );
  BUF_X4 U13136 ( .A(n11458), .Z(n17853) );
  AOI22_X1 U13137 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17833), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11423) );
  NAND4_X1 U13138 ( .A1(n11426), .A2(n11425), .A3(n11424), .A4(n11423), .ZN(
        n11436) );
  AOI22_X1 U13139 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11434) );
  NOR2_X1 U13140 ( .A1(n11428), .A2(n20824), .ZN(n11507) );
  CLKBUF_X3 U13141 ( .A(n11507), .Z(n17849) );
  AOI22_X1 U13142 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U13144 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U13146 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11431) );
  NAND4_X1 U13147 ( .A1(n11434), .A2(n11433), .A3(n11432), .A4(n11431), .ZN(
        n11435) );
  AOI22_X1 U13148 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U13149 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U13150 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U13151 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11438) );
  NAND4_X1 U13152 ( .A1(n11441), .A2(n11440), .A3(n11439), .A4(n11438), .ZN(
        n11447) );
  AOI22_X1 U13153 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17849), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U13154 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U13155 ( .A1(n17861), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11443) );
  BUF_X4 U13156 ( .A(n17859), .Z(n17718) );
  AOI22_X1 U13157 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11442) );
  NAND4_X1 U13158 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11446) );
  AOI22_X1 U13159 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U13160 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U13161 ( .A1(n17832), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U13162 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17833), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11448) );
  NAND4_X1 U13163 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(
        n11457) );
  AOI22_X1 U13164 ( .A1(n17848), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U13165 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17849), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U13166 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17838), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U13167 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11452) );
  NAND4_X1 U13168 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n11456) );
  NOR2_X1 U13169 ( .A1(n11457), .A2(n11456), .ZN(n20642) );
  INV_X1 U13170 ( .A(n20642), .ZN(n11526) );
  AOI22_X1 U13171 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U13172 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11517), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11467) );
  INV_X1 U13173 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17706) );
  AOI22_X1 U13174 ( .A1(n11437), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11469), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11459) );
  OAI21_X1 U13175 ( .B1(n11506), .B2(n17706), .A(n11459), .ZN(n11465) );
  AOI22_X1 U13176 ( .A1(n11510), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11508), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U13177 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U13178 ( .A1(n11560), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11507), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U13179 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11473), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11460) );
  NAND4_X1 U13180 ( .A1(n11463), .A2(n11462), .A3(n11461), .A4(n11460), .ZN(
        n11464) );
  AOI211_X1 U13181 ( .C1(n17853), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n11465), .B(n11464), .ZN(n11466) );
  NAND3_X1 U13182 ( .A1(n11468), .A2(n11467), .A3(n11466), .ZN(n11667) );
  INV_X1 U13183 ( .A(n11667), .ZN(n20651) );
  INV_X1 U13184 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17873) );
  AOI22_X1 U13185 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11437), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n11469), .ZN(n11470) );
  OAI21_X1 U13186 ( .B1(n17873), .B2(n11506), .A(n11470), .ZN(n11471) );
  AOI22_X1 U13187 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11507), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U13188 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11509), .B1(
        n11510), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11472) );
  INV_X1 U13189 ( .A(n11472), .ZN(n11478) );
  AOI22_X1 U13190 ( .A1(n11566), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n11508), .ZN(n11476) );
  AOI22_X1 U13191 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10971), .B1(
        n11473), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11475) );
  NAND3_X1 U13192 ( .A1(n11476), .A2(n11475), .A3(n11474), .ZN(n11477) );
  AOI22_X1 U13193 ( .A1(n11560), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11517), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U13194 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17859), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11482) );
  NAND3_X1 U13195 ( .A1(n11484), .A2(n11483), .A3(n11482), .ZN(n20774) );
  AOI22_X1 U13196 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11494) );
  AOI22_X1 U13197 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17838), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11493) );
  INV_X1 U13198 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17717) );
  AOI22_X1 U13199 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11485) );
  OAI21_X1 U13200 ( .B1(n11506), .B2(n17717), .A(n11485), .ZN(n11491) );
  AOI22_X1 U13201 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U13202 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U13203 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U13204 ( .A1(n17718), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11486) );
  NAND4_X1 U13205 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11490) );
  AOI211_X1 U13206 ( .C1(n17853), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n11491), .B(n11490), .ZN(n11492) );
  NAND3_X1 U13207 ( .A1(n11494), .A2(n11493), .A3(n11492), .ZN(n11673) );
  INV_X1 U13208 ( .A(n11673), .ZN(n20638) );
  AOI22_X1 U13209 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U13210 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U13211 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11495) );
  OAI21_X1 U13212 ( .B1(n11506), .B2(n17730), .A(n11495), .ZN(n11501) );
  AOI22_X1 U13213 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17838), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U13214 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U13215 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11497) );
  AOI22_X1 U13216 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11496) );
  NAND4_X1 U13217 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n11500) );
  AOI211_X1 U13218 ( .C1(n17853), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n11501), .B(n11500), .ZN(n11502) );
  NAND3_X1 U13219 ( .A1(n11504), .A2(n11503), .A3(n11502), .ZN(n20629) );
  INV_X1 U13220 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17902) );
  NAND2_X1 U13221 ( .A1(n18190), .A2(n17902), .ZN(n17900) );
  INV_X1 U13222 ( .A(n17900), .ZN(n17987) );
  NOR2_X1 U13223 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17972) );
  INV_X1 U13224 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n20999) );
  NAND3_X1 U13225 ( .A1(n17987), .A2(n17972), .A3(n20999), .ZN(n17956) );
  NOR2_X1 U13226 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17956), .ZN(
        n18007) );
  INV_X1 U13227 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20891) );
  INV_X1 U13228 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20864) );
  INV_X1 U13229 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17684) );
  AOI22_X1 U13230 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11469), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11505) );
  OAI21_X1 U13231 ( .B1(n11506), .B2(n17684), .A(n11505), .ZN(n11516) );
  AOI22_X1 U13232 ( .A1(n11473), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U13233 ( .A1(n11507), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U13234 ( .A1(n11508), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U13235 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11510), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11511) );
  NAND4_X1 U13236 ( .A1(n11514), .A2(n11513), .A3(n11512), .A4(n11511), .ZN(
        n11515) );
  AOI211_X1 U13237 ( .C1(n17853), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n11516), .B(n11515), .ZN(n11520) );
  AOI22_X1 U13238 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11517), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U13239 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17850), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11518) );
  NOR2_X1 U13240 ( .A1(n18270), .A2(n18278), .ZN(n18269) );
  NOR2_X1 U13241 ( .A1(n20774), .A2(n20864), .ZN(n11521) );
  XNOR2_X1 U13242 ( .A(n11667), .B(n20774), .ZN(n11523) );
  NOR2_X1 U13243 ( .A1(n11522), .A2(n11523), .ZN(n11524) );
  XNOR2_X1 U13244 ( .A(n11526), .B(n11676), .ZN(n18249) );
  XOR2_X1 U13245 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11529), .Z(
        n18234) );
  NOR2_X1 U13246 ( .A1(n18235), .A2(n18234), .ZN(n18233) );
  INV_X1 U13247 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20883) );
  NOR2_X1 U13248 ( .A1(n20883), .A2(n11529), .ZN(n11530) );
  XNOR2_X1 U13249 ( .A(n20633), .B(n11531), .ZN(n11532) );
  NOR2_X1 U13250 ( .A1(n11533), .A2(n11532), .ZN(n11534) );
  INV_X1 U13251 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11698) );
  XOR2_X1 U13252 ( .A(n20629), .B(n11535), .Z(n11536) );
  XOR2_X1 U13253 ( .A(n11698), .B(n11536), .Z(n18213) );
  NOR2_X1 U13254 ( .A1(n18212), .A2(n11537), .ZN(n11539) );
  OAI21_X1 U13255 ( .B1(n11538), .B2(n17893), .A(n18190), .ZN(n11540) );
  XNOR2_X1 U13256 ( .A(n11539), .B(n11540), .ZN(n18202) );
  NOR2_X1 U13257 ( .A1(n11539), .A2(n11540), .ZN(n11541) );
  NAND2_X1 U13258 ( .A1(n21199), .A2(n21177), .ZN(n18162) );
  NOR2_X1 U13259 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18162), .ZN(
        n17936) );
  INV_X1 U13260 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n20952) );
  NOR2_X1 U13261 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11546) );
  NOR2_X1 U13262 ( .A1(n21199), .A2(n21177), .ZN(n20934) );
  NAND3_X1 U13263 ( .A1(n20934), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17941) );
  INV_X1 U13264 ( .A(n17941), .ZN(n20959) );
  NAND2_X1 U13265 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n20959), .ZN(
        n20962) );
  NAND2_X1 U13266 ( .A1(n20958), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n20982) );
  INV_X1 U13267 ( .A(n20982), .ZN(n20979) );
  NAND2_X1 U13268 ( .A1(n20979), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21148) );
  NOR2_X1 U13269 ( .A1(n11547), .A2(n21148), .ZN(n11552) );
  INV_X1 U13270 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21087) );
  NAND2_X1 U13271 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21135) );
  NOR2_X1 U13272 ( .A1(n21135), .A2(n17902), .ZN(n11700) );
  NAND2_X1 U13273 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n20837) );
  NOR2_X1 U13274 ( .A1(n20999), .A2(n20837), .ZN(n17960) );
  NAND2_X1 U13275 ( .A1(n11700), .A2(n17960), .ZN(n11752) );
  NOR2_X1 U13276 ( .A1(n21087), .A2(n11752), .ZN(n20993) );
  INV_X1 U13277 ( .A(n20993), .ZN(n11750) );
  OAI21_X1 U13278 ( .B1(n17920), .B2(n11750), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11548) );
  INV_X1 U13279 ( .A(n11548), .ZN(n11549) );
  NOR2_X1 U13280 ( .A1(n11550), .A2(n11549), .ZN(n11555) );
  INV_X1 U13281 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11551) );
  OAI22_X1 U13282 ( .A1(n11552), .A2(n11551), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18190), .ZN(n11553) );
  INV_X1 U13283 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21147) );
  NAND2_X1 U13284 ( .A1(n18123), .A2(n21147), .ZN(n18122) );
  NAND2_X1 U13285 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21093) );
  NAND2_X1 U13286 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11754) );
  INV_X1 U13287 ( .A(n11754), .ZN(n11558) );
  INV_X1 U13288 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18070) );
  INV_X1 U13289 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21025) );
  AOI21_X1 U13290 ( .B1(n18070), .B2(n21025), .A(n18189), .ZN(n11557) );
  INV_X1 U13291 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21036) );
  NAND2_X1 U13292 ( .A1(n11559), .A2(n21036), .ZN(n11765) );
  NOR2_X1 U13293 ( .A1(n11559), .A2(n21036), .ZN(n11743) );
  NAND2_X1 U13294 ( .A1(n18053), .A2(n18189), .ZN(n18052) );
  NAND2_X1 U13295 ( .A1(n18052), .A2(n11765), .ZN(n18045) );
  NOR2_X1 U13296 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18189), .ZN(
        n18098) );
  AOI21_X1 U13297 ( .B1(n18189), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18098), .ZN(n18046) );
  NAND2_X1 U13298 ( .A1(n18045), .A2(n18046), .ZN(n18044) );
  AOI22_X1 U13299 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17838), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U13300 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U13301 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U13302 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11562) );
  NAND4_X1 U13303 ( .A1(n11565), .A2(n11564), .A3(n11563), .A4(n11562), .ZN(
        n11572) );
  AOI22_X1 U13304 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U13305 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U13306 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U13307 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11567) );
  NAND4_X1 U13308 ( .A1(n11570), .A2(n11569), .A3(n11568), .A4(n11567), .ZN(
        n11571) );
  AOI22_X1 U13309 ( .A1(n17848), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11573) );
  OAI21_X1 U13310 ( .B1(n11641), .B2(n17873), .A(n11573), .ZN(n11579) );
  AOI22_X1 U13311 ( .A1(n17838), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U13312 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U13313 ( .A1(n17832), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11469), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U13314 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17833), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11574) );
  NAND4_X1 U13315 ( .A1(n11577), .A2(n11576), .A3(n11575), .A4(n11574), .ZN(
        n11578) );
  NAND2_X1 U13316 ( .A1(n18997), .A2(n20596), .ZN(n11731) );
  AOI22_X1 U13317 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U13318 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U13319 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11469), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U13320 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11583) );
  NAND4_X1 U13321 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11583), .ZN(
        n11592) );
  AOI22_X1 U13322 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U13323 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U13324 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U13325 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11587) );
  NAND4_X1 U13326 ( .A1(n11590), .A2(n11589), .A3(n11588), .A4(n11587), .ZN(
        n11591) );
  INV_X1 U13327 ( .A(n18957), .ZN(n11653) );
  AOI22_X1 U13328 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17838), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U13329 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U13330 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U13331 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11593) );
  NAND4_X1 U13332 ( .A1(n11596), .A2(n11595), .A3(n11594), .A4(n11593), .ZN(
        n11602) );
  AOI22_X1 U13333 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U13334 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U13335 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U13336 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11509), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11597) );
  NAND4_X1 U13337 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(
        n11601) );
  NAND2_X1 U13338 ( .A1(n11634), .A2(n18997), .ZN(n11732) );
  AND2_X1 U13339 ( .A1(n11653), .A2(n11732), .ZN(n11638) );
  AOI22_X1 U13340 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U13341 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U13342 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11469), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U13343 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11603) );
  NAND4_X1 U13344 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11612) );
  AOI22_X1 U13345 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U13346 ( .A1(n17861), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U13347 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17725), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U13348 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11607) );
  NAND4_X1 U13349 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n11611) );
  NAND2_X1 U13350 ( .A1(n18997), .A2(n18916), .ZN(n11714) );
  INV_X1 U13351 ( .A(n11714), .ZN(n11623) );
  AOI22_X1 U13352 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U13353 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U13354 ( .A1(n17838), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11613) );
  OAI21_X1 U13355 ( .B1(n11641), .B2(n17730), .A(n11613), .ZN(n11619) );
  AOI22_X1 U13356 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U13357 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U13358 ( .A1(n17832), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U13359 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10977), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11614) );
  NAND4_X1 U13360 ( .A1(n11617), .A2(n11616), .A3(n11615), .A4(n11614), .ZN(
        n11618) );
  AOI211_X1 U13361 ( .C1(n17849), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n11619), .B(n11618), .ZN(n11620) );
  NAND3_X1 U13362 ( .A1(n11622), .A2(n11621), .A3(n11620), .ZN(n11635) );
  NAND2_X1 U13363 ( .A1(n20653), .A2(n11635), .ZN(n11706) );
  NAND2_X1 U13364 ( .A1(n11623), .A2(n11706), .ZN(n11637) );
  AOI22_X1 U13365 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U13366 ( .A1(n17838), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U13367 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17833), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U13368 ( .A1(n17832), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11624) );
  NAND4_X1 U13369 ( .A1(n11627), .A2(n11626), .A3(n11625), .A4(n11624), .ZN(
        n11633) );
  AOI22_X1 U13370 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U13371 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U13372 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U13373 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11628) );
  NAND4_X1 U13374 ( .A1(n11631), .A2(n11630), .A3(n11629), .A4(n11628), .ZN(
        n11632) );
  NOR2_X1 U13375 ( .A1(n18916), .A2(n11635), .ZN(n11664) );
  INV_X1 U13376 ( .A(n11736), .ZN(n11652) );
  INV_X1 U13377 ( .A(n18997), .ZN(n11639) );
  OR2_X1 U13378 ( .A1(n11639), .A2(n11662), .ZN(n11711) );
  AOI22_X1 U13379 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17849), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U13380 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17838), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U13381 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11640) );
  OAI21_X1 U13382 ( .B1(n11641), .B2(n17695), .A(n11640), .ZN(n11647) );
  AOI22_X1 U13383 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U13384 ( .A1(n17861), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U13385 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U13386 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11469), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11642) );
  NAND4_X1 U13387 ( .A1(n11645), .A2(n11644), .A3(n11643), .A4(n11642), .ZN(
        n11646) );
  AOI21_X1 U13388 ( .B1(n20622), .B2(n11652), .A(n18916), .ZN(n11651) );
  AOI21_X1 U13389 ( .B1(n11652), .B2(n11711), .A(n11651), .ZN(n11656) );
  NAND2_X1 U13390 ( .A1(n20622), .A2(n20788), .ZN(n20600) );
  NOR2_X1 U13391 ( .A1(n20596), .A2(n19087), .ZN(n11663) );
  NAND2_X1 U13392 ( .A1(n20600), .A2(n11663), .ZN(n11713) );
  AOI21_X1 U13393 ( .B1(n11713), .B2(n11653), .A(n11660), .ZN(n11654) );
  INV_X1 U13394 ( .A(n11654), .ZN(n11655) );
  NAND3_X1 U13395 ( .A1(n11657), .A2(n11656), .A3(n11655), .ZN(n20820) );
  NAND4_X1 U13396 ( .A1(n18916), .A2(n18957), .A3(n11660), .A4(n11736), .ZN(
        n11702) );
  OR2_X1 U13397 ( .A1(n11702), .A2(n18997), .ZN(n11709) );
  NAND3_X1 U13398 ( .A1(n20653), .A2(n11707), .A3(n11657), .ZN(n11658) );
  NAND2_X1 U13399 ( .A1(n11709), .A2(n11658), .ZN(n17881) );
  NAND2_X1 U13400 ( .A1(n18997), .A2(n18957), .ZN(n20800) );
  NOR2_X1 U13401 ( .A1(n11706), .A2(n20800), .ZN(n15624) );
  NAND3_X1 U13402 ( .A1(n20106), .A2(n11660), .A3(n15624), .ZN(n11703) );
  NAND3_X1 U13403 ( .A1(n17125), .A2(n11703), .A3(n20114), .ZN(n20802) );
  NAND2_X1 U13404 ( .A1(n11701), .A2(n11702), .ZN(n20819) );
  INV_X1 U13405 ( .A(n11707), .ZN(n11665) );
  NAND2_X1 U13406 ( .A1(n20596), .A2(n11665), .ZN(n20798) );
  NAND2_X1 U13407 ( .A1(n20800), .A2(n20798), .ZN(n11749) );
  INV_X1 U13408 ( .A(n11664), .ZN(n20801) );
  NAND2_X1 U13409 ( .A1(n18044), .A2(n20856), .ZN(n11746) );
  INV_X1 U13410 ( .A(n11746), .ZN(n11705) );
  INV_X1 U13411 ( .A(n11700), .ZN(n17898) );
  NOR2_X1 U13412 ( .A1(n21148), .A2(n17898), .ZN(n17897) );
  INV_X1 U13413 ( .A(n20780), .ZN(n11678) );
  NOR2_X1 U13414 ( .A1(n20642), .A2(n11675), .ZN(n11672) );
  NAND2_X1 U13415 ( .A1(n11672), .A2(n11673), .ZN(n11670) );
  NOR2_X1 U13416 ( .A1(n20633), .A2(n11670), .ZN(n11669) );
  NAND2_X1 U13417 ( .A1(n11669), .A2(n20629), .ZN(n11668) );
  NOR2_X1 U13418 ( .A1(n20625), .A2(n11668), .ZN(n11695) );
  XOR2_X1 U13419 ( .A(n20625), .B(n11668), .Z(n18204) );
  XOR2_X1 U13420 ( .A(n20629), .B(n11669), .Z(n11689) );
  XOR2_X1 U13421 ( .A(n20633), .B(n11670), .Z(n11671) );
  NAND2_X1 U13422 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11671), .ZN(
        n11688) );
  XOR2_X1 U13423 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11671), .Z(
        n18224) );
  XOR2_X1 U13424 ( .A(n11673), .B(n11672), .Z(n11684) );
  XOR2_X1 U13425 ( .A(n20642), .B(n11675), .Z(n11674) );
  NAND2_X1 U13426 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11674), .ZN(
        n11683) );
  XOR2_X1 U13427 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11674), .Z(
        n18247) );
  NAND2_X1 U13428 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11677), .ZN(
        n11682) );
  XNOR2_X1 U13429 ( .A(n11522), .B(n11677), .ZN(n18260) );
  INV_X1 U13430 ( .A(n18270), .ZN(n18272) );
  INV_X1 U13431 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20994) );
  NAND2_X1 U13432 ( .A1(n11678), .A2(n20994), .ZN(n18277) );
  NOR2_X1 U13433 ( .A1(n18272), .A2(n18277), .ZN(n18271) );
  AOI211_X1 U13434 ( .C1(n11680), .C2(n20864), .A(n11679), .B(n18271), .ZN(
        n18261) );
  NAND2_X1 U13435 ( .A1(n18260), .A2(n18261), .ZN(n11681) );
  NAND2_X1 U13436 ( .A1(n11682), .A2(n11681), .ZN(n18246) );
  NAND2_X1 U13437 ( .A1(n18247), .A2(n18246), .ZN(n18245) );
  NAND2_X1 U13438 ( .A1(n11683), .A2(n18245), .ZN(n11685) );
  NAND2_X1 U13439 ( .A1(n11684), .A2(n11685), .ZN(n11686) );
  XNOR2_X1 U13440 ( .A(n11685), .B(n11684), .ZN(n18232) );
  NAND2_X1 U13441 ( .A1(n11686), .A2(n18237), .ZN(n18223) );
  NAND2_X1 U13442 ( .A1(n18224), .A2(n18223), .ZN(n11687) );
  NAND2_X1 U13443 ( .A1(n11688), .A2(n11687), .ZN(n11690) );
  NAND2_X1 U13444 ( .A1(n11689), .A2(n11690), .ZN(n11691) );
  XOR2_X1 U13445 ( .A(n11690), .B(n11689), .Z(n18217) );
  NAND2_X1 U13446 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18217), .ZN(
        n18216) );
  NAND2_X1 U13447 ( .A1(n11695), .A2(n11692), .ZN(n11696) );
  NAND2_X1 U13448 ( .A1(n18204), .A2(n18205), .ZN(n18203) );
  NAND2_X1 U13449 ( .A1(n11695), .A2(n11694), .ZN(n11693) );
  OAI211_X1 U13450 ( .C1(n11695), .C2(n11694), .A(n18203), .B(n11693), .ZN(
        n18194) );
  NAND2_X1 U13451 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18194), .ZN(
        n18193) );
  INV_X1 U13452 ( .A(n18149), .ZN(n20936) );
  INV_X1 U13453 ( .A(n21138), .ZN(n11697) );
  OAI22_X1 U13454 ( .A1(n20936), .A2(n21050), .B1(n21137), .B2(n11697), .ZN(
        n20929) );
  NAND2_X1 U13455 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20928) );
  NAND3_X1 U13456 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20901) );
  NOR2_X1 U13457 ( .A1(n11698), .A2(n20901), .ZN(n20908) );
  AOI21_X1 U13458 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20873) );
  INV_X1 U13459 ( .A(n20873), .ZN(n20876) );
  NAND2_X1 U13460 ( .A1(n20908), .A2(n20876), .ZN(n20910) );
  NOR2_X1 U13461 ( .A1(n20928), .A2(n20910), .ZN(n20978) );
  INV_X1 U13462 ( .A(n20978), .ZN(n11699) );
  NOR2_X1 U13463 ( .A1(n21148), .A2(n11699), .ZN(n21139) );
  NAND2_X1 U13464 ( .A1(n11700), .A2(n21139), .ZN(n20836) );
  NAND2_X1 U13465 ( .A1(n21207), .A2(n11703), .ZN(n21007) );
  NAND2_X1 U13466 ( .A1(n21192), .A2(n20994), .ZN(n20853) );
  NAND2_X1 U13467 ( .A1(n21187), .A2(n20853), .ZN(n20872) );
  NAND3_X1 U13468 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n20908), .ZN(n20909) );
  NOR2_X1 U13469 ( .A1(n20918), .A2(n20909), .ZN(n21191) );
  NAND2_X1 U13470 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21191), .ZN(
        n20932) );
  INV_X1 U13471 ( .A(n20932), .ZN(n11747) );
  NAND2_X1 U13472 ( .A1(n17897), .A2(n11747), .ZN(n11756) );
  OAI22_X1 U13473 ( .A1(n21172), .A2(n20836), .B1(n20872), .B2(n11756), .ZN(
        n21053) );
  AOI21_X1 U13474 ( .B1(n17897), .B2(n20929), .A(n21053), .ZN(n21089) );
  INV_X1 U13475 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21105) );
  NOR2_X1 U13476 ( .A1(n21105), .A2(n21093), .ZN(n11753) );
  NAND2_X1 U13477 ( .A1(n17960), .A2(n11753), .ZN(n21010) );
  OR2_X1 U13478 ( .A1(n21010), .A2(n11754), .ZN(n18090) );
  NOR2_X1 U13479 ( .A1(n21089), .A2(n18090), .ZN(n21034) );
  AND2_X1 U13480 ( .A1(n21034), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11704) );
  AOI21_X1 U13481 ( .B1(n11705), .B2(n18189), .A(n11704), .ZN(n11742) );
  OAI211_X1 U13482 ( .C1(n11708), .C2(n18916), .A(n11707), .B(n11706), .ZN(
        n11710) );
  OAI21_X1 U13483 ( .B1(n11711), .B2(n11710), .A(n11709), .ZN(n11712) );
  OAI211_X1 U13484 ( .C1(n11715), .C2(n11714), .A(n11713), .B(n11712), .ZN(
        n15642) );
  INV_X1 U13485 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18795) );
  AOI22_X1 U13486 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18795), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20813), .ZN(n11723) );
  OAI22_X1 U13487 ( .A1(n11420), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18796), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11726) );
  NAND2_X1 U13488 ( .A1(n18802), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11727) );
  OR2_X1 U13489 ( .A1(n11726), .A2(n11727), .ZN(n11716) );
  NAND2_X1 U13490 ( .A1(n11723), .A2(n11724), .ZN(n11717) );
  OAI22_X1 U13491 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17124), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11718), .ZN(n11720) );
  NOR2_X1 U13492 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17124), .ZN(
        n11719) );
  NAND2_X1 U13493 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11718), .ZN(
        n11721) );
  AOI22_X1 U13494 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11720), .B1(
        n11719), .B2(n11721), .ZN(n11725) );
  OAI211_X1 U13495 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18802), .A(
        n11725), .B(n11727), .ZN(n11733) );
  AOI21_X1 U13496 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11721), .A(
        n11720), .ZN(n11722) );
  XOR2_X1 U13497 ( .A(n11724), .B(n11723), .Z(n11734) );
  NAND2_X1 U13498 ( .A1(n11725), .A2(n11734), .ZN(n11730) );
  OAI211_X1 U13499 ( .C1(n11733), .C2(n11726), .A(n11728), .B(n11730), .ZN(
        n11740) );
  NAND2_X1 U13500 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n21652) );
  XNOR2_X1 U13501 ( .A(n11727), .B(n11726), .ZN(n11729) );
  NOR2_X1 U13502 ( .A1(n21607), .A2(n21226), .ZN(n15645) );
  INV_X2 U13503 ( .A(n21651), .ZN(n18364) );
  NOR2_X1 U13504 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n21654), .ZN(n21648) );
  NOR2_X1 U13505 ( .A1(n21654), .A2(n21651), .ZN(n18360) );
  INV_X2 U13506 ( .A(n18360), .ZN(n18363) );
  OAI211_X1 U13507 ( .C1(n18997), .C2(n20596), .A(n20105), .B(n11731), .ZN(
        n21228) );
  NAND3_X1 U13508 ( .A1(n15645), .A2(n11732), .A3(n21228), .ZN(n11739) );
  INV_X1 U13509 ( .A(n11733), .ZN(n11735) );
  AOI21_X1 U13510 ( .B1(n11735), .B2(n11734), .A(n21226), .ZN(n21209) );
  AND2_X1 U13511 ( .A1(n21209), .A2(n20596), .ZN(n11737) );
  OAI211_X1 U13512 ( .C1(n11737), .C2(n21205), .A(n11736), .B(n18997), .ZN(
        n11738) );
  OAI211_X1 U13513 ( .C1(n18916), .C2(n11740), .A(n11739), .B(n11738), .ZN(
        n11741) );
  NOR2_X1 U13514 ( .A1(n11742), .A2(n21194), .ZN(n11763) );
  INV_X1 U13515 ( .A(n11743), .ZN(n11745) );
  NAND2_X1 U13516 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18189), .ZN(
        n11744) );
  AOI221_X1 U13517 ( .B1(n20625), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), 
        .C1(n11746), .C2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n18097), .ZN(
        n11761) );
  NAND2_X1 U13518 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n11747), .ZN(
        n21186) );
  INV_X1 U13519 ( .A(n21186), .ZN(n20944) );
  NAND2_X1 U13520 ( .A1(n17897), .A2(n20944), .ZN(n20840) );
  INV_X1 U13521 ( .A(n20802), .ZN(n11748) );
  AOI21_X1 U13522 ( .B1(n11749), .B2(n11748), .A(n20820), .ZN(n20943) );
  NOR2_X1 U13523 ( .A1(n18090), .A2(n21036), .ZN(n21054) );
  INV_X1 U13524 ( .A(n21054), .ZN(n11755) );
  NAND3_X1 U13525 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21028) );
  NOR2_X1 U13526 ( .A1(n18070), .A2(n21028), .ZN(n21039) );
  INV_X1 U13527 ( .A(n21139), .ZN(n11751) );
  OAI21_X1 U13528 ( .B1(n11751), .B2(n11750), .A(n21204), .ZN(n21099) );
  OAI21_X1 U13529 ( .B1(n21039), .B2(n21172), .A(n21099), .ZN(n21035) );
  AOI221_X1 U13530 ( .B1(n20840), .B2(n21188), .C1(n11755), .C2(n21188), .A(
        n21035), .ZN(n21047) );
  INV_X1 U13531 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18140) );
  NAND2_X1 U13532 ( .A1(n21138), .A2(n20958), .ZN(n18139) );
  NAND2_X1 U13533 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n20976), .ZN(
        n20984) );
  NAND2_X1 U13534 ( .A1(n11753), .A2(n20839), .ZN(n18017) );
  NOR2_X1 U13535 ( .A1(n11754), .A2(n18017), .ZN(n21022) );
  NAND3_X1 U13536 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n21022), .ZN(n21055) );
  INV_X1 U13537 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18042) );
  AOI22_X1 U13538 ( .A1(n21114), .A2(n21055), .B1(n21203), .B2(n18100), .ZN(
        n11759) );
  NOR2_X1 U13539 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21248) );
  NAND2_X1 U13540 ( .A1(n21248), .A2(n21246), .ZN(n17884) );
  NOR2_X2 U13541 ( .A1(n10979), .A2(n21171), .ZN(n21080) );
  INV_X1 U13542 ( .A(n21080), .ZN(n21094) );
  NOR2_X1 U13543 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21172), .ZN(
        n21052) );
  NOR2_X1 U13544 ( .A1(n11756), .A2(n11755), .ZN(n21048) );
  INV_X1 U13545 ( .A(n21048), .ZN(n11757) );
  OAI21_X1 U13546 ( .B1(n21052), .B2(n21007), .A(n11757), .ZN(n11758) );
  NAND4_X1 U13547 ( .A1(n21047), .A2(n11759), .A3(n21094), .A4(n11758), .ZN(
        n11760) );
  OR2_X1 U13548 ( .A1(n11761), .A2(n11760), .ZN(n11762) );
  OAI211_X1 U13549 ( .C1(n11763), .C2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11762), .B(n11764), .ZN(n11767) );
  INV_X1 U13550 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n20539) );
  NOR2_X1 U13551 ( .A1(n11764), .A2(n20539), .ZN(n18037) );
  NAND2_X1 U13552 ( .A1(n11767), .A2(n11766), .ZN(P3_U2834) );
  AOI22_X1 U13553 ( .A1(n10963), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U13554 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U13555 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11770) );
  AND2_X4 U13556 ( .A1(n14939), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11975) );
  AND2_X4 U13557 ( .A1(n14939), .A2(n17066), .ZN(n11977) );
  AOI22_X1 U13558 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11769) );
  NAND4_X1 U13559 ( .A1(n11772), .A2(n11771), .A3(n11770), .A4(n11769), .ZN(
        n11773) );
  AOI22_X1 U13560 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U13561 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U13562 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U13563 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11774) );
  NAND4_X1 U13564 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n11778) );
  NAND2_X1 U13565 ( .A1(n11778), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11779) );
  AOI22_X1 U13566 ( .A1(n10963), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U13567 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U13568 ( .A1(n15776), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U13569 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11781) );
  NAND4_X1 U13570 ( .A1(n11784), .A2(n11783), .A3(n11782), .A4(n11781), .ZN(
        n11785) );
  NAND2_X1 U13571 ( .A1(n11785), .A2(n11832), .ZN(n11792) );
  AOI22_X1 U13572 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U13573 ( .A1(n10963), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U13574 ( .A1(n10967), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U13575 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11786) );
  NAND4_X1 U13576 ( .A1(n11789), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n11790) );
  NAND2_X1 U13577 ( .A1(n11790), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11791) );
  AOI22_X1 U13578 ( .A1(n10963), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11797) );
  INV_X4 U13579 ( .A(n15785), .ZN(n15777) );
  AOI22_X1 U13580 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U13581 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U13582 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11794) );
  NAND4_X1 U13583 ( .A1(n11797), .A2(n11796), .A3(n11795), .A4(n11794), .ZN(
        n11798) );
  AOI22_X1 U13584 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U13585 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U13586 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U13587 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11799) );
  NAND4_X1 U13588 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11803) );
  NAND2_X1 U13589 ( .A1(n11886), .A2(n12894), .ZN(n12601) );
  AOI22_X1 U13590 ( .A1(n10963), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U13591 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U13592 ( .A1(n15776), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U13593 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U13594 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U13595 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U13596 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U13597 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11810) );
  NAND3_X1 U13598 ( .A1(n11812), .A2(n11811), .A3(n11810), .ZN(n11813) );
  AOI22_X1 U13599 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11818) );
  AOI22_X1 U13600 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U13601 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U13602 ( .A1(n10966), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10964), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11814) );
  NAND2_X1 U13603 ( .A1(n11818), .A2(n11817), .ZN(n11824) );
  AOI22_X1 U13604 ( .A1(n10963), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U13605 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U13606 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U13607 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11819) );
  NAND4_X1 U13608 ( .A1(n11822), .A2(n11821), .A3(n11820), .A4(n11819), .ZN(
        n11823) );
  MUX2_X2 U13609 ( .A(n11824), .B(n11823), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12901) );
  NAND2_X1 U13610 ( .A1(n12899), .A2(n12901), .ZN(n11827) );
  NOR2_X1 U13611 ( .A1(n12635), .A2(n10969), .ZN(n11825) );
  NAND2_X1 U13612 ( .A1(n12892), .A2(n11880), .ZN(n11826) );
  NAND2_X1 U13613 ( .A1(n11827), .A2(n11826), .ZN(n11907) );
  AOI22_X1 U13614 ( .A1(n10962), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U13615 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U13616 ( .A1(n10967), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U13617 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11828) );
  NAND4_X1 U13618 ( .A1(n11831), .A2(n11830), .A3(n11829), .A4(n11828), .ZN(
        n11833) );
  NAND2_X1 U13619 ( .A1(n11833), .A2(n11832), .ZN(n11841) );
  AOI22_X1 U13620 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U13621 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U13622 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11834) );
  NAND3_X1 U13623 ( .A1(n11836), .A2(n11835), .A3(n11834), .ZN(n11839) );
  AOI22_X1 U13624 ( .A1(n10963), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11837) );
  NAND2_X1 U13625 ( .A1(n11841), .A2(n11840), .ZN(n11869) );
  AOI22_X1 U13626 ( .A1(n10963), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11010), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U13627 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U13628 ( .A1(n15776), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U13629 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11843) );
  NAND4_X1 U13630 ( .A1(n11846), .A2(n11845), .A3(n11844), .A4(n11843), .ZN(
        n11852) );
  AOI22_X1 U13631 ( .A1(n10963), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11010), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U13632 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U13633 ( .A1(n10967), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U13634 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11847) );
  NAND4_X1 U13635 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11851) );
  MUX2_X2 U13636 ( .A(n11852), .B(n11851), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12641) );
  NAND2_X2 U13637 ( .A1(n19703), .A2(n12641), .ZN(n15000) );
  NAND2_X1 U13638 ( .A1(n11907), .A2(n15291), .ZN(n11872) );
  NAND2_X1 U13639 ( .A1(n11853), .A2(n11884), .ZN(n11855) );
  NAND2_X1 U13640 ( .A1(n11886), .A2(n12901), .ZN(n11854) );
  NAND2_X1 U13641 ( .A1(n19376), .A2(n10969), .ZN(n11866) );
  AOI22_X1 U13642 ( .A1(n10963), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U13643 ( .A1(n15793), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U13644 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U13645 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11856) );
  NAND4_X1 U13646 ( .A1(n11859), .A2(n11858), .A3(n11857), .A4(n11856), .ZN(
        n11865) );
  AOI22_X1 U13647 ( .A1(n10963), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15793), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U13648 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U13649 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U13650 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11860) );
  NAND4_X1 U13651 ( .A1(n11863), .A2(n11862), .A3(n11861), .A4(n11860), .ZN(
        n11864) );
  MUX2_X2 U13652 ( .A(n11865), .B(n11864), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n17083) );
  INV_X2 U13653 ( .A(n17083), .ZN(n12600) );
  NAND3_X1 U13654 ( .A1(n11870), .A2(n18657), .A3(n12627), .ZN(n12905) );
  AND2_X1 U13655 ( .A1(n11886), .A2(n12633), .ZN(n12891) );
  NAND2_X1 U13656 ( .A1(n12891), .A2(n12892), .ZN(n11906) );
  NAND2_X1 U13657 ( .A1(n11906), .A2(n12627), .ZN(n11871) );
  NAND2_X1 U13658 ( .A1(n11872), .A2(n11904), .ZN(n11873) );
  AND3_X2 U13659 ( .A1(n12600), .A2(n12901), .A3(n12635), .ZN(n11877) );
  NAND2_X1 U13660 ( .A1(n12641), .A2(n11875), .ZN(n11878) );
  NAND2_X1 U13661 ( .A1(n11878), .A2(n11881), .ZN(n12883) );
  INV_X1 U13662 ( .A(n12883), .ZN(n11879) );
  NAND2_X1 U13663 ( .A1(n18711), .A2(n17057), .ZN(n18695) );
  NAND2_X1 U13664 ( .A1(n12633), .A2(n12627), .ZN(n18656) );
  INV_X1 U13665 ( .A(n18656), .ZN(n15019) );
  AND2_X1 U13666 ( .A1(n19376), .A2(n12635), .ZN(n13272) );
  OAI211_X1 U13667 ( .C1(n18695), .C2(n14986), .A(n11887), .B(n11889), .ZN(
        n11882) );
  INV_X1 U13668 ( .A(n11882), .ZN(n11883) );
  INV_X1 U13669 ( .A(n11896), .ZN(n11894) );
  INV_X1 U13670 ( .A(n11884), .ZN(n11885) );
  NAND2_X1 U13671 ( .A1(n11915), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11893) );
  NOR2_X1 U13672 ( .A1(n11897), .A2(n15000), .ZN(n11888) );
  AND2_X2 U13673 ( .A1(n12890), .A2(n11888), .ZN(n12906) );
  AOI22_X1 U13674 ( .A1(n11899), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11892) );
  INV_X1 U13675 ( .A(n11889), .ZN(n11890) );
  NAND3_X1 U13676 ( .A1(n11893), .A2(n11892), .A3(n11891), .ZN(n11895) );
  NAND2_X1 U13677 ( .A1(n15291), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11898) );
  NOR2_X1 U13678 ( .A1(n11898), .A2(n11897), .ZN(n11900) );
  INV_X1 U13679 ( .A(n18695), .ZN(n11932) );
  NAND2_X1 U13680 ( .A1(n11932), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11901) );
  INV_X1 U13681 ( .A(n11904), .ZN(n11905) );
  AOI21_X1 U13682 ( .B1(n11907), .B2(n11906), .A(n11905), .ZN(n11913) );
  NAND2_X1 U13683 ( .A1(n11915), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11912) );
  INV_X1 U13684 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n12645) );
  OAI21_X1 U13685 ( .B1(n12282), .B2(n12645), .A(n11908), .ZN(n11911) );
  NAND2_X1 U13686 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11909) );
  OAI211_X1 U13687 ( .C1(n12274), .C2(n14843), .A(n18695), .B(n11909), .ZN(
        n11910) );
  INV_X4 U13688 ( .A(n11916), .ZN(n12337) );
  INV_X1 U13689 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n11919) );
  NAND2_X1 U13690 ( .A1(n10980), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11918) );
  NAND2_X1 U13691 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11917) );
  OAI211_X1 U13692 ( .C1(n12274), .C2(n11919), .A(n11918), .B(n11917), .ZN(
        n11920) );
  AOI21_X2 U13693 ( .B1(n12346), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11920), .ZN(n11924) );
  NAND2_X1 U13694 ( .A1(n11921), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11923) );
  AOI21_X1 U13695 ( .B1(n18711), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11922) );
  INV_X1 U13696 ( .A(n11924), .ZN(n11925) );
  INV_X1 U13697 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n15338) );
  NAND2_X1 U13698 ( .A1(n10980), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11930) );
  NAND2_X1 U13699 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11929) );
  OAI211_X1 U13700 ( .C1(n12274), .C2(n15338), .A(n11930), .B(n11929), .ZN(
        n11931) );
  NAND2_X1 U13701 ( .A1(n11921), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11934) );
  NAND2_X1 U13702 ( .A1(n11932), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11933) );
  INV_X1 U13703 ( .A(n11937), .ZN(n11939) );
  INV_X1 U13704 ( .A(n11942), .ZN(n11938) );
  XNOR2_X2 U13705 ( .A(n11939), .B(n11938), .ZN(n14681) );
  OR2_X1 U13706 ( .A1(n11941), .A2(n11940), .ZN(n11945) );
  INV_X1 U13707 ( .A(n12950), .ZN(n18393) );
  INV_X1 U13708 ( .A(n12944), .ZN(n11943) );
  INV_X1 U13709 ( .A(n11944), .ZN(n11946) );
  NAND2_X1 U13710 ( .A1(n11946), .A2(n11945), .ZN(n11959) );
  INV_X1 U13711 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11947) );
  OAI21_X1 U13712 ( .B1(n12025), .B2(n11947), .A(n12651), .ZN(n11948) );
  NOR2_X1 U13713 ( .A1(n11949), .A2(n11948), .ZN(n11954) );
  NAND2_X1 U13714 ( .A1(n14681), .A2(n12950), .ZN(n11955) );
  AOI22_X1 U13715 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12105), .B1(
        n12104), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11953) );
  INV_X1 U13716 ( .A(n11955), .ZN(n11950) );
  AOI22_X1 U13717 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n12099), .B1(
        n19273), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11952) );
  NOR2_X1 U13718 ( .A1(n12950), .A2(n11937), .ZN(n11957) );
  INV_X1 U13719 ( .A(n11957), .ZN(n11958) );
  NOR2_X2 U13720 ( .A1(n11009), .A2(n11958), .ZN(n19360) );
  AOI22_X1 U13721 ( .A1(n15231), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n19360), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11951) );
  NOR2_X2 U13722 ( .A1(n11009), .A2(n11955), .ZN(n19344) );
  AOI22_X1 U13723 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19344), .B1(
        n19288), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11968) );
  NOR2_X2 U13724 ( .A1(n11009), .A2(n11959), .ZN(n19333) );
  INV_X1 U13725 ( .A(n11959), .ZN(n11963) );
  AOI22_X1 U13726 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12097), .B1(
        n19259), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11965) );
  NAND2_X1 U13727 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11974) );
  AOI22_X1 U13728 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11973) );
  AND2_X2 U13729 ( .A1(n14978), .A2(n13083), .ZN(n13103) );
  AOI22_X1 U13730 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11972) );
  NAND2_X1 U13731 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11971) );
  AND4_X1 U13732 ( .A1(n11974), .A2(n11973), .A3(n11972), .A4(n11971), .ZN(
        n11989) );
  NAND3_X1 U13733 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12246) );
  AOI211_X1 U13734 ( .C1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .C2(n13118), .A(
        n11401), .B(n11404), .ZN(n11988) );
  INV_X1 U13735 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11976) );
  INV_X1 U13736 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12701) );
  OAI22_X1 U13737 ( .A1(n12046), .A2(n11976), .B1(n13030), .B2(n12701), .ZN(
        n11980) );
  INV_X1 U13738 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12696) );
  INV_X1 U13739 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11978) );
  OAI22_X1 U13740 ( .A1(n13033), .A2(n12696), .B1(n13032), .B2(n11978), .ZN(
        n11979) );
  NOR2_X1 U13741 ( .A1(n11980), .A2(n11979), .ZN(n11987) );
  INV_X1 U13742 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11984) );
  NAND2_X1 U13743 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11983) );
  INV_X1 U13744 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11981) );
  NAND2_X1 U13745 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11982) );
  OAI211_X1 U13746 ( .C1(n11984), .C2(n13026), .A(n11983), .B(n11982), .ZN(
        n11985) );
  INV_X1 U13747 ( .A(n11985), .ZN(n11986) );
  NAND4_X1 U13748 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n12059) );
  INV_X1 U13749 ( .A(n12059), .ZN(n14675) );
  INV_X1 U13750 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12721) );
  INV_X1 U13751 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13137) );
  OAI22_X1 U13752 ( .A1(n13033), .A2(n12721), .B1(n13032), .B2(n13137), .ZN(
        n11990) );
  INV_X1 U13753 ( .A(n11990), .ZN(n11995) );
  AOI22_X1 U13754 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n13118), .ZN(n11994) );
  AOI22_X1 U13755 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13108), .B1(
        n11991), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U13756 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12763), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11992) );
  NAND4_X1 U13757 ( .A1(n11995), .A2(n11994), .A3(n11993), .A4(n11992), .ZN(
        n12002) );
  AOI22_X1 U13758 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U13759 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13103), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U13760 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n13022), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U13761 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12012), .B1(
        n13115), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11997) );
  NAND4_X1 U13762 ( .A1(n12000), .A2(n11999), .A3(n11998), .A4(n11997), .ZN(
        n12001) );
  NOR2_X1 U13763 ( .A1(n14675), .A2(n12060), .ZN(n12003) );
  NAND2_X1 U13764 ( .A1(n12633), .A2(n12003), .ZN(n12063) );
  INV_X1 U13765 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13011) );
  INV_X1 U13766 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13007) );
  OAI22_X1 U13767 ( .A1(n12046), .A2(n13011), .B1(n13030), .B2(n13007), .ZN(
        n12006) );
  INV_X1 U13768 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12738) );
  INV_X1 U13769 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12004) );
  OAI22_X1 U13770 ( .A1(n13033), .A2(n12738), .B1(n13032), .B2(n12004), .ZN(
        n12005) );
  OR2_X1 U13771 ( .A1(n12006), .A2(n12005), .ZN(n12011) );
  INV_X1 U13772 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12009) );
  NAND2_X1 U13773 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12008) );
  NAND2_X1 U13774 ( .A1(n13117), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12007) );
  OAI211_X1 U13775 ( .C1(n12009), .C2(n12191), .A(n12008), .B(n12007), .ZN(
        n12010) );
  NOR2_X1 U13776 ( .A1(n12011), .A2(n12010), .ZN(n12023) );
  NAND2_X1 U13777 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12016) );
  AOI22_X1 U13778 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U13779 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12014) );
  NAND2_X1 U13780 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12013) );
  NAND4_X1 U13781 ( .A1(n12016), .A2(n12015), .A3(n12014), .A4(n12013), .ZN(
        n12021) );
  INV_X1 U13782 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12019) );
  NAND2_X1 U13783 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12018) );
  NAND2_X1 U13784 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12017) );
  OAI211_X1 U13785 ( .C1(n12019), .C2(n13026), .A(n12018), .B(n12017), .ZN(
        n12020) );
  NOR2_X1 U13786 ( .A1(n12021), .A2(n12020), .ZN(n12022) );
  NAND2_X1 U13787 ( .A1(n12063), .A2(n12663), .ZN(n12024) );
  AOI22_X1 U13788 ( .A1(n12096), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__3__SCAN_IN), .B2(n19288), .ZN(n12029) );
  AOI22_X1 U13789 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19344), .B1(
        n19333), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U13790 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12098), .B1(
        n15140), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U13791 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n15231), .B1(
        n19273), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U13792 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12105), .B1(
        n12106), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U13793 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19360), .B1(
        n12097), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U13794 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12104), .B1(
        n12099), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12030) );
  INV_X1 U13795 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12756) );
  INV_X1 U13796 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13025) );
  OAI22_X1 U13797 ( .A1(n13033), .A2(n12756), .B1(n13030), .B2(n13025), .ZN(
        n12037) );
  NAND2_X1 U13798 ( .A1(n13117), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12035) );
  NAND2_X1 U13799 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12034) );
  NAND2_X1 U13800 ( .A1(n12035), .A2(n12034), .ZN(n12036) );
  NOR2_X1 U13801 ( .A1(n12037), .A2(n12036), .ZN(n12053) );
  INV_X1 U13802 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12040) );
  NAND2_X1 U13803 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12039) );
  NAND2_X1 U13804 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12038) );
  OAI211_X1 U13805 ( .C1(n12040), .C2(n13026), .A(n12039), .B(n12038), .ZN(
        n12041) );
  INV_X1 U13806 ( .A(n12041), .ZN(n12052) );
  NAND2_X1 U13807 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12045) );
  AOI22_X1 U13808 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U13809 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12043) );
  NAND2_X1 U13810 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12042) );
  AND4_X1 U13811 ( .A1(n12045), .A2(n12044), .A3(n12043), .A4(n12042), .ZN(
        n12051) );
  INV_X1 U13812 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13031) );
  NAND2_X1 U13813 ( .A1(n13113), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12048) );
  NAND2_X1 U13814 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12047) );
  OAI211_X1 U13815 ( .C1(n12046), .C2(n13031), .A(n12048), .B(n12047), .ZN(
        n12049) );
  INV_X1 U13816 ( .A(n12049), .ZN(n12050) );
  NAND4_X1 U13817 ( .A1(n12053), .A2(n12052), .A3(n12051), .A4(n12050), .ZN(
        n12668) );
  INV_X1 U13818 ( .A(n12668), .ZN(n12054) );
  NAND2_X1 U13819 ( .A1(n12054), .A2(n12633), .ZN(n12055) );
  NAND2_X1 U13820 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14675), .ZN(
        n14674) );
  NOR2_X1 U13821 ( .A1(n12060), .A2(n14674), .ZN(n12062) );
  INV_X1 U13822 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15284) );
  NOR2_X1 U13823 ( .A1(n12059), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12061) );
  XNOR2_X1 U13824 ( .A(n12061), .B(n12060), .ZN(n14686) );
  NOR2_X1 U13825 ( .A1(n15284), .A2(n14686), .ZN(n14685) );
  NOR2_X1 U13826 ( .A1(n12062), .A2(n14685), .ZN(n12065) );
  XOR2_X1 U13827 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12065), .Z(
        n15666) );
  INV_X1 U13828 ( .A(n15666), .ZN(n12064) );
  XNOR2_X1 U13829 ( .A(n12063), .B(n12663), .ZN(n15664) );
  NAND2_X1 U13830 ( .A1(n12064), .A2(n15664), .ZN(n15677) );
  INV_X1 U13831 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15670) );
  OR2_X1 U13832 ( .A1(n12065), .A2(n15670), .ZN(n12066) );
  NAND2_X1 U13833 ( .A1(n15677), .A2(n12066), .ZN(n12067) );
  INV_X1 U13834 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15212) );
  XNOR2_X1 U13835 ( .A(n12067), .B(n15212), .ZN(n15160) );
  NAND2_X1 U13836 ( .A1(n12067), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12068) );
  INV_X1 U13837 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12069) );
  INV_X1 U13838 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12776) );
  OAI22_X1 U13839 ( .A1(n12046), .A2(n12069), .B1(n13030), .B2(n12776), .ZN(
        n12073) );
  INV_X1 U13840 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12071) );
  INV_X1 U13841 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12070) );
  OAI22_X1 U13842 ( .A1(n13033), .A2(n12071), .B1(n13032), .B2(n12070), .ZN(
        n12072) );
  NOR2_X1 U13843 ( .A1(n12073), .A2(n12072), .ZN(n12089) );
  INV_X1 U13844 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12780) );
  NAND2_X1 U13845 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12075) );
  NAND2_X1 U13846 ( .A1(n13117), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12074) );
  OAI211_X1 U13847 ( .C1(n12191), .C2(n12780), .A(n12075), .B(n12074), .ZN(
        n12076) );
  INV_X1 U13848 ( .A(n12076), .ZN(n12088) );
  NAND2_X1 U13849 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12081) );
  AOI22_X1 U13850 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12077), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U13851 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13103), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12079) );
  NAND2_X1 U13852 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12078) );
  AND4_X1 U13853 ( .A1(n12081), .A2(n12080), .A3(n12079), .A4(n12078), .ZN(
        n12087) );
  INV_X1 U13854 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12084) );
  NAND2_X1 U13855 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12083) );
  NAND2_X1 U13856 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12082) );
  OAI211_X1 U13857 ( .C1(n13026), .C2(n12084), .A(n12083), .B(n12082), .ZN(
        n12085) );
  INV_X1 U13858 ( .A(n12085), .ZN(n12086) );
  NAND4_X1 U13859 ( .A1(n12089), .A2(n12088), .A3(n12087), .A4(n12086), .ZN(
        n12233) );
  NAND2_X1 U13860 ( .A1(n12090), .A2(n12675), .ZN(n12091) );
  INV_X1 U13861 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18678) );
  INV_X1 U13862 ( .A(n12092), .ZN(n12094) );
  NAND2_X1 U13863 ( .A1(n12094), .A2(n12093), .ZN(n12095) );
  AOI22_X1 U13864 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19344), .B1(
        n12096), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U13865 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19360), .B1(
        n12097), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U13866 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n12098), .B1(
        n19259), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U13867 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n12099), .B1(
        n19273), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U13868 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19333), .B1(
        n19288), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U13869 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19226), .B1(
        n15140), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U13870 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n12104), .B1(
        n15231), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U13871 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n12105), .B1(
        n12106), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12107) );
  NAND2_X1 U13872 ( .A1(n11416), .A2(n11415), .ZN(n12132) );
  INV_X1 U13873 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12112) );
  INV_X1 U13874 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12111) );
  OAI22_X1 U13875 ( .A1(n12046), .A2(n12112), .B1(n13030), .B2(n12111), .ZN(
        n12115) );
  INV_X1 U13876 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12800) );
  INV_X1 U13877 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12113) );
  OAI22_X1 U13878 ( .A1(n13033), .A2(n12800), .B1(n13032), .B2(n12113), .ZN(
        n12114) );
  OR2_X1 U13879 ( .A1(n12115), .A2(n12114), .ZN(n12120) );
  INV_X1 U13880 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12118) );
  NAND2_X1 U13881 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12117) );
  NAND2_X1 U13882 ( .A1(n13117), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12116) );
  OAI211_X1 U13883 ( .C1(n12118), .C2(n12191), .A(n12117), .B(n12116), .ZN(
        n12119) );
  NOR2_X1 U13884 ( .A1(n12120), .A2(n12119), .ZN(n12130) );
  NAND2_X1 U13885 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12124) );
  AOI22_X1 U13886 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U13887 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12122) );
  NAND2_X1 U13888 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12121) );
  NAND4_X1 U13889 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12128) );
  INV_X1 U13890 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13213) );
  NAND2_X1 U13891 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12126) );
  INV_X1 U13892 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19479) );
  NAND2_X1 U13893 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12125) );
  OAI211_X1 U13894 ( .C1(n13213), .C2(n13026), .A(n12126), .B(n12125), .ZN(
        n12127) );
  NOR2_X1 U13895 ( .A1(n12128), .A2(n12127), .ZN(n12129) );
  NAND2_X1 U13896 ( .A1(n19642), .A2(n12682), .ZN(n12131) );
  INV_X1 U13897 ( .A(n12135), .ZN(n12133) );
  NAND2_X1 U13898 ( .A1(n12134), .A2(n12133), .ZN(n12136) );
  INV_X1 U13899 ( .A(n10991), .ZN(n12172) );
  AOI22_X1 U13900 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12096), .B1(
        n19288), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U13901 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19344), .B1(
        n19333), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U13902 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n15231), .B1(
        n19226), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U13903 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12105), .B1(
        n12106), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12138) );
  NAND4_X1 U13904 ( .A1(n12141), .A2(n12140), .A3(n12139), .A4(n12138), .ZN(
        n12147) );
  AOI22_X1 U13905 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12098), .B1(
        n15140), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U13906 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19360), .B1(
        n19259), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U13907 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12097), .B1(
        n19273), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U13908 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12104), .B1(
        n12099), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12142) );
  NAND4_X1 U13909 ( .A1(n12145), .A2(n12144), .A3(n12143), .A4(n12142), .ZN(
        n12146) );
  INV_X1 U13910 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12149) );
  INV_X1 U13911 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12148) );
  OAI22_X1 U13912 ( .A1(n12046), .A2(n12149), .B1(n13030), .B2(n12148), .ZN(
        n12153) );
  INV_X1 U13913 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12151) );
  INV_X1 U13914 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12150) );
  OAI22_X1 U13915 ( .A1(n13033), .A2(n12151), .B1(n13032), .B2(n12150), .ZN(
        n12152) );
  OR2_X1 U13916 ( .A1(n12153), .A2(n12152), .ZN(n12157) );
  INV_X1 U13917 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13236) );
  NAND2_X1 U13918 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12155) );
  NAND2_X1 U13919 ( .A1(n13117), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12154) );
  OAI211_X1 U13920 ( .C1(n12191), .C2(n13236), .A(n12155), .B(n12154), .ZN(
        n12156) );
  NOR2_X1 U13921 ( .A1(n12157), .A2(n12156), .ZN(n12167) );
  NAND2_X1 U13922 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12161) );
  AOI22_X1 U13923 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12077), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U13924 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13103), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12159) );
  NAND2_X1 U13925 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12158) );
  NAND4_X1 U13926 ( .A1(n12161), .A2(n12160), .A3(n12159), .A4(n12158), .ZN(
        n12165) );
  INV_X1 U13927 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13239) );
  NAND2_X1 U13928 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12163) );
  NAND2_X1 U13929 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12162) );
  OAI211_X1 U13930 ( .C1(n13026), .C2(n13239), .A(n12163), .B(n12162), .ZN(
        n12164) );
  NOR2_X1 U13931 ( .A1(n12165), .A2(n12164), .ZN(n12166) );
  NAND2_X1 U13932 ( .A1(n19642), .A2(n12684), .ZN(n12168) );
  OAI21_X1 U13933 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n11354), .A(
        n12170), .ZN(n12176) );
  INV_X1 U13934 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18693) );
  MUX2_X1 U13935 ( .A(n12183), .B(n18693), .S(n12389), .Z(n12174) );
  OAI21_X1 U13936 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12393), .A(
        n12174), .ZN(n12175) );
  INV_X1 U13937 ( .A(n12177), .ZN(n12178) );
  NAND2_X1 U13938 ( .A1(n12181), .A2(n12393), .ZN(n12182) );
  INV_X1 U13939 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12185) );
  INV_X1 U13940 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15786) );
  OAI22_X1 U13941 ( .A1(n12046), .A2(n12185), .B1(n13030), .B2(n15786), .ZN(
        n12188) );
  INV_X1 U13942 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12833) );
  INV_X1 U13943 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12186) );
  OAI22_X1 U13944 ( .A1(n13033), .A2(n12833), .B1(n13032), .B2(n12186), .ZN(
        n12187) );
  OR2_X1 U13945 ( .A1(n12188), .A2(n12187), .ZN(n12193) );
  INV_X1 U13946 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15783) );
  NAND2_X1 U13947 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12190) );
  NAND2_X1 U13948 ( .A1(n13117), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12189) );
  OAI211_X1 U13949 ( .C1(n12191), .C2(n15783), .A(n12190), .B(n12189), .ZN(
        n12192) );
  NOR2_X1 U13950 ( .A1(n12193), .A2(n12192), .ZN(n12203) );
  NAND2_X1 U13951 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12197) );
  AOI22_X1 U13952 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12077), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U13953 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13103), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12195) );
  NAND2_X1 U13954 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12194) );
  NAND4_X1 U13955 ( .A1(n12197), .A2(n12196), .A3(n12195), .A4(n12194), .ZN(
        n12201) );
  INV_X1 U13956 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15788) );
  NAND2_X1 U13957 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12199) );
  NAND2_X1 U13958 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12198) );
  OAI211_X1 U13959 ( .C1(n15788), .C2(n13026), .A(n12199), .B(n12198), .ZN(
        n12200) );
  NOR2_X1 U13960 ( .A1(n12201), .A2(n12200), .ZN(n12202) );
  XNOR2_X1 U13961 ( .A(n12209), .B(n12535), .ZN(n12204) );
  XNOR2_X1 U13962 ( .A(n12204), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17021) );
  INV_X1 U13963 ( .A(n12204), .ZN(n12205) );
  NAND2_X1 U13964 ( .A1(n12205), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12206) );
  NAND2_X1 U13965 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12408) );
  INV_X1 U13966 ( .A(n12408), .ZN(n12207) );
  INV_X1 U13967 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17000) );
  OAI21_X1 U13968 ( .B1(n12209), .B2(n12535), .A(n17000), .ZN(n12210) );
  AND2_X1 U13969 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16912) );
  AND2_X1 U13970 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16921) );
  AND2_X1 U13971 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12212) );
  NAND3_X1 U13972 ( .A1(n16912), .A2(n16921), .A3(n12212), .ZN(n16857) );
  AND2_X1 U13973 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13338) );
  INV_X1 U13974 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16905) );
  INV_X1 U13975 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15693) );
  INV_X1 U13976 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16907) );
  NOR3_X1 U13977 ( .A1(n16905), .A2(n15693), .A3(n16907), .ZN(n16858) );
  NAND2_X1 U13978 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16858), .ZN(
        n13340) );
  INV_X1 U13979 ( .A(n13340), .ZN(n12213) );
  NAND3_X1 U13980 ( .A1(n13338), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n12213), .ZN(n12214) );
  NOR2_X1 U13981 ( .A1(n16857), .A2(n12214), .ZN(n16833) );
  INV_X1 U13982 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16847) );
  INV_X1 U13983 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16812) );
  INV_X1 U13984 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16597) );
  NOR2_X1 U13985 ( .A1(n16812), .A2(n16597), .ZN(n12215) );
  INV_X1 U13986 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16799) );
  NAND2_X1 U13987 ( .A1(n11144), .A2(n11399), .ZN(n13300) );
  INV_X1 U13988 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15704) );
  NAND2_X1 U13989 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13314) );
  NAND2_X1 U13990 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12216) );
  NOR2_X1 U13991 ( .A1(n13314), .A2(n12216), .ZN(n12923) );
  INV_X1 U13992 ( .A(n12242), .ZN(n12218) );
  NAND2_X1 U13993 ( .A1(n14972), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12217) );
  INV_X1 U13994 ( .A(n12579), .ZN(n12576) );
  MUX2_X1 U13995 ( .A(n12576), .B(n14675), .S(n15291), .Z(n12366) );
  MUX2_X1 U13996 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14986), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12577) );
  INV_X1 U13997 ( .A(n12577), .ZN(n12219) );
  NAND2_X1 U13998 ( .A1(n12219), .A2(n12242), .ZN(n12221) );
  NAND2_X1 U13999 ( .A1(n14986), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12220) );
  NAND2_X1 U14000 ( .A1(n12221), .A2(n12220), .ZN(n12225) );
  XNOR2_X1 U14001 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12224) );
  XNOR2_X1 U14002 ( .A(n12225), .B(n12224), .ZN(n12586) );
  OAI21_X1 U14003 ( .B1(n15291), .B2(n12223), .A(n12222), .ZN(n12356) );
  OAI21_X1 U14004 ( .B1(n12366), .B2(n12577), .A(n12356), .ZN(n12234) );
  NAND2_X1 U14005 ( .A1(n12225), .A2(n12224), .ZN(n12227) );
  NAND2_X1 U14006 ( .A1(n19257), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12226) );
  INV_X1 U14007 ( .A(n12230), .ZN(n12228) );
  XNOR2_X1 U14008 ( .A(n12231), .B(n12228), .ZN(n12240) );
  MUX2_X1 U14009 ( .A(n12240), .B(n12668), .S(n15291), .Z(n12360) );
  NOR2_X1 U14010 ( .A1(n11832), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12229) );
  NOR2_X1 U14011 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17137), .ZN(
        n12232) );
  NAND2_X1 U14012 ( .A1(n12236), .A2(n12232), .ZN(n12241) );
  MUX2_X1 U14013 ( .A(n12241), .B(n12233), .S(n15291), .Z(n12378) );
  NAND3_X1 U14014 ( .A1(n12234), .A2(n12360), .A3(n12378), .ZN(n12239) );
  NAND2_X1 U14015 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17137), .ZN(
        n12235) );
  NAND2_X1 U14016 ( .A1(n12236), .A2(n12235), .ZN(n12238) );
  NAND2_X1 U14017 ( .A1(n18660), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12237) );
  AND2_X1 U14018 ( .A1(n12239), .A2(n12594), .ZN(n15003) );
  AND2_X1 U14019 ( .A1(n19642), .A2(n19703), .ZN(n15030) );
  NAND2_X1 U14020 ( .A1(n15003), .A2(n15030), .ZN(n12597) );
  XNOR2_X1 U14021 ( .A(n12577), .B(n12242), .ZN(n12578) );
  NAND2_X1 U14022 ( .A1(n12244), .A2(n12578), .ZN(n12243) );
  NAND2_X1 U14023 ( .A1(n12244), .A2(n12579), .ZN(n12245) );
  NAND2_X1 U14024 ( .A1(n15004), .A2(n12245), .ZN(n12249) );
  AND2_X1 U14025 ( .A1(n12246), .A2(n18660), .ZN(n18655) );
  INV_X1 U14026 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12247) );
  NAND2_X1 U14027 ( .A1(n12247), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12248) );
  AOI21_X1 U14028 ( .B1(n12046), .B2(n18655), .A(n12248), .ZN(n17420) );
  AOI21_X1 U14029 ( .B1(n12249), .B2(n17057), .A(n17420), .ZN(n17134) );
  NAND2_X1 U14030 ( .A1(n17134), .A2(n15291), .ZN(n12250) );
  NAND2_X1 U14031 ( .A1(n12597), .A2(n12250), .ZN(n12252) );
  INV_X1 U14032 ( .A(n12251), .ZN(n15008) );
  NAND2_X1 U14033 ( .A1(n12252), .A2(n15008), .ZN(n15022) );
  NOR2_X2 U14034 ( .A1(n18721), .A2(n12651), .ZN(n16766) );
  INV_X1 U14035 ( .A(n17419), .ZN(n12253) );
  NOR2_X1 U14036 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n12253), .ZN(n18372) );
  NAND2_X1 U14037 ( .A1(n18372), .A2(n18711), .ZN(n12254) );
  NAND2_X1 U14038 ( .A1(n21597), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12255) );
  NAND2_X1 U14039 ( .A1(n15129), .A2(n12255), .ZN(n14678) );
  NAND2_X1 U14040 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16399), .ZN(
        n16401) );
  INV_X1 U14041 ( .A(n16401), .ZN(n12256) );
  INV_X1 U14042 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16628) );
  INV_X1 U14043 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16407) );
  INV_X1 U14044 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16413) );
  INV_X1 U14045 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15750) );
  INV_X1 U14046 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15276) );
  XNOR2_X1 U14047 ( .A(n15277), .B(n15276), .ZN(n18649) );
  INV_X1 U14048 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n18626) );
  AOI22_X1 U14049 ( .A1(n12622), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12257) );
  OAI21_X1 U14050 ( .B1(n12349), .B2(n18626), .A(n12257), .ZN(n12258) );
  AOI21_X1 U14051 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12337), .A(
        n12258), .ZN(n12351) );
  INV_X1 U14052 ( .A(n12260), .ZN(n12262) );
  NAND2_X1 U14053 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  INV_X1 U14054 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12266) );
  NAND2_X1 U14055 ( .A1(n12622), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12265) );
  NAND2_X1 U14056 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12264) );
  OAI211_X1 U14057 ( .C1(n12349), .C2(n12266), .A(n12265), .B(n12264), .ZN(
        n12267) );
  AOI21_X1 U14058 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n12267), .ZN(n14834) );
  INV_X1 U14059 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U14060 ( .A1(n12337), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12269) );
  AOI22_X1 U14061 ( .A1(n12622), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12268) );
  OAI211_X1 U14062 ( .C1(n12270), .C2(n12349), .A(n12269), .B(n12268), .ZN(
        n14824) );
  INV_X1 U14063 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n12688) );
  NAND2_X1 U14064 ( .A1(n12622), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12272) );
  NAND2_X1 U14065 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12271) );
  OAI211_X1 U14066 ( .C1(n12349), .C2(n12688), .A(n12272), .B(n12271), .ZN(
        n12273) );
  AOI21_X1 U14067 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n12273), .ZN(n15046) );
  INV_X1 U14068 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12710) );
  NAND2_X1 U14069 ( .A1(n12622), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12276) );
  NAND2_X1 U14070 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12275) );
  OAI211_X1 U14071 ( .C1(n12349), .C2(n12710), .A(n12276), .B(n12275), .ZN(
        n12277) );
  AOI21_X1 U14072 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n12277), .ZN(n12278) );
  INV_X1 U14073 ( .A(n12278), .ZN(n15083) );
  NAND2_X1 U14074 ( .A1(n12337), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12285) );
  INV_X1 U14075 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n12281) );
  NAND2_X1 U14076 ( .A1(n12622), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n12280) );
  NAND2_X1 U14077 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12279) );
  OAI211_X1 U14078 ( .C1(n12349), .C2(n12281), .A(n12280), .B(n12279), .ZN(
        n12283) );
  INV_X1 U14079 ( .A(n12283), .ZN(n12284) );
  NAND2_X1 U14080 ( .A1(n12285), .A2(n12284), .ZN(n14897) );
  AND2_X1 U14081 ( .A1(n15083), .A2(n14897), .ZN(n12286) );
  NAND2_X1 U14082 ( .A1(n14896), .A2(n12286), .ZN(n15040) );
  INV_X1 U14083 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n16767) );
  NAND2_X1 U14084 ( .A1(n12622), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12288) );
  NAND2_X1 U14085 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12287) );
  OAI211_X1 U14086 ( .C1(n12349), .C2(n16767), .A(n12288), .B(n12287), .ZN(
        n12289) );
  AOI21_X1 U14087 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12289), .ZN(n15041) );
  INV_X1 U14088 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n16747) );
  NAND2_X1 U14089 ( .A1(n12622), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12292) );
  NAND2_X1 U14090 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12291) );
  OAI211_X1 U14091 ( .C1(n12349), .C2(n16747), .A(n12292), .B(n12291), .ZN(
        n12293) );
  AOI21_X1 U14092 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n12293), .ZN(n15059) );
  INV_X1 U14093 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n18433) );
  NAND2_X1 U14094 ( .A1(n12337), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12295) );
  AOI22_X1 U14095 ( .A1(n12622), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12294) );
  OAI211_X1 U14096 ( .C1(n12349), .C2(n18433), .A(n12295), .B(n12294), .ZN(
        n15108) );
  INV_X1 U14097 ( .A(n15072), .ZN(n12300) );
  INV_X1 U14098 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n17484) );
  NAND2_X1 U14099 ( .A1(n12622), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12297) );
  NAND2_X1 U14100 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12296) );
  OAI211_X1 U14101 ( .C1(n12349), .C2(n17484), .A(n12297), .B(n12296), .ZN(
        n12298) );
  AOI21_X1 U14102 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12298), .ZN(n15073) );
  INV_X1 U14103 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n17485) );
  NAND2_X1 U14104 ( .A1(n12622), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12302) );
  NAND2_X1 U14105 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12301) );
  OAI211_X1 U14106 ( .C1(n12349), .C2(n17485), .A(n12302), .B(n12301), .ZN(
        n12303) );
  AOI21_X1 U14107 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n12303), .ZN(n15119) );
  INV_X1 U14108 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n16697) );
  NAND2_X1 U14109 ( .A1(n12337), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12305) );
  AOI22_X1 U14110 ( .A1(n12622), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12304) );
  OAI211_X1 U14111 ( .C1(n12349), .C2(n16697), .A(n12305), .B(n12304), .ZN(
        n15184) );
  INV_X1 U14112 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n12844) );
  NAND2_X1 U14113 ( .A1(n12622), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12307) );
  NAND2_X1 U14114 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12306) );
  OAI211_X1 U14115 ( .C1(n12349), .C2(n12844), .A(n12307), .B(n12306), .ZN(
        n12308) );
  AOI21_X1 U14116 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12308), .ZN(n12559) );
  INV_X1 U14117 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n17486) );
  NAND2_X1 U14118 ( .A1(n12622), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12311) );
  NAND2_X1 U14119 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12310) );
  OAI211_X1 U14120 ( .C1(n12349), .C2(n17486), .A(n12311), .B(n12310), .ZN(
        n12312) );
  AOI21_X1 U14121 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12312), .ZN(n15315) );
  INV_X1 U14122 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n18498) );
  NAND2_X1 U14123 ( .A1(n12337), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12314) );
  AOI22_X1 U14124 ( .A1(n12622), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12313) );
  OAI211_X1 U14125 ( .C1(n12349), .C2(n18498), .A(n12314), .B(n12313), .ZN(
        n15396) );
  INV_X1 U14126 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n18512) );
  NAND2_X1 U14127 ( .A1(n12337), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12316) );
  AOI22_X1 U14128 ( .A1(n12622), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n12315) );
  OAI211_X1 U14129 ( .C1(n12349), .C2(n18512), .A(n12316), .B(n12315), .ZN(
        n15371) );
  INV_X1 U14130 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n17487) );
  NAND2_X1 U14131 ( .A1(n12622), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U14132 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12317) );
  OAI211_X1 U14133 ( .C1(n12349), .C2(n17487), .A(n12318), .B(n12317), .ZN(
        n12319) );
  AOI21_X1 U14134 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12319), .ZN(n15488) );
  INV_X1 U14135 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n17488) );
  NAND2_X1 U14136 ( .A1(n12622), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12322) );
  NAND2_X1 U14137 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12321) );
  OAI211_X1 U14138 ( .C1(n12349), .C2(n17488), .A(n12322), .B(n12321), .ZN(
        n12323) );
  AOI21_X1 U14139 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12323), .ZN(n15502) );
  INV_X1 U14140 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n13296) );
  NAND2_X1 U14141 ( .A1(n12622), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12325) );
  NAND2_X1 U14142 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12324) );
  OAI211_X1 U14143 ( .C1(n12349), .C2(n13296), .A(n12325), .B(n12324), .ZN(
        n12326) );
  AOI21_X1 U14144 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12326), .ZN(n13294) );
  INV_X1 U14145 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n17489) );
  NAND2_X1 U14146 ( .A1(n12337), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12328) );
  AOI22_X1 U14147 ( .A1(n12622), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n12327) );
  OAI211_X1 U14148 ( .C1(n12349), .C2(n17489), .A(n12328), .B(n12327), .ZN(
        n16519) );
  NAND2_X1 U14149 ( .A1(n16520), .A2(n16519), .ZN(n16522) );
  INV_X1 U14150 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n12331) );
  NAND2_X1 U14151 ( .A1(n12622), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12330) );
  NAND2_X1 U14152 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12329) );
  OAI211_X1 U14153 ( .C1(n12349), .C2(n12331), .A(n12330), .B(n12329), .ZN(
        n12332) );
  AOI21_X1 U14154 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12332), .ZN(n16509) );
  INV_X1 U14155 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n17490) );
  NAND2_X1 U14156 ( .A1(n12622), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12334) );
  NAND2_X1 U14157 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12333) );
  OAI211_X1 U14158 ( .C1(n12349), .C2(n17490), .A(n12334), .B(n12333), .ZN(
        n12335) );
  AOI21_X1 U14159 ( .B1(n12337), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12335), .ZN(n16433) );
  INV_X1 U14160 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n16603) );
  NAND2_X1 U14161 ( .A1(n12337), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12339) );
  AOI22_X1 U14162 ( .A1(n12622), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12338) );
  OAI211_X1 U14163 ( .C1(n12349), .C2(n16603), .A(n12339), .B(n12338), .ZN(
        n16498) );
  INV_X1 U14164 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n17491) );
  NAND2_X1 U14165 ( .A1(n12337), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12341) );
  AOI22_X1 U14166 ( .A1(n12622), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12340) );
  OAI211_X1 U14167 ( .C1(n12349), .C2(n17491), .A(n12341), .B(n12340), .ZN(
        n16491) );
  INV_X1 U14168 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n17492) );
  NAND2_X1 U14169 ( .A1(n12346), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12343) );
  AOI22_X1 U14170 ( .A1(n12622), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12342) );
  OAI211_X1 U14171 ( .C1(n12349), .C2(n17492), .A(n12343), .B(n12342), .ZN(
        n16419) );
  INV_X1 U14172 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n17493) );
  AOI22_X1 U14173 ( .A1(n12622), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12344) );
  OAI21_X1 U14174 ( .B1(n12349), .B2(n17493), .A(n12344), .ZN(n12345) );
  AOI21_X1 U14175 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n12337), .A(
        n12345), .ZN(n13359) );
  INV_X1 U14176 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n17494) );
  NAND2_X1 U14177 ( .A1(n12346), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12348) );
  AOI22_X1 U14178 ( .A1(n12622), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12347) );
  OAI211_X1 U14179 ( .C1(n12349), .C2(n17494), .A(n12348), .B(n12347), .ZN(
        n13303) );
  NAND2_X1 U14180 ( .A1(n13304), .A2(n13303), .ZN(n12350) );
  AOI21_X1 U14181 ( .B1(n12351), .B2(n12350), .A(n12626), .ZN(n18624) );
  AND2_X1 U14182 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12352) );
  NAND2_X2 U14183 ( .A1(n17417), .A2(n12352), .ZN(n17410) );
  INV_X1 U14184 ( .A(n17410), .ZN(n16711) );
  NAND2_X1 U14185 ( .A1(n18624), .A2(n16711), .ZN(n12354) );
  OR2_X1 U14186 ( .A1(n19355), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17394) );
  INV_X2 U14187 ( .A(n18500), .ZN(n18680) );
  NOR2_X1 U14188 ( .A1(n18680), .A2(n18626), .ZN(n15706) );
  AOI21_X1 U14189 ( .B1(n16750), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15706), .ZN(n12353) );
  OAI211_X1 U14190 ( .C1(n16782), .C2(n18649), .A(n12354), .B(n12353), .ZN(
        n12355) );
  AOI21_X1 U14191 ( .B1(n15713), .B2(n16766), .A(n12355), .ZN(n12547) );
  MUX2_X1 U14192 ( .A(n12356), .B(P2_EBX_REG_2__SCAN_IN), .S(n12539), .Z(
        n12370) );
  INV_X1 U14193 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14814) );
  NAND3_X1 U14194 ( .A1(n12539), .A2(n14814), .A3(n14843), .ZN(n12359) );
  NOR2_X2 U14195 ( .A1(n12370), .A2(n11036), .ZN(n12361) );
  MUX2_X1 U14196 ( .A(n12360), .B(n15338), .S(n12539), .Z(n12362) );
  INV_X1 U14197 ( .A(n12382), .ZN(n12365) );
  INV_X1 U14198 ( .A(n12361), .ZN(n12372) );
  INV_X1 U14199 ( .A(n12362), .ZN(n12363) );
  NAND2_X1 U14200 ( .A1(n12372), .A2(n12363), .ZN(n12364) );
  NAND2_X1 U14201 ( .A1(n12365), .A2(n12364), .ZN(n15343) );
  XNOR2_X1 U14202 ( .A(n12376), .B(n15212), .ZN(n15155) );
  MUX2_X1 U14203 ( .A(n12366), .B(n14843), .S(n12539), .Z(n18390) );
  INV_X1 U14204 ( .A(n18390), .ZN(n12367) );
  NAND2_X1 U14205 ( .A1(n12367), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14673) );
  OR3_X1 U14206 ( .A1(n12357), .A2(n14814), .A3(n14843), .ZN(n12368) );
  NAND2_X1 U14207 ( .A1(n11036), .A2(n12368), .ZN(n16468) );
  AND2_X1 U14208 ( .A1(n14673), .A2(n16468), .ZN(n14682) );
  NOR2_X1 U14209 ( .A1(n14673), .A2(n16468), .ZN(n14683) );
  NOR2_X1 U14210 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14683), .ZN(
        n12369) );
  NOR2_X1 U14211 ( .A1(n14682), .A2(n12369), .ZN(n15663) );
  NAND2_X1 U14212 ( .A1(n12370), .A2(n11036), .ZN(n12371) );
  NAND2_X1 U14213 ( .A1(n12372), .A2(n12371), .ZN(n15329) );
  XNOR2_X1 U14214 ( .A(n15329), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15662) );
  NAND2_X1 U14215 ( .A1(n15663), .A2(n15662), .ZN(n12375) );
  INV_X1 U14216 ( .A(n15329), .ZN(n12373) );
  NAND2_X1 U14217 ( .A1(n12373), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12374) );
  NAND2_X1 U14218 ( .A1(n12375), .A2(n12374), .ZN(n15156) );
  NAND2_X1 U14219 ( .A1(n12376), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12377) );
  INV_X1 U14220 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n18396) );
  MUX2_X1 U14221 ( .A(n12378), .B(n18396), .S(n12539), .Z(n12381) );
  XNOR2_X1 U14222 ( .A(n12382), .B(n12381), .ZN(n12379) );
  XNOR2_X1 U14223 ( .A(n12379), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15209) );
  INV_X1 U14224 ( .A(n12379), .ZN(n18398) );
  NAND2_X1 U14225 ( .A1(n18398), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12380) );
  AND2_X2 U14226 ( .A1(n12382), .A2(n12381), .ZN(n12384) );
  INV_X1 U14227 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n15418) );
  INV_X1 U14228 ( .A(n12682), .ZN(n12383) );
  MUX2_X1 U14229 ( .A(n15418), .B(n12383), .S(n12357), .Z(n12385) );
  NAND2_X1 U14230 ( .A1(n12384), .A2(n12385), .ZN(n12396) );
  INV_X1 U14231 ( .A(n12384), .ZN(n12387) );
  INV_X1 U14232 ( .A(n12385), .ZN(n12386) );
  NAND2_X1 U14233 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  NAND2_X1 U14234 ( .A1(n12396), .A2(n12388), .ZN(n15424) );
  NAND2_X1 U14235 ( .A1(n17398), .A2(n17397), .ZN(n12392) );
  NAND2_X1 U14236 ( .A1(n12390), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12391) );
  NAND2_X1 U14237 ( .A1(n12393), .A2(n12535), .ZN(n12394) );
  MUX2_X1 U14238 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n12684), .S(n12357), .Z(
        n12397) );
  XNOR2_X1 U14239 ( .A(n12396), .B(n12397), .ZN(n15366) );
  NAND2_X1 U14240 ( .A1(n12394), .A2(n15366), .ZN(n12409) );
  INV_X1 U14241 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12395) );
  INV_X1 U14242 ( .A(n12396), .ZN(n12399) );
  INV_X1 U14243 ( .A(n12397), .ZN(n12398) );
  NAND2_X1 U14244 ( .A1(n12399), .A2(n12398), .ZN(n12402) );
  INV_X1 U14245 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12401) );
  MUX2_X1 U14246 ( .A(n12401), .B(n12689), .S(n12357), .Z(n12403) );
  XNOR2_X1 U14247 ( .A(n12402), .B(n12403), .ZN(n18414) );
  AND2_X1 U14248 ( .A1(n18414), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17017) );
  INV_X1 U14249 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12404) );
  NOR2_X1 U14250 ( .A1(n12357), .A2(n12404), .ZN(n12406) );
  NAND2_X1 U14251 ( .A1(n12405), .A2(n12406), .ZN(n12407) );
  NAND2_X1 U14252 ( .A1(n12412), .A2(n12407), .ZN(n18422) );
  OR2_X1 U14253 ( .A1(n18422), .A2(n12408), .ZN(n16777) );
  INV_X1 U14254 ( .A(n16777), .ZN(n12417) );
  OR2_X1 U14255 ( .A1(n17017), .A2(n12417), .ZN(n16759) );
  INV_X1 U14256 ( .A(n16759), .ZN(n12410) );
  NAND2_X1 U14257 ( .A1(n12409), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16757) );
  AND2_X1 U14258 ( .A1(n12410), .A2(n16757), .ZN(n12411) );
  NAND2_X1 U14259 ( .A1(n12539), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12413) );
  NAND2_X1 U14260 ( .A1(n12539), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12421) );
  XNOR2_X1 U14261 ( .A(n12423), .B(n12421), .ZN(n15303) );
  NAND2_X1 U14262 ( .A1(n15303), .A2(n12689), .ZN(n12437) );
  INV_X1 U14263 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16977) );
  AND2_X1 U14264 ( .A1(n12437), .A2(n16977), .ZN(n16742) );
  XNOR2_X1 U14265 ( .A(n12412), .B(n12413), .ZN(n15433) );
  AOI21_X1 U14266 ( .B1(n15433), .B2(n12689), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16756) );
  INV_X1 U14267 ( .A(n16756), .ZN(n12418) );
  INV_X1 U14268 ( .A(n18414), .ZN(n12414) );
  INV_X1 U14269 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16999) );
  NAND2_X1 U14270 ( .A1(n12414), .A2(n16999), .ZN(n17016) );
  OR2_X1 U14271 ( .A1(n18422), .A2(n12535), .ZN(n12415) );
  NAND2_X1 U14272 ( .A1(n12415), .A2(n17000), .ZN(n16778) );
  AND2_X1 U14273 ( .A1(n17016), .A2(n16778), .ZN(n12416) );
  OR2_X1 U14274 ( .A1(n12417), .A2(n12416), .ZN(n16760) );
  NAND2_X1 U14275 ( .A1(n12418), .A2(n16760), .ZN(n16740) );
  OR2_X1 U14276 ( .A1(n16742), .A2(n16740), .ZN(n12419) );
  INV_X1 U14277 ( .A(n12419), .ZN(n12420) );
  INV_X1 U14278 ( .A(n12421), .ZN(n12422) );
  NOR2_X2 U14279 ( .A1(n12423), .A2(n12422), .ZN(n12424) );
  NAND2_X1 U14280 ( .A1(n12539), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12425) );
  NAND2_X1 U14281 ( .A1(n12424), .A2(n12425), .ZN(n12432) );
  INV_X1 U14282 ( .A(n12424), .ZN(n12427) );
  INV_X1 U14283 ( .A(n12425), .ZN(n12426) );
  NAND2_X1 U14284 ( .A1(n12427), .A2(n12426), .ZN(n12428) );
  NAND2_X1 U14285 ( .A1(n12432), .A2(n12428), .ZN(n18437) );
  OR2_X1 U14286 ( .A1(n18437), .A2(n12535), .ZN(n12429) );
  INV_X1 U14287 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16965) );
  NAND2_X1 U14288 ( .A1(n12429), .A2(n16965), .ZN(n16730) );
  INV_X1 U14289 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12430) );
  NOR2_X1 U14290 ( .A1(n12357), .A2(n12430), .ZN(n12431) );
  NOR2_X2 U14291 ( .A1(n12432), .A2(n12431), .ZN(n12440) );
  INV_X1 U14292 ( .A(n12440), .ZN(n12473) );
  NAND2_X1 U14293 ( .A1(n12432), .A2(n12431), .ZN(n12433) );
  AND2_X1 U14294 ( .A1(n12473), .A2(n12433), .ZN(n12439) );
  AND2_X1 U14295 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12434) );
  NAND2_X1 U14296 ( .A1(n12439), .A2(n12434), .ZN(n16718) );
  NAND2_X1 U14297 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12435) );
  OR2_X1 U14298 ( .A1(n18437), .A2(n12435), .ZN(n16729) );
  INV_X1 U14299 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16991) );
  NOR2_X1 U14300 ( .A1(n12535), .A2(n16991), .ZN(n12436) );
  NAND2_X1 U14301 ( .A1(n15433), .A2(n12436), .ZN(n16754) );
  OR2_X1 U14302 ( .A1(n12437), .A2(n16977), .ZN(n16743) );
  NAND2_X1 U14303 ( .A1(n16754), .A2(n16743), .ZN(n16731) );
  INV_X1 U14304 ( .A(n16731), .ZN(n12438) );
  AND2_X1 U14305 ( .A1(n16729), .A2(n12438), .ZN(n16716) );
  NAND2_X1 U14306 ( .A1(n16718), .A2(n16716), .ZN(n13277) );
  INV_X1 U14307 ( .A(n12439), .ZN(n18447) );
  INV_X1 U14308 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16714) );
  OAI21_X1 U14309 ( .B1(n18447), .B2(n12535), .A(n16714), .ZN(n16719) );
  NAND2_X1 U14310 ( .A1(n12539), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12471) );
  INV_X1 U14311 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12441) );
  NOR2_X1 U14312 ( .A1(n12357), .A2(n12441), .ZN(n12468) );
  INV_X1 U14313 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12442) );
  NAND2_X1 U14314 ( .A1(n12539), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12458) );
  AND2_X2 U14315 ( .A1(n12457), .A2(n12458), .ZN(n12456) );
  NAND2_X1 U14316 ( .A1(n12539), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12462) );
  NAND2_X1 U14317 ( .A1(n12456), .A2(n12462), .ZN(n12466) );
  INV_X1 U14318 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n12443) );
  NOR2_X1 U14319 ( .A1(n12357), .A2(n12443), .ZN(n12453) );
  OR2_X2 U14320 ( .A1(n12466), .A2(n12453), .ZN(n12455) );
  INV_X1 U14321 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12444) );
  NOR2_X1 U14322 ( .A1(n12357), .A2(n12444), .ZN(n12449) );
  NAND2_X1 U14323 ( .A1(n12539), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12445) );
  INV_X1 U14324 ( .A(n12445), .ZN(n12446) );
  NAND2_X1 U14325 ( .A1(n11041), .A2(n12446), .ZN(n12447) );
  NAND2_X1 U14326 ( .A1(n11038), .A2(n11080), .ZN(n12448) );
  NAND2_X1 U14327 ( .A1(n11026), .A2(n12448), .ZN(n16454) );
  NOR2_X1 U14328 ( .A1(n16454), .A2(n12535), .ZN(n12478) );
  OR2_X1 U14329 ( .A1(n12478), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13288) );
  NAND2_X1 U14330 ( .A1(n12455), .A2(n12449), .ZN(n12450) );
  NAND2_X1 U14331 ( .A1(n11041), .A2(n12450), .ZN(n18530) );
  OR2_X1 U14332 ( .A1(n18530), .A2(n12535), .ZN(n12452) );
  INV_X1 U14333 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12451) );
  NAND2_X1 U14334 ( .A1(n12452), .A2(n12451), .ZN(n16653) );
  NAND2_X1 U14335 ( .A1(n12466), .A2(n12453), .ZN(n12454) );
  AND2_X1 U14336 ( .A1(n12455), .A2(n12454), .ZN(n18511) );
  NAND2_X1 U14337 ( .A1(n18511), .A2(n12689), .ZN(n12481) );
  INV_X1 U14338 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16891) );
  NAND2_X1 U14339 ( .A1(n12481), .A2(n16891), .ZN(n16663) );
  NAND2_X1 U14340 ( .A1(n16653), .A2(n16663), .ZN(n13285) );
  XNOR2_X1 U14341 ( .A(n12470), .B(n11078), .ZN(n15463) );
  AOI21_X1 U14342 ( .B1(n15463), .B2(n12689), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12555) );
  INV_X1 U14343 ( .A(n12456), .ZN(n12464) );
  INV_X1 U14344 ( .A(n12457), .ZN(n12460) );
  INV_X1 U14345 ( .A(n12458), .ZN(n12459) );
  NAND2_X1 U14346 ( .A1(n12460), .A2(n12459), .ZN(n12461) );
  NAND2_X1 U14347 ( .A1(n18482), .A2(n12689), .ZN(n12489) );
  XNOR2_X1 U14348 ( .A(n12489), .B(n16905), .ZN(n15697) );
  INV_X1 U14349 ( .A(n12462), .ZN(n12463) );
  NAND2_X1 U14350 ( .A1(n12464), .A2(n12463), .ZN(n12465) );
  NAND2_X1 U14351 ( .A1(n12466), .A2(n12465), .ZN(n18502) );
  OR2_X1 U14352 ( .A1(n18502), .A2(n12535), .ZN(n12467) );
  NAND2_X1 U14353 ( .A1(n12467), .A2(n16907), .ZN(n16671) );
  NAND2_X1 U14354 ( .A1(n12475), .A2(n12468), .ZN(n12469) );
  NAND2_X1 U14355 ( .A1(n12470), .A2(n12469), .ZN(n18471) );
  INV_X1 U14356 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16920) );
  OAI21_X1 U14357 ( .B1(n18471), .B2(n12535), .A(n16920), .ZN(n12554) );
  INV_X1 U14358 ( .A(n12471), .ZN(n12472) );
  NAND2_X1 U14359 ( .A1(n12473), .A2(n12472), .ZN(n12474) );
  NAND2_X1 U14360 ( .A1(n12475), .A2(n12474), .ZN(n18462) );
  OR2_X1 U14361 ( .A1(n18462), .A2(n12535), .ZN(n12485) );
  INV_X1 U14362 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16938) );
  NAND2_X1 U14363 ( .A1(n12485), .A2(n16938), .ZN(n16702) );
  AND2_X1 U14364 ( .A1(n12554), .A2(n16702), .ZN(n13276) );
  NAND2_X1 U14365 ( .A1(n16671), .A2(n13276), .ZN(n12476) );
  NOR4_X1 U14366 ( .A1(n13285), .A2(n12555), .A3(n15697), .A4(n12476), .ZN(
        n12477) );
  OAI211_X1 U14367 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n13286), .A(
        n13288), .B(n12477), .ZN(n12494) );
  INV_X1 U14368 ( .A(n12478), .ZN(n12480) );
  INV_X1 U14369 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12479) );
  INV_X1 U14370 ( .A(n12481), .ZN(n12482) );
  NAND2_X1 U14371 ( .A1(n12482), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16661) );
  NAND2_X1 U14372 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12483) );
  OR2_X2 U14373 ( .A1(n18530), .A2(n12483), .ZN(n16652) );
  AND2_X1 U14374 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12484) );
  NAND2_X1 U14375 ( .A1(n15463), .A2(n12484), .ZN(n12556) );
  INV_X1 U14376 ( .A(n12485), .ZN(n12486) );
  NAND2_X1 U14377 ( .A1(n12486), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16703) );
  INV_X1 U14378 ( .A(n18471), .ZN(n12488) );
  AND2_X1 U14379 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12487) );
  NAND2_X1 U14380 ( .A1(n12488), .A2(n12487), .ZN(n12553) );
  AND3_X1 U14381 ( .A1(n12556), .A2(n16703), .A3(n12553), .ZN(n13279) );
  INV_X1 U14382 ( .A(n12489), .ZN(n12490) );
  NAND2_X1 U14383 ( .A1(n12490), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16672) );
  NAND2_X1 U14384 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12491) );
  OR2_X1 U14385 ( .A1(n18502), .A2(n12491), .ZN(n16670) );
  AND2_X1 U14386 ( .A1(n16672), .A2(n16670), .ZN(n13283) );
  NAND4_X1 U14387 ( .A1(n16661), .A2(n16652), .A3(n13279), .A4(n13283), .ZN(
        n12492) );
  AOI21_X1 U14388 ( .B1(n13286), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12492), .ZN(n12493) );
  INV_X1 U14389 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n12495) );
  NOR2_X1 U14390 ( .A1(n12357), .A2(n12495), .ZN(n12496) );
  NAND2_X1 U14391 ( .A1(n11026), .A2(n12496), .ZN(n12497) );
  NAND2_X1 U14392 ( .A1(n12499), .A2(n12497), .ZN(n18551) );
  OR2_X1 U14393 ( .A1(n18551), .A2(n12535), .ZN(n12498) );
  NOR2_X1 U14394 ( .A1(n12498), .A2(n16847), .ZN(n16637) );
  NAND2_X1 U14395 ( .A1(n12498), .A2(n16847), .ZN(n16635) );
  NAND2_X1 U14396 ( .A1(n12539), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12502) );
  XNOR2_X1 U14397 ( .A(n12499), .B(n12502), .ZN(n18563) );
  NAND2_X1 U14398 ( .A1(n18563), .A2(n12689), .ZN(n12500) );
  INV_X1 U14399 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16834) );
  AND2_X1 U14400 ( .A1(n12500), .A2(n16834), .ZN(n16625) );
  INV_X1 U14401 ( .A(n12500), .ZN(n12501) );
  NAND2_X1 U14402 ( .A1(n12501), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16624) );
  NAND2_X1 U14403 ( .A1(n12503), .A2(n12502), .ZN(n12506) );
  INV_X1 U14404 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n12504) );
  NOR2_X1 U14405 ( .A1(n12357), .A2(n12504), .ZN(n12505) );
  NAND2_X1 U14406 ( .A1(n12506), .A2(n12505), .ZN(n12507) );
  NAND2_X1 U14407 ( .A1(n12511), .A2(n12507), .ZN(n16442) );
  OR2_X1 U14408 ( .A1(n16442), .A2(n12535), .ZN(n12508) );
  NOR2_X1 U14409 ( .A1(n12508), .A2(n16597), .ZN(n16614) );
  NAND2_X1 U14410 ( .A1(n12508), .A2(n16597), .ZN(n16612) );
  INV_X1 U14411 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n12509) );
  NAND2_X1 U14412 ( .A1(n12539), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12513) );
  XNOR2_X1 U14413 ( .A(n12515), .B(n12513), .ZN(n18584) );
  NAND2_X1 U14414 ( .A1(n18584), .A2(n12689), .ZN(n12510) );
  XOR2_X1 U14415 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n12510), .Z(
        n16587) );
  XNOR2_X1 U14416 ( .A(n12511), .B(n11091), .ZN(n18573) );
  AOI21_X1 U14417 ( .B1(n18573), .B2(n12689), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16601) );
  INV_X1 U14418 ( .A(n12513), .ZN(n12514) );
  NAND2_X1 U14419 ( .A1(n12539), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12519) );
  INV_X1 U14420 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n18597) );
  NOR2_X1 U14421 ( .A1(n12357), .A2(n18597), .ZN(n12516) );
  NAND2_X1 U14422 ( .A1(n12523), .A2(n12516), .ZN(n12517) );
  NAND2_X1 U14423 ( .A1(n12533), .A2(n12517), .ZN(n18595) );
  INV_X1 U14424 ( .A(n12518), .ZN(n12521) );
  INV_X1 U14425 ( .A(n12519), .ZN(n12520) );
  NAND2_X1 U14426 ( .A1(n12521), .A2(n12520), .ZN(n12522) );
  NAND2_X1 U14427 ( .A1(n12523), .A2(n12522), .ZN(n16429) );
  NOR2_X1 U14428 ( .A1(n16429), .A2(n12535), .ZN(n13352) );
  NAND2_X1 U14429 ( .A1(n13351), .A2(n12524), .ZN(n12525) );
  INV_X1 U14430 ( .A(n12526), .ZN(n12527) );
  OAI21_X1 U14431 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n12527), .ZN(n12530) );
  NAND3_X1 U14432 ( .A1(n18584), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n12689), .ZN(n12529) );
  AND2_X1 U14433 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12528) );
  NAND2_X1 U14434 ( .A1(n18573), .A2(n12528), .ZN(n16599) );
  AND2_X1 U14435 ( .A1(n12529), .A2(n16599), .ZN(n13350) );
  NAND2_X1 U14436 ( .A1(n12539), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12537) );
  XNOR2_X1 U14437 ( .A(n12538), .B(n12537), .ZN(n12536) );
  INV_X1 U14438 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12534) );
  OAI21_X1 U14439 ( .B1(n12536), .B2(n12535), .A(n12534), .ZN(n13308) );
  NAND2_X1 U14440 ( .A1(n13310), .A2(n13308), .ZN(n12570) );
  INV_X1 U14441 ( .A(n12536), .ZN(n18612) );
  NAND3_X1 U14442 ( .A1(n18612), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12689), .ZN(n13309) );
  NAND2_X1 U14443 ( .A1(n12570), .A2(n13309), .ZN(n12544) );
  NAND2_X1 U14444 ( .A1(n12538), .A2(n12537), .ZN(n12571) );
  NAND2_X1 U14445 ( .A1(n12539), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12540) );
  XNOR2_X1 U14446 ( .A(n12571), .B(n12540), .ZN(n18633) );
  AOI21_X1 U14447 ( .B1(n18633), .B2(n12689), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12569) );
  AND2_X1 U14448 ( .A1(n12689), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12541) );
  NAND2_X1 U14449 ( .A1(n18633), .A2(n12541), .ZN(n12568) );
  INV_X1 U14450 ( .A(n12568), .ZN(n12542) );
  NOR2_X1 U14451 ( .A1(n12569), .A2(n12542), .ZN(n12543) );
  INV_X1 U14452 ( .A(n18721), .ZN(n12545) );
  INV_X1 U14453 ( .A(n16912), .ZN(n16914) );
  INV_X1 U14454 ( .A(n16921), .ZN(n12548) );
  NOR2_X2 U14455 ( .A1(n16705), .A2(n12548), .ZN(n16692) );
  NOR2_X1 U14456 ( .A1(n15716), .A2(n17408), .ZN(n12567) );
  INV_X1 U14457 ( .A(n12550), .ZN(n12552) );
  INV_X1 U14458 ( .A(n16703), .ZN(n12551) );
  OAI21_X1 U14459 ( .B1(n12552), .B2(n12551), .A(n16702), .ZN(n16696) );
  AND2_X1 U14460 ( .A1(n12554), .A2(n12553), .ZN(n16695) );
  NAND2_X1 U14461 ( .A1(n16696), .A2(n16695), .ZN(n16694) );
  NAND2_X1 U14462 ( .A1(n16694), .A2(n12554), .ZN(n12558) );
  INV_X1 U14463 ( .A(n12555), .ZN(n13281) );
  NAND2_X1 U14464 ( .A1(n13281), .A2(n12556), .ZN(n12557) );
  XNOR2_X1 U14465 ( .A(n12558), .B(n12557), .ZN(n15728) );
  NAND2_X1 U14466 ( .A1(n15186), .A2(n12559), .ZN(n12560) );
  NOR2_X1 U14467 ( .A1(n12561), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12562) );
  OR2_X1 U14468 ( .A1(n16398), .A2(n12562), .ZN(n15466) );
  NAND2_X1 U14469 ( .A1(n18532), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15718) );
  NAND2_X1 U14470 ( .A1(n16750), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12563) );
  OAI211_X1 U14471 ( .C1(n16782), .C2(n15466), .A(n15718), .B(n12563), .ZN(
        n12564) );
  AOI21_X1 U14472 ( .B1(n15717), .B2(n16711), .A(n12564), .ZN(n12565) );
  OAI21_X1 U14473 ( .B1(n12570), .B2(n12569), .A(n11410), .ZN(n12575) );
  NOR2_X1 U14474 ( .A1(n12571), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12572) );
  MUX2_X1 U14475 ( .A(n12405), .B(n12572), .S(n12539), .Z(n18643) );
  NAND2_X1 U14476 ( .A1(n18643), .A2(n12689), .ZN(n12573) );
  XNOR2_X1 U14477 ( .A(n12573), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12574) );
  XNOR2_X1 U14478 ( .A(n12575), .B(n12574), .ZN(n15767) );
  NAND2_X1 U14479 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n18716) );
  NAND2_X2 U14480 ( .A1(n17495), .A2(n21640), .ZN(n17496) );
  NOR2_X1 U14481 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n17129) );
  NAND2_X1 U14482 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17129), .ZN(n17477) );
  NAND2_X1 U14483 ( .A1(n18716), .A2(n21630), .ZN(n15029) );
  INV_X1 U14484 ( .A(n15029), .ZN(n15014) );
  NAND2_X1 U14485 ( .A1(n17083), .A2(n15014), .ZN(n12619) );
  NOR2_X1 U14486 ( .A1(n12577), .A2(n12576), .ZN(n12581) );
  OAI211_X1 U14487 ( .C1(n12651), .C2(n12579), .A(n12627), .B(n12578), .ZN(
        n12580) );
  OAI21_X1 U14488 ( .B1(n15000), .B2(n12581), .A(n12580), .ZN(n12583) );
  NAND2_X1 U14489 ( .A1(n12583), .A2(n12582), .ZN(n12584) );
  OAI21_X1 U14490 ( .B1(n12585), .B2(n18656), .A(n12584), .ZN(n12592) );
  NAND2_X1 U14491 ( .A1(n18377), .A2(n12651), .ZN(n12587) );
  MUX2_X1 U14492 ( .A(n12587), .B(n15000), .S(n12223), .Z(n12591) );
  NAND2_X1 U14493 ( .A1(n15291), .A2(n12588), .ZN(n12589) );
  NAND2_X1 U14494 ( .A1(n12589), .A2(n12594), .ZN(n12590) );
  AOI21_X1 U14495 ( .B1(n12592), .B2(n12591), .A(n12590), .ZN(n12593) );
  MUX2_X1 U14496 ( .A(n18660), .B(n12593), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n12614) );
  OR2_X1 U14497 ( .A1(n15128), .A2(n19642), .ZN(n14949) );
  NAND2_X1 U14498 ( .A1(n17134), .A2(n12651), .ZN(n12596) );
  NAND2_X1 U14499 ( .A1(n12597), .A2(n12596), .ZN(n12598) );
  NAND2_X1 U14500 ( .A1(n12598), .A2(n15008), .ZN(n12613) );
  NAND2_X1 U14501 ( .A1(n12601), .A2(n12600), .ZN(n12602) );
  NAND2_X1 U14502 ( .A1(n12599), .A2(n12602), .ZN(n12608) );
  AOI21_X1 U14503 ( .B1(n19703), .B2(n12635), .A(n17083), .ZN(n12603) );
  OR2_X1 U14504 ( .A1(n11884), .A2(n12651), .ZN(n12887) );
  AOI21_X1 U14505 ( .B1(n12603), .B2(n12887), .A(n12895), .ZN(n12607) );
  NAND2_X1 U14506 ( .A1(n12604), .A2(n12635), .ZN(n12605) );
  NAND2_X1 U14507 ( .A1(n12605), .A2(n15030), .ZN(n12900) );
  NAND4_X1 U14508 ( .A1(n12608), .A2(n12607), .A3(n12900), .A4(n12606), .ZN(
        n12888) );
  NOR2_X1 U14509 ( .A1(n11881), .A2(n15029), .ZN(n12609) );
  AND2_X1 U14510 ( .A1(n15004), .A2(n12609), .ZN(n12610) );
  NOR2_X1 U14511 ( .A1(n12888), .A2(n12610), .ZN(n14953) );
  MUX2_X1 U14512 ( .A(n15031), .B(n17083), .S(n19642), .Z(n12611) );
  NAND3_X1 U14513 ( .A1(n12611), .A2(n15004), .A3(n18716), .ZN(n12612) );
  OAI21_X1 U14514 ( .B1(n12614), .B2(n19703), .A(n12894), .ZN(n12615) );
  INV_X1 U14515 ( .A(n12615), .ZN(n12616) );
  NAND2_X1 U14516 ( .A1(n14949), .A2(n12616), .ZN(n12617) );
  OAI211_X1 U14517 ( .C1(n12619), .C2(n14949), .A(n12618), .B(n12617), .ZN(
        n12620) );
  NOR2_X1 U14518 ( .A1(n12251), .A2(n15000), .ZN(n12621) );
  INV_X1 U14519 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15280) );
  AOI22_X1 U14520 ( .A1(n12622), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12624) );
  NAND2_X1 U14521 ( .A1(n10980), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12623) );
  OAI211_X1 U14522 ( .C1(n11916), .C2(n15280), .A(n12624), .B(n12623), .ZN(
        n12625) );
  XNOR2_X1 U14523 ( .A(n12626), .B(n12625), .ZN(n16472) );
  INV_X1 U14524 ( .A(n12884), .ZN(n14568) );
  OR2_X1 U14525 ( .A1(n12628), .A2(n14568), .ZN(n14981) );
  NAND2_X1 U14526 ( .A1(n14981), .A2(n19642), .ZN(n12631) );
  INV_X1 U14527 ( .A(n12629), .ZN(n12630) );
  NAND2_X1 U14528 ( .A1(n12631), .A2(n12630), .ZN(n12632) );
  NOR2_X1 U14529 ( .A1(n12635), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12638) );
  AOI22_X1 U14530 ( .A1(n12875), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12636) );
  OAI21_X1 U14531 ( .B1(n12878), .B2(n18512), .A(n12636), .ZN(n15403) );
  AND2_X1 U14532 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12639) );
  NOR2_X1 U14533 ( .A1(n12638), .A2(n12639), .ZN(n12640) );
  INV_X1 U14534 ( .A(n11886), .ZN(n13259) );
  NAND2_X1 U14535 ( .A1(n13259), .A2(n12647), .ZN(n12661) );
  INV_X1 U14536 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19685) );
  NAND2_X1 U14537 ( .A1(n12641), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12642) );
  OAI211_X1 U14538 ( .C1(n12635), .C2(n19685), .A(n12642), .B(n12654), .ZN(
        n12643) );
  INV_X1 U14539 ( .A(n12643), .ZN(n12644) );
  OAI21_X1 U14540 ( .B1(n12878), .B2(n12645), .A(n12644), .ZN(n18385) );
  NAND2_X1 U14541 ( .A1(n18386), .A2(n18385), .ZN(n12658) );
  INV_X1 U14542 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U14543 ( .A1(n12638), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12647), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12648) );
  INV_X1 U14544 ( .A(n12659), .ZN(n12650) );
  XNOR2_X1 U14545 ( .A(n12658), .B(n12650), .ZN(n16461) );
  INV_X1 U14546 ( .A(n12635), .ZN(n14813) );
  OAI22_X1 U14547 ( .A1(n12652), .A2(n12651), .B1(n14813), .B2(n13259), .ZN(
        n12653) );
  INV_X1 U14548 ( .A(n12653), .ZN(n12655) );
  NAND2_X1 U14549 ( .A1(n16461), .A2(n16460), .ZN(n16465) );
  NAND2_X1 U14550 ( .A1(n12659), .A2(n12658), .ZN(n12660) );
  NAND2_X1 U14551 ( .A1(n16465), .A2(n12660), .ZN(n12665) );
  NAND2_X1 U14552 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12662) );
  OAI211_X1 U14553 ( .C1(n12826), .C2(n12663), .A(n12662), .B(n12661), .ZN(
        n12664) );
  XNOR2_X1 U14554 ( .A(n12665), .B(n12664), .ZN(n15325) );
  AOI222_X1 U14555 ( .A1(n12870), .A2(P2_REIP_REG_2__SCAN_IN), .B1(n12875), 
        .B2(P2_EAX_REG_2__SCAN_IN), .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), 
        .C2(n12647), .ZN(n15324) );
  INV_X1 U14556 ( .A(n12664), .ZN(n12666) );
  NAND2_X1 U14557 ( .A1(n12666), .A2(n12665), .ZN(n12667) );
  NAND2_X1 U14558 ( .A1(n12870), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12674) );
  NAND2_X1 U14559 ( .A1(n12846), .A2(n12668), .ZN(n12673) );
  INV_X1 U14560 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17436) );
  NAND2_X1 U14561 ( .A1(n12875), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12670) );
  NAND2_X1 U14562 ( .A1(n12647), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12669) );
  OAI211_X1 U14563 ( .C1(n17436), .C2(n12654), .A(n12670), .B(n12669), .ZN(
        n12671) );
  INV_X1 U14564 ( .A(n12671), .ZN(n12672) );
  AOI22_X1 U14565 ( .A1(n12870), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n12875), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12678) );
  OAI22_X1 U14566 ( .A1(n12826), .A2(n12675), .B1(n12679), .B2(n18678), .ZN(
        n12676) );
  INV_X1 U14567 ( .A(n12676), .ZN(n12677) );
  NAND2_X1 U14568 ( .A1(n12678), .A2(n12677), .ZN(n15215) );
  INV_X1 U14569 ( .A(n15412), .ZN(n12683) );
  NAND2_X1 U14570 ( .A1(n12870), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U14571 ( .A1(n12875), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12647), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12680) );
  OAI211_X1 U14572 ( .C1(n12682), .C2(n12826), .A(n12681), .B(n12680), .ZN(
        n15410) );
  NAND2_X1 U14573 ( .A1(n12683), .A2(n15410), .ZN(n15414) );
  INV_X1 U14574 ( .A(n12684), .ZN(n12685) );
  NAND2_X1 U14575 ( .A1(n12846), .A2(n12685), .ZN(n12686) );
  NAND2_X1 U14576 ( .A1(n15414), .A2(n12686), .ZN(n15353) );
  AOI22_X1 U14577 ( .A1(n12875), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12647), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12687) );
  OAI21_X1 U14578 ( .B1(n12878), .B2(n12688), .A(n12687), .ZN(n15352) );
  AOI21_X1 U14579 ( .B1(n12846), .B2(n12689), .A(n15355), .ZN(n17030) );
  AOI222_X1 U14580 ( .A1(n12870), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n12875), 
        .B2(P2_EAX_REG_7__SCAN_IN), .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), 
        .C2(n12647), .ZN(n17029) );
  NAND2_X1 U14581 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12693) );
  AOI22_X1 U14582 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12692) );
  AOI22_X1 U14583 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12691) );
  NAND2_X1 U14584 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12690) );
  NAND4_X1 U14585 ( .A1(n12693), .A2(n12692), .A3(n12691), .A4(n12690), .ZN(
        n12698) );
  NAND2_X1 U14586 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12695) );
  NAND2_X1 U14587 ( .A1(n13117), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12694) );
  OAI211_X1 U14588 ( .C1(n12696), .C2(n13026), .A(n12695), .B(n12694), .ZN(
        n12697) );
  NOR2_X1 U14589 ( .A1(n12698), .A2(n12697), .ZN(n12707) );
  INV_X1 U14590 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12699) );
  INV_X1 U14591 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13093) );
  OAI22_X1 U14592 ( .A1(n12046), .A2(n12699), .B1(n13030), .B2(n13093), .ZN(
        n12703) );
  INV_X1 U14593 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12700) );
  OAI22_X1 U14594 ( .A1(n13033), .A2(n12701), .B1(n13032), .B2(n12700), .ZN(
        n12702) );
  NOR2_X1 U14595 ( .A1(n12703), .A2(n12702), .ZN(n12706) );
  AOI22_X1 U14596 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13022), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12705) );
  NAND2_X1 U14597 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12704) );
  NAND4_X1 U14598 ( .A1(n12707), .A2(n12706), .A3(n12705), .A4(n12704), .ZN(
        n15086) );
  NAND2_X1 U14599 ( .A1(n12846), .A2(n15086), .ZN(n12709) );
  AOI22_X1 U14600 ( .A1(n12875), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12647), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12708) );
  OAI211_X1 U14601 ( .C1(n12878), .C2(n12710), .A(n12709), .B(n12708), .ZN(
        n17006) );
  AOI22_X1 U14602 ( .A1(n13114), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U14603 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n13115), .ZN(n12713) );
  AOI22_X1 U14604 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12712) );
  NAND2_X1 U14605 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12711) );
  AND4_X1 U14606 ( .A1(n12714), .A2(n12713), .A3(n12712), .A4(n12711), .ZN(
        n12725) );
  NAND2_X1 U14607 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12718) );
  AOI22_X1 U14608 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12077), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U14609 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13103), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12716) );
  NAND2_X1 U14610 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12715) );
  NAND4_X1 U14611 ( .A1(n12718), .A2(n12717), .A3(n12716), .A4(n12715), .ZN(
        n12723) );
  NAND2_X1 U14612 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12720) );
  NAND2_X1 U14613 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12719) );
  OAI211_X1 U14614 ( .C1(n13026), .C2(n12721), .A(n12720), .B(n12719), .ZN(
        n12722) );
  NOR2_X1 U14615 ( .A1(n12723), .A2(n12722), .ZN(n12724) );
  NAND2_X1 U14616 ( .A1(n12870), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U14617 ( .A1(n12875), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12647), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12726) );
  OAI211_X1 U14618 ( .C1(n15054), .C2(n12826), .A(n12727), .B(n12726), .ZN(
        n15427) );
  NAND2_X1 U14619 ( .A1(n12870), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12745) );
  AOI22_X1 U14620 ( .A1(n13114), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12731) );
  AOI22_X1 U14621 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13115), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U14622 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U14623 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12728) );
  AND4_X1 U14624 ( .A1(n12731), .A2(n12730), .A3(n12729), .A4(n12728), .ZN(
        n12742) );
  NAND2_X1 U14625 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12735) );
  AOI22_X1 U14626 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U14627 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12733) );
  NAND2_X1 U14628 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12732) );
  NAND4_X1 U14629 ( .A1(n12735), .A2(n12734), .A3(n12733), .A4(n12732), .ZN(
        n12740) );
  NAND2_X1 U14630 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12737) );
  NAND2_X1 U14631 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12736) );
  OAI211_X1 U14632 ( .C1(n12738), .C2(n13026), .A(n12737), .B(n12736), .ZN(
        n12739) );
  NOR2_X1 U14633 ( .A1(n12740), .A2(n12739), .ZN(n12741) );
  AND2_X1 U14634 ( .A1(n12742), .A2(n12741), .ZN(n12967) );
  INV_X1 U14635 ( .A(n12967), .ZN(n15056) );
  NAND2_X1 U14636 ( .A1(n12846), .A2(n15056), .ZN(n12744) );
  AOI22_X1 U14637 ( .A1(n12875), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U14638 ( .A1(n13114), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U14639 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13115), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U14640 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12747) );
  NAND2_X1 U14641 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12746) );
  AND4_X1 U14642 ( .A1(n12749), .A2(n12748), .A3(n12747), .A4(n12746), .ZN(
        n12760) );
  NAND2_X1 U14643 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12753) );
  AOI22_X1 U14644 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U14645 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12751) );
  NAND2_X1 U14646 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12750) );
  NAND4_X1 U14647 ( .A1(n12753), .A2(n12752), .A3(n12751), .A4(n12750), .ZN(
        n12758) );
  NAND2_X1 U14648 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12755) );
  NAND2_X1 U14649 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12754) );
  OAI211_X1 U14650 ( .C1(n12756), .C2(n13026), .A(n12755), .B(n12754), .ZN(
        n12757) );
  NOR2_X1 U14651 ( .A1(n12758), .A2(n12757), .ZN(n12759) );
  NAND2_X1 U14652 ( .A1(n12870), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U14653 ( .A1(n12875), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12761) );
  OAI211_X1 U14654 ( .C1(n15112), .C2(n12826), .A(n12762), .B(n12761), .ZN(
        n16957) );
  NAND2_X1 U14655 ( .A1(n12870), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12788) );
  INV_X1 U14656 ( .A(n12763), .ZN(n12819) );
  INV_X1 U14657 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12764) );
  INV_X1 U14658 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13200) );
  OAI22_X1 U14659 ( .A1(n12819), .A2(n12764), .B1(n13030), .B2(n13200), .ZN(
        n12769) );
  INV_X1 U14660 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12767) );
  INV_X1 U14661 ( .A(n13117), .ZN(n12766) );
  INV_X1 U14662 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12765) );
  OAI22_X1 U14663 ( .A1(n12767), .A2(n13112), .B1(n12766), .B2(n12765), .ZN(
        n12768) );
  NOR2_X1 U14664 ( .A1(n12769), .A2(n12768), .ZN(n12785) );
  NAND2_X1 U14665 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12773) );
  AOI22_X1 U14666 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12077), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12772) );
  AOI22_X1 U14667 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n13103), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12771) );
  NAND2_X1 U14668 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12770) );
  AND4_X1 U14669 ( .A1(n12773), .A2(n12772), .A3(n12771), .A4(n12770), .ZN(
        n12784) );
  NAND2_X1 U14670 ( .A1(n13108), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12775) );
  NAND2_X1 U14671 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12774) );
  OAI211_X1 U14672 ( .C1(n13033), .C2(n12776), .A(n12775), .B(n12774), .ZN(
        n12777) );
  INV_X1 U14673 ( .A(n12777), .ZN(n12783) );
  NAND2_X1 U14674 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12779) );
  NAND2_X1 U14675 ( .A1(n13113), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12778) );
  OAI211_X1 U14676 ( .C1(n12046), .C2(n12780), .A(n12779), .B(n12778), .ZN(
        n12781) );
  INV_X1 U14677 ( .A(n12781), .ZN(n12782) );
  NAND4_X1 U14678 ( .A1(n12785), .A2(n12784), .A3(n12783), .A4(n12782), .ZN(
        n15079) );
  NAND2_X1 U14679 ( .A1(n12846), .A2(n15079), .ZN(n12787) );
  AOI22_X1 U14680 ( .A1(n12875), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12786) );
  NAND2_X1 U14681 ( .A1(n12789), .A2(n11411), .ZN(n16931) );
  NAND2_X1 U14682 ( .A1(n12870), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U14683 ( .A1(n13114), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U14684 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13115), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U14685 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12791) );
  NAND2_X1 U14686 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12790) );
  AND4_X1 U14687 ( .A1(n12793), .A2(n12792), .A3(n12791), .A4(n12790), .ZN(
        n12804) );
  NAND2_X1 U14688 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12797) );
  AOI22_X1 U14689 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12796) );
  AOI22_X1 U14690 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12795) );
  NAND2_X1 U14691 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12794) );
  NAND4_X1 U14692 ( .A1(n12797), .A2(n12796), .A3(n12795), .A4(n12794), .ZN(
        n12802) );
  NAND2_X1 U14693 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12799) );
  NAND2_X1 U14694 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12798) );
  OAI211_X1 U14695 ( .C1(n12800), .C2(n13026), .A(n12799), .B(n12798), .ZN(
        n12801) );
  NOR2_X1 U14696 ( .A1(n12802), .A2(n12801), .ZN(n12803) );
  INV_X1 U14697 ( .A(n12974), .ZN(n15116) );
  NAND2_X1 U14698 ( .A1(n12846), .A2(n15116), .ZN(n12806) );
  AOI22_X1 U14699 ( .A1(n12875), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U14700 ( .A1(n13114), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13022), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U14701 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12810) );
  AOI22_X1 U14702 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n13113), .B1(
        n13115), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12809) );
  NAND2_X1 U14703 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12808) );
  AND4_X1 U14704 ( .A1(n12811), .A2(n12810), .A3(n12809), .A4(n12808), .ZN(
        n12823) );
  NAND2_X1 U14705 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12815) );
  AOI22_X1 U14706 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12077), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U14707 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13103), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12813) );
  NAND2_X1 U14708 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12812) );
  NAND4_X1 U14709 ( .A1(n12815), .A2(n12814), .A3(n12813), .A4(n12812), .ZN(
        n12821) );
  INV_X1 U14710 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12818) );
  NAND2_X1 U14711 ( .A1(n13108), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12817) );
  NAND2_X1 U14712 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12816) );
  OAI211_X1 U14713 ( .C1(n12819), .C2(n12818), .A(n12817), .B(n12816), .ZN(
        n12820) );
  NOR2_X1 U14714 ( .A1(n12821), .A2(n12820), .ZN(n12822) );
  NAND2_X1 U14715 ( .A1(n12870), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12825) );
  AOI22_X1 U14716 ( .A1(n12875), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12824) );
  OAI211_X1 U14717 ( .C1(n15189), .C2(n12826), .A(n12825), .B(n12824), .ZN(
        n16916) );
  NAND2_X1 U14718 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12830) );
  AOI22_X1 U14719 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12077), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12829) );
  AOI22_X1 U14720 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n13103), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12828) );
  NAND2_X1 U14721 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12827) );
  NAND4_X1 U14722 ( .A1(n12830), .A2(n12829), .A3(n12828), .A4(n12827), .ZN(
        n12835) );
  NAND2_X1 U14723 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12832) );
  NAND2_X1 U14724 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12831) );
  OAI211_X1 U14725 ( .C1(n12833), .C2(n13026), .A(n12832), .B(n12831), .ZN(
        n12834) );
  NOR2_X1 U14726 ( .A1(n12835), .A2(n12834), .ZN(n12842) );
  INV_X1 U14727 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12836) );
  OAI22_X1 U14728 ( .A1(n12046), .A2(n15783), .B1(n13030), .B2(n12836), .ZN(
        n12838) );
  INV_X1 U14729 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15237) );
  OAI22_X1 U14730 ( .A1(n13033), .A2(n15786), .B1(n13032), .B2(n15237), .ZN(
        n12837) );
  NOR2_X1 U14731 ( .A1(n12838), .A2(n12837), .ZN(n12841) );
  AOI22_X1 U14732 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12840) );
  NAND2_X1 U14733 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12839) );
  NAND4_X1 U14734 ( .A1(n12842), .A2(n12841), .A3(n12840), .A4(n12839), .ZN(
        n15148) );
  AOI22_X1 U14735 ( .A1(n12875), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12843) );
  OAI21_X1 U14736 ( .B1(n12878), .B2(n12844), .A(n12843), .ZN(n12845) );
  AOI21_X1 U14737 ( .B1(n12846), .B2(n15148), .A(n12845), .ZN(n15465) );
  AOI22_X1 U14738 ( .A1(n12875), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12847) );
  OAI21_X1 U14739 ( .B1(n12878), .B2(n17486), .A(n12847), .ZN(n15239) );
  NAND2_X1 U14740 ( .A1(n12870), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12849) );
  AOI22_X1 U14741 ( .A1(n12875), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12848) );
  NAND2_X1 U14742 ( .A1(n12870), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U14743 ( .A1(n12875), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12850) );
  NAND2_X1 U14744 ( .A1(n12870), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U14745 ( .A1(n12875), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U14746 ( .A1(n12875), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12854) );
  OAI21_X1 U14747 ( .B1(n12878), .B2(n13296), .A(n12854), .ZN(n13336) );
  NAND2_X1 U14748 ( .A1(n13335), .A2(n13336), .ZN(n13334) );
  NAND2_X1 U14749 ( .A1(n12870), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12856) );
  AOI22_X1 U14750 ( .A1(n12875), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12855) );
  NAND2_X1 U14751 ( .A1(n12870), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12858) );
  AOI22_X1 U14752 ( .A1(n12875), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12857) );
  INV_X1 U14753 ( .A(n16562), .ZN(n12859) );
  AOI22_X1 U14754 ( .A1(n12875), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12860) );
  OAI21_X1 U14755 ( .B1(n12878), .B2(n17490), .A(n12860), .ZN(n16436) );
  AOI22_X1 U14756 ( .A1(n12875), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12861) );
  OAI21_X1 U14757 ( .B1(n12878), .B2(n16603), .A(n12861), .ZN(n16545) );
  INV_X1 U14758 ( .A(n16548), .ZN(n12865) );
  NAND2_X1 U14759 ( .A1(n12870), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12863) );
  AOI22_X1 U14760 ( .A1(n12875), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12862) );
  AND2_X1 U14761 ( .A1(n12863), .A2(n12862), .ZN(n16536) );
  INV_X1 U14762 ( .A(n16536), .ZN(n12864) );
  NAND2_X1 U14763 ( .A1(n12865), .A2(n12864), .ZN(n16538) );
  NAND2_X1 U14764 ( .A1(n12870), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12867) );
  AOI22_X1 U14765 ( .A1(n12875), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12866) );
  AND2_X1 U14766 ( .A1(n12867), .A2(n12866), .ZN(n16421) );
  AOI22_X1 U14767 ( .A1(n12875), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12868) );
  OAI21_X1 U14768 ( .B1(n12878), .B2(n17493), .A(n12868), .ZN(n13362) );
  AOI22_X1 U14769 ( .A1(n12875), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12869) );
  OAI21_X1 U14770 ( .B1(n12878), .B2(n17494), .A(n12869), .ZN(n13260) );
  INV_X1 U14771 ( .A(n15703), .ZN(n12874) );
  NAND2_X1 U14772 ( .A1(n12870), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12872) );
  AOI22_X1 U14773 ( .A1(n12875), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12871) );
  AND2_X1 U14774 ( .A1(n12872), .A2(n12871), .ZN(n15702) );
  INV_X1 U14775 ( .A(n15702), .ZN(n12873) );
  INV_X1 U14776 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n12877) );
  AOI22_X1 U14777 ( .A1(n12875), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12647), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12876) );
  OAI21_X1 U14778 ( .B1(n12878), .B2(n12877), .A(n12876), .ZN(n12879) );
  INV_X1 U14779 ( .A(n12879), .ZN(n12880) );
  AND2_X1 U14780 ( .A1(n12883), .A2(n12882), .ZN(n14810) );
  INV_X1 U14781 ( .A(n14810), .ZN(n15013) );
  NAND2_X1 U14782 ( .A1(n12599), .A2(n12884), .ZN(n15006) );
  NAND2_X1 U14783 ( .A1(n15006), .A2(n12651), .ZN(n12885) );
  NAND2_X1 U14784 ( .A1(n15013), .A2(n12885), .ZN(n12886) );
  NAND2_X1 U14785 ( .A1(n12890), .A2(n12889), .ZN(n13254) );
  INV_X1 U14786 ( .A(n12891), .ZN(n12893) );
  NAND3_X1 U14787 ( .A1(n12893), .A2(n12895), .A3(n12892), .ZN(n12898) );
  NAND2_X1 U14788 ( .A1(n19703), .A2(n17083), .ZN(n12897) );
  INV_X1 U14789 ( .A(n13256), .ZN(n14572) );
  OAI21_X1 U14790 ( .B1(n12895), .B2(n12894), .A(n14572), .ZN(n12896) );
  AND4_X1 U14791 ( .A1(n13254), .A2(n12898), .A3(n12897), .A4(n12896), .ZN(
        n12904) );
  NAND2_X1 U14792 ( .A1(n12899), .A2(n12651), .ZN(n14971) );
  NAND2_X1 U14793 ( .A1(n14971), .A2(n12900), .ZN(n12902) );
  NAND2_X1 U14794 ( .A1(n12902), .A2(n12901), .ZN(n12903) );
  AND3_X1 U14795 ( .A1(n12905), .A2(n12904), .A3(n12903), .ZN(n14970) );
  INV_X1 U14796 ( .A(n12906), .ZN(n14811) );
  NAND2_X1 U14797 ( .A1(n14970), .A2(n14811), .ZN(n12907) );
  NAND2_X1 U14798 ( .A1(n17005), .A2(n17002), .ZN(n18671) );
  INV_X1 U14799 ( .A(n18671), .ZN(n12921) );
  NAND2_X1 U14800 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12920) );
  NAND2_X1 U14801 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17052) );
  NAND2_X1 U14802 ( .A1(n15670), .A2(n17052), .ZN(n15660) );
  NAND2_X1 U14803 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18675) );
  NOR2_X1 U14804 ( .A1(n15212), .A2(n18675), .ZN(n12908) );
  AND2_X1 U14805 ( .A1(n15660), .A2(n12908), .ZN(n17003) );
  NOR2_X1 U14806 ( .A1(n17000), .A2(n16999), .ZN(n16998) );
  NAND3_X1 U14807 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17003), .A3(
        n16998), .ZN(n12912) );
  NOR2_X1 U14808 ( .A1(n17005), .A2(n12912), .ZN(n12910) );
  OR2_X1 U14809 ( .A1(n15670), .A2(n17052), .ZN(n15659) );
  NAND2_X1 U14810 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12908), .ZN(
        n16995) );
  NOR2_X1 U14811 ( .A1(n15659), .A2(n16995), .ZN(n17001) );
  NAND2_X1 U14812 ( .A1(n16998), .A2(n17001), .ZN(n12915) );
  NOR2_X1 U14813 ( .A1(n17002), .A2(n12915), .ZN(n12909) );
  AND2_X1 U14814 ( .A1(n16833), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12911) );
  NAND2_X1 U14815 ( .A1(n16990), .A2(n12911), .ZN(n16837) );
  NOR2_X1 U14816 ( .A1(n16837), .A2(n16834), .ZN(n12922) );
  AND2_X1 U14817 ( .A1(n12922), .A2(n16597), .ZN(n16820) );
  INV_X1 U14818 ( .A(n12912), .ZN(n12913) );
  NOR2_X1 U14819 ( .A1(n17005), .A2(n12913), .ZN(n12914) );
  NOR2_X1 U14820 ( .A1(n12933), .A2(n18500), .ZN(n18665) );
  OR2_X1 U14821 ( .A1(n12914), .A2(n18665), .ZN(n15691) );
  INV_X1 U14822 ( .A(n12915), .ZN(n16856) );
  NOR2_X1 U14823 ( .A1(n17002), .A2(n16856), .ZN(n12916) );
  NOR2_X1 U14824 ( .A1(n15691), .A2(n12916), .ZN(n16987) );
  INV_X1 U14825 ( .A(n16833), .ZN(n12917) );
  NAND2_X1 U14826 ( .A1(n18671), .A2(n12917), .ZN(n12918) );
  AND2_X1 U14827 ( .A1(n16987), .A2(n12918), .ZN(n16848) );
  OAI21_X1 U14828 ( .B1(n16847), .B2(n16834), .A(n18671), .ZN(n12919) );
  NAND2_X1 U14829 ( .A1(n16848), .A2(n12919), .ZN(n16823) );
  OR2_X1 U14830 ( .A1(n16820), .A2(n16823), .ZN(n16816) );
  AOI21_X1 U14831 ( .B1(n12920), .B2(n18671), .A(n16816), .ZN(n16787) );
  OAI21_X1 U14832 ( .B1(n12921), .B2(n12923), .A(n16787), .ZN(n15709) );
  AND2_X1 U14833 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n12922), .ZN(
        n16811) );
  NAND3_X1 U14834 ( .A1(n12923), .A2(n13323), .A3(n15280), .ZN(n12924) );
  NAND2_X1 U14835 ( .A1(n18532), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n15760) );
  NAND2_X1 U14836 ( .A1(n12924), .A2(n15760), .ZN(n12925) );
  AOI21_X1 U14837 ( .B1(n15709), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12925), .ZN(n12926) );
  OAI21_X1 U14838 ( .B1(n16472), .B2(n18666), .A(n12929), .ZN(n12930) );
  INV_X1 U14839 ( .A(n12930), .ZN(n12935) );
  INV_X1 U14840 ( .A(n15030), .ZN(n15002) );
  NOR2_X1 U14841 ( .A1(n12251), .A2(n15002), .ZN(n12932) );
  OAI211_X1 U14842 ( .C1(n15767), .C2(n18664), .A(n12935), .B(n12934), .ZN(
        P2_U3015) );
  NAND2_X1 U14843 ( .A1(n14819), .A2(n12956), .ZN(n12940) );
  NAND2_X1 U14844 ( .A1(n19376), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12936) );
  NAND2_X1 U14845 ( .A1(n19327), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12946) );
  AOI21_X1 U14846 ( .B1(n12946), .B2(n17436), .A(n19355), .ZN(n12938) );
  INV_X1 U14847 ( .A(n12946), .ZN(n12937) );
  NAND2_X1 U14848 ( .A1(n12937), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n17079) );
  AOI22_X1 U14849 ( .A1(n12953), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n12938), .B2(n17079), .ZN(n12939) );
  NAND2_X1 U14850 ( .A1(n12940), .A2(n12939), .ZN(n12943) );
  INV_X1 U14851 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13172) );
  NAND2_X1 U14852 ( .A1(n12943), .A2(n12942), .ZN(n12965) );
  NAND2_X1 U14853 ( .A1(n12944), .A2(n12956), .ZN(n12949) );
  INV_X1 U14854 ( .A(n19327), .ZN(n19302) );
  NAND2_X1 U14855 ( .A1(n19302), .A2(n19257), .ZN(n12945) );
  NAND2_X1 U14856 ( .A1(n12946), .A2(n12945), .ZN(n17100) );
  NOR2_X1 U14857 ( .A1(n17100), .A2(n19355), .ZN(n12947) );
  AOI21_X1 U14858 ( .B1(n12953), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12947), .ZN(n12948) );
  NOR2_X1 U14859 ( .A1(n19355), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12951) );
  NAND2_X1 U14860 ( .A1(n12953), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12954) );
  NOR2_X1 U14861 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17101) );
  INV_X1 U14862 ( .A(n17101), .ZN(n19301) );
  NAND3_X1 U14863 ( .A1(n19346), .A2(n19302), .A3(n19301), .ZN(n19339) );
  NAND2_X1 U14864 ( .A1(n12954), .A2(n19339), .ZN(n12955) );
  INV_X1 U14865 ( .A(n14842), .ZN(n12958) );
  NAND2_X1 U14866 ( .A1(n12958), .A2(n12957), .ZN(n12959) );
  INV_X1 U14867 ( .A(n12960), .ZN(n12961) );
  NAND2_X1 U14868 ( .A1(n12962), .A2(n12961), .ZN(n12963) );
  NAND2_X1 U14869 ( .A1(n19376), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12964) );
  AND2_X1 U14870 ( .A1(n12965), .A2(n12964), .ZN(n12966) );
  INV_X1 U14871 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17095) );
  NAND2_X1 U14872 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14895) );
  NOR2_X1 U14873 ( .A1(n17095), .A2(n14895), .ZN(n12971) );
  INV_X1 U14874 ( .A(n15112), .ZN(n12969) );
  NOR2_X1 U14875 ( .A1(n12967), .A2(n15054), .ZN(n12968) );
  AND2_X1 U14876 ( .A1(n12968), .A2(n15086), .ZN(n15055) );
  AND2_X1 U14877 ( .A1(n12969), .A2(n15055), .ZN(n12970) );
  AND2_X1 U14878 ( .A1(n12971), .A2(n12970), .ZN(n15076) );
  AND2_X1 U14879 ( .A1(n15079), .A2(n15076), .ZN(n12972) );
  INV_X1 U14880 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19530) );
  NOR2_X1 U14881 ( .A1(n13149), .A2(n19530), .ZN(n15075) );
  AND2_X1 U14882 ( .A1(n12972), .A2(n15075), .ZN(n12973) );
  NAND2_X1 U14883 ( .A1(n14822), .A2(n12973), .ZN(n15078) );
  OR2_X1 U14884 ( .A1(n15078), .A2(n12974), .ZN(n15188) );
  INV_X1 U14885 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12981) );
  NAND2_X1 U14886 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12978) );
  AOI22_X1 U14887 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12977) );
  AOI22_X1 U14888 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12976) );
  NAND2_X1 U14889 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12975) );
  AND4_X1 U14890 ( .A1(n12978), .A2(n12977), .A3(n12976), .A4(n12975), .ZN(
        n12980) );
  AOI22_X1 U14891 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13108), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12979) );
  OAI211_X1 U14892 ( .C1(n13112), .C2(n12981), .A(n12980), .B(n12979), .ZN(
        n12987) );
  AOI22_X1 U14893 ( .A1(n13114), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U14894 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13115), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U14895 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12983) );
  NAND2_X1 U14896 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12982) );
  NAND4_X1 U14897 ( .A1(n12985), .A2(n12984), .A3(n12983), .A4(n12982), .ZN(
        n12986) );
  INV_X1 U14898 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12994) );
  NAND2_X1 U14899 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12991) );
  AOI22_X1 U14900 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12077), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12990) );
  AOI22_X1 U14901 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13103), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12989) );
  NAND2_X1 U14902 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12988) );
  AND4_X1 U14903 ( .A1(n12991), .A2(n12990), .A3(n12989), .A4(n12988), .ZN(
        n12993) );
  AOI22_X1 U14904 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13108), .B1(
        n11991), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12992) );
  OAI211_X1 U14905 ( .C1(n12994), .C2(n13112), .A(n12993), .B(n12992), .ZN(
        n13000) );
  AOI22_X1 U14906 ( .A1(n13114), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U14907 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n13115), .ZN(n12997) );
  AOI22_X1 U14908 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12996) );
  NAND2_X1 U14909 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12995) );
  NAND4_X1 U14910 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n12995), .ZN(
        n12999) );
  NOR2_X1 U14911 ( .A1(n13000), .A2(n12999), .ZN(n15195) );
  NAND2_X1 U14912 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13004) );
  AOI22_X1 U14913 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U14914 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13002) );
  NAND2_X1 U14915 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13001) );
  NAND4_X1 U14916 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        n13009) );
  NAND2_X1 U14917 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13006) );
  NAND2_X1 U14918 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n13005) );
  OAI211_X1 U14919 ( .C1(n13026), .C2(n13007), .A(n13006), .B(n13005), .ZN(
        n13008) );
  NOR2_X1 U14920 ( .A1(n13009), .A2(n13008), .ZN(n13017) );
  INV_X1 U14921 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17090) );
  INV_X1 U14922 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13010) );
  OAI22_X1 U14923 ( .A1(n12046), .A2(n17090), .B1(n13030), .B2(n13010), .ZN(
        n13013) );
  INV_X1 U14924 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13159) );
  OAI22_X1 U14925 ( .A1(n13033), .A2(n13159), .B1(n13032), .B2(n13011), .ZN(
        n13012) );
  NOR2_X1 U14926 ( .A1(n13013), .A2(n13012), .ZN(n13016) );
  AOI22_X1 U14927 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13015) );
  NAND2_X1 U14928 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13014) );
  NAND4_X1 U14929 ( .A1(n13017), .A2(n13016), .A3(n13015), .A4(n13014), .ZN(
        n15369) );
  NAND2_X1 U14930 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13021) );
  AOI22_X1 U14931 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13020) );
  AOI22_X1 U14932 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13019) );
  NAND2_X1 U14933 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13018) );
  NAND4_X1 U14934 ( .A1(n13021), .A2(n13020), .A3(n13019), .A4(n13018), .ZN(
        n13028) );
  NAND2_X1 U14935 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13024) );
  NAND2_X1 U14936 ( .A1(n13022), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n13023) );
  OAI211_X1 U14937 ( .C1(n13026), .C2(n13025), .A(n13024), .B(n13023), .ZN(
        n13027) );
  NOR2_X1 U14938 ( .A1(n13028), .A2(n13027), .ZN(n13039) );
  INV_X1 U14939 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13029) );
  OAI22_X1 U14940 ( .A1(n12046), .A2(n13172), .B1(n13030), .B2(n13029), .ZN(
        n13035) );
  INV_X1 U14941 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13179) );
  OAI22_X1 U14942 ( .A1(n13033), .A2(n13179), .B1(n13032), .B2(n13031), .ZN(
        n13034) );
  NOR2_X1 U14943 ( .A1(n13035), .A2(n13034), .ZN(n13038) );
  AOI22_X1 U14944 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13037) );
  NAND2_X1 U14945 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13036) );
  NAND4_X1 U14946 ( .A1(n13039), .A2(n13038), .A3(n13037), .A4(n13036), .ZN(
        n15450) );
  INV_X1 U14947 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13046) );
  NAND2_X1 U14948 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13043) );
  AOI22_X1 U14949 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12077), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U14950 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n13103), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13041) );
  NAND2_X1 U14951 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13040) );
  AND4_X1 U14952 ( .A1(n13043), .A2(n13042), .A3(n13041), .A4(n13040), .ZN(
        n13045) );
  AOI22_X1 U14953 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13108), .B1(
        n11991), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13044) );
  OAI211_X1 U14954 ( .C1(n13046), .C2(n13112), .A(n13045), .B(n13044), .ZN(
        n13052) );
  AOI22_X1 U14955 ( .A1(n13114), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U14956 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__4__SCAN_IN), .B2(n13115), .ZN(n13049) );
  AOI22_X1 U14957 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13048) );
  NAND2_X1 U14958 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13047) );
  NAND4_X1 U14959 ( .A1(n13050), .A2(n13049), .A3(n13048), .A4(n13047), .ZN(
        n13051) );
  INV_X1 U14960 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13060) );
  NAND2_X1 U14961 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13057) );
  AOI22_X1 U14962 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U14963 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13055) );
  NAND2_X1 U14964 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13054) );
  AND4_X1 U14965 ( .A1(n13057), .A2(n13056), .A3(n13055), .A4(n13054), .ZN(
        n13059) );
  AOI22_X1 U14966 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13108), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13058) );
  OAI211_X1 U14967 ( .C1(n13112), .C2(n13060), .A(n13059), .B(n13058), .ZN(
        n13066) );
  AOI22_X1 U14968 ( .A1(n13114), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U14969 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13115), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U14970 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13062) );
  NAND2_X1 U14971 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13061) );
  NAND4_X1 U14972 ( .A1(n13064), .A2(n13063), .A3(n13062), .A4(n13061), .ZN(
        n13065) );
  NOR2_X1 U14973 ( .A1(n13066), .A2(n13065), .ZN(n15518) );
  INV_X1 U14974 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13073) );
  NAND2_X1 U14975 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13070) );
  AOI22_X1 U14976 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12077), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13069) );
  AOI22_X1 U14977 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n13103), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13068) );
  NAND2_X1 U14978 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n13067) );
  AND4_X1 U14979 ( .A1(n13070), .A2(n13069), .A3(n13068), .A4(n13067), .ZN(
        n13072) );
  AOI22_X1 U14980 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n13108), .B1(
        n11991), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13071) );
  OAI211_X1 U14981 ( .C1(n13073), .C2(n13112), .A(n13072), .B(n13071), .ZN(
        n13079) );
  AOI22_X1 U14982 ( .A1(n13114), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U14983 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__6__SCAN_IN), .B2(n13115), .ZN(n13076) );
  AOI22_X1 U14984 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13075) );
  NAND2_X1 U14985 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n13074) );
  NAND4_X1 U14986 ( .A1(n13077), .A2(n13076), .A3(n13075), .A4(n13074), .ZN(
        n13078) );
  NOR2_X1 U14987 ( .A1(n13079), .A2(n13078), .ZN(n16517) );
  INV_X1 U14988 ( .A(n16517), .ZN(n13080) );
  AOI22_X1 U14989 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10967), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U14990 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U14991 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13089) );
  NAND2_X1 U14992 ( .A1(n11977), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13086) );
  INV_X1 U14993 ( .A(n13083), .ZN(n13085) );
  NAND2_X1 U14994 ( .A1(n10990), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13084) );
  NAND2_X1 U14995 ( .A1(n13085), .A2(n13084), .ZN(n15784) );
  OAI211_X1 U14996 ( .C1(n13082), .C2(n11981), .A(n13086), .B(n15784), .ZN(
        n13087) );
  INV_X1 U14997 ( .A(n13087), .ZN(n13088) );
  NAND4_X1 U14998 ( .A1(n13091), .A2(n13090), .A3(n13089), .A4(n13088), .ZN(
        n13100) );
  AOI22_X1 U14999 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U15000 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13097) );
  AOI22_X1 U15001 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13096) );
  NAND2_X1 U15002 ( .A1(n11977), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13092) );
  INV_X1 U15003 ( .A(n15784), .ZN(n13219) );
  OAI211_X1 U15004 ( .C1(n13082), .C2(n13093), .A(n13092), .B(n13219), .ZN(
        n13094) );
  INV_X1 U15005 ( .A(n13094), .ZN(n13095) );
  NAND4_X1 U15006 ( .A1(n13098), .A2(n13097), .A3(n13096), .A4(n13095), .ZN(
        n13099) );
  NAND2_X1 U15007 ( .A1(n13100), .A2(n13099), .ZN(n13126) );
  INV_X1 U15008 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13111) );
  NAND2_X1 U15009 ( .A1(n13101), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13107) );
  AOI22_X1 U15010 ( .A1(n12077), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13102), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U15011 ( .A1(n13103), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11996), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13105) );
  NAND2_X1 U15012 ( .A1(n12012), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n13104) );
  AND4_X1 U15013 ( .A1(n13107), .A2(n13106), .A3(n13105), .A4(n13104), .ZN(
        n13110) );
  AOI22_X1 U15014 ( .A1(n11991), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13108), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13109) );
  OAI211_X1 U15015 ( .C1(n13112), .C2(n13111), .A(n13110), .B(n13109), .ZN(
        n13124) );
  AOI22_X1 U15016 ( .A1(n13114), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13113), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U15017 ( .A1(n13116), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13115), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U15018 ( .A1(n12763), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13117), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13120) );
  NAND2_X1 U15019 ( .A1(n13118), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13119) );
  NAND4_X1 U15020 ( .A1(n13122), .A2(n13121), .A3(n13120), .A4(n13119), .ZN(
        n13123) );
  NOR2_X1 U15021 ( .A1(n13124), .A2(n13123), .ZN(n13125) );
  XOR2_X1 U15022 ( .A(n13126), .B(n13125), .Z(n16508) );
  INV_X1 U15023 ( .A(n13125), .ZN(n13128) );
  INV_X1 U15024 ( .A(n13126), .ZN(n13127) );
  AOI22_X1 U15025 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11842), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U15026 ( .A1(n15792), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10964), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13134) );
  AOI22_X1 U15027 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13133) );
  INV_X1 U15028 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13130) );
  NAND2_X1 U15029 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13129) );
  OAI211_X1 U15030 ( .C1(n10968), .C2(n13130), .A(n13129), .B(n15784), .ZN(
        n13131) );
  INV_X1 U15031 ( .A(n13131), .ZN(n13132) );
  NAND4_X1 U15032 ( .A1(n13135), .A2(n13134), .A3(n13133), .A4(n13132), .ZN(
        n13144) );
  AOI22_X1 U15033 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11842), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13142) );
  AOI22_X1 U15034 ( .A1(n15792), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13141) );
  AOI22_X1 U15035 ( .A1(n15776), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13140) );
  NAND2_X1 U15036 ( .A1(n11975), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13136) );
  OAI211_X1 U15037 ( .C1(n10968), .C2(n13137), .A(n13136), .B(n13219), .ZN(
        n13138) );
  INV_X1 U15038 ( .A(n13138), .ZN(n13139) );
  NAND4_X1 U15039 ( .A1(n13142), .A2(n13141), .A3(n13140), .A4(n13139), .ZN(
        n13143) );
  NAND2_X1 U15040 ( .A1(n13144), .A2(n13143), .ZN(n13147) );
  INV_X1 U15041 ( .A(n13147), .ZN(n13145) );
  NAND2_X1 U15042 ( .A1(n13146), .A2(n13145), .ZN(n13151) );
  INV_X1 U15043 ( .A(n13146), .ZN(n13148) );
  OAI21_X1 U15044 ( .B1(n13149), .B2(n13148), .A(n13147), .ZN(n13150) );
  OAI21_X1 U15045 ( .B1(n19642), .B2(n13151), .A(n13150), .ZN(n16504) );
  INV_X1 U15046 ( .A(n13151), .ZN(n13167) );
  AOI22_X1 U15047 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10967), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U15048 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13156) );
  AOI22_X1 U15049 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13155) );
  NAND2_X1 U15050 ( .A1(n11977), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13152) );
  OAI211_X1 U15051 ( .C1(n13082), .C2(n17090), .A(n13152), .B(n15784), .ZN(
        n13153) );
  INV_X1 U15052 ( .A(n13153), .ZN(n13154) );
  NAND4_X1 U15053 ( .A1(n13157), .A2(n13156), .A3(n13155), .A4(n13154), .ZN(
        n13166) );
  AOI22_X1 U15054 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10966), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13164) );
  AOI22_X1 U15055 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13163) );
  AOI22_X1 U15056 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13162) );
  NAND2_X1 U15057 ( .A1(n11977), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13158) );
  OAI211_X1 U15058 ( .C1(n13082), .C2(n13159), .A(n13158), .B(n13219), .ZN(
        n13160) );
  INV_X1 U15059 ( .A(n13160), .ZN(n13161) );
  NAND4_X1 U15060 ( .A1(n13164), .A2(n13163), .A3(n13162), .A4(n13161), .ZN(
        n13165) );
  AND2_X1 U15061 ( .A1(n13166), .A2(n13165), .ZN(n13168) );
  NAND2_X1 U15062 ( .A1(n13167), .A2(n13168), .ZN(n13192) );
  OAI211_X1 U15063 ( .C1(n13167), .C2(n13168), .A(n13208), .B(n13192), .ZN(
        n13170) );
  INV_X1 U15064 ( .A(n13168), .ZN(n13169) );
  NOR2_X1 U15065 ( .A1(n12651), .A2(n13169), .ZN(n16497) );
  NAND2_X1 U15066 ( .A1(n16495), .A2(n16497), .ZN(n16496) );
  AOI22_X1 U15067 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10966), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13177) );
  AOI22_X1 U15068 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13176) );
  AOI22_X1 U15069 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13175) );
  NAND2_X1 U15070 ( .A1(n11977), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13171) );
  OAI211_X1 U15071 ( .C1(n13082), .C2(n13172), .A(n13171), .B(n15784), .ZN(
        n13173) );
  INV_X1 U15072 ( .A(n13173), .ZN(n13174) );
  NAND4_X1 U15073 ( .A1(n13177), .A2(n13176), .A3(n13175), .A4(n13174), .ZN(
        n13186) );
  AOI22_X1 U15074 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13184) );
  AOI22_X1 U15075 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13183) );
  AOI22_X1 U15076 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13182) );
  NAND2_X1 U15077 ( .A1(n11977), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13178) );
  OAI211_X1 U15078 ( .C1(n13082), .C2(n13179), .A(n13178), .B(n13219), .ZN(
        n13180) );
  INV_X1 U15079 ( .A(n13180), .ZN(n13181) );
  NAND4_X1 U15080 ( .A1(n13184), .A2(n13183), .A3(n13182), .A4(n13181), .ZN(
        n13185) );
  AND2_X1 U15081 ( .A1(n13186), .A2(n13185), .ZN(n13190) );
  XNOR2_X1 U15082 ( .A(n13192), .B(n13190), .ZN(n13187) );
  NAND2_X1 U15083 ( .A1(n19642), .A2(n13190), .ZN(n16488) );
  INV_X1 U15084 ( .A(n13190), .ZN(n13191) );
  NOR2_X1 U15085 ( .A1(n13192), .A2(n13191), .ZN(n13209) );
  AOI22_X1 U15086 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11008), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13198) );
  AOI22_X1 U15087 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13197) );
  AOI22_X1 U15088 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13196) );
  NAND2_X1 U15089 ( .A1(n11977), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13193) );
  OAI211_X1 U15090 ( .C1(n13082), .C2(n19530), .A(n13193), .B(n15784), .ZN(
        n13194) );
  INV_X1 U15091 ( .A(n13194), .ZN(n13195) );
  NAND4_X1 U15092 ( .A1(n13198), .A2(n13197), .A3(n13196), .A4(n13195), .ZN(
        n13207) );
  AOI22_X1 U15093 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15776), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U15094 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10964), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13204) );
  AOI22_X1 U15095 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13203) );
  NAND2_X1 U15096 ( .A1(n11977), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13199) );
  OAI211_X1 U15097 ( .C1(n13082), .C2(n13200), .A(n13199), .B(n13219), .ZN(
        n13201) );
  INV_X1 U15098 ( .A(n13201), .ZN(n13202) );
  NAND4_X1 U15099 ( .A1(n13205), .A2(n13204), .A3(n13203), .A4(n13202), .ZN(
        n13206) );
  AND2_X1 U15100 ( .A1(n13207), .A2(n13206), .ZN(n13210) );
  NAND2_X1 U15101 ( .A1(n13209), .A2(n13210), .ZN(n16475) );
  OAI211_X1 U15102 ( .C1(n13209), .C2(n13210), .A(n13208), .B(n16475), .ZN(
        n13230) );
  INV_X1 U15103 ( .A(n13210), .ZN(n13211) );
  OAI21_X1 U15104 ( .B1(n13082), .B2(n19479), .A(n15784), .ZN(n13215) );
  INV_X1 U15105 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13212) );
  OAI22_X1 U15106 ( .A1(n11793), .A2(n13213), .B1(n13081), .B2(n13212), .ZN(
        n13214) );
  AOI211_X1 U15107 ( .C1(n11977), .C2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n13215), .B(n13214), .ZN(n13218) );
  AOI22_X1 U15108 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10964), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13217) );
  AOI22_X1 U15109 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10967), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13216) );
  NAND3_X1 U15110 ( .A1(n13218), .A2(n13217), .A3(n13216), .ZN(n13229) );
  INV_X1 U15111 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13220) );
  OAI21_X1 U15112 ( .B1(n13082), .B2(n13220), .A(n13219), .ZN(n13224) );
  INV_X1 U15113 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13222) );
  INV_X1 U15114 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13221) );
  OAI22_X1 U15115 ( .A1(n11793), .A2(n13222), .B1(n13081), .B2(n13221), .ZN(
        n13223) );
  AOI211_X1 U15116 ( .C1(n11977), .C2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n13224), .B(n13223), .ZN(n13227) );
  AOI22_X1 U15117 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13226) );
  AOI22_X1 U15118 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10966), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13225) );
  NAND3_X1 U15119 ( .A1(n13227), .A2(n13226), .A3(n13225), .ZN(n13228) );
  AND2_X1 U15120 ( .A1(n13229), .A2(n13228), .ZN(n13251) );
  NAND2_X1 U15121 ( .A1(n13231), .A2(n13230), .ZN(n16481) );
  AOI22_X1 U15122 ( .A1(n11008), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n15792), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13233) );
  AOI22_X1 U15123 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13232) );
  NAND2_X1 U15124 ( .A1(n13233), .A2(n13232), .ZN(n13247) );
  AOI22_X1 U15125 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13235) );
  AOI21_X1 U15126 ( .B1(n15777), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n15784), .ZN(n13234) );
  OAI211_X1 U15127 ( .C1(n15787), .C2(n13236), .A(n13235), .B(n13234), .ZN(
        n13246) );
  INV_X1 U15128 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19418) );
  OAI21_X1 U15129 ( .B1(n13082), .B2(n19418), .A(n15784), .ZN(n13241) );
  INV_X1 U15130 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13237) );
  OAI22_X1 U15131 ( .A1(n11793), .A2(n13239), .B1(n11011), .B2(n13237), .ZN(
        n13240) );
  AOI211_X1 U15132 ( .C1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .C2(n11977), .A(
        n13241), .B(n13240), .ZN(n13244) );
  AOI22_X1 U15133 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15791), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U15134 ( .A1(n10966), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13242) );
  NAND3_X1 U15135 ( .A1(n13244), .A2(n13243), .A3(n13242), .ZN(n13245) );
  OAI21_X1 U15136 ( .B1(n13247), .B2(n13246), .A(n13245), .ZN(n13248) );
  NAND2_X1 U15137 ( .A1(n13249), .A2(n13248), .ZN(n15772) );
  INV_X1 U15138 ( .A(n15772), .ZN(n13250) );
  NOR2_X1 U15139 ( .A1(n13249), .A2(n13248), .ZN(n15773) );
  NOR2_X1 U15140 ( .A1(n13250), .A2(n15773), .ZN(n13252) );
  INV_X1 U15141 ( .A(n13251), .ZN(n16477) );
  NOR3_X1 U15142 ( .A1(n16475), .A2(n19642), .A3(n16477), .ZN(n15771) );
  XNOR2_X1 U15143 ( .A(n13252), .B(n15771), .ZN(n15770) );
  INV_X1 U15144 ( .A(n15128), .ZN(n13253) );
  NAND2_X1 U15145 ( .A1(n13253), .A2(n15010), .ZN(n14954) );
  NAND2_X1 U15146 ( .A1(n14954), .A2(n13254), .ZN(n13255) );
  NAND2_X1 U15147 ( .A1(n18371), .A2(n15015), .ZN(n13257) );
  OAI21_X1 U15148 ( .B1(n13360), .B2(n13260), .A(n15703), .ZN(n13317) );
  INV_X1 U15149 ( .A(n13317), .ZN(n18614) );
  NOR4_X1 U15150 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13264) );
  NOR4_X1 U15151 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n13263) );
  NOR4_X1 U15152 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13262) );
  NOR4_X1 U15153 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n13261) );
  NAND4_X1 U15154 ( .A1(n13264), .A2(n13263), .A3(n13262), .A4(n13261), .ZN(
        n13269) );
  NOR4_X1 U15155 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n13267) );
  NOR4_X1 U15156 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13266) );
  NOR4_X1 U15157 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13265) );
  NAND4_X1 U15158 ( .A1(n13267), .A2(n13266), .A3(n13265), .A4(n19821), .ZN(
        n13268) );
  INV_X1 U15159 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20075) );
  NOR2_X1 U15160 ( .A1(n15131), .A2(n20075), .ZN(n13270) );
  AOI21_X1 U15161 ( .B1(n15131), .B2(BUF2_REG_13__SCAN_IN), .A(n13270), .ZN(
        n19199) );
  INV_X1 U15162 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14859) );
  OAI22_X1 U15163 ( .A1(n19189), .A2(n19199), .B1(n19686), .B2(n14859), .ZN(
        n13271) );
  AOI21_X1 U15164 ( .B1(n18614), .B2(n19633), .A(n13271), .ZN(n13274) );
  AOI22_X1 U15165 ( .A1(n19185), .A2(BUF2_REG_29__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n13273) );
  OAI21_X1 U15166 ( .B1(n15770), .B2(n19636), .A(n13275), .ZN(P2_U2890) );
  NAND3_X1 U15167 ( .A1(n16715), .A2(n13276), .A3(n16719), .ZN(n13280) );
  INV_X1 U15168 ( .A(n13277), .ZN(n13278) );
  NAND3_X1 U15169 ( .A1(n13280), .A2(n13279), .A3(n13278), .ZN(n13282) );
  NAND2_X1 U15170 ( .A1(n13288), .A2(n13287), .ZN(n13289) );
  XNOR2_X1 U15171 ( .A(n13290), .B(n13289), .ZN(n13349) );
  AND2_X1 U15172 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16664) );
  NAND2_X1 U15173 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16664), .ZN(
        n16649) );
  NOR2_X1 U15174 ( .A1(n16649), .A2(n12451), .ZN(n13291) );
  OAI21_X1 U15175 ( .B1(n13293), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n13292), .ZN(n13332) );
  AOI21_X1 U15176 ( .B1(n13294), .B2(n15505), .A(n16520), .ZN(n16451) );
  AND2_X1 U15177 ( .A1(n16402), .A2(n16447), .ZN(n13295) );
  OR2_X1 U15178 ( .A1(n13295), .A2(n11079), .ZN(n16444) );
  NOR2_X1 U15179 ( .A1(n18680), .A2(n13296), .ZN(n13343) );
  AOI21_X1 U15180 ( .B1(n16750), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n13343), .ZN(n13297) );
  OAI21_X1 U15181 ( .B1(n16782), .B2(n16444), .A(n13297), .ZN(n13298) );
  OAI211_X1 U15182 ( .C1(n13349), .C2(n17411), .A(n11400), .B(n13299), .ZN(
        P2_U2993) );
  AOI21_X1 U15183 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13302) );
  INV_X1 U15184 ( .A(n13300), .ZN(n13301) );
  NOR2_X1 U15185 ( .A1(n13302), .A2(n13301), .ZN(n13328) );
  OAI21_X1 U15186 ( .B1(n13304), .B2(n13303), .A(n12350), .ZN(n18613) );
  NOR2_X1 U15187 ( .A1(n18680), .A2(n17494), .ZN(n13316) );
  OAI21_X1 U15188 ( .B1(n11016), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15277), .ZN(n18619) );
  NOR2_X1 U15189 ( .A1(n16782), .A2(n18619), .ZN(n13305) );
  AOI211_X1 U15190 ( .C1(n16750), .C2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n13316), .B(n13305), .ZN(n13306) );
  OAI21_X1 U15191 ( .B1(n18613), .B2(n17410), .A(n13306), .ZN(n13307) );
  AOI21_X1 U15192 ( .B1(n13328), .B2(n16766), .A(n13307), .ZN(n13313) );
  NAND2_X1 U15193 ( .A1(n13309), .A2(n13308), .ZN(n13311) );
  NAND2_X1 U15194 ( .A1(n13313), .A2(n13312), .ZN(P2_U2985) );
  INV_X1 U15195 ( .A(n13323), .ZN(n13315) );
  NOR2_X1 U15196 ( .A1(n13315), .A2(n13314), .ZN(n15705) );
  INV_X1 U15197 ( .A(n15705), .ZN(n13319) );
  INV_X1 U15198 ( .A(n13316), .ZN(n13318) );
  INV_X1 U15199 ( .A(n13320), .ZN(n13326) );
  NAND2_X1 U15200 ( .A1(n13323), .A2(n12524), .ZN(n16790) );
  NAND2_X1 U15201 ( .A1(n16787), .A2(n16790), .ZN(n13366) );
  INV_X1 U15202 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13321) );
  AND2_X1 U15203 ( .A1(n13321), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13322) );
  NAND2_X1 U15204 ( .A1(n13323), .A2(n13322), .ZN(n13363) );
  INV_X1 U15205 ( .A(n13363), .ZN(n13324) );
  OAI21_X1 U15206 ( .B1(n13366), .B2(n13324), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13325) );
  OAI211_X1 U15207 ( .C1(n18613), .C2(n18666), .A(n13326), .B(n13325), .ZN(
        n13327) );
  AOI21_X1 U15208 ( .B1(n13328), .B2(n15725), .A(n13327), .ZN(n13331) );
  NAND2_X1 U15209 ( .A1(n13331), .A2(n13330), .ZN(P2_U3017) );
  INV_X1 U15210 ( .A(n16451), .ZN(n13333) );
  NOR2_X1 U15211 ( .A1(n13333), .A2(n18666), .ZN(n13347) );
  OR2_X1 U15212 ( .A1(n13335), .A2(n13336), .ZN(n13337) );
  NAND2_X1 U15213 ( .A1(n13334), .A2(n13337), .ZN(n16448) );
  INV_X1 U15214 ( .A(n16857), .ZN(n15689) );
  NAND2_X1 U15215 ( .A1(n16990), .A2(n15689), .ZN(n16855) );
  INV_X1 U15216 ( .A(n13338), .ZN(n13339) );
  NOR3_X1 U15217 ( .A1(n16855), .A2(n13340), .A3(n13339), .ZN(n13342) );
  INV_X1 U15218 ( .A(n16848), .ZN(n13341) );
  OAI21_X1 U15219 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13342), .A(
        n13341), .ZN(n13345) );
  INV_X1 U15220 ( .A(n13343), .ZN(n13344) );
  OAI211_X1 U15221 ( .C1(n18662), .C2(n16448), .A(n13345), .B(n13344), .ZN(
        n13346) );
  OAI211_X1 U15222 ( .C1(n13349), .C2(n18664), .A(n11398), .B(n13348), .ZN(
        P2_U3025) );
  INV_X1 U15223 ( .A(n13354), .ZN(n13355) );
  XNOR2_X1 U15224 ( .A(n13357), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15756) );
  XNOR2_X1 U15225 ( .A(n13358), .B(n13359), .ZN(n18602) );
  INV_X1 U15226 ( .A(n13360), .ZN(n13361) );
  OAI21_X1 U15227 ( .B1(n16422), .B2(n13362), .A(n13361), .ZN(n18611) );
  NOR2_X1 U15228 ( .A1(n18680), .A2(n17493), .ZN(n15753) );
  INV_X1 U15229 ( .A(n15753), .ZN(n13364) );
  OAI211_X1 U15230 ( .C1(n18611), .C2(n18662), .A(n13364), .B(n13363), .ZN(
        n13365) );
  AOI21_X1 U15231 ( .B1(n13366), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n13365), .ZN(n13367) );
  OAI21_X1 U15232 ( .B1(n18602), .B2(n18666), .A(n13367), .ZN(n13368) );
  AOI21_X1 U15233 ( .B1(n15756), .B2(n15725), .A(n13368), .ZN(n13369) );
  OAI21_X1 U15234 ( .B1(n15758), .B2(n18664), .A(n13369), .ZN(P2_U3018) );
  INV_X1 U15235 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13797) );
  AND2_X4 U15236 ( .A1(n14764), .A2(n14762), .ZN(n13438) );
  AOI22_X1 U15238 ( .A1(n13519), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10975), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13372) );
  NOR2_X4 U15239 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14763) );
  AND2_X4 U15240 ( .A1(n13381), .A2(n14764), .ZN(n13444) );
  AND2_X4 U15241 ( .A1(n14762), .A2(n14763), .ZN(n13560) );
  AOI22_X1 U15242 ( .A1(n13514), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13377) );
  AOI22_X1 U15243 ( .A1(n13451), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13376) );
  AND2_X4 U15244 ( .A1(n13381), .A2(n14763), .ZN(n13534) );
  AOI22_X1 U15245 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13450), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13385) );
  AOI22_X1 U15246 ( .A1(n13431), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13383) );
  AOI22_X1 U15247 ( .A1(n13432), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13604), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13389) );
  AOI22_X1 U15248 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10975), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13386) );
  AOI22_X1 U15249 ( .A1(n13432), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13431), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13395) );
  AOI22_X1 U15250 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13450), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13394) );
  AOI22_X1 U15251 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13451), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13393) );
  AOI22_X1 U15252 ( .A1(n13443), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13399) );
  AOI22_X1 U15253 ( .A1(n13514), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13398) );
  AOI22_X1 U15254 ( .A1(n11417), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10975), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13397) );
  NAND2_X2 U15255 ( .A1(n13401), .A2(n13400), .ZN(n13475) );
  AOI22_X1 U15256 ( .A1(n13514), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13405) );
  AOI22_X1 U15257 ( .A1(n13458), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13404) );
  AOI22_X1 U15258 ( .A1(n11417), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10975), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U15259 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13406) );
  NAND2_X2 U15260 ( .A1(n13410), .A2(n11039), .ZN(n13504) );
  INV_X2 U15261 ( .A(n13504), .ZN(n13844) );
  AOI22_X1 U15262 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13414) );
  AOI22_X1 U15263 ( .A1(n13514), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13443), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U15264 ( .A1(n13432), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13431), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13412) );
  AOI22_X1 U15265 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13451), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13411) );
  AND4_X2 U15266 ( .A1(n13414), .A2(n13411), .A3(n13412), .A4(n13413), .ZN(
        n13419) );
  AOI22_X1 U15267 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13450), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13418) );
  AOI22_X1 U15268 ( .A1(n13458), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U15269 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U15270 ( .A1(n11417), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10975), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13415) );
  NAND2_X1 U15271 ( .A1(n13844), .A2(n13473), .ZN(n13495) );
  AOI22_X1 U15272 ( .A1(n13432), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13422) );
  AOI22_X1 U15273 ( .A1(n13458), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13421) );
  AOI22_X1 U15274 ( .A1(n11417), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13420) );
  AOI22_X1 U15275 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10975), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13427) );
  AOI22_X1 U15276 ( .A1(n13431), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13604), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13425) );
  AOI22_X1 U15277 ( .A1(n13450), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13451), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13424) );
  NAND2_X2 U15278 ( .A1(n13428), .A2(n11419), .ZN(n13968) );
  AND2_X2 U15279 ( .A1(n14661), .A2(n13430), .ZN(n13845) );
  NAND2_X1 U15280 ( .A1(n13431), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13437) );
  NAND2_X1 U15281 ( .A1(n13432), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13436) );
  NAND2_X1 U15282 ( .A1(n10974), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13435) );
  NAND2_X1 U15283 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13434) );
  NAND2_X1 U15284 ( .A1(n13458), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13442) );
  NAND2_X1 U15285 ( .A1(n13560), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13441) );
  NAND2_X1 U15286 ( .A1(n13514), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13440) );
  NAND2_X1 U15287 ( .A1(n13438), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13439) );
  NAND2_X1 U15288 ( .A1(n11417), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13449) );
  NAND2_X1 U15289 ( .A1(n13443), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13448) );
  NAND2_X1 U15290 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13447) );
  NAND2_X1 U15291 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13446) );
  NAND2_X1 U15292 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13454) );
  NAND2_X1 U15293 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13453) );
  NAND2_X1 U15294 ( .A1(n13451), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13452) );
  NAND2_X1 U15295 ( .A1(n21611), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21619) );
  INV_X1 U15296 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n13456) );
  NAND2_X1 U15297 ( .A1(n13456), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U15298 ( .A1(n13443), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13462) );
  AOI22_X1 U15299 ( .A1(n13519), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10975), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13461) );
  AOI22_X1 U15300 ( .A1(n13514), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13460) );
  AOI22_X1 U15301 ( .A1(n13458), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13459) );
  AOI22_X1 U15302 ( .A1(n13432), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13431), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13465) );
  AOI22_X1 U15303 ( .A1(n13604), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13464) );
  AOI22_X1 U15304 ( .A1(n14419), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13450), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13463) );
  NAND3_X4 U15305 ( .A1(n11042), .A2(n13466), .A3(n11020), .ZN(n13491) );
  NOR2_X1 U15306 ( .A1(n13491), .A2(n13786), .ZN(n13467) );
  NAND2_X1 U15307 ( .A1(n13506), .A2(n13467), .ZN(n14753) );
  INV_X1 U15308 ( .A(n14753), .ZN(n13469) );
  NAND2_X1 U15309 ( .A1(n13968), .A2(n13831), .ZN(n14889) );
  INV_X1 U15310 ( .A(n14889), .ZN(n13468) );
  NAND2_X1 U15311 ( .A1(n13470), .A2(n13484), .ZN(n13487) );
  INV_X1 U15312 ( .A(n13487), .ZN(n13472) );
  NAND2_X1 U15313 ( .A1(n13472), .A2(n13471), .ZN(n13489) );
  NAND2_X1 U15314 ( .A1(n13489), .A2(n13473), .ZN(n13481) );
  INV_X1 U15315 ( .A(n13475), .ZN(n13474) );
  NAND2_X1 U15316 ( .A1(n13484), .A2(n13486), .ZN(n13482) );
  NAND2_X1 U15317 ( .A1(n13484), .A2(n13476), .ZN(n13477) );
  NAND2_X1 U15318 ( .A1(n13477), .A2(n13844), .ZN(n13478) );
  OAI21_X1 U15319 ( .B1(n13482), .B2(n13844), .A(n13478), .ZN(n13479) );
  NOR2_X1 U15320 ( .A1(n13482), .A2(n13860), .ZN(n13483) );
  NAND2_X1 U15321 ( .A1(n22117), .A2(n13831), .ZN(n13485) );
  AND2_X1 U15322 ( .A1(n13485), .A2(n13968), .ZN(n13832) );
  NAND2_X1 U15323 ( .A1(n13832), .A2(n13474), .ZN(n13492) );
  INV_X1 U15324 ( .A(n13492), .ZN(n13488) );
  NAND2_X1 U15326 ( .A1(n13836), .A2(n13490), .ZN(n13493) );
  OR2_X1 U15327 ( .A1(n13482), .A2(n13865), .ZN(n14754) );
  AND3_X1 U15328 ( .A1(n13493), .A2(n14754), .A3(n13508), .ZN(n13498) );
  INV_X1 U15329 ( .A(n10997), .ZN(n13496) );
  MUX2_X1 U15330 ( .A(n14533), .B(n13841), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n13499) );
  INV_X1 U15331 ( .A(n13865), .ZN(n15733) );
  AOI21_X1 U15332 ( .B1(n13473), .B2(n13487), .A(n15733), .ZN(n13501) );
  MUX2_X1 U15333 ( .A(n13502), .B(n13501), .S(n15814), .Z(n13503) );
  INV_X1 U15334 ( .A(n13503), .ZN(n13511) );
  NAND3_X1 U15335 ( .A1(n13836), .A2(n13490), .A3(n13491), .ZN(n13509) );
  CLKBUF_X1 U15336 ( .A(n13504), .Z(n13505) );
  NAND2_X1 U15337 ( .A1(n16385), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20046) );
  AOI21_X1 U15338 ( .B1(n13505), .B2(n13860), .A(n20046), .ZN(n13507) );
  NAND2_X1 U15339 ( .A1(n13506), .A2(n22167), .ZN(n13977) );
  AND4_X1 U15340 ( .A1(n13509), .A2(n13508), .A3(n13507), .A4(n13977), .ZN(
        n13510) );
  NAND2_X1 U15341 ( .A1(n13511), .A2(n13510), .ZN(n13557) );
  INV_X1 U15342 ( .A(n13557), .ZN(n13512) );
  NAND2_X1 U15343 ( .A1(n14037), .A2(n17186), .ZN(n13543) );
  AOI22_X1 U15344 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13513), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13518) );
  AOI22_X1 U15345 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13517) );
  AOI22_X1 U15346 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13516) );
  AOI22_X1 U15347 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13451), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13515) );
  NAND4_X1 U15348 ( .A1(n13518), .A2(n13517), .A3(n13516), .A4(n13515), .ZN(
        n13528) );
  AOI22_X1 U15349 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14478), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13526) );
  INV_X1 U15350 ( .A(n14770), .ZN(n13521) );
  AOI22_X1 U15351 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13525) );
  AOI22_X1 U15352 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13524) );
  AOI22_X1 U15353 ( .A1(n13560), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13523) );
  NAND4_X1 U15354 ( .A1(n13526), .A2(n13525), .A3(n13524), .A4(n13523), .ZN(
        n13527) );
  AOI22_X1 U15355 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13529), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13533) );
  AOI22_X1 U15356 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14478), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13532) );
  AOI22_X1 U15357 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13531) );
  AOI22_X1 U15358 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n14484), .B1(
        n13451), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13530) );
  NAND4_X1 U15359 ( .A1(n13533), .A2(n13532), .A3(n13531), .A4(n13530), .ZN(
        n13540) );
  AOI22_X1 U15360 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n13534), .B1(
        n13513), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13538) );
  AOI22_X1 U15361 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13537) );
  AOI22_X1 U15362 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13536) );
  AOI22_X1 U15363 ( .A1(n13560), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13535) );
  NAND4_X1 U15364 ( .A1(n13538), .A2(n13537), .A3(n13536), .A4(n13535), .ZN(
        n13539) );
  XNOR2_X1 U15365 ( .A(n13723), .B(n13572), .ZN(n13541) );
  NAND2_X1 U15366 ( .A1(n13541), .A2(n13583), .ZN(n13542) );
  INV_X1 U15367 ( .A(n13572), .ZN(n13546) );
  NAND2_X1 U15368 ( .A1(n13814), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13545) );
  AOI21_X1 U15369 ( .B1(n13474), .B2(n13739), .A(n17186), .ZN(n13544) );
  XNOR2_X2 U15370 ( .A(n13580), .B(n13579), .ZN(n14035) );
  INV_X1 U15371 ( .A(n13821), .ZN(n13550) );
  INV_X1 U15372 ( .A(n13547), .ZN(n17177) );
  NAND2_X1 U15373 ( .A1(n21737), .A2(n13473), .ZN(n13619) );
  OAI21_X1 U15374 ( .B1(n17177), .B2(n13572), .A(n13619), .ZN(n13548) );
  INV_X1 U15375 ( .A(n13548), .ZN(n13549) );
  XNOR2_X1 U15376 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21762) );
  NAND2_X1 U15377 ( .A1(n17179), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13592) );
  OAI21_X1 U15378 ( .B1(n14533), .B2(n21762), .A(n13592), .ZN(n13552) );
  INV_X1 U15379 ( .A(n13552), .ZN(n13553) );
  INV_X1 U15380 ( .A(n13555), .ZN(n13556) );
  NAND2_X1 U15381 ( .A1(n13558), .A2(n13557), .ZN(n13559) );
  OR2_X2 U15382 ( .A1(n21771), .A2(n13559), .ZN(n13596) );
  NAND2_X1 U15383 ( .A1(n13559), .A2(n21771), .ZN(n21752) );
  AOI22_X1 U15384 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13534), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13564) );
  AOI22_X1 U15385 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13563) );
  AOI22_X1 U15386 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13562) );
  AOI22_X1 U15387 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13561) );
  NAND4_X1 U15388 ( .A1(n13564), .A2(n13563), .A3(n13562), .A4(n13561), .ZN(
        n13570) );
  AOI22_X1 U15389 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13568) );
  AOI22_X1 U15390 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13451), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U15391 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13566) );
  AOI22_X1 U15392 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13565) );
  NAND4_X1 U15393 ( .A1(n13568), .A2(n13567), .A3(n13566), .A4(n13565), .ZN(
        n13569) );
  NAND2_X1 U15394 ( .A1(n13583), .A2(n13584), .ZN(n13571) );
  NAND2_X1 U15395 ( .A1(n13572), .A2(n13584), .ZN(n13646) );
  OAI21_X1 U15396 ( .B1(n13584), .B2(n13572), .A(n13646), .ZN(n13573) );
  OAI211_X1 U15397 ( .C1(n13573), .C2(n17177), .A(n13496), .B(n13786), .ZN(
        n13574) );
  INV_X1 U15398 ( .A(n13574), .ZN(n13575) );
  INV_X1 U15399 ( .A(n13576), .ZN(n13577) );
  OR2_X1 U15400 ( .A1(n11005), .A2(n13577), .ZN(n13578) );
  INV_X1 U15401 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21301) );
  NAND2_X1 U15402 ( .A1(n13580), .A2(n13579), .ZN(n13581) );
  NAND2_X1 U15403 ( .A1(n13583), .A2(n13739), .ZN(n13735) );
  NAND2_X1 U15404 ( .A1(n13581), .A2(n13735), .ZN(n13589) );
  INV_X1 U15405 ( .A(n13589), .ZN(n13582) );
  XNOR2_X1 U15406 ( .A(n13582), .B(n13590), .ZN(n13588) );
  NAND2_X1 U15407 ( .A1(n13583), .A2(n13723), .ZN(n13586) );
  NAND3_X1 U15408 ( .A1(n21737), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n13584), 
        .ZN(n13585) );
  NAND2_X1 U15409 ( .A1(n13586), .A2(n13585), .ZN(n14028) );
  INV_X1 U15410 ( .A(n13592), .ZN(n13594) );
  OAI21_X1 U15411 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13594), .A(
        n13593), .ZN(n13595) );
  NAND2_X1 U15412 ( .A1(n13597), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13601) );
  INV_X1 U15413 ( .A(n14533), .ZN(n13627) );
  NAND2_X1 U15414 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13598) );
  NAND2_X1 U15415 ( .A1(n21875), .A2(n13598), .ZN(n13599) );
  NOR2_X1 U15416 ( .A1(n21875), .A2(n21763), .ZN(n21916) );
  NAND2_X1 U15417 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21916), .ZN(
        n13625) );
  AOI22_X1 U15418 ( .A1(n13627), .A2(n21738), .B1(n17179), .B2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13600) );
  AOI22_X1 U15419 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13608) );
  AOI22_X1 U15420 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13607) );
  AOI22_X1 U15421 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13606) );
  AOI22_X1 U15422 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13605) );
  NAND4_X1 U15423 ( .A1(n13608), .A2(n13607), .A3(n13606), .A4(n13605), .ZN(
        n13614) );
  AOI22_X1 U15424 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13612) );
  AOI22_X1 U15425 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13611) );
  AOI22_X1 U15426 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13610) );
  AOI22_X1 U15427 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13609) );
  NAND4_X1 U15428 ( .A1(n13612), .A2(n13611), .A3(n13610), .A4(n13609), .ZN(
        n13613) );
  AOI22_X1 U15429 ( .A1(n13814), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13794), .B2(n13618), .ZN(n13615) );
  INV_X1 U15430 ( .A(n13618), .ZN(n13645) );
  XNOR2_X1 U15431 ( .A(n13646), .B(n13645), .ZN(n13621) );
  INV_X1 U15432 ( .A(n13619), .ZN(n13620) );
  AOI21_X1 U15433 ( .B1(n13621), .B2(n13547), .A(n13620), .ZN(n13622) );
  NAND2_X1 U15434 ( .A1(n13623), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13624) );
  INV_X1 U15435 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21317) );
  INV_X1 U15436 ( .A(n13643), .ZN(n13642) );
  NAND2_X1 U15437 ( .A1(n13597), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13629) );
  INV_X1 U15438 ( .A(n13625), .ZN(n21913) );
  NAND2_X1 U15439 ( .A1(n21913), .A2(n13778), .ZN(n21811) );
  NAND2_X1 U15440 ( .A1(n13625), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13626) );
  NAND2_X1 U15441 ( .A1(n21811), .A2(n13626), .ZN(n21824) );
  AOI22_X1 U15442 ( .A1(n13627), .A2(n21824), .B1(n17179), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13628) );
  XNOR2_X2 U15443 ( .A(n14748), .B(n21784), .ZN(n21823) );
  AOI22_X1 U15444 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13513), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13633) );
  AOI22_X1 U15445 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13632) );
  AOI22_X1 U15446 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13631) );
  AOI22_X1 U15447 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13630) );
  NAND4_X1 U15448 ( .A1(n13633), .A2(n13632), .A3(n13631), .A4(n13630), .ZN(
        n13639) );
  AOI22_X1 U15449 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13637) );
  AOI22_X1 U15450 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13636) );
  AOI22_X1 U15451 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13635) );
  INV_X1 U15452 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U15453 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13634) );
  NAND4_X1 U15454 ( .A1(n13637), .A2(n13636), .A3(n13635), .A4(n13634), .ZN(
        n13638) );
  AOI22_X1 U15455 ( .A1(n13814), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13794), .B2(n13664), .ZN(n13640) );
  INV_X1 U15456 ( .A(n14927), .ZN(n14928) );
  NAND2_X1 U15457 ( .A1(n13643), .A2(n14928), .ZN(n13644) );
  OR2_X1 U15458 ( .A1(n21821), .A2(n13550), .ZN(n13650) );
  NAND2_X1 U15459 ( .A1(n13646), .A2(n13645), .ZN(n13665) );
  INV_X1 U15460 ( .A(n13664), .ZN(n13647) );
  XNOR2_X1 U15461 ( .A(n13665), .B(n13647), .ZN(n13648) );
  NAND2_X1 U15462 ( .A1(n13648), .A2(n13547), .ZN(n13649) );
  NAND2_X1 U15463 ( .A1(n13650), .A2(n13649), .ZN(n15093) );
  NAND2_X1 U15464 ( .A1(n13651), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13652) );
  INV_X1 U15465 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21311) );
  INV_X1 U15466 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U15467 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13513), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13656) );
  AOI22_X1 U15468 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13655) );
  AOI22_X1 U15469 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13654) );
  AOI22_X1 U15470 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13653) );
  NAND4_X1 U15471 ( .A1(n13656), .A2(n13655), .A3(n13654), .A4(n13653), .ZN(
        n13662) );
  AOI22_X1 U15472 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13660) );
  AOI22_X1 U15473 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13659) );
  AOI22_X1 U15474 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U15475 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13657) );
  NAND4_X1 U15476 ( .A1(n13660), .A2(n13659), .A3(n13658), .A4(n13657), .ZN(
        n13661) );
  NAND2_X1 U15477 ( .A1(n14065), .A2(n13821), .ZN(n13669) );
  NAND2_X1 U15478 ( .A1(n13665), .A2(n13664), .ZN(n13688) );
  XNOR2_X1 U15479 ( .A(n13688), .B(n13666), .ZN(n13667) );
  NAND2_X1 U15480 ( .A1(n13667), .A2(n13547), .ZN(n13668) );
  NAND2_X1 U15481 ( .A1(n13669), .A2(n13668), .ZN(n19992) );
  NAND2_X1 U15482 ( .A1(n13670), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13671) );
  INV_X1 U15483 ( .A(n13672), .ZN(n13674) );
  NAND2_X1 U15484 ( .A1(n13674), .A2(n13673), .ZN(n13694) );
  INV_X1 U15485 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13686) );
  AOI22_X1 U15486 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13678) );
  AOI22_X1 U15487 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13677) );
  AOI22_X1 U15488 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13676) );
  AOI22_X1 U15489 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13675) );
  NAND4_X1 U15490 ( .A1(n13678), .A2(n13677), .A3(n13676), .A4(n13675), .ZN(
        n13684) );
  AOI22_X1 U15491 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13682) );
  AOI22_X1 U15492 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13681) );
  AOI22_X1 U15493 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13680) );
  AOI22_X1 U15494 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13679) );
  NAND4_X1 U15495 ( .A1(n13682), .A2(n13681), .A3(n13680), .A4(n13679), .ZN(
        n13683) );
  INV_X1 U15496 ( .A(n13715), .ZN(n13685) );
  XNOR2_X1 U15497 ( .A(n13694), .B(n13695), .ZN(n14072) );
  NAND2_X1 U15498 ( .A1(n14072), .A2(n13821), .ZN(n13691) );
  OR2_X1 U15499 ( .A1(n13688), .A2(n13687), .ZN(n13714) );
  XNOR2_X1 U15500 ( .A(n13714), .B(n13715), .ZN(n13689) );
  NAND2_X1 U15501 ( .A1(n13689), .A2(n13547), .ZN(n13690) );
  NAND2_X1 U15502 ( .A1(n13691), .A2(n13690), .ZN(n13692) );
  INV_X1 U15503 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13984) );
  XNOR2_X1 U15504 ( .A(n13692), .B(n13984), .ZN(n19998) );
  NAND2_X1 U15505 ( .A1(n13692), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13693) );
  INV_X1 U15506 ( .A(n13694), .ZN(n13696) );
  NAND2_X1 U15507 ( .A1(n13814), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13709) );
  AOI22_X1 U15508 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13513), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U15509 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13699) );
  AOI22_X1 U15510 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13698) );
  AOI22_X1 U15511 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13697) );
  NAND4_X1 U15512 ( .A1(n13700), .A2(n13699), .A3(n13698), .A4(n13697), .ZN(
        n13706) );
  AOI22_X1 U15513 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13704) );
  AOI22_X1 U15514 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13703) );
  AOI22_X1 U15515 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U15516 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13701) );
  NAND4_X1 U15517 ( .A1(n13704), .A2(n13703), .A3(n13702), .A4(n13701), .ZN(
        n13705) );
  INV_X1 U15518 ( .A(n13727), .ZN(n13707) );
  NAND2_X1 U15519 ( .A1(n13713), .A2(n13712), .ZN(n14073) );
  NAND3_X1 U15520 ( .A1(n13737), .A2(n13821), .A3(n14073), .ZN(n13719) );
  INV_X1 U15521 ( .A(n13714), .ZN(n13716) );
  NAND2_X1 U15522 ( .A1(n13716), .A2(n13715), .ZN(n13726) );
  XNOR2_X1 U15523 ( .A(n13726), .B(n13727), .ZN(n13717) );
  NAND2_X1 U15524 ( .A1(n13717), .A2(n13547), .ZN(n13718) );
  NAND2_X1 U15525 ( .A1(n13719), .A2(n13718), .ZN(n13721) );
  XNOR2_X1 U15526 ( .A(n13721), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n20004) );
  INV_X1 U15527 ( .A(n20004), .ZN(n13720) );
  OR2_X1 U15528 ( .A1(n13721), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13722) );
  INV_X1 U15529 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13724) );
  OAI22_X1 U15530 ( .A1(n14027), .A2(n13724), .B1(n13806), .B2(n13723), .ZN(
        n13725) );
  NAND2_X1 U15531 ( .A1(n14020), .A2(n13821), .ZN(n13731) );
  INV_X1 U15532 ( .A(n13726), .ZN(n13728) );
  NAND2_X1 U15533 ( .A1(n13728), .A2(n13727), .ZN(n13738) );
  XNOR2_X1 U15534 ( .A(n13738), .B(n13739), .ZN(n13729) );
  NAND2_X1 U15535 ( .A1(n13729), .A2(n13547), .ZN(n13730) );
  NAND2_X1 U15536 ( .A1(n13731), .A2(n13730), .ZN(n13733) );
  XNOR2_X1 U15537 ( .A(n13733), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n20010) );
  INV_X1 U15538 ( .A(n20010), .ZN(n13732) );
  NAND2_X1 U15539 ( .A1(n13733), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13734) );
  NOR2_X1 U15540 ( .A1(n13735), .A2(n13550), .ZN(n13736) );
  INV_X1 U15541 ( .A(n13738), .ZN(n13740) );
  NAND3_X1 U15542 ( .A1(n13740), .A2(n13547), .A3(n13739), .ZN(n13741) );
  NAND2_X1 U15543 ( .A1(n13755), .A2(n13741), .ZN(n13742) );
  XNOR2_X1 U15544 ( .A(n13742), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15530) );
  OR2_X1 U15545 ( .A1(n13742), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13743) );
  XNOR2_X1 U15546 ( .A(n13755), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15553) );
  INV_X1 U15547 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13893) );
  NAND2_X1 U15548 ( .A1(n16336), .A2(n13893), .ZN(n13744) );
  INV_X1 U15549 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16134) );
  XNOR2_X1 U15550 ( .A(n13755), .B(n16134), .ZN(n16162) );
  NAND2_X1 U15551 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13745) );
  AND2_X1 U15552 ( .A1(n13755), .A2(n13745), .ZN(n16158) );
  INV_X1 U15553 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16133) );
  INV_X1 U15554 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16149) );
  AND2_X1 U15555 ( .A1(n16336), .A2(n16149), .ZN(n13746) );
  AND2_X1 U15556 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16302) );
  NAND2_X1 U15557 ( .A1(n16302), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16241) );
  INV_X1 U15558 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13981) );
  INV_X1 U15559 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16342) );
  AND2_X1 U15560 ( .A1(n13981), .A2(n16342), .ZN(n13748) );
  OR2_X1 U15561 ( .A1(n13755), .A2(n16133), .ZN(n16159) );
  INV_X1 U15562 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16138) );
  NAND3_X1 U15563 ( .A1(n16149), .A2(n16134), .A3(n16138), .ZN(n16296) );
  INV_X1 U15564 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13917) );
  NAND2_X1 U15565 ( .A1(n21353), .A2(n13917), .ZN(n13749) );
  NAND2_X1 U15566 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16242) );
  NAND2_X1 U15567 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13750) );
  NOR2_X1 U15568 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13752) );
  INV_X1 U15569 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16232) );
  AND2_X1 U15570 ( .A1(n13752), .A2(n16232), .ZN(n13761) );
  NAND2_X1 U15571 ( .A1(n13759), .A2(n13761), .ZN(n13756) );
  XNOR2_X1 U15572 ( .A(n13755), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16127) );
  INV_X1 U15573 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13923) );
  INV_X1 U15574 ( .A(n16113), .ZN(n13754) );
  INV_X1 U15575 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16276) );
  INV_X1 U15576 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16122) );
  INV_X1 U15577 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16253) );
  OAI22_X1 U15578 ( .A1(n13760), .A2(n13756), .B1(n13759), .B2(n16337), .ZN(
        n13757) );
  AND2_X1 U15579 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16201) );
  NAND2_X1 U15580 ( .A1(n16201), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13998) );
  NAND2_X1 U15581 ( .A1(n16336), .A2(n13998), .ZN(n16057) );
  NAND2_X1 U15582 ( .A1(n13757), .A2(n16057), .ZN(n16081) );
  INV_X1 U15583 ( .A(n16081), .ZN(n13758) );
  INV_X1 U15584 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16202) );
  INV_X1 U15585 ( .A(n13761), .ZN(n16058) );
  NAND2_X1 U15586 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16181) );
  INV_X1 U15587 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16194) );
  INV_X1 U15588 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16063) );
  NAND2_X1 U15589 ( .A1(n16194), .A2(n16063), .ZN(n16180) );
  INV_X1 U15590 ( .A(n16180), .ZN(n13763) );
  NOR2_X1 U15591 ( .A1(n16337), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14006) );
  XNOR2_X1 U15592 ( .A(n13755), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13768) );
  INV_X1 U15593 ( .A(n13768), .ZN(n13766) );
  NOR2_X1 U15594 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13764) );
  OR2_X1 U15595 ( .A1(n13764), .A2(n16336), .ZN(n13765) );
  NAND2_X1 U15596 ( .A1(n13767), .A2(n11069), .ZN(n13775) );
  INV_X1 U15597 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16049) );
  NAND2_X1 U15598 ( .A1(n16336), .A2(n16049), .ZN(n13770) );
  NAND3_X1 U15599 ( .A1(n13769), .A2(n13768), .A3(n13770), .ZN(n13774) );
  INV_X1 U15600 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14000) );
  NOR2_X1 U15601 ( .A1(n16336), .A2(n14000), .ZN(n16042) );
  INV_X1 U15602 ( .A(n13770), .ZN(n13771) );
  AOI211_X1 U15603 ( .C1(n16337), .C2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16042), .B(n13771), .ZN(n13772) );
  NAND3_X1 U15604 ( .A1(n13775), .A2(n13774), .A3(n13773), .ZN(n14541) );
  MUX2_X1 U15605 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n21875), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13789) );
  NAND2_X1 U15606 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21885), .ZN(
        n13798) );
  NOR2_X1 U15607 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21763), .ZN(
        n13776) );
  NOR2_X1 U15608 ( .A1(n13798), .A2(n13776), .ZN(n13777) );
  NAND2_X1 U15609 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14922), .ZN(
        n13780) );
  INV_X1 U15610 ( .A(n13818), .ZN(n13785) );
  MUX2_X1 U15611 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n13778), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13781) );
  XNOR2_X1 U15612 ( .A(n13782), .B(n13781), .ZN(n13784) );
  AOI22_X1 U15613 ( .A1(n13785), .A2(n13823), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17186), .ZN(n13816) );
  INV_X1 U15614 ( .A(n13823), .ZN(n13813) );
  NAND2_X1 U15615 ( .A1(n21935), .A2(n13786), .ZN(n13787) );
  NAND2_X1 U15616 ( .A1(n15814), .A2(n13787), .ZN(n13807) );
  XNOR2_X1 U15617 ( .A(n13789), .B(n13788), .ZN(n13822) );
  NOR3_X1 U15618 ( .A1(n11174), .A2(n13822), .A3(n13806), .ZN(n13812) );
  XNOR2_X1 U15619 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n13798), .ZN(
        n13790) );
  XNOR2_X1 U15620 ( .A(n13790), .B(n21763), .ZN(n13824) );
  INV_X1 U15621 ( .A(n13824), .ZN(n13791) );
  OAI211_X1 U15622 ( .C1(n21935), .C2(n13806), .A(n13791), .B(n13800), .ZN(
        n13796) );
  INV_X1 U15623 ( .A(n13792), .ZN(n13793) );
  OAI21_X1 U15624 ( .B1(n13794), .B2(n13793), .A(n13824), .ZN(n13795) );
  NAND2_X1 U15625 ( .A1(n13796), .A2(n13795), .ZN(n13810) );
  INV_X1 U15626 ( .A(n13798), .ZN(n13799) );
  AOI21_X1 U15627 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n13797), .A(
        n13799), .ZN(n13801) );
  OAI21_X1 U15628 ( .B1(n21737), .B2(n13482), .A(n13801), .ZN(n13805) );
  NAND3_X1 U15629 ( .A1(n21935), .A2(n13800), .A3(n13824), .ZN(n13804) );
  INV_X1 U15630 ( .A(n13801), .ZN(n13802) );
  OAI21_X1 U15631 ( .B1(n13806), .B2(n13802), .A(n13818), .ZN(n13803) );
  OAI211_X1 U15632 ( .C1(n13807), .C2(n13805), .A(n13804), .B(n13803), .ZN(
        n13809) );
  AOI21_X1 U15633 ( .B1(n13810), .B2(n13809), .A(n13808), .ZN(n13811) );
  OAI22_X1 U15634 ( .A1(n13814), .A2(n13813), .B1(n13812), .B2(n13811), .ZN(
        n13815) );
  NAND2_X1 U15635 ( .A1(n13816), .A2(n13815), .ZN(n13817) );
  NAND2_X1 U15636 ( .A1(n13821), .A2(n22167), .ZN(n13840) );
  NOR3_X1 U15637 ( .A1(n13824), .A2(n13823), .A3(n13822), .ZN(n13827) );
  INV_X1 U15638 ( .A(n13825), .ZN(n13826) );
  NAND2_X1 U15639 ( .A1(n13491), .A2(n21617), .ZN(n13829) );
  NAND4_X1 U15640 ( .A1(n14738), .A2(n13505), .A3(n21667), .A4(n13829), .ZN(
        n13839) );
  INV_X1 U15641 ( .A(n13830), .ZN(n14666) );
  OR2_X1 U15642 ( .A1(n13482), .A2(n13831), .ZN(n13833) );
  AND2_X1 U15643 ( .A1(n13833), .A2(n13832), .ZN(n13973) );
  NAND2_X1 U15644 ( .A1(n13490), .A2(n21737), .ZN(n13834) );
  NAND3_X1 U15645 ( .A1(n13973), .A2(n13496), .A3(n13834), .ZN(n13851) );
  INV_X1 U15646 ( .A(n13851), .ZN(n13837) );
  AND2_X1 U15647 ( .A1(n13840), .A2(n13860), .ZN(n13835) );
  NAND2_X1 U15648 ( .A1(n13836), .A2(n13835), .ZN(n13975) );
  NAND2_X1 U15649 ( .A1(n13837), .A2(n13975), .ZN(n13838) );
  NAND2_X1 U15650 ( .A1(n14666), .A2(n13838), .ZN(n14743) );
  OAI211_X1 U15651 ( .C1(n13843), .C2(n13840), .A(n13839), .B(n14743), .ZN(
        n13842) );
  NAND2_X1 U15652 ( .A1(n13842), .A2(n14880), .ZN(n13850) );
  INV_X1 U15653 ( .A(n21617), .ZN(n14695) );
  OAI21_X1 U15654 ( .B1(n13491), .B2(n14695), .A(n21667), .ZN(n14517) );
  INV_X1 U15655 ( .A(n14517), .ZN(n13846) );
  NAND2_X1 U15656 ( .A1(n10996), .A2(n13846), .ZN(n13847) );
  NAND3_X1 U15657 ( .A1(n13847), .A2(n13860), .A3(n14889), .ZN(n13848) );
  NAND3_X1 U15658 ( .A1(n11017), .A2(n13844), .A3(n13848), .ZN(n13849) );
  NOR2_X1 U15659 ( .A1(n13851), .A2(n13482), .ZN(n17168) );
  AND2_X1 U15660 ( .A1(n11315), .A2(n13496), .ZN(n13852) );
  NAND2_X1 U15661 ( .A1(n13852), .A2(n14152), .ZN(n14767) );
  INV_X1 U15662 ( .A(n14767), .ZN(n13853) );
  NOR2_X1 U15663 ( .A1(n17168), .A2(n13853), .ZN(n14663) );
  OR2_X1 U15664 ( .A1(n13857), .A2(n13474), .ZN(n13858) );
  NAND4_X1 U15665 ( .A1(n14663), .A2(n13855), .A3(n13856), .A4(n13858), .ZN(
        n13859) );
  INV_X1 U15666 ( .A(n13473), .ZN(n22025) );
  NAND2_X1 U15667 ( .A1(n22025), .A2(n13860), .ZN(n13881) );
  NAND2_X2 U15668 ( .A1(n13881), .A2(n10981), .ZN(n14704) );
  OAI22_X1 U15669 ( .A1(n14704), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n14721), .ZN(n15735) );
  AND2_X1 U15670 ( .A1(n14721), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13861) );
  AOI21_X1 U15671 ( .B1(n14704), .B2(P1_EBX_REG_31__SCAN_IN), .A(n13861), .ZN(
        n13862) );
  XNOR2_X1 U15672 ( .A(n15735), .B(n13862), .ZN(n13966) );
  INV_X1 U15673 ( .A(n13862), .ZN(n13863) );
  NAND2_X1 U15674 ( .A1(n13863), .A2(n10981), .ZN(n13965) );
  MUX2_X1 U15675 ( .A(n13869), .B(n10981), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n13867) );
  OR2_X1 U15676 ( .A1(n14704), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13866) );
  INV_X1 U15677 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13868) );
  OAI22_X1 U15678 ( .A1(n13881), .A2(n13868), .B1(n10981), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n14705) );
  MUX2_X1 U15679 ( .A(n13869), .B(n10981), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13870) );
  OAI21_X1 U15680 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14704), .A(
        n13870), .ZN(n13871) );
  INV_X1 U15681 ( .A(n13871), .ZN(n14863) );
  INV_X1 U15682 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13872) );
  NAND2_X1 U15683 ( .A1(n13957), .A2(n13872), .ZN(n13876) );
  NAND2_X1 U15684 ( .A1(n13881), .A2(n21317), .ZN(n13874) );
  NAND2_X1 U15685 ( .A1(n13864), .A2(n13872), .ZN(n13873) );
  NAND3_X1 U15686 ( .A1(n13874), .A2(n10981), .A3(n13873), .ZN(n13875) );
  AND2_X1 U15687 ( .A1(n13876), .A2(n13875), .ZN(n15069) );
  MUX2_X1 U15688 ( .A(n13869), .B(n10981), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13877) );
  OAI21_X1 U15689 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n14704), .A(
        n13877), .ZN(n17193) );
  INV_X1 U15690 ( .A(n13957), .ZN(n13964) );
  NAND2_X1 U15691 ( .A1(n10981), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13878) );
  NAND2_X1 U15692 ( .A1(n13881), .A2(n13878), .ZN(n13879) );
  OAI21_X1 U15693 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(n14721), .A(n13879), .ZN(
        n13880) );
  OAI21_X1 U15694 ( .B1(n13964), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13880), .ZN(
        n15151) );
  INV_X1 U15695 ( .A(n19973), .ZN(n13885) );
  NAND2_X1 U15696 ( .A1(n10981), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13882) );
  OAI211_X1 U15697 ( .C1(n14721), .C2(P1_EBX_REG_6__SCAN_IN), .A(n13881), .B(
        n13882), .ZN(n13883) );
  OAI21_X1 U15698 ( .B1(n13869), .B2(P1_EBX_REG_6__SCAN_IN), .A(n13883), .ZN(
        n19972) );
  INV_X1 U15699 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13886) );
  NAND2_X1 U15700 ( .A1(n13957), .A2(n13886), .ZN(n13890) );
  INV_X1 U15701 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21337) );
  NAND2_X1 U15702 ( .A1(n13881), .A2(n21337), .ZN(n13888) );
  NAND2_X1 U15703 ( .A1(n13864), .A2(n13886), .ZN(n13887) );
  NAND3_X1 U15704 ( .A1(n13888), .A2(n10981), .A3(n13887), .ZN(n13889) );
  AND2_X1 U15705 ( .A1(n13890), .A2(n13889), .ZN(n15206) );
  MUX2_X1 U15706 ( .A(n13869), .B(n10981), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13891) );
  OAI21_X1 U15707 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n14704), .A(
        n13891), .ZN(n13892) );
  INV_X1 U15708 ( .A(n13892), .ZN(n15375) );
  INV_X1 U15709 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15388) );
  NAND2_X1 U15710 ( .A1(n13957), .A2(n15388), .ZN(n13897) );
  NAND2_X1 U15711 ( .A1(n13881), .A2(n13893), .ZN(n13895) );
  NAND2_X1 U15712 ( .A1(n13864), .A2(n15388), .ZN(n13894) );
  NAND3_X1 U15713 ( .A1(n13895), .A2(n10981), .A3(n13894), .ZN(n13896) );
  NAND2_X1 U15714 ( .A1(n13897), .A2(n13896), .ZN(n15385) );
  NAND2_X1 U15715 ( .A1(n10981), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13898) );
  OAI211_X1 U15716 ( .C1(n14721), .C2(P1_EBX_REG_10__SCAN_IN), .A(n13881), .B(
        n13898), .ZN(n13899) );
  OAI21_X1 U15717 ( .B1(n13869), .B2(P1_EBX_REG_10__SCAN_IN), .A(n13899), .ZN(
        n16351) );
  INV_X1 U15718 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15514) );
  NAND2_X1 U15719 ( .A1(n13957), .A2(n15514), .ZN(n13903) );
  NAND2_X1 U15720 ( .A1(n13881), .A2(n16342), .ZN(n13901) );
  NAND2_X1 U15721 ( .A1(n13864), .A2(n15514), .ZN(n13900) );
  NAND3_X1 U15722 ( .A1(n13901), .A2(n10981), .A3(n13900), .ZN(n13902) );
  AND2_X1 U15723 ( .A1(n13903), .A2(n13902), .ZN(n15512) );
  NAND2_X1 U15724 ( .A1(n10981), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13904) );
  OAI211_X1 U15725 ( .C1(n14721), .C2(P1_EBX_REG_12__SCAN_IN), .A(n13881), .B(
        n13904), .ZN(n13905) );
  OAI21_X1 U15726 ( .B1(n13869), .B2(P1_EBX_REG_12__SCAN_IN), .A(n13905), .ZN(
        n16330) );
  INV_X1 U15727 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15744) );
  NAND2_X1 U15728 ( .A1(n13957), .A2(n15744), .ZN(n13909) );
  NAND2_X1 U15729 ( .A1(n13881), .A2(n16134), .ZN(n13907) );
  NAND2_X1 U15730 ( .A1(n13864), .A2(n15744), .ZN(n13906) );
  NAND3_X1 U15731 ( .A1(n13907), .A2(n10981), .A3(n13906), .ZN(n13908) );
  NAND2_X1 U15732 ( .A1(n13909), .A2(n13908), .ZN(n15739) );
  MUX2_X1 U15733 ( .A(n13869), .B(n10981), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n13910) );
  OAI21_X1 U15734 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14704), .A(
        n13910), .ZN(n15601) );
  INV_X1 U15735 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15977) );
  NAND2_X1 U15736 ( .A1(n13957), .A2(n15977), .ZN(n13914) );
  NAND2_X1 U15737 ( .A1(n13881), .A2(n16138), .ZN(n13912) );
  NAND2_X1 U15738 ( .A1(n13864), .A2(n15977), .ZN(n13911) );
  NAND3_X1 U15739 ( .A1(n13912), .A2(n10981), .A3(n13911), .ZN(n13913) );
  MUX2_X1 U15740 ( .A(n13869), .B(n10981), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n13915) );
  OAI21_X1 U15741 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n14704), .A(
        n13915), .ZN(n13916) );
  INV_X1 U15742 ( .A(n13916), .ZN(n15883) );
  INV_X1 U15743 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n19988) );
  NAND2_X1 U15744 ( .A1(n13957), .A2(n19988), .ZN(n13921) );
  NAND2_X1 U15745 ( .A1(n13881), .A2(n13917), .ZN(n13919) );
  NAND2_X1 U15746 ( .A1(n13864), .A2(n19988), .ZN(n13918) );
  NAND3_X1 U15747 ( .A1(n13919), .A2(n10981), .A3(n13918), .ZN(n13920) );
  NAND2_X1 U15748 ( .A1(n13921), .A2(n13920), .ZN(n15873) );
  INV_X1 U15749 ( .A(n14704), .ZN(n13922) );
  NAND2_X1 U15750 ( .A1(n13923), .A2(n13922), .ZN(n13925) );
  MUX2_X1 U15751 ( .A(n13869), .B(n10981), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n13924) );
  NAND2_X1 U15752 ( .A1(n13925), .A2(n13924), .ZN(n15960) );
  INV_X1 U15753 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15959) );
  NAND2_X1 U15754 ( .A1(n13957), .A2(n15959), .ZN(n13929) );
  NAND2_X1 U15755 ( .A1(n10981), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13926) );
  NAND2_X1 U15756 ( .A1(n13881), .A2(n13926), .ZN(n13927) );
  OAI21_X1 U15757 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(n14721), .A(n13927), .ZN(
        n13928) );
  MUX2_X1 U15758 ( .A(n13869), .B(n10981), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n13930) );
  OAI21_X1 U15759 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14704), .A(
        n13930), .ZN(n13931) );
  INV_X1 U15760 ( .A(n13931), .ZN(n15949) );
  INV_X1 U15761 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n13932) );
  NAND2_X1 U15762 ( .A1(n13957), .A2(n13932), .ZN(n13936) );
  NAND2_X1 U15763 ( .A1(n13881), .A2(n16253), .ZN(n13934) );
  NAND2_X1 U15764 ( .A1(n13864), .A2(n13932), .ZN(n13933) );
  NAND3_X1 U15765 ( .A1(n13934), .A2(n10981), .A3(n13933), .ZN(n13935) );
  NAND2_X1 U15766 ( .A1(n13936), .A2(n13935), .ZN(n15944) );
  NAND2_X1 U15767 ( .A1(n10981), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13937) );
  OAI211_X1 U15768 ( .C1(n14721), .C2(P1_EBX_REG_22__SCAN_IN), .A(n13881), .B(
        n13937), .ZN(n13938) );
  OAI21_X1 U15769 ( .B1(n13869), .B2(P1_EBX_REG_22__SCAN_IN), .A(n13938), .ZN(
        n15939) );
  OR2_X2 U15770 ( .A1(n15943), .A2(n15939), .ZN(n15937) );
  INV_X1 U15771 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n13939) );
  NAND2_X1 U15772 ( .A1(n13957), .A2(n13939), .ZN(n13943) );
  NAND2_X1 U15773 ( .A1(n13881), .A2(n16232), .ZN(n13941) );
  NAND2_X1 U15774 ( .A1(n13864), .A2(n13939), .ZN(n13940) );
  NAND3_X1 U15775 ( .A1(n13941), .A2(n10981), .A3(n13940), .ZN(n13942) );
  NOR2_X2 U15776 ( .A1(n15937), .A2(n15928), .ZN(n15929) );
  INV_X1 U15777 ( .A(n13869), .ZN(n13945) );
  INV_X1 U15778 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n13944) );
  NAND2_X1 U15779 ( .A1(n13945), .A2(n13944), .ZN(n13948) );
  NAND2_X1 U15780 ( .A1(n10981), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13946) );
  OAI211_X1 U15781 ( .C1(n14721), .C2(P1_EBX_REG_24__SCAN_IN), .A(n13881), .B(
        n13946), .ZN(n13947) );
  INV_X1 U15782 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n21561) );
  NAND2_X1 U15783 ( .A1(n13957), .A2(n21561), .ZN(n13952) );
  INV_X1 U15784 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16212) );
  NAND2_X1 U15785 ( .A1(n13881), .A2(n16212), .ZN(n13950) );
  NAND2_X1 U15786 ( .A1(n13864), .A2(n21561), .ZN(n13949) );
  NAND3_X1 U15787 ( .A1(n13950), .A2(n10981), .A3(n13949), .ZN(n13951) );
  NAND2_X1 U15788 ( .A1(n13952), .A2(n13951), .ZN(n15911) );
  MUX2_X1 U15789 ( .A(n13869), .B(n10981), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n13953) );
  OAI21_X1 U15790 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14704), .A(
        n13953), .ZN(n15860) );
  MUX2_X1 U15791 ( .A(n13869), .B(n10981), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13954) );
  OAI21_X1 U15792 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14704), .A(
        n13954), .ZN(n13955) );
  INV_X1 U15793 ( .A(n13955), .ZN(n15834) );
  INV_X1 U15794 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n13956) );
  NAND2_X1 U15795 ( .A1(n13957), .A2(n13956), .ZN(n13960) );
  NAND2_X1 U15796 ( .A1(n13881), .A2(n16194), .ZN(n13958) );
  OAI211_X1 U15797 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n14721), .A(n13958), .B(
        n10981), .ZN(n13959) );
  NAND2_X1 U15798 ( .A1(n13960), .A2(n13959), .ZN(n15848) );
  NAND2_X1 U15799 ( .A1(n15834), .A2(n15848), .ZN(n13961) );
  OR2_X1 U15800 ( .A1(n14704), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13963) );
  INV_X1 U15801 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15904) );
  NAND2_X1 U15802 ( .A1(n13864), .A2(n15904), .ZN(n13962) );
  NAND2_X1 U15803 ( .A1(n13963), .A2(n13962), .ZN(n15731) );
  OAI22_X1 U15804 ( .A1(n15731), .A2(n15733), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n13964), .ZN(n14007) );
  NAND2_X1 U15805 ( .A1(n15836), .A2(n14007), .ZN(n15734) );
  MUX2_X1 U15806 ( .A(n13966), .B(n13965), .S(n15734), .Z(n15902) );
  NAND2_X1 U15807 ( .A1(n10996), .A2(n13547), .ZN(n14692) );
  OAI21_X1 U15808 ( .B1(n13857), .B2(n13475), .A(n14692), .ZN(n13967) );
  NOR2_X1 U15809 ( .A1(n15902), .A2(n21338), .ZN(n14003) );
  INV_X1 U15810 ( .A(n16201), .ZN(n16085) );
  NAND2_X1 U15811 ( .A1(n13482), .A2(n21737), .ZN(n13969) );
  OAI211_X1 U15812 ( .C1(n13844), .C2(n13831), .A(n13969), .B(n14882), .ZN(
        n13970) );
  OAI21_X1 U15813 ( .B1(n13506), .B2(n13970), .A(n13491), .ZN(n13972) );
  NAND2_X1 U15814 ( .A1(n10997), .A2(n13860), .ZN(n13971) );
  OAI211_X1 U15815 ( .C1(n13973), .C2(n10981), .A(n13972), .B(n13971), .ZN(
        n13974) );
  INV_X1 U15816 ( .A(n13974), .ZN(n13976) );
  OAI21_X1 U15817 ( .B1(n14754), .B2(n13860), .A(n13977), .ZN(n13978) );
  OR2_X1 U15818 ( .A1(n14757), .A2(n13978), .ZN(n13979) );
  NAND2_X1 U15819 ( .A1(n13986), .A2(n13979), .ZN(n16312) );
  INV_X1 U15820 ( .A(n21285), .ZN(n21299) );
  AND2_X1 U15821 ( .A1(n13496), .A2(n13864), .ZN(n13980) );
  NAND2_X1 U15822 ( .A1(n14152), .A2(n13980), .ZN(n14766) );
  INV_X1 U15823 ( .A(n14766), .ZN(n14664) );
  NOR2_X1 U15824 ( .A1(n21289), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13990) );
  INV_X1 U15825 ( .A(n16241), .ZN(n16287) );
  AND2_X1 U15826 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16282) );
  NAND3_X1 U15827 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16287), .A3(
        n16282), .ZN(n13985) );
  NAND3_X1 U15828 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15560) );
  INV_X1 U15829 ( .A(n15560), .ZN(n15558) );
  NAND2_X1 U15830 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15558), .ZN(
        n16357) );
  NOR2_X1 U15831 ( .A1(n13981), .A2(n16357), .ZN(n16343) );
  NAND2_X1 U15832 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16343), .ZN(
        n16326) );
  NOR2_X1 U15833 ( .A1(n16133), .A2(n16326), .ZN(n21275) );
  NOR2_X1 U15834 ( .A1(n21311), .A2(n21317), .ZN(n21306) );
  INV_X1 U15835 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21283) );
  INV_X1 U15836 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21300) );
  OAI21_X1 U15837 ( .B1(n21283), .B2(n21300), .A(n21301), .ZN(n21304) );
  NAND2_X1 U15838 ( .A1(n21306), .A2(n21304), .ZN(n21327) );
  NOR2_X1 U15839 ( .A1(n13984), .A2(n21327), .ZN(n15538) );
  NAND2_X1 U15840 ( .A1(n21275), .A2(n15538), .ZN(n16262) );
  NOR2_X1 U15841 ( .A1(n13985), .A2(n16262), .ZN(n16237) );
  NAND3_X1 U15842 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n13982) );
  NOR2_X1 U15843 ( .A1(n13982), .A2(n16242), .ZN(n13983) );
  AND2_X1 U15844 ( .A1(n16237), .A2(n13983), .ZN(n13989) );
  NAND3_X1 U15845 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21306), .ZN(n15555) );
  NOR2_X1 U15846 ( .A1(n13984), .A2(n15555), .ZN(n15535) );
  NAND2_X1 U15847 ( .A1(n15535), .A2(n21275), .ZN(n16316) );
  OR2_X1 U15848 ( .A1(n16316), .A2(n13985), .ZN(n16235) );
  NOR2_X1 U15849 ( .A1(n16242), .A2(n16253), .ZN(n16245) );
  NAND2_X1 U15850 ( .A1(n16245), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13995) );
  NOR2_X1 U15851 ( .A1(n16235), .A2(n13995), .ZN(n13994) );
  OR2_X1 U15852 ( .A1(n21285), .A2(n13994), .ZN(n13988) );
  OR2_X1 U15853 ( .A1(n16312), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13987) );
  INV_X2 U15854 ( .A(n21288), .ZN(n21348) );
  OR2_X1 U15855 ( .A1(n13986), .A2(n21348), .ZN(n16366) );
  OAI211_X1 U15856 ( .C1(n13989), .C2(n21289), .A(n13988), .B(n21284), .ZN(
        n16219) );
  AOI211_X1 U15857 ( .C1(n16085), .C2(n21299), .A(n13990), .B(n16219), .ZN(
        n16213) );
  NAND3_X1 U15858 ( .A1(n16213), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16189) );
  NOR2_X1 U15859 ( .A1(n16189), .A2(n16181), .ZN(n14009) );
  NAND2_X1 U15860 ( .A1(n21285), .A2(n21289), .ZN(n16286) );
  NOR2_X1 U15861 ( .A1(n16328), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16171) );
  NOR2_X1 U15862 ( .A1(n16171), .A2(n16049), .ZN(n13992) );
  INV_X1 U15863 ( .A(n16213), .ZN(n13991) );
  NOR2_X1 U15864 ( .A1(n13991), .A2(n16286), .ZN(n16190) );
  INV_X1 U15865 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16378) );
  AOI211_X1 U15866 ( .C1(n14009), .C2(n13992), .A(n16190), .B(n16378), .ZN(
        n14002) );
  INV_X1 U15867 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n19947) );
  NOR2_X1 U15868 ( .A1(n21288), .A2(n19947), .ZN(n14537) );
  INV_X1 U15869 ( .A(n16365), .ZN(n13993) );
  NOR2_X1 U15870 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13993), .ZN(
        n14725) );
  NAND2_X1 U15871 ( .A1(n21302), .A2(n13994), .ZN(n16220) );
  INV_X1 U15872 ( .A(n13995), .ZN(n13996) );
  NAND3_X1 U15873 ( .A1(n21305), .A2(n13996), .A3(n16237), .ZN(n13997) );
  NAND2_X1 U15874 ( .A1(n16220), .A2(n13997), .ZN(n16231) );
  INV_X1 U15875 ( .A(n13998), .ZN(n13999) );
  NAND2_X1 U15876 ( .A1(n16231), .A2(n13999), .ZN(n16204) );
  NOR2_X1 U15877 ( .A1(n16204), .A2(n16202), .ZN(n16195) );
  NOR2_X1 U15878 ( .A1(n16181), .A2(n14000), .ZN(n16043) );
  NAND2_X1 U15879 ( .A1(n16195), .A2(n16043), .ZN(n16175) );
  NOR3_X1 U15880 ( .A1(n16175), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16049), .ZN(n14001) );
  NOR4_X1 U15881 ( .A1(n14003), .A2(n14002), .A3(n14537), .A4(n14001), .ZN(
        n14004) );
  OAI21_X1 U15882 ( .B1(n14541), .B2(n21339), .A(n14004), .ZN(P1_U3000) );
  XNOR2_X1 U15883 ( .A(n14005), .B(n11406), .ZN(n15653) );
  OAI21_X1 U15884 ( .B1(n15836), .B2(n14007), .A(n15734), .ZN(n15903) );
  INV_X1 U15885 ( .A(n15903), .ZN(n14008) );
  NAND2_X1 U15886 ( .A1(n14008), .A2(n21345), .ZN(n14013) );
  NOR2_X1 U15887 ( .A1(n14009), .A2(n16190), .ZN(n16172) );
  INV_X1 U15888 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n19943) );
  NOR2_X1 U15889 ( .A1(n21288), .A2(n19943), .ZN(n15649) );
  INV_X1 U15890 ( .A(n16195), .ZN(n14010) );
  NOR3_X1 U15891 ( .A1(n14010), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n16181), .ZN(n14011) );
  AOI211_X1 U15892 ( .C1(n16172), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15649), .B(n14011), .ZN(n14012) );
  OAI21_X1 U15893 ( .B1(n15653), .B2(n21339), .A(n14014), .ZN(P1_U3002) );
  NOR2_X2 U15894 ( .A1(n14882), .A2(n21917), .ZN(n14038) );
  INV_X1 U15895 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n14018) );
  NAND2_X1 U15896 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14047) );
  NAND2_X1 U15897 ( .A1(n14060), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14059) );
  INV_X1 U15898 ( .A(n14059), .ZN(n14068) );
  OAI21_X1 U15899 ( .B1(n14074), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n14097), .ZN(n21420) );
  AOI22_X1 U15900 ( .A1(n21420), .A2(n14497), .B1(n14501), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14017) );
  OAI21_X1 U15901 ( .B1(n14081), .B2(n14018), .A(n14017), .ZN(n14019) );
  NAND2_X1 U15902 ( .A1(n13468), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14052) );
  XNOR2_X1 U15903 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21361) );
  AOI21_X1 U15904 ( .B1(n14497), .B2(n21361), .A(n14501), .ZN(n14022) );
  NAND2_X1 U15905 ( .A1(n14502), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n14021) );
  OAI211_X1 U15906 ( .C1(n14052), .C2(n13370), .A(n14022), .B(n14021), .ZN(
        n14023) );
  INV_X1 U15907 ( .A(n14023), .ZN(n14024) );
  NAND2_X1 U15908 ( .A1(n14501), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14044) );
  INV_X1 U15909 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14026) );
  NOR2_X1 U15910 ( .A1(n14027), .A2(n14026), .ZN(n14029) );
  NOR2_X1 U15911 ( .A1(n14029), .A2(n14028), .ZN(n14030) );
  NAND2_X1 U15912 ( .A1(n21759), .A2(n14229), .ZN(n14034) );
  AOI22_X1 U15913 ( .A1(n14502), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21917), .ZN(n14032) );
  INV_X1 U15914 ( .A(n14052), .ZN(n14056) );
  NAND2_X1 U15915 ( .A1(n14056), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14031) );
  AND2_X1 U15916 ( .A1(n14032), .A2(n14031), .ZN(n14033) );
  NAND2_X1 U15917 ( .A1(n14035), .A2(n22167), .ZN(n14036) );
  NAND2_X1 U15918 ( .A1(n14036), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14710) );
  NAND2_X1 U15919 ( .A1(n14038), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n14040) );
  NAND2_X1 U15920 ( .A1(n21917), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14039) );
  OAI211_X1 U15921 ( .C1(n14052), .C2(n13797), .A(n14040), .B(n14039), .ZN(
        n14041) );
  AOI21_X1 U15922 ( .B1(n21772), .B2(n14229), .A(n14041), .ZN(n14042) );
  OR2_X1 U15923 ( .A1(n14710), .A2(n14042), .ZN(n14711) );
  INV_X1 U15924 ( .A(n14042), .ZN(n14712) );
  OR2_X1 U15925 ( .A1(n14712), .A2(n17185), .ZN(n14043) );
  NAND2_X1 U15926 ( .A1(n14711), .A2(n14043), .ZN(n14779) );
  INV_X1 U15927 ( .A(n21821), .ZN(n14046) );
  NAND2_X1 U15928 ( .A1(n14046), .A2(n14229), .ZN(n14055) );
  INV_X1 U15929 ( .A(n14047), .ZN(n14049) );
  INV_X1 U15930 ( .A(n14060), .ZN(n14048) );
  OAI21_X1 U15931 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n14049), .A(
        n14048), .ZN(n15259) );
  AOI22_X1 U15932 ( .A1(n14497), .A2(n15259), .B1(n14501), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14051) );
  NAND2_X1 U15933 ( .A1(n14038), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n14050) );
  OAI211_X1 U15934 ( .C1(n14052), .C2(n14776), .A(n14051), .B(n14050), .ZN(
        n14053) );
  INV_X1 U15935 ( .A(n14053), .ZN(n14054) );
  NAND2_X1 U15936 ( .A1(n15065), .A2(n15066), .ZN(n15103) );
  NAND2_X1 U15937 ( .A1(n14056), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14063) );
  INV_X1 U15938 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14057) );
  AOI21_X1 U15939 ( .B1(n14057), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14058) );
  AOI21_X1 U15940 ( .B1(n14038), .B2(P1_EAX_REG_4__SCAN_IN), .A(n14058), .ZN(
        n14062) );
  OAI21_X1 U15941 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n14060), .A(
        n14059), .ZN(n21382) );
  NOR2_X1 U15942 ( .A1(n21382), .A2(n17185), .ZN(n14061) );
  AOI21_X1 U15943 ( .B1(n14063), .B2(n14062), .A(n14061), .ZN(n14064) );
  AOI21_X1 U15944 ( .B1(n14065), .B2(n14229), .A(n14064), .ZN(n15102) );
  INV_X1 U15945 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n14070) );
  OAI21_X1 U15946 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n14068), .A(
        n14075), .ZN(n21396) );
  AOI22_X1 U15947 ( .A1(n14497), .A2(n21396), .B1(n14501), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n14069) );
  OAI21_X1 U15948 ( .B1(n14081), .B2(n14070), .A(n14069), .ZN(n14071) );
  INV_X1 U15949 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n14080) );
  NAND2_X1 U15950 ( .A1(n14073), .A2(n14229), .ZN(n14079) );
  INV_X1 U15951 ( .A(n14074), .ZN(n14077) );
  INV_X1 U15952 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21397) );
  NAND2_X1 U15953 ( .A1(n21397), .A2(n14075), .ZN(n14076) );
  NAND2_X1 U15954 ( .A1(n14077), .A2(n14076), .ZN(n21408) );
  AOI22_X1 U15955 ( .A1(n21408), .A2(n14497), .B1(n14501), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n14078) );
  OAI211_X1 U15956 ( .C1(n14081), .C2(n14080), .A(n14079), .B(n14078), .ZN(
        n15178) );
  NAND2_X1 U15957 ( .A1(n14083), .A2(n14082), .ZN(n15203) );
  XNOR2_X1 U15958 ( .A(n14097), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n21425) );
  INV_X1 U15959 ( .A(n14501), .ZN(n14203) );
  OAI22_X1 U15960 ( .A1(n21425), .A2(n17185), .B1(n14203), .B2(n15532), .ZN(
        n14084) );
  AOI21_X1 U15961 ( .B1(n14038), .B2(P1_EAX_REG_8__SCAN_IN), .A(n14084), .ZN(
        n14096) );
  AOI22_X1 U15962 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n14484), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14088) );
  AOI22_X1 U15963 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14087) );
  AOI22_X1 U15964 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n14770), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14086) );
  AOI22_X1 U15965 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14085) );
  NAND4_X1 U15966 ( .A1(n14088), .A2(n14087), .A3(n14086), .A4(n14085), .ZN(
        n14094) );
  AOI22_X1 U15967 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13529), .B1(
        n13534), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U15968 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n13513), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14091) );
  AOI22_X1 U15969 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14090) );
  AOI22_X1 U15970 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14089) );
  NAND4_X1 U15971 ( .A1(n14092), .A2(n14091), .A3(n14090), .A4(n14089), .ZN(
        n14093) );
  OAI21_X1 U15972 ( .B1(n14094), .B2(n14093), .A(n14229), .ZN(n14095) );
  NOR2_X2 U15973 ( .A1(n15203), .A2(n15348), .ZN(n15379) );
  XOR2_X1 U15974 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n14111), .Z(n15579) );
  AOI22_X1 U15975 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14101) );
  AOI22_X1 U15976 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14100) );
  AOI22_X1 U15977 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14099) );
  AOI22_X1 U15978 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14098) );
  NAND4_X1 U15979 ( .A1(n14101), .A2(n14100), .A3(n14099), .A4(n14098), .ZN(
        n14107) );
  AOI22_X1 U15980 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14770), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14105) );
  AOI22_X1 U15981 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U15982 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14103) );
  AOI22_X1 U15983 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14102) );
  NAND4_X1 U15984 ( .A1(n14105), .A2(n14104), .A3(n14103), .A4(n14102), .ZN(
        n14106) );
  OR2_X1 U15985 ( .A1(n14107), .A2(n14106), .ZN(n14108) );
  AOI22_X1 U15986 ( .A1(n14229), .A2(n14108), .B1(n14501), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14110) );
  NAND2_X1 U15987 ( .A1(n14038), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n14109) );
  OAI211_X1 U15988 ( .C1(n15579), .C2(n17185), .A(n14110), .B(n14109), .ZN(
        n15383) );
  NAND2_X1 U15989 ( .A1(n15379), .A2(n15383), .ZN(n15381) );
  XNOR2_X1 U15990 ( .A(n14128), .B(n21436), .ZN(n21439) );
  NAND2_X1 U15991 ( .A1(n21439), .A2(n14497), .ZN(n14126) );
  AOI22_X1 U15992 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14770), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14115) );
  AOI22_X1 U15993 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U15994 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14113) );
  AOI22_X1 U15995 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14112) );
  NAND4_X1 U15996 ( .A1(n14115), .A2(n14114), .A3(n14113), .A4(n14112), .ZN(
        n14121) );
  AOI22_X1 U15997 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14119) );
  AOI22_X1 U15998 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14118) );
  AOI22_X1 U15999 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14117) );
  AOI22_X1 U16000 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14116) );
  NAND4_X1 U16001 ( .A1(n14119), .A2(n14118), .A3(n14117), .A4(n14116), .ZN(
        n14120) );
  OAI21_X1 U16002 ( .B1(n14121), .B2(n14120), .A(n14229), .ZN(n14123) );
  NAND2_X1 U16003 ( .A1(n14038), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n14122) );
  OAI211_X1 U16004 ( .C1(n14203), .C2(n21436), .A(n14123), .B(n14122), .ZN(
        n14124) );
  INV_X1 U16005 ( .A(n14124), .ZN(n14125) );
  NAND2_X1 U16006 ( .A1(n14126), .A2(n14125), .ZN(n15458) );
  NAND2_X1 U16007 ( .A1(n14038), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n14131) );
  OAI21_X1 U16008 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n14129), .A(
        n14219), .ZN(n21448) );
  AOI22_X1 U16009 ( .A1(n14497), .A2(n21448), .B1(n14501), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n14130) );
  NAND2_X1 U16010 ( .A1(n14131), .A2(n14130), .ZN(n15509) );
  AOI22_X1 U16011 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13534), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14135) );
  AOI22_X1 U16012 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14134) );
  AOI22_X1 U16013 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14133) );
  AOI22_X1 U16014 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14132) );
  NAND4_X1 U16015 ( .A1(n14135), .A2(n14134), .A3(n14133), .A4(n14132), .ZN(
        n14141) );
  AOI22_X1 U16016 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14770), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14139) );
  AOI22_X1 U16017 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14138) );
  AOI22_X1 U16018 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14137) );
  AOI22_X1 U16019 ( .A1(n13560), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14136) );
  NAND4_X1 U16020 ( .A1(n14139), .A2(n14138), .A3(n14137), .A4(n14136), .ZN(
        n14140) );
  OR2_X1 U16021 ( .A1(n14141), .A2(n14140), .ZN(n14142) );
  NAND2_X1 U16022 ( .A1(n15457), .A2(n15511), .ZN(n14143) );
  XOR2_X1 U16023 ( .A(n15875), .B(n14237), .Z(n20032) );
  AOI22_X1 U16024 ( .A1(n14502), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n14501), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14156) );
  AOI22_X1 U16025 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13513), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U16026 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14146) );
  AOI22_X1 U16027 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14145) );
  AOI22_X1 U16028 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14144) );
  NAND4_X1 U16029 ( .A1(n14147), .A2(n14146), .A3(n14145), .A4(n14144), .ZN(
        n14154) );
  AOI22_X1 U16030 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14151) );
  AOI22_X1 U16031 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14150) );
  AOI22_X1 U16032 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14149) );
  AOI22_X1 U16033 ( .A1(n13560), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14148) );
  NAND4_X1 U16034 ( .A1(n14151), .A2(n14150), .A3(n14149), .A4(n14148), .ZN(
        n14153) );
  OAI21_X1 U16035 ( .B1(n14154), .B2(n14153), .A(n14493), .ZN(n14155) );
  OAI211_X1 U16036 ( .C1(n20032), .C2(n17185), .A(n14156), .B(n14155), .ZN(
        n14157) );
  INV_X1 U16037 ( .A(n14157), .ZN(n15871) );
  XNOR2_X1 U16038 ( .A(n14158), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16140) );
  NAND2_X1 U16039 ( .A1(n16140), .A2(n14497), .ZN(n14174) );
  AOI22_X1 U16040 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13534), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U16041 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14161) );
  AOI22_X1 U16042 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14160) );
  AOI22_X1 U16043 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14159) );
  NAND4_X1 U16044 ( .A1(n14162), .A2(n14161), .A3(n14160), .A4(n14159), .ZN(
        n14170) );
  AOI22_X1 U16045 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n13513), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14168) );
  AOI22_X1 U16046 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14167) );
  NAND2_X1 U16047 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n14164) );
  NAND2_X1 U16048 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14163) );
  AND3_X1 U16049 ( .A1(n14164), .A2(n14163), .A3(n17185), .ZN(n14166) );
  AOI22_X1 U16050 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14165) );
  NAND4_X1 U16051 ( .A1(n14168), .A2(n14167), .A3(n14166), .A4(n14165), .ZN(
        n14169) );
  NAND2_X1 U16052 ( .A1(n14472), .A2(n17185), .ZN(n14322) );
  OAI21_X1 U16053 ( .B1(n14170), .B2(n14169), .A(n14322), .ZN(n14172) );
  AOI22_X1 U16054 ( .A1(n14502), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21917), .ZN(n14171) );
  NAND2_X1 U16055 ( .A1(n14172), .A2(n14171), .ZN(n14173) );
  NAND2_X1 U16056 ( .A1(n14174), .A2(n14173), .ZN(n15882) );
  XOR2_X1 U16057 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n14175), .Z(
        n20029) );
  INV_X1 U16058 ( .A(n20029), .ZN(n21466) );
  AOI22_X1 U16059 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14179) );
  AOI22_X1 U16060 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14178) );
  AOI22_X1 U16061 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14177) );
  AOI22_X1 U16062 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14176) );
  NAND4_X1 U16063 ( .A1(n14179), .A2(n14178), .A3(n14177), .A4(n14176), .ZN(
        n14185) );
  AOI22_X1 U16064 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14183) );
  AOI22_X1 U16065 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14182) );
  AOI22_X1 U16066 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14181) );
  AOI22_X1 U16067 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14180) );
  NAND4_X1 U16068 ( .A1(n14183), .A2(n14182), .A3(n14181), .A4(n14180), .ZN(
        n14184) );
  OAI21_X1 U16069 ( .B1(n14185), .B2(n14184), .A(n14229), .ZN(n14188) );
  NAND2_X1 U16070 ( .A1(n14038), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n14187) );
  NAND2_X1 U16071 ( .A1(n14501), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14186) );
  NAND3_X1 U16072 ( .A1(n14188), .A2(n14187), .A3(n14186), .ZN(n14189) );
  AOI21_X1 U16073 ( .B1(n21466), .B2(n14497), .A(n14189), .ZN(n15971) );
  OR2_X1 U16074 ( .A1(n15882), .A2(n15971), .ZN(n15869) );
  XNOR2_X1 U16075 ( .A(n14190), .B(n15607), .ZN(n16153) );
  AOI22_X1 U16076 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14194) );
  AOI22_X1 U16077 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14193) );
  AOI22_X1 U16078 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14192) );
  AOI22_X1 U16079 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14191) );
  NAND4_X1 U16080 ( .A1(n14194), .A2(n14193), .A3(n14192), .A4(n14191), .ZN(
        n14200) );
  AOI22_X1 U16081 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13534), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14198) );
  AOI22_X1 U16082 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14197) );
  AOI22_X1 U16083 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14196) );
  AOI22_X1 U16084 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14195) );
  NAND4_X1 U16085 ( .A1(n14198), .A2(n14197), .A3(n14196), .A4(n14195), .ZN(
        n14199) );
  OAI21_X1 U16086 ( .B1(n14200), .B2(n14199), .A(n14229), .ZN(n14202) );
  NAND2_X1 U16087 ( .A1(n14038), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n14201) );
  OAI211_X1 U16088 ( .C1(n14203), .C2(n15607), .A(n14202), .B(n14201), .ZN(
        n14204) );
  AOI21_X1 U16089 ( .B1(n16153), .B2(n14497), .A(n14204), .ZN(n15600) );
  XOR2_X1 U16090 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n14206), .Z(
        n16168) );
  AOI22_X1 U16091 ( .A1(n14502), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n14501), 
        .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14218) );
  AOI22_X1 U16092 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14210) );
  AOI22_X1 U16093 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14209) );
  AOI22_X1 U16094 ( .A1(n11006), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14208) );
  AOI22_X1 U16095 ( .A1(n13560), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14207) );
  NAND4_X1 U16096 ( .A1(n14210), .A2(n14209), .A3(n14208), .A4(n14207), .ZN(
        n14216) );
  AOI22_X1 U16097 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14478), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14214) );
  AOI22_X1 U16098 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14213) );
  AOI22_X1 U16099 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14770), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14212) );
  AOI22_X1 U16100 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14211) );
  NAND4_X1 U16101 ( .A1(n14214), .A2(n14213), .A3(n14212), .A4(n14211), .ZN(
        n14215) );
  OAI21_X1 U16102 ( .B1(n14216), .B2(n14215), .A(n14229), .ZN(n14217) );
  OAI211_X1 U16103 ( .C1(n16168), .C2(n17185), .A(n14218), .B(n14217), .ZN(
        n15587) );
  XOR2_X1 U16104 ( .A(n14220), .B(n14219), .Z(n21461) );
  AOI22_X1 U16105 ( .A1(n14502), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n14501), 
        .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14233) );
  AOI22_X1 U16106 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14224) );
  AOI22_X1 U16107 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14223) );
  AOI22_X1 U16108 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14222) );
  AOI22_X1 U16109 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14221) );
  NAND4_X1 U16110 ( .A1(n14224), .A2(n14223), .A3(n14222), .A4(n14221), .ZN(
        n14231) );
  AOI22_X1 U16111 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14228) );
  AOI22_X1 U16112 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14227) );
  AOI22_X1 U16113 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14226) );
  AOI22_X1 U16114 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14225) );
  NAND4_X1 U16115 ( .A1(n14228), .A2(n14227), .A3(n14226), .A4(n14225), .ZN(
        n14230) );
  OAI21_X1 U16116 ( .B1(n14231), .B2(n14230), .A(n14229), .ZN(n14232) );
  OAI211_X1 U16117 ( .C1(n21461), .C2(n17185), .A(n14233), .B(n14232), .ZN(
        n15591) );
  AND2_X1 U16118 ( .A1(n15587), .A2(n15591), .ZN(n15585) );
  XNOR2_X1 U16119 ( .A(n14265), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n21482) );
  AOI21_X1 U16120 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n21478), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14238) );
  AOI21_X1 U16121 ( .B1(n14038), .B2(P1_EAX_REG_18__SCAN_IN), .A(n14238), .ZN(
        n14250) );
  AOI22_X1 U16122 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13534), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14242) );
  AOI22_X1 U16123 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14241) );
  AOI22_X1 U16124 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14240) );
  AOI22_X1 U16125 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14239) );
  NAND4_X1 U16126 ( .A1(n14242), .A2(n14241), .A3(n14240), .A4(n14239), .ZN(
        n14248) );
  AOI22_X1 U16127 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14246) );
  AOI22_X1 U16128 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14245) );
  AOI22_X1 U16129 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14244) );
  AOI22_X1 U16130 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14243) );
  NAND4_X1 U16131 ( .A1(n14246), .A2(n14245), .A3(n14244), .A4(n14243), .ZN(
        n14247) );
  OAI21_X1 U16132 ( .B1(n14248), .B2(n14247), .A(n14493), .ZN(n14249) );
  AOI22_X1 U16133 ( .A1(n21482), .A2(n14497), .B1(n14250), .B2(n14249), .ZN(
        n15614) );
  AOI22_X1 U16134 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14254) );
  AOI22_X1 U16135 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14253) );
  AOI22_X1 U16136 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14252) );
  AOI22_X1 U16137 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14251) );
  NAND4_X1 U16138 ( .A1(n14254), .A2(n14253), .A3(n14252), .A4(n14251), .ZN(
        n14260) );
  AOI22_X1 U16139 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14258) );
  AOI22_X1 U16140 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14257) );
  AOI22_X1 U16141 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14256) );
  AOI22_X1 U16142 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14255) );
  NAND4_X1 U16143 ( .A1(n14258), .A2(n14257), .A3(n14256), .A4(n14255), .ZN(
        n14259) );
  NOR2_X1 U16144 ( .A1(n14260), .A2(n14259), .ZN(n14264) );
  NAND2_X1 U16145 ( .A1(n21917), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14261) );
  NAND2_X1 U16146 ( .A1(n17185), .A2(n14261), .ZN(n14262) );
  AOI21_X1 U16147 ( .B1(n14038), .B2(P1_EAX_REG_19__SCAN_IN), .A(n14262), .ZN(
        n14263) );
  OAI21_X1 U16148 ( .B1(n14472), .B2(n14264), .A(n14263), .ZN(n14272) );
  INV_X1 U16149 ( .A(n14304), .ZN(n14270) );
  INV_X1 U16150 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14268) );
  INV_X1 U16151 ( .A(n14266), .ZN(n14267) );
  NAND2_X1 U16152 ( .A1(n14268), .A2(n14267), .ZN(n14269) );
  NAND2_X1 U16153 ( .A1(n14270), .A2(n14269), .ZN(n21491) );
  AOI22_X1 U16154 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14276) );
  AOI22_X1 U16155 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14770), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14275) );
  AOI22_X1 U16156 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14274) );
  AOI22_X1 U16157 ( .A1(n10976), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14273) );
  NAND4_X1 U16158 ( .A1(n14276), .A2(n14275), .A3(n14274), .A4(n14273), .ZN(
        n14284) );
  NAND2_X1 U16159 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n14278) );
  NAND2_X1 U16160 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14277) );
  AND3_X1 U16161 ( .A1(n14278), .A2(n14277), .A3(n17185), .ZN(n14282) );
  AOI22_X1 U16162 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14484), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14281) );
  AOI22_X1 U16163 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14478), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14280) );
  AOI22_X1 U16164 ( .A1(n11006), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14279) );
  NAND4_X1 U16165 ( .A1(n14282), .A2(n14281), .A3(n14280), .A4(n14279), .ZN(
        n14283) );
  OAI21_X1 U16166 ( .B1(n14284), .B2(n14283), .A(n14322), .ZN(n14286) );
  AOI22_X1 U16167 ( .A1(n14502), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n21917), .ZN(n14285) );
  NAND2_X1 U16168 ( .A1(n14286), .A2(n14285), .ZN(n14288) );
  INV_X1 U16169 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21509) );
  XNOR2_X1 U16170 ( .A(n14304), .B(n21509), .ZN(n21502) );
  NAND2_X1 U16171 ( .A1(n21502), .A2(n14497), .ZN(n14287) );
  NAND2_X1 U16172 ( .A1(n14288), .A2(n14287), .ZN(n15947) );
  AOI22_X1 U16173 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14294) );
  AOI22_X1 U16174 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14293) );
  AOI22_X1 U16175 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14292) );
  AOI22_X1 U16176 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14291) );
  NAND4_X1 U16177 ( .A1(n14294), .A2(n14293), .A3(n14292), .A4(n14291), .ZN(
        n14300) );
  AOI22_X1 U16178 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13513), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14298) );
  AOI22_X1 U16179 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14297) );
  AOI22_X1 U16180 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14296) );
  AOI22_X1 U16181 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14295) );
  NAND4_X1 U16182 ( .A1(n14298), .A2(n14297), .A3(n14296), .A4(n14295), .ZN(
        n14299) );
  NOR2_X1 U16183 ( .A1(n14300), .A2(n14299), .ZN(n14303) );
  OAI21_X1 U16184 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n16117), .A(n17185), 
        .ZN(n14301) );
  AOI21_X1 U16185 ( .B1(n14038), .B2(P1_EAX_REG_21__SCAN_IN), .A(n14301), .ZN(
        n14302) );
  OAI21_X1 U16186 ( .B1(n14472), .B2(n14303), .A(n14302), .ZN(n14308) );
  AND2_X1 U16187 ( .A1(n14305), .A2(n16117), .ZN(n14306) );
  NOR2_X1 U16188 ( .A1(n14350), .A2(n14306), .ZN(n21510) );
  NAND2_X1 U16189 ( .A1(n21510), .A2(n14497), .ZN(n14307) );
  NAND2_X1 U16190 ( .A1(n14308), .A2(n14307), .ZN(n15942) );
  NOR2_X2 U16191 ( .A1(n15941), .A2(n15942), .ZN(n15933) );
  NAND2_X1 U16192 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n14310) );
  NAND2_X1 U16193 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14309) );
  AND3_X1 U16194 ( .A1(n14310), .A2(n14309), .A3(n17185), .ZN(n14314) );
  AOI22_X1 U16195 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13534), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14313) );
  AOI22_X1 U16196 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14312) );
  AOI22_X1 U16197 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14311) );
  NAND4_X1 U16198 ( .A1(n14314), .A2(n14313), .A3(n14312), .A4(n14311), .ZN(
        n14320) );
  AOI22_X1 U16199 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U16200 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14317) );
  AOI22_X1 U16201 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14316) );
  AOI22_X1 U16202 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14315) );
  NAND4_X1 U16203 ( .A1(n14318), .A2(n14317), .A3(n14316), .A4(n14315), .ZN(
        n14319) );
  OR2_X1 U16204 ( .A1(n14320), .A2(n14319), .ZN(n14321) );
  NAND2_X1 U16205 ( .A1(n14322), .A2(n14321), .ZN(n14325) );
  AOI22_X1 U16206 ( .A1(n14502), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21917), .ZN(n14324) );
  INV_X1 U16207 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16109) );
  XNOR2_X1 U16208 ( .A(n14350), .B(n16109), .ZN(n21522) );
  AND2_X1 U16209 ( .A1(n21522), .A2(n14497), .ZN(n14323) );
  AOI21_X1 U16210 ( .B1(n14325), .B2(n14324), .A(n14323), .ZN(n15936) );
  AOI22_X1 U16211 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14329) );
  AOI22_X1 U16212 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n14484), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14328) );
  AOI22_X1 U16213 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14327) );
  AOI22_X1 U16214 ( .A1(n13560), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14326) );
  NAND4_X1 U16215 ( .A1(n14329), .A2(n14328), .A3(n14327), .A4(n14326), .ZN(
        n14335) );
  AOI22_X1 U16216 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n13513), .B1(
        n14770), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14333) );
  AOI22_X1 U16217 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14332) );
  AOI22_X1 U16218 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14331) );
  AOI22_X1 U16219 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n13534), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14330) );
  NAND4_X1 U16220 ( .A1(n14333), .A2(n14332), .A3(n14331), .A4(n14330), .ZN(
        n14334) );
  NOR2_X1 U16221 ( .A1(n14335), .A2(n14334), .ZN(n14357) );
  AOI22_X1 U16222 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13534), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14339) );
  AOI22_X1 U16223 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14338) );
  AOI22_X1 U16224 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14337) );
  AOI22_X1 U16225 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14336) );
  NAND4_X1 U16226 ( .A1(n14339), .A2(n14338), .A3(n14337), .A4(n14336), .ZN(
        n14345) );
  AOI22_X1 U16227 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14343) );
  AOI22_X1 U16228 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14342) );
  AOI22_X1 U16229 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14341) );
  AOI22_X1 U16230 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14340) );
  NAND4_X1 U16231 ( .A1(n14343), .A2(n14342), .A3(n14341), .A4(n14340), .ZN(
        n14344) );
  NOR2_X1 U16232 ( .A1(n14345), .A2(n14344), .ZN(n14356) );
  XNOR2_X1 U16233 ( .A(n14357), .B(n14356), .ZN(n14349) );
  NAND2_X1 U16234 ( .A1(n21917), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14346) );
  NAND2_X1 U16235 ( .A1(n17185), .A2(n14346), .ZN(n14347) );
  AOI21_X1 U16236 ( .B1(n14038), .B2(P1_EAX_REG_23__SCAN_IN), .A(n14347), .ZN(
        n14348) );
  OAI21_X1 U16237 ( .B1(n14472), .B2(n14349), .A(n14348), .ZN(n14355) );
  INV_X1 U16238 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14351) );
  NAND2_X1 U16239 ( .A1(n14352), .A2(n14351), .ZN(n14353) );
  NAND2_X1 U16240 ( .A1(n14374), .A2(n14353), .ZN(n21543) );
  NOR2_X1 U16241 ( .A1(n14357), .A2(n14356), .ZN(n14380) );
  AOI22_X1 U16242 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13513), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14361) );
  AOI22_X1 U16243 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14360) );
  AOI22_X1 U16244 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14359) );
  AOI22_X1 U16245 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14358) );
  NAND4_X1 U16246 ( .A1(n14361), .A2(n14360), .A3(n14359), .A4(n14358), .ZN(
        n14367) );
  AOI22_X1 U16247 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14365) );
  AOI22_X1 U16248 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14364) );
  AOI22_X1 U16249 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14363) );
  AOI22_X1 U16250 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14362) );
  NAND4_X1 U16251 ( .A1(n14365), .A2(n14364), .A3(n14363), .A4(n14362), .ZN(
        n14366) );
  OR2_X1 U16252 ( .A1(n14367), .A2(n14366), .ZN(n14379) );
  XNOR2_X1 U16253 ( .A(n14380), .B(n14379), .ZN(n14371) );
  NAND2_X1 U16254 ( .A1(n21917), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14368) );
  NAND2_X1 U16255 ( .A1(n17185), .A2(n14368), .ZN(n14369) );
  AOI21_X1 U16256 ( .B1(n14038), .B2(P1_EAX_REG_24__SCAN_IN), .A(n14369), .ZN(
        n14370) );
  OAI21_X1 U16257 ( .B1(n14371), .B2(n14472), .A(n14370), .ZN(n14373) );
  XNOR2_X1 U16258 ( .A(n14374), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n21544) );
  NAND2_X1 U16259 ( .A1(n21544), .A2(n14497), .ZN(n14372) );
  NAND2_X1 U16260 ( .A1(n14373), .A2(n14372), .ZN(n15917) );
  INV_X1 U16261 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14376) );
  NAND2_X1 U16262 ( .A1(n14377), .A2(n14376), .ZN(n14378) );
  NAND2_X1 U16263 ( .A1(n14415), .A2(n14378), .ZN(n21559) );
  NAND2_X1 U16264 ( .A1(n14380), .A2(n14379), .ZN(n14409) );
  AOI22_X1 U16265 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14384) );
  AOI22_X1 U16266 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14383) );
  AOI22_X1 U16267 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14770), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14382) );
  AOI22_X1 U16268 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14381) );
  NAND4_X1 U16269 ( .A1(n14384), .A2(n14383), .A3(n14382), .A4(n14381), .ZN(
        n14390) );
  AOI22_X1 U16270 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U16271 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14387) );
  AOI22_X1 U16272 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14386) );
  AOI22_X1 U16273 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14385) );
  NAND4_X1 U16274 ( .A1(n14388), .A2(n14387), .A3(n14386), .A4(n14385), .ZN(
        n14389) );
  NOR2_X1 U16275 ( .A1(n14390), .A2(n14389), .ZN(n14410) );
  XNOR2_X1 U16276 ( .A(n14409), .B(n14410), .ZN(n14393) );
  AOI21_X1 U16277 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n21917), .A(
        n14497), .ZN(n14392) );
  NAND2_X1 U16278 ( .A1(n14038), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n14391) );
  OAI211_X1 U16279 ( .C1(n14393), .C2(n14472), .A(n14392), .B(n14391), .ZN(
        n14394) );
  OAI21_X1 U16280 ( .B1(n17185), .B2(n21559), .A(n14394), .ZN(n15910) );
  INV_X1 U16281 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14395) );
  NOR2_X1 U16282 ( .A1(n14396), .A2(n14395), .ZN(n14400) );
  INV_X1 U16283 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14398) );
  OAI22_X1 U16284 ( .A1(n13520), .A2(n14398), .B1(n13522), .B2(n14397), .ZN(
        n14399) );
  AOI211_X1 U16285 ( .C1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .C2(n14478), .A(
        n14400), .B(n14399), .ZN(n14408) );
  AOI22_X1 U16286 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14484), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14404) );
  AOI22_X1 U16287 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14403) );
  AOI22_X1 U16288 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14402) );
  AOI22_X1 U16289 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14401) );
  AND4_X1 U16290 ( .A1(n14404), .A2(n14403), .A3(n14402), .A4(n14401), .ZN(
        n14407) );
  AOI22_X1 U16291 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14406) );
  AOI22_X1 U16292 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14405) );
  NAND4_X1 U16293 ( .A1(n14408), .A2(n14407), .A3(n14406), .A4(n14405), .ZN(
        n14430) );
  NOR2_X1 U16294 ( .A1(n14410), .A2(n14409), .ZN(n14431) );
  XOR2_X1 U16295 ( .A(n14430), .B(n14431), .Z(n14411) );
  NAND2_X1 U16296 ( .A1(n14411), .A2(n14493), .ZN(n14414) );
  INV_X1 U16297 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16077) );
  AOI21_X1 U16298 ( .B1(n16077), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n14412) );
  AOI21_X1 U16299 ( .B1(n14038), .B2(P1_EAX_REG_26__SCAN_IN), .A(n14412), .ZN(
        n14413) );
  XNOR2_X1 U16300 ( .A(n14415), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16079) );
  AOI22_X1 U16301 ( .A1(n14414), .A2(n14413), .B1(n14497), .B2(n16079), .ZN(
        n15856) );
  INV_X1 U16302 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15847) );
  NAND2_X1 U16303 ( .A1(n14417), .A2(n15847), .ZN(n14418) );
  NAND2_X1 U16304 ( .A1(n14453), .A2(n14418), .ZN(n16073) );
  AOI22_X1 U16305 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14419), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14423) );
  AOI22_X1 U16306 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14422) );
  AOI22_X1 U16307 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14421) );
  AOI22_X1 U16308 ( .A1(n13560), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14420) );
  NAND4_X1 U16309 ( .A1(n14423), .A2(n14422), .A3(n14421), .A4(n14420), .ZN(
        n14429) );
  AOI22_X1 U16310 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U16311 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14478), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14426) );
  AOI22_X1 U16312 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14461), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14425) );
  AOI22_X1 U16313 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14424) );
  NAND4_X1 U16314 ( .A1(n14427), .A2(n14426), .A3(n14425), .A4(n14424), .ZN(
        n14428) );
  NOR2_X1 U16315 ( .A1(n14429), .A2(n14428), .ZN(n14448) );
  NAND2_X1 U16316 ( .A1(n14431), .A2(n14430), .ZN(n14447) );
  XNOR2_X1 U16317 ( .A(n14448), .B(n14447), .ZN(n14434) );
  OAI21_X1 U16318 ( .B1(n21900), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n21917), .ZN(n14433) );
  NAND2_X1 U16319 ( .A1(n14502), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n14432) );
  OAI211_X1 U16320 ( .C1(n14434), .C2(n14472), .A(n14433), .B(n14432), .ZN(
        n14435) );
  OAI21_X1 U16321 ( .B1(n17185), .B2(n16073), .A(n14435), .ZN(n15846) );
  INV_X1 U16322 ( .A(n14453), .ZN(n14436) );
  XOR2_X1 U16323 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B(n14436), .Z(
        n16069) );
  AOI22_X1 U16324 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13513), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14440) );
  AOI22_X1 U16325 ( .A1(n13529), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14439) );
  AOI22_X1 U16326 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U16327 ( .A1(n14770), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14437) );
  NAND4_X1 U16328 ( .A1(n14440), .A2(n14439), .A3(n14438), .A4(n14437), .ZN(
        n14446) );
  AOI22_X1 U16329 ( .A1(n14478), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13444), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14444) );
  AOI22_X1 U16330 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14443) );
  AOI22_X1 U16331 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14442) );
  AOI22_X1 U16332 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14441) );
  NAND4_X1 U16333 ( .A1(n14444), .A2(n14443), .A3(n14442), .A4(n14441), .ZN(
        n14445) );
  OR2_X1 U16334 ( .A1(n14446), .A2(n14445), .ZN(n14468) );
  NOR2_X1 U16335 ( .A1(n14448), .A2(n14447), .ZN(n14469) );
  XOR2_X1 U16336 ( .A(n14468), .B(n14469), .Z(n14451) );
  INV_X1 U16337 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16065) );
  NAND2_X1 U16338 ( .A1(n14502), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n14449) );
  OAI211_X1 U16339 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n16065), .A(n14449), 
        .B(n17185), .ZN(n14450) );
  AOI21_X1 U16340 ( .B1(n14451), .B2(n14493), .A(n14450), .ZN(n14452) );
  AOI21_X1 U16341 ( .B1(n14497), .B2(n16069), .A(n14452), .ZN(n15833) );
  INV_X1 U16342 ( .A(n14454), .ZN(n14455) );
  INV_X1 U16343 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15824) );
  NAND2_X1 U16344 ( .A1(n14455), .A2(n15824), .ZN(n14456) );
  NAND2_X1 U16345 ( .A1(n14509), .A2(n14456), .ZN(n15823) );
  AOI22_X1 U16346 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14478), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14460) );
  AOI22_X1 U16347 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14459) );
  AOI22_X1 U16348 ( .A1(n14477), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14458) );
  AOI22_X1 U16349 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14457) );
  NAND4_X1 U16350 ( .A1(n14460), .A2(n14459), .A3(n14458), .A4(n14457), .ZN(
        n14467) );
  AOI22_X1 U16351 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14770), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14465) );
  AOI22_X1 U16352 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14464) );
  AOI22_X1 U16353 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11006), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14463) );
  AOI22_X1 U16354 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14462) );
  NAND4_X1 U16355 ( .A1(n14465), .A2(n14464), .A3(n14463), .A4(n14462), .ZN(
        n14466) );
  NOR2_X1 U16356 ( .A1(n14467), .A2(n14466), .ZN(n14476) );
  NAND2_X1 U16357 ( .A1(n14469), .A2(n14468), .ZN(n14475) );
  XNOR2_X1 U16358 ( .A(n14476), .B(n14475), .ZN(n14473) );
  AOI21_X1 U16359 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n21917), .A(
        n14497), .ZN(n14471) );
  NAND2_X1 U16360 ( .A1(n14502), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n14470) );
  OAI211_X1 U16361 ( .C1(n14473), .C2(n14472), .A(n14471), .B(n14470), .ZN(
        n14474) );
  OAI21_X1 U16362 ( .B1(n17185), .B2(n15823), .A(n14474), .ZN(n15648) );
  NOR2_X1 U16363 ( .A1(n14476), .A2(n14475), .ZN(n14492) );
  AOI22_X1 U16364 ( .A1(n13534), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14477), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14483) );
  AOI22_X1 U16365 ( .A1(n14479), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14478), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14482) );
  AOI22_X1 U16366 ( .A1(n11006), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10974), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14481) );
  AOI22_X1 U16367 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10976), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14480) );
  NAND4_X1 U16368 ( .A1(n14483), .A2(n14482), .A3(n14481), .A4(n14480), .ZN(
        n14490) );
  AOI22_X1 U16369 ( .A1(n14484), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13529), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14488) );
  AOI22_X1 U16370 ( .A1(n13513), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14770), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14487) );
  AOI22_X1 U16371 ( .A1(n13444), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13438), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14486) );
  AOI22_X1 U16372 ( .A1(n14461), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14485) );
  NAND4_X1 U16373 ( .A1(n14488), .A2(n14487), .A3(n14486), .A4(n14485), .ZN(
        n14489) );
  NOR2_X1 U16374 ( .A1(n14490), .A2(n14489), .ZN(n14491) );
  XNOR2_X1 U16375 ( .A(n14492), .B(n14491), .ZN(n14494) );
  NAND2_X1 U16376 ( .A1(n14494), .A2(n14493), .ZN(n14500) );
  NAND2_X1 U16377 ( .A1(n21917), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14495) );
  NAND2_X1 U16378 ( .A1(n17185), .A2(n14495), .ZN(n14496) );
  AOI21_X1 U16379 ( .B1(n14038), .B2(P1_EAX_REG_30__SCAN_IN), .A(n14496), .ZN(
        n14499) );
  XNOR2_X1 U16380 ( .A(n14509), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16051) );
  AND2_X1 U16381 ( .A1(n16051), .A2(n14497), .ZN(n14498) );
  AOI21_X1 U16382 ( .B1(n14500), .B2(n14499), .A(n14498), .ZN(n15730) );
  AOI22_X1 U16383 ( .A1(n14502), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n14501), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14503) );
  INV_X1 U16384 ( .A(n14503), .ZN(n14504) );
  INV_X1 U16385 ( .A(n15654), .ZN(n14531) );
  NAND2_X1 U16386 ( .A1(n14659), .A2(n14880), .ZN(n14627) );
  NAND2_X1 U16387 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n21586), .ZN(n17183) );
  NOR2_X1 U16388 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n16379), .ZN(n14506) );
  NOR2_X1 U16389 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21581) );
  NAND2_X1 U16390 ( .A1(n14506), .A2(n21581), .ZN(n14507) );
  OAI211_X1 U16391 ( .C1(n17183), .C2(n17186), .A(n21288), .B(n14507), .ZN(
        n14508) );
  INV_X1 U16392 ( .A(n14509), .ZN(n14510) );
  NAND2_X1 U16393 ( .A1(n14510), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14512) );
  INV_X1 U16394 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14511) );
  NAND2_X1 U16395 ( .A1(n13491), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14520) );
  AND2_X1 U16396 ( .A1(n21667), .A2(n21900), .ZN(n14515) );
  NOR2_X1 U16397 ( .A1(n14520), .A2(n14515), .ZN(n14516) );
  NOR2_X1 U16398 ( .A1(n14517), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14522) );
  NAND3_X1 U16399 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .ZN(n21377) );
  INV_X1 U16400 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21376) );
  NOR2_X1 U16401 ( .A1(n21377), .A2(n21376), .ZN(n21385) );
  NAND2_X1 U16402 ( .A1(n21385), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n21402) );
  INV_X1 U16403 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21401) );
  NOR2_X1 U16404 ( .A1(n21402), .A2(n21401), .ZN(n21409) );
  NAND3_X1 U16405 ( .A1(n21409), .A2(P1_REIP_REG_7__SCAN_IN), .A3(
        P1_REIP_REG_8__SCAN_IN), .ZN(n15742) );
  INV_X1 U16406 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21453) );
  NAND2_X1 U16407 ( .A1(n21460), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n15747) );
  INV_X1 U16408 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n19922) );
  NAND2_X1 U16409 ( .A1(n15605), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n21475) );
  INV_X1 U16410 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21474) );
  NOR2_X2 U16411 ( .A1(n21475), .A2(n21474), .ZN(n15879) );
  INV_X1 U16412 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n19927) );
  INV_X1 U16413 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21487) );
  INV_X1 U16414 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21527) );
  NOR2_X2 U16415 ( .A1(n21518), .A2(n21527), .ZN(n21525) );
  NAND2_X1 U16416 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n21525), .ZN(n21536) );
  INV_X1 U16417 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21535) );
  NOR2_X2 U16418 ( .A1(n21536), .A2(n21535), .ZN(n21556) );
  NAND2_X1 U16419 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14518) );
  NOR2_X2 U16420 ( .A1(n21565), .A2(n14518), .ZN(n15857) );
  INV_X1 U16421 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14519) );
  NAND3_X1 U16422 ( .A1(n14527), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n21567), 
        .ZN(n14526) );
  INV_X1 U16423 ( .A(n14520), .ZN(n14521) );
  NOR2_X1 U16424 ( .A1(n14522), .A2(n14521), .ZN(n14523) );
  AND2_X2 U16425 ( .A1(n14524), .A2(n14523), .ZN(n21551) );
  AOI22_X1 U16426 ( .A1(n21551), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n21564), .ZN(n14525) );
  OAI211_X1 U16427 ( .C1(n15902), .C2(n21572), .A(n14526), .B(n14525), .ZN(
        n14529) );
  NOR2_X1 U16428 ( .A1(n14527), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14528) );
  OAI21_X1 U16429 ( .B1(n14531), .B2(n21553), .A(n14530), .ZN(P1_U2809) );
  NAND3_X1 U16430 ( .A1(n17186), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n21579) );
  INV_X1 U16431 ( .A(n21579), .ZN(n14532) );
  NAND2_X1 U16432 ( .A1(n21923), .A2(n14533), .ZN(n21263) );
  NAND2_X1 U16433 ( .A1(n21263), .A2(n17186), .ZN(n14534) );
  NAND2_X1 U16434 ( .A1(n17186), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17180) );
  NAND2_X1 U16435 ( .A1(n21900), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14535) );
  AND2_X1 U16436 ( .A1(n17180), .A2(n14535), .ZN(n14730) );
  INV_X1 U16437 ( .A(n14730), .ZN(n14536) );
  AOI21_X1 U16438 ( .B1(n20038), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14537), .ZN(n14538) );
  OAI21_X1 U16439 ( .B1(n20043), .B2(n15250), .A(n14538), .ZN(n14539) );
  AOI21_X1 U16440 ( .B1(n15654), .B2(n21732), .A(n14539), .ZN(n14540) );
  OAI21_X1 U16441 ( .B1(n14541), .B2(n21574), .A(n14540), .ZN(P1_U2968) );
  NOR2_X1 U16442 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14543) );
  NOR4_X1 U16443 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14542) );
  NAND4_X1 U16444 ( .A1(n14543), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14542), .ZN(n14556) );
  NOR4_X1 U16445 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n14547) );
  NOR4_X1 U16446 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n14546) );
  NOR4_X1 U16447 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n14545) );
  NOR4_X1 U16448 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n14544) );
  AND4_X1 U16449 ( .A1(n14547), .A2(n14546), .A3(n14545), .A4(n14544), .ZN(
        n14552) );
  NOR4_X1 U16450 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n14550) );
  NOR4_X1 U16451 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n14549) );
  NOR4_X1 U16452 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n14548) );
  AND4_X1 U16453 ( .A1(n14550), .A2(n14549), .A3(n14548), .A4(n19909), .ZN(
        n14551) );
  NAND2_X1 U16454 ( .A1(n14552), .A2(n14551), .ZN(n14553) );
  INV_X1 U16455 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n17356) );
  INV_X1 U16456 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20100) );
  NOR4_X1 U16457 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n17356), .A4(n20100), .ZN(n14555) );
  NOR4_X1 U16458 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14554) );
  NAND3_X1 U16459 ( .A1(n21730), .A2(n14555), .A3(n14554), .ZN(U214) );
  INV_X1 U16460 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18357) );
  INV_X1 U16461 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17117) );
  NAND4_X1 U16462 ( .A1(n17883), .A2(n17117), .A3(n21602), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n21243) );
  NOR2_X2 U16463 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21246), .ZN(n21239) );
  NAND2_X1 U16464 ( .A1(n21202), .A2(n21239), .ZN(n21253) );
  NAND2_X1 U16465 ( .A1(n14558), .A2(n14557), .ZN(n20792) );
  NOR2_X1 U16466 ( .A1(n20595), .A2(n20101), .ZN(n20584) );
  INV_X1 U16467 ( .A(n20584), .ZN(n20197) );
  OAI22_X1 U16468 ( .A1(n18357), .A2(n20586), .B1(n20792), .B2(n20197), .ZN(
        n14566) );
  INV_X1 U16469 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17875) );
  AOI211_X1 U16470 ( .C1(n20106), .C2(n20105), .A(n21607), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n14561) );
  AOI211_X4 U16471 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n20596), .A(n14561), .B(
        n14562), .ZN(n20588) );
  INV_X1 U16472 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n20583) );
  INV_X1 U16473 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20549) );
  INV_X1 U16474 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20517) );
  NAND2_X1 U16475 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18034) );
  NAND2_X1 U16476 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17997) );
  NAND2_X1 U16477 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20378) );
  NAND2_X1 U16478 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20322) );
  NOR2_X1 U16479 ( .A1(n20322), .A2(n18135), .ZN(n20348) );
  NAND2_X1 U16480 ( .A1(n18241), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20196) );
  NAND3_X1 U16481 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20269) );
  NAND2_X1 U16482 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18108), .ZN(
        n14559) );
  INV_X1 U16483 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20229) );
  OAI21_X1 U16484 ( .B1(n20556), .B2(n20229), .A(n20561), .ZN(n20324) );
  OAI22_X1 U16485 ( .A1(n17875), .A2(n20516), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20324), .ZN(n14565) );
  NAND2_X1 U16486 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20596), .ZN(n14560) );
  AOI211_X4 U16487 ( .C1(n21652), .C2(n21602), .A(n14562), .B(n14560), .ZN(
        n20587) );
  INV_X1 U16488 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17505) );
  NAND2_X1 U16489 ( .A1(n17505), .A2(n17875), .ZN(n20176) );
  OAI21_X1 U16490 ( .B1(n17875), .B2(n17505), .A(n20176), .ZN(n17876) );
  INV_X1 U16491 ( .A(n14561), .ZN(n21237) );
  OAI22_X1 U16492 ( .A1(n20564), .A2(n17876), .B1(n20450), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n14564) );
  NAND2_X1 U16493 ( .A1(n20523), .A2(n20561), .ZN(n20571) );
  AOI221_X1 U16494 ( .B1(n20582), .B2(n20571), .C1(n20582), .C2(n20229), .A(
        n20169), .ZN(n14563) );
  OR4_X1 U16495 ( .A1(n14566), .A2(n14565), .A3(n14564), .A4(n14563), .ZN(
        P3_U2670) );
  INV_X1 U16496 ( .A(n12599), .ZN(n14567) );
  NAND2_X1 U16497 ( .A1(n14567), .A2(n14569), .ZN(n18400) );
  INV_X1 U16498 ( .A(n18400), .ZN(n14571) );
  INV_X1 U16499 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n14570) );
  OAI211_X1 U16500 ( .C1(n14571), .C2(n14570), .A(n17394), .B(n14574), .ZN(
        P2_U2814) );
  NOR2_X1 U16501 ( .A1(n18371), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n14573)
         );
  AOI22_X1 U16502 ( .A1(n14573), .A2(n17394), .B1(n14572), .B2(n18371), .ZN(
        P2_U3612) );
  INV_X1 U16503 ( .A(n18716), .ZN(n21624) );
  INV_X1 U16504 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n14576) );
  NAND3_X1 U16505 ( .A1(n15298), .A2(n12651), .A3(n18716), .ZN(n14625) );
  AOI22_X1 U16506 ( .A1(n15130), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n15131), .ZN(n19701) );
  NOR2_X1 U16507 ( .A1(n14625), .A2(n19701), .ZN(n14581) );
  AOI21_X1 U16508 ( .B1(n14622), .B2(P2_EAX_REG_16__SCAN_IN), .A(n14581), .ZN(
        n14575) );
  OAI21_X1 U16509 ( .B1(n14630), .B2(n14576), .A(n14575), .ZN(P2_U2952) );
  INV_X1 U16510 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n14578) );
  AOI22_X1 U16511 ( .A1(n15130), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14617), .ZN(n19584) );
  NOR2_X1 U16512 ( .A1(n14625), .A2(n19584), .ZN(n14586) );
  AOI21_X1 U16513 ( .B1(n14622), .B2(P2_EAX_REG_18__SCAN_IN), .A(n14586), .ZN(
        n14577) );
  OAI21_X1 U16514 ( .B1(n14630), .B2(n14578), .A(n14577), .ZN(P2_U2954) );
  INV_X1 U16515 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n14580) );
  AOI22_X1 U16516 ( .A1(n15130), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14617), .ZN(n19538) );
  NOR2_X1 U16517 ( .A1(n14625), .A2(n19538), .ZN(n14596) );
  AOI21_X1 U16518 ( .B1(n14622), .B2(P2_EAX_REG_3__SCAN_IN), .A(n14596), .ZN(
        n14579) );
  OAI21_X1 U16519 ( .B1(n14630), .B2(n14580), .A(n14579), .ZN(P2_U2970) );
  INV_X1 U16520 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n14583) );
  AOI21_X1 U16521 ( .B1(n14622), .B2(P2_EAX_REG_0__SCAN_IN), .A(n14581), .ZN(
        n14582) );
  OAI21_X1 U16522 ( .B1(n14630), .B2(n14583), .A(n14582), .ZN(P2_U2967) );
  INV_X1 U16523 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n14585) );
  AOI22_X1 U16524 ( .A1(n15130), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14617), .ZN(n19218) );
  NOR2_X1 U16525 ( .A1(n14625), .A2(n19218), .ZN(n14589) );
  AOI21_X1 U16526 ( .B1(n14622), .B2(P2_EAX_REG_7__SCAN_IN), .A(n14589), .ZN(
        n14584) );
  OAI21_X1 U16527 ( .B1(n14630), .B2(n14585), .A(n14584), .ZN(P2_U2974) );
  INV_X1 U16528 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n14588) );
  AOI21_X1 U16529 ( .B1(n14622), .B2(P2_EAX_REG_2__SCAN_IN), .A(n14586), .ZN(
        n14587) );
  OAI21_X1 U16530 ( .B1(n14630), .B2(n14588), .A(n14587), .ZN(P2_U2969) );
  INV_X1 U16531 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n14591) );
  AOI21_X1 U16532 ( .B1(n14622), .B2(P2_EAX_REG_23__SCAN_IN), .A(n14589), .ZN(
        n14590) );
  OAI21_X1 U16533 ( .B1(n14630), .B2(n14591), .A(n14590), .ZN(P2_U2959) );
  INV_X1 U16534 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n14593) );
  AOI22_X1 U16535 ( .A1(n15130), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14617), .ZN(n19436) );
  NOR2_X1 U16536 ( .A1(n14625), .A2(n19436), .ZN(n14602) );
  AOI21_X1 U16537 ( .B1(n14622), .B2(P2_EAX_REG_5__SCAN_IN), .A(n14602), .ZN(
        n14592) );
  OAI21_X1 U16538 ( .B1(n14630), .B2(n14593), .A(n14592), .ZN(P2_U2972) );
  INV_X1 U16539 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n14595) );
  AOI22_X1 U16540 ( .A1(n15130), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14617), .ZN(n19640) );
  NOR2_X1 U16541 ( .A1(n14625), .A2(n19640), .ZN(n14599) );
  AOI21_X1 U16542 ( .B1(n14622), .B2(P2_EAX_REG_17__SCAN_IN), .A(n14599), .ZN(
        n14594) );
  OAI21_X1 U16543 ( .B1(n14630), .B2(n14595), .A(n14594), .ZN(P2_U2953) );
  INV_X1 U16544 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n14598) );
  AOI21_X1 U16545 ( .B1(n14622), .B2(P2_EAX_REG_19__SCAN_IN), .A(n14596), .ZN(
        n14597) );
  OAI21_X1 U16546 ( .B1(n14630), .B2(n14598), .A(n14597), .ZN(P2_U2955) );
  INV_X1 U16547 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n14601) );
  AOI21_X1 U16548 ( .B1(n14622), .B2(P2_EAX_REG_1__SCAN_IN), .A(n14599), .ZN(
        n14600) );
  OAI21_X1 U16549 ( .B1(n14630), .B2(n14601), .A(n14600), .ZN(P2_U2968) );
  INV_X1 U16550 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n14604) );
  AOI21_X1 U16551 ( .B1(n14622), .B2(P2_EAX_REG_21__SCAN_IN), .A(n14602), .ZN(
        n14603) );
  OAI21_X1 U16552 ( .B1(n14630), .B2(n14604), .A(n14603), .ZN(P2_U2957) );
  INV_X1 U16553 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n14606) );
  INV_X1 U16554 ( .A(n14625), .ZN(n14645) );
  AOI22_X1 U16555 ( .A1(n15130), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14617), .ZN(n19374) );
  INV_X1 U16556 ( .A(n19374), .ZN(n16573) );
  NAND2_X1 U16557 ( .A1(n14645), .A2(n16573), .ZN(n14643) );
  NAND2_X1 U16558 ( .A1(n14622), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n14605) );
  OAI211_X1 U16559 ( .C1(n14630), .C2(n14606), .A(n14643), .B(n14605), .ZN(
        P2_U2973) );
  INV_X1 U16560 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n14610) );
  INV_X1 U16561 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n14607) );
  NOR2_X1 U16562 ( .A1(n15130), .A2(n14607), .ZN(n14608) );
  AOI21_X1 U16563 ( .B1(BUF1_REG_10__SCAN_IN), .B2(n15130), .A(n14608), .ZN(
        n19209) );
  INV_X1 U16564 ( .A(n19209), .ZN(n16541) );
  NAND2_X1 U16565 ( .A1(n14645), .A2(n16541), .ZN(n14638) );
  NAND2_X1 U16566 ( .A1(n14622), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n14609) );
  OAI211_X1 U16567 ( .C1(n14630), .C2(n14610), .A(n14638), .B(n14609), .ZN(
        P2_U2977) );
  INV_X1 U16568 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n14613) );
  AOI22_X1 U16569 ( .A1(n15130), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n14617), .ZN(n19194) );
  INV_X1 U16570 ( .A(n19194), .ZN(n14611) );
  NAND2_X1 U16571 ( .A1(n14645), .A2(n14611), .ZN(n14653) );
  NAND2_X1 U16572 ( .A1(n14622), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n14612) );
  OAI211_X1 U16573 ( .C1(n14630), .C2(n14613), .A(n14653), .B(n14612), .ZN(
        P2_U2981) );
  INV_X1 U16574 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n14616) );
  INV_X1 U16575 ( .A(n19199), .ZN(n14614) );
  NAND2_X1 U16576 ( .A1(n14645), .A2(n14614), .ZN(n14631) );
  NAND2_X1 U16577 ( .A1(n14622), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n14615) );
  OAI211_X1 U16578 ( .C1(n14630), .C2(n14616), .A(n14631), .B(n14615), .ZN(
        P2_U2980) );
  INV_X1 U16579 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n14620) );
  AOI22_X1 U16580 ( .A1(n15130), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n14617), .ZN(n19215) );
  INV_X1 U16581 ( .A(n19215), .ZN(n14618) );
  NAND2_X1 U16582 ( .A1(n14645), .A2(n14618), .ZN(n14633) );
  NAND2_X1 U16583 ( .A1(n14622), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n14619) );
  OAI211_X1 U16584 ( .C1(n14630), .C2(n14620), .A(n14633), .B(n14619), .ZN(
        P2_U2975) );
  INV_X1 U16585 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n14624) );
  NOR2_X1 U16586 ( .A1(n15130), .A2(n20608), .ZN(n14621) );
  AOI21_X1 U16587 ( .B1(BUF1_REG_12__SCAN_IN), .B2(n15130), .A(n14621), .ZN(
        n19200) );
  INV_X1 U16588 ( .A(n19200), .ZN(n16527) );
  NAND2_X1 U16589 ( .A1(n14645), .A2(n16527), .ZN(n14651) );
  NAND2_X1 U16590 ( .A1(n14622), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n14623) );
  OAI211_X1 U16591 ( .C1(n14630), .C2(n14624), .A(n14651), .B(n14623), .ZN(
        P2_U2979) );
  INV_X1 U16592 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14626) );
  AOI22_X1 U16593 ( .A1(n15130), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15131), .ZN(n19193) );
  INV_X1 U16594 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n17476) );
  OAI222_X1 U16595 ( .A1(n14630), .A2(n14626), .B1(n14625), .B2(n19193), .C1(
        n14714), .C2(n17476), .ZN(P2_U2982) );
  INV_X1 U16596 ( .A(n14627), .ZN(n14629) );
  INV_X1 U16597 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14628) );
  AND2_X1 U16598 ( .A1(n21896), .A2(n16379), .ZN(n15391) );
  INV_X1 U16599 ( .A(n15391), .ZN(n15813) );
  OAI211_X1 U16600 ( .C1(n14629), .C2(n14628), .A(n15813), .B(n21665), .ZN(
        P1_U2801) );
  NAND2_X1 U16601 ( .A1(n14655), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14632) );
  OAI211_X1 U16602 ( .C1(n14714), .C2(n14859), .A(n14632), .B(n14631), .ZN(
        P2_U2965) );
  INV_X1 U16603 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n16557) );
  NAND2_X1 U16604 ( .A1(n14655), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n14634) );
  OAI211_X1 U16605 ( .C1(n14714), .C2(n16557), .A(n14634), .B(n14633), .ZN(
        P2_U2960) );
  INV_X1 U16606 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19206) );
  NAND2_X1 U16607 ( .A1(n14655), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n14637) );
  NAND2_X1 U16608 ( .A1(n15131), .A2(BUF2_REG_11__SCAN_IN), .ZN(n14636) );
  INV_X1 U16609 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20071) );
  OR2_X1 U16610 ( .A1(n15131), .A2(n20071), .ZN(n14635) );
  NAND2_X1 U16611 ( .A1(n14636), .A2(n14635), .ZN(n19203) );
  NAND2_X1 U16612 ( .A1(n14645), .A2(n19203), .ZN(n14649) );
  OAI211_X1 U16613 ( .C1(n19206), .C2(n14714), .A(n14637), .B(n14649), .ZN(
        P2_U2978) );
  INV_X1 U16614 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n16539) );
  NAND2_X1 U16615 ( .A1(n14655), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14639) );
  OAI211_X1 U16616 ( .C1(n14714), .C2(n16539), .A(n14639), .B(n14638), .ZN(
        P2_U2962) );
  INV_X1 U16617 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19214) );
  NAND2_X1 U16618 ( .A1(n14655), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n14642) );
  NAND2_X1 U16619 ( .A1(n15131), .A2(BUF2_REG_9__SCAN_IN), .ZN(n14641) );
  INV_X1 U16620 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20067) );
  OR2_X1 U16621 ( .A1(n15131), .A2(n20067), .ZN(n14640) );
  NAND2_X1 U16622 ( .A1(n14641), .A2(n14640), .ZN(n19211) );
  NAND2_X1 U16623 ( .A1(n14645), .A2(n19211), .ZN(n14656) );
  OAI211_X1 U16624 ( .C1(n19214), .C2(n14714), .A(n14642), .B(n14656), .ZN(
        P2_U2976) );
  INV_X1 U16625 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n16571) );
  NAND2_X1 U16626 ( .A1(n14655), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n14644) );
  OAI211_X1 U16627 ( .C1(n14714), .C2(n16571), .A(n14644), .B(n14643), .ZN(
        P2_U2958) );
  INV_X1 U16628 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19480) );
  NAND2_X1 U16629 ( .A1(n14655), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n14646) );
  AOI22_X1 U16630 ( .A1(n15130), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14617), .ZN(n19488) );
  INV_X1 U16631 ( .A(n19488), .ZN(n15499) );
  NAND2_X1 U16632 ( .A1(n14645), .A2(n15499), .ZN(n14647) );
  OAI211_X1 U16633 ( .C1(n19480), .C2(n14714), .A(n14646), .B(n14647), .ZN(
        P2_U2971) );
  INV_X1 U16634 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n15497) );
  NAND2_X1 U16635 ( .A1(n14655), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n14648) );
  OAI211_X1 U16636 ( .C1(n14714), .C2(n15497), .A(n14648), .B(n14647), .ZN(
        P2_U2956) );
  INV_X1 U16637 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14855) );
  NAND2_X1 U16638 ( .A1(n14655), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14650) );
  OAI211_X1 U16639 ( .C1(n14855), .C2(n14714), .A(n14650), .B(n14649), .ZN(
        P2_U2963) );
  INV_X1 U16640 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n16525) );
  NAND2_X1 U16641 ( .A1(n14655), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14652) );
  OAI211_X1 U16642 ( .C1(n14714), .C2(n16525), .A(n14652), .B(n14651), .ZN(
        P2_U2964) );
  INV_X1 U16643 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n15804) );
  NAND2_X1 U16644 ( .A1(n14655), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14654) );
  OAI211_X1 U16645 ( .C1(n14714), .C2(n15804), .A(n14654), .B(n14653), .ZN(
        P2_U2966) );
  INV_X1 U16646 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14852) );
  NAND2_X1 U16647 ( .A1(n14655), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14657) );
  OAI211_X1 U16648 ( .C1(n14852), .C2(n14714), .A(n14657), .B(n14656), .ZN(
        P2_U2961) );
  OAI22_X1 U16649 ( .A1(n14659), .A2(n14658), .B1(n11315), .B2(n13843), .ZN(
        n20044) );
  NAND3_X1 U16650 ( .A1(n14721), .A2(n15814), .A3(n21617), .ZN(n21266) );
  AND2_X1 U16651 ( .A1(n21266), .A2(n21667), .ZN(n14660) );
  NOR2_X1 U16652 ( .A1(n20044), .A2(n14660), .ZN(n17167) );
  OR2_X1 U16653 ( .A1(n17167), .A2(n21592), .ZN(n14669) );
  INV_X1 U16654 ( .A(n14669), .ZN(n21576) );
  INV_X1 U16655 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n14671) );
  NAND3_X1 U16656 ( .A1(n14661), .A2(n13496), .A3(n13860), .ZN(n14662) );
  NAND2_X1 U16657 ( .A1(n14663), .A2(n14662), .ZN(n14665) );
  MUX2_X1 U16658 ( .A(n14665), .B(n14664), .S(n13843), .Z(n14668) );
  NOR2_X1 U16659 ( .A1(n14738), .A2(n14666), .ZN(n14667) );
  OAI21_X1 U16660 ( .B1(n14668), .B2(n14667), .A(n14882), .ZN(n17171) );
  OR2_X1 U16661 ( .A1(n14669), .A2(n17171), .ZN(n14670) );
  OAI21_X1 U16662 ( .B1(n21576), .B2(n14671), .A(n14670), .ZN(P1_U3484) );
  INV_X1 U16663 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18667) );
  NAND2_X1 U16664 ( .A1(n18390), .A2(n18667), .ZN(n14672) );
  NAND2_X1 U16665 ( .A1(n14673), .A2(n14672), .ZN(n18663) );
  INV_X1 U16666 ( .A(n18663), .ZN(n14677) );
  OAI21_X1 U16667 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14675), .A(
        n14674), .ZN(n18674) );
  NAND2_X1 U16668 ( .A1(n18500), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n18672) );
  OAI21_X1 U16669 ( .B1(n17408), .B2(n18674), .A(n18672), .ZN(n14676) );
  AOI21_X1 U16670 ( .B1(n12546), .B2(n14677), .A(n14676), .ZN(n14680) );
  OAI21_X1 U16671 ( .B1(n16750), .B2(n14678), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14679) );
  OAI211_X1 U16672 ( .C1(n17410), .C2(n12950), .A(n14680), .B(n14679), .ZN(
        P2_U3014) );
  INV_X1 U16673 ( .A(n14681), .ZN(n14691) );
  NOR2_X1 U16674 ( .A1(n14683), .A2(n14682), .ZN(n14684) );
  XOR2_X1 U16675 ( .A(n14684), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n17050) );
  AOI21_X1 U16676 ( .B1(n15284), .B2(n14686), .A(n14685), .ZN(n17051) );
  INV_X1 U16677 ( .A(n17051), .ZN(n14688) );
  MUX2_X1 U16678 ( .A(n16782), .B(n17417), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14687) );
  NAND2_X1 U16679 ( .A1(n18500), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n17048) );
  OAI211_X1 U16680 ( .C1(n17408), .C2(n14688), .A(n14687), .B(n17048), .ZN(
        n14689) );
  AOI21_X1 U16681 ( .B1(n12546), .B2(n17050), .A(n14689), .ZN(n14690) );
  OAI21_X1 U16682 ( .B1(n14691), .B2(n17410), .A(n14690), .ZN(P2_U3013) );
  INV_X1 U16683 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14698) );
  INV_X1 U16684 ( .A(n14692), .ZN(n14693) );
  NAND2_X1 U16685 ( .A1(n17152), .A2(n11017), .ZN(n14694) );
  NAND2_X1 U16686 ( .A1(n21720), .A2(n14694), .ZN(n14696) );
  NAND2_X1 U16687 ( .A1(n19882), .A2(n13860), .ZN(n14803) );
  NOR2_X1 U16688 ( .A1(n21917), .A2(n16379), .ZN(n14924) );
  INV_X1 U16689 ( .A(n14924), .ZN(n15035) );
  AOI22_X1 U16690 ( .A1(n19897), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19894), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14697) );
  OAI21_X1 U16691 ( .B1(n14698), .B2(n14803), .A(n14697), .ZN(P1_U2913) );
  AOI22_X1 U16692 ( .A1(n21264), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n19894), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14699) );
  OAI21_X1 U16693 ( .B1(n16008), .B2(n14803), .A(n14699), .ZN(P1_U2914) );
  INV_X1 U16694 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14701) );
  AOI22_X1 U16695 ( .A1(n21264), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n19894), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14700) );
  OAI21_X1 U16696 ( .B1(n14701), .B2(n14803), .A(n14700), .ZN(P1_U2915) );
  INV_X1 U16697 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21691) );
  AOI22_X1 U16698 ( .A1(n21264), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19894), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14702) );
  OAI21_X1 U16699 ( .B1(n21691), .B2(n14803), .A(n14702), .ZN(P1_U2911) );
  INV_X1 U16700 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n21686) );
  AOI22_X1 U16701 ( .A1(n21264), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n19894), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14703) );
  OAI21_X1 U16702 ( .B1(n21686), .B2(n14803), .A(n14703), .ZN(P1_U2912) );
  NOR2_X1 U16703 ( .A1(n14704), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14706) );
  OR2_X1 U16704 ( .A1(n14706), .A2(n14705), .ZN(n15895) );
  NAND4_X1 U16705 ( .A1(n14707), .A2(n14708), .A3(n13429), .A4(n13831), .ZN(
        n14877) );
  OAI22_X1 U16706 ( .A1(n13843), .A2(n14766), .B1(n14877), .B2(n14721), .ZN(
        n14709) );
  INV_X1 U16707 ( .A(n14710), .ZN(n14713) );
  OAI21_X1 U16708 ( .B1(n14713), .B2(n14712), .A(n14711), .ZN(n15892) );
  OAI222_X1 U16709 ( .A1(n15895), .A2(n19979), .B1(n13868), .B2(n19989), .C1(
        n15892), .C2(n15965), .ZN(P1_U2872) );
  INV_X1 U16710 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n15404) );
  OR2_X1 U16711 ( .A1(n12599), .A2(n18718), .ZN(n14715) );
  OAI21_X1 U16712 ( .B1(n14949), .B2(n14715), .A(n14714), .ZN(n14716) );
  INV_X1 U16713 ( .A(n18377), .ZN(n14717) );
  NOR2_X1 U16714 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17419), .ZN(n17465) );
  NOR2_X4 U16715 ( .A1(n17448), .A2(n17473), .ZN(n17464) );
  AOI22_X1 U16716 ( .A1(n17465), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14718) );
  OAI21_X1 U16717 ( .B1(n15404), .B2(n14862), .A(n14718), .ZN(P2_U2933) );
  INV_X1 U16718 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n15199) );
  AOI22_X1 U16719 ( .A1(n17465), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14719) );
  OAI21_X1 U16720 ( .B1(n15199), .B2(n14862), .A(n14719), .ZN(P2_U2934) );
  XNOR2_X1 U16721 ( .A(n14720), .B(n14721), .ZN(n14781) );
  OR2_X1 U16722 ( .A1(n14722), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14785) );
  NAND3_X1 U16723 ( .A1(n14785), .A2(n14723), .A3(n21346), .ZN(n14729) );
  INV_X1 U16724 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n15268) );
  NOR2_X1 U16725 ( .A1(n21288), .A2(n15268), .ZN(n14784) );
  NAND2_X1 U16726 ( .A1(n21289), .A2(n16312), .ZN(n14724) );
  NAND2_X1 U16727 ( .A1(n14724), .A2(n21283), .ZN(n16369) );
  AOI21_X1 U16728 ( .B1(n16366), .B2(n16369), .A(n21300), .ZN(n14727) );
  NOR3_X1 U16729 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16328), .A3(
        n14725), .ZN(n14726) );
  NOR3_X1 U16730 ( .A1(n14784), .A2(n14727), .A3(n14726), .ZN(n14728) );
  OAI211_X1 U16731 ( .C1(n21338), .C2(n14781), .A(n14729), .B(n14728), .ZN(
        P1_U3030) );
  NAND2_X1 U16732 ( .A1(n14730), .A2(n16164), .ZN(n14735) );
  INV_X1 U16733 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14731) );
  NOR2_X1 U16734 ( .A1(n21288), .A2(n14731), .ZN(n16363) );
  OAI21_X1 U16735 ( .B1(n14732), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11005), .ZN(n16362) );
  NOR2_X1 U16736 ( .A1(n16362), .A2(n21574), .ZN(n14734) );
  AOI211_X1 U16737 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n14735), .A(
        n16363), .B(n14734), .ZN(n14736) );
  OAI21_X1 U16738 ( .B1(n20022), .B2(n15892), .A(n14736), .ZN(P1_U2999) );
  NOR2_X1 U16739 ( .A1(n17186), .A2(n15035), .ZN(n21582) );
  INV_X1 U16740 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21881) );
  NOR2_X1 U16741 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21881), .ZN(n21736) );
  INV_X1 U16742 ( .A(n21667), .ZN(n21616) );
  NOR2_X1 U16743 ( .A1(n21617), .A2(n21616), .ZN(n17178) );
  OAI21_X1 U16744 ( .B1(n17152), .B2(n10996), .A(n17178), .ZN(n14737) );
  MUX2_X1 U16745 ( .A(n14766), .B(n14737), .S(n13843), .Z(n14746) );
  INV_X1 U16746 ( .A(n13855), .ZN(n14750) );
  NAND3_X1 U16747 ( .A1(n14750), .A2(n14738), .A3(n21667), .ZN(n14741) );
  NAND2_X1 U16748 ( .A1(n21663), .A2(n14767), .ZN(n14739) );
  NAND2_X1 U16749 ( .A1(n14739), .A2(n13843), .ZN(n14740) );
  NAND2_X1 U16750 ( .A1(n14741), .A2(n14740), .ZN(n14879) );
  NAND3_X1 U16751 ( .A1(n13844), .A2(n21737), .A3(n13491), .ZN(n14742) );
  NAND2_X1 U16752 ( .A1(n14743), .A2(n14742), .ZN(n14744) );
  NOR2_X1 U16753 ( .A1(n14879), .A2(n14744), .ZN(n14745) );
  NOR2_X1 U16754 ( .A1(n17161), .A2(n21592), .ZN(n14747) );
  AOI211_X1 U16755 ( .C1(P1_FLUSH_REG_SCAN_IN), .C2(n21582), .A(n21736), .B(
        n14747), .ZN(n16393) );
  INV_X1 U16756 ( .A(n16393), .ZN(n14752) );
  INV_X1 U16757 ( .A(n21784), .ZN(n21871) );
  NOR2_X1 U16758 ( .A1(n14748), .A2(n21871), .ZN(n14749) );
  XOR2_X1 U16759 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n14749), .Z(
        n14917) );
  NAND4_X1 U16760 ( .A1(n14752), .A2(n16385), .A3(n14750), .A4(n14917), .ZN(
        n14751) );
  OAI21_X1 U16761 ( .B1(n14752), .B2(n14922), .A(n14751), .ZN(P1_U3468) );
  INV_X1 U16762 ( .A(n21823), .ZN(n15263) );
  INV_X1 U16763 ( .A(n13845), .ZN(n14755) );
  NAND3_X1 U16764 ( .A1(n14755), .A2(n14753), .A3(n14754), .ZN(n14756) );
  NOR2_X1 U16765 ( .A1(n14757), .A2(n14756), .ZN(n14758) );
  AND2_X1 U16766 ( .A1(n14758), .A2(n13855), .ZN(n16375) );
  NAND2_X1 U16767 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14760) );
  INV_X1 U16768 ( .A(n14760), .ZN(n14759) );
  MUX2_X1 U16769 ( .A(n14760), .B(n14759), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14761) );
  INV_X1 U16770 ( .A(n14761), .ZN(n14769) );
  MUX2_X1 U16771 ( .A(n14763), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14762), .Z(n14765) );
  NOR2_X1 U16772 ( .A1(n14765), .A2(n14764), .ZN(n14768) );
  NAND2_X1 U16773 ( .A1(n14767), .A2(n14766), .ZN(n14903) );
  AOI22_X1 U16774 ( .A1(n17152), .A2(n14769), .B1(n14768), .B2(n14903), .ZN(
        n14774) );
  INV_X1 U16775 ( .A(n14771), .ZN(n14772) );
  OAI211_X1 U16776 ( .C1(n14762), .C2(n14776), .A(n13521), .B(n14772), .ZN(
        n14775) );
  NAND3_X1 U16777 ( .A1(n16375), .A2(n14708), .A3(n14775), .ZN(n14773) );
  OAI211_X1 U16778 ( .C1(n15263), .C2(n16375), .A(n14774), .B(n14773), .ZN(
        n14912) );
  INV_X1 U16779 ( .A(n16380), .ZN(n21587) );
  AOI22_X1 U16780 ( .A1(n14912), .A2(n16385), .B1(n14775), .B2(n21587), .ZN(
        n14777) );
  MUX2_X1 U16781 ( .A(n14777), .B(n14776), .S(n16393), .Z(n14778) );
  INV_X1 U16782 ( .A(n14778), .ZN(P1_U3469) );
  OAI21_X1 U16783 ( .B1(n14780), .B2(n14779), .A(n14867), .ZN(n15275) );
  INV_X1 U16784 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14782) );
  OAI222_X1 U16785 ( .A1(n15275), .A2(n15965), .B1(n14782), .B2(n19989), .C1(
        n14781), .C2(n19979), .ZN(P1_U2871) );
  NOR2_X1 U16786 ( .A1(n20043), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14783) );
  AOI211_X1 U16787 ( .C1(n20038), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14784), .B(n14783), .ZN(n14787) );
  NAND3_X1 U16788 ( .A1(n14785), .A2(n14723), .A3(n20039), .ZN(n14786) );
  OAI211_X1 U16789 ( .C1(n15275), .C2(n20022), .A(n14787), .B(n14786), .ZN(
        P1_U2998) );
  INV_X1 U16790 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14789) );
  AOI22_X1 U16791 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n19905), .B1(n19897), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14788) );
  OAI21_X1 U16792 ( .B1(n14789), .B2(n14803), .A(n14788), .ZN(P1_U2920) );
  INV_X1 U16793 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14791) );
  AOI22_X1 U16794 ( .A1(n19897), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14790) );
  OAI21_X1 U16795 ( .B1(n14791), .B2(n14803), .A(n14790), .ZN(P1_U2919) );
  INV_X1 U16796 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14793) );
  AOI22_X1 U16797 ( .A1(n21264), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14792) );
  OAI21_X1 U16798 ( .B1(n14793), .B2(n14803), .A(n14792), .ZN(P1_U2916) );
  INV_X1 U16799 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21696) );
  AOI22_X1 U16800 ( .A1(n21264), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14794) );
  OAI21_X1 U16801 ( .B1(n21696), .B2(n14803), .A(n14794), .ZN(P1_U2910) );
  INV_X1 U16802 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n21706) );
  AOI22_X1 U16803 ( .A1(n21264), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14795) );
  OAI21_X1 U16804 ( .B1(n21706), .B2(n14803), .A(n14795), .ZN(P1_U2908) );
  INV_X1 U16805 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14797) );
  AOI22_X1 U16806 ( .A1(n21264), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14796) );
  OAI21_X1 U16807 ( .B1(n14797), .B2(n14803), .A(n14796), .ZN(P1_U2917) );
  INV_X1 U16808 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n21711) );
  AOI22_X1 U16809 ( .A1(n21264), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14798) );
  OAI21_X1 U16810 ( .B1(n21711), .B2(n14803), .A(n14798), .ZN(P1_U2907) );
  INV_X1 U16811 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n21716) );
  AOI22_X1 U16812 ( .A1(n21264), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14799) );
  OAI21_X1 U16813 ( .B1(n21716), .B2(n14803), .A(n14799), .ZN(P1_U2906) );
  INV_X1 U16814 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U16815 ( .A1(n21264), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14800) );
  OAI21_X1 U16816 ( .B1(n14801), .B2(n14803), .A(n14800), .ZN(P1_U2918) );
  INV_X1 U16817 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n21701) );
  AOI22_X1 U16818 ( .A1(n21264), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14802) );
  OAI21_X1 U16819 ( .B1(n21701), .B2(n14803), .A(n14802), .ZN(P1_U2909) );
  INV_X1 U16820 ( .A(n14804), .ZN(n14807) );
  INV_X1 U16821 ( .A(n14805), .ZN(n14806) );
  NAND2_X1 U16822 ( .A1(n14807), .A2(n14806), .ZN(n14808) );
  NAND2_X1 U16823 ( .A1(n15128), .A2(n14810), .ZN(n14955) );
  NAND2_X1 U16824 ( .A1(n14955), .A2(n14811), .ZN(n14812) );
  NOR2_X1 U16825 ( .A1(n16473), .A2(n14814), .ZN(n14815) );
  AOI21_X1 U16826 ( .B1(n14681), .B2(n16473), .A(n14815), .ZN(n14816) );
  OAI21_X1 U16827 ( .B1(n19424), .B2(n16524), .A(n14816), .ZN(P2_U2886) );
  INV_X1 U16828 ( .A(n14819), .ZN(n15157) );
  NOR2_X1 U16829 ( .A1(n15157), .A2(n16513), .ZN(n14820) );
  AOI21_X1 U16830 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n16513), .A(n14820), .ZN(
        n14821) );
  OAI21_X1 U16831 ( .B1(n19431), .B2(n16524), .A(n14821), .ZN(P2_U2884) );
  NAND2_X1 U16832 ( .A1(n14822), .A2(n15075), .ZN(n15049) );
  XOR2_X1 U16833 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n15049), .Z(n14827)
         );
  OR2_X1 U16834 ( .A1(n14824), .A2(n14823), .ZN(n14825) );
  NAND2_X1 U16835 ( .A1(n14825), .A2(n15045), .ZN(n17402) );
  MUX2_X1 U16836 ( .A(n15418), .B(n17402), .S(n16473), .Z(n14826) );
  OAI21_X1 U16837 ( .B1(n14827), .B2(n16524), .A(n14826), .ZN(P2_U2882) );
  MUX2_X1 U16838 ( .A(n11919), .B(n11943), .S(n16473), .Z(n14832) );
  OAI21_X1 U16839 ( .B1(n19579), .B2(n16524), .A(n14832), .ZN(P2_U2885) );
  OR2_X1 U16840 ( .A1(n14822), .A2(n15075), .ZN(n14833) );
  NAND2_X1 U16841 ( .A1(n15049), .A2(n14833), .ZN(n19484) );
  NAND2_X1 U16842 ( .A1(n14835), .A2(n14834), .ZN(n14837) );
  INV_X1 U16843 ( .A(n14823), .ZN(n14836) );
  NAND2_X1 U16844 ( .A1(n14837), .A2(n14836), .ZN(n18399) );
  MUX2_X1 U16845 ( .A(n18396), .B(n18399), .S(n16473), .Z(n14838) );
  OAI21_X1 U16846 ( .B1(n19484), .B2(n16524), .A(n14838), .ZN(P2_U2883) );
  NAND2_X1 U16847 ( .A1(n12651), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14839) );
  AND4_X1 U16848 ( .A1(n14840), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n14839), 
        .A4(n12654), .ZN(n14841) );
  MUX2_X1 U16849 ( .A(n12950), .B(n14843), .S(n16513), .Z(n14844) );
  OAI21_X1 U16850 ( .B1(n19425), .B2(n16524), .A(n14844), .ZN(P2_U2887) );
  INV_X1 U16851 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n15240) );
  AOI22_X1 U16852 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17464), .B1(n17473), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14845) );
  OAI21_X1 U16853 ( .B1(n15240), .B2(n14862), .A(n14845), .ZN(P2_U2935) );
  AOI22_X1 U16854 ( .A1(n17473), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14846) );
  OAI21_X1 U16855 ( .B1(n16525), .B2(n14862), .A(n14846), .ZN(P2_U2923) );
  AOI22_X1 U16856 ( .A1(n17473), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14847) );
  OAI21_X1 U16857 ( .B1(n16571), .B2(n14862), .A(n14847), .ZN(P2_U2929) );
  AOI22_X1 U16858 ( .A1(n17473), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14848) );
  OAI21_X1 U16859 ( .B1(n16557), .B2(n14862), .A(n14848), .ZN(P2_U2927) );
  INV_X1 U16860 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14850) );
  AOI22_X1 U16861 ( .A1(n17473), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14849) );
  OAI21_X1 U16862 ( .B1(n14850), .B2(n14862), .A(n14849), .ZN(P2_U2928) );
  AOI22_X1 U16863 ( .A1(n17473), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14851) );
  OAI21_X1 U16864 ( .B1(n14852), .B2(n14862), .A(n14851), .ZN(P2_U2926) );
  AOI22_X1 U16865 ( .A1(n17473), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14853) );
  OAI21_X1 U16866 ( .B1(n15497), .B2(n14862), .A(n14853), .ZN(P2_U2931) );
  AOI22_X1 U16867 ( .A1(n17473), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14854) );
  OAI21_X1 U16868 ( .B1(n14855), .B2(n14862), .A(n14854), .ZN(P2_U2924) );
  AOI22_X1 U16869 ( .A1(n17473), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14856) );
  OAI21_X1 U16870 ( .B1(n16539), .B2(n14862), .A(n14856), .ZN(P2_U2925) );
  INV_X1 U16871 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15522) );
  AOI22_X1 U16872 ( .A1(n17473), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14857) );
  OAI21_X1 U16873 ( .B1(n15522), .B2(n14862), .A(n14857), .ZN(P2_U2930) );
  AOI22_X1 U16874 ( .A1(n17473), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14858) );
  OAI21_X1 U16875 ( .B1(n14859), .B2(n14862), .A(n14858), .ZN(P2_U2922) );
  INV_X1 U16876 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15452) );
  AOI22_X1 U16877 ( .A1(n17465), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14860) );
  OAI21_X1 U16878 ( .B1(n15452), .B2(n14862), .A(n14860), .ZN(P2_U2932) );
  AOI22_X1 U16879 ( .A1(n17465), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14861) );
  OAI21_X1 U16880 ( .B1(n15804), .B2(n14862), .A(n14861), .ZN(P2_U2921) );
  OAI21_X1 U16881 ( .B1(n14864), .B2(n14863), .A(n15068), .ZN(n21287) );
  INV_X1 U16882 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14869) );
  NAND2_X1 U16883 ( .A1(n14866), .A2(n14867), .ZN(n14868) );
  AND2_X1 U16884 ( .A1(n14865), .A2(n14868), .ZN(n21366) );
  INV_X1 U16885 ( .A(n21366), .ZN(n14894) );
  OAI222_X1 U16886 ( .A1(n21287), .A2(n19979), .B1(n14869), .B2(n19989), .C1(
        n14894), .C2(n15965), .ZN(P1_U2870) );
  OAI21_X1 U16887 ( .B1(n14870), .B2(n14871), .A(n14873), .ZN(n21291) );
  AOI22_X1 U16888 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n21348), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14874) );
  OAI21_X1 U16889 ( .B1(n20043), .B2(n21361), .A(n14874), .ZN(n14875) );
  AOI21_X1 U16890 ( .B1(n21366), .B2(n21732), .A(n14875), .ZN(n14876) );
  OAI21_X1 U16891 ( .B1(n21574), .B2(n21291), .A(n14876), .ZN(P1_U2997) );
  NOR2_X1 U16892 ( .A1(n14877), .A2(n15814), .ZN(n14878) );
  AND2_X1 U16893 ( .A1(n22117), .A2(n14882), .ZN(n14888) );
  INV_X1 U16894 ( .A(n14888), .ZN(n14883) );
  AND2_X1 U16895 ( .A1(n14883), .A2(n14889), .ZN(n14884) );
  INV_X1 U16896 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n14885) );
  OR2_X1 U16897 ( .A1(n21731), .A2(n14885), .ZN(n14887) );
  NAND2_X1 U16898 ( .A1(n21731), .A2(DATAI_0_), .ZN(n14886) );
  INV_X1 U16899 ( .A(n16027), .ZN(n14890) );
  NOR2_X1 U16900 ( .A1(n15655), .A2(n14889), .ZN(n15616) );
  INV_X1 U16901 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19884) );
  OAI222_X1 U16902 ( .A1(n16033), .A2(n15892), .B1(n21729), .B2(n16040), .C1(
        n16039), .C2(n19884), .ZN(P1_U2904) );
  INV_X1 U16903 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n14891) );
  OR2_X1 U16904 ( .A1(n21731), .A2(n14891), .ZN(n14893) );
  NAND2_X1 U16905 ( .A1(n21731), .A2(DATAI_2_), .ZN(n14892) );
  AND2_X1 U16906 ( .A1(n14893), .A2(n14892), .ZN(n21976) );
  INV_X1 U16907 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19888) );
  OAI222_X1 U16908 ( .A1(n16033), .A2(n14894), .B1(n21976), .B2(n16040), .C1(
        n16039), .C2(n19888), .ZN(P1_U2902) );
  XOR2_X1 U16909 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n15050), .Z(n14900)
         );
  NAND2_X1 U16910 ( .A1(n14897), .A2(n14896), .ZN(n15082) );
  OR2_X1 U16911 ( .A1(n14897), .A2(n14896), .ZN(n14898) );
  NAND2_X1 U16912 ( .A1(n15082), .A2(n14898), .ZN(n18416) );
  MUX2_X1 U16913 ( .A(n12401), .B(n18416), .S(n16473), .Z(n14899) );
  OAI21_X1 U16914 ( .B1(n14900), .B2(n16524), .A(n14899), .ZN(P2_U2880) );
  INV_X1 U16915 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19886) );
  OR2_X1 U16916 ( .A1(n21731), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14902) );
  INV_X1 U16917 ( .A(DATAI_1_), .ZN(n17290) );
  NAND2_X1 U16918 ( .A1(n21731), .A2(n17290), .ZN(n14901) );
  NAND2_X1 U16919 ( .A1(n14902), .A2(n14901), .ZN(n21933) );
  OAI222_X1 U16920 ( .A1(n15275), .A2(n16033), .B1(n16039), .B2(n19886), .C1(
        n21933), .C2(n16040), .ZN(P1_U2903) );
  INV_X1 U16921 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21575) );
  NAND2_X1 U16922 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21575), .ZN(n14923) );
  INV_X1 U16923 ( .A(n14764), .ZN(n14914) );
  OR2_X1 U16924 ( .A1(n21872), .A2(n16375), .ZN(n14911) );
  INV_X1 U16925 ( .A(n16375), .ZN(n14908) );
  XNOR2_X1 U16926 ( .A(n14762), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14904) );
  INV_X1 U16927 ( .A(n14904), .ZN(n16390) );
  NAND2_X1 U16928 ( .A1(n14708), .A2(n16390), .ZN(n14907) );
  XNOR2_X1 U16929 ( .A(n13370), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14905) );
  AOI22_X1 U16930 ( .A1(n17152), .A2(n14905), .B1(n14904), .B2(n14903), .ZN(
        n14906) );
  OAI21_X1 U16931 ( .B1(n14908), .B2(n14907), .A(n14906), .ZN(n14909) );
  INV_X1 U16932 ( .A(n14909), .ZN(n14910) );
  NAND2_X1 U16933 ( .A1(n14911), .A2(n14910), .ZN(n16386) );
  MUX2_X1 U16934 ( .A(n16386), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n17161), .Z(n17163) );
  MUX2_X1 U16935 ( .A(n14912), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n17161), .Z(n17164) );
  NAND3_X1 U16936 ( .A1(n17163), .A2(n17164), .A3(n16379), .ZN(n14913) );
  OAI21_X1 U16937 ( .B1(n14923), .B2(n14914), .A(n14913), .ZN(n17175) );
  INV_X1 U16938 ( .A(n17175), .ZN(n14916) );
  NOR2_X1 U16939 ( .A1(n14916), .A2(n14915), .ZN(n15036) );
  INV_X1 U16940 ( .A(n14917), .ZN(n21374) );
  NOR2_X1 U16941 ( .A1(n13855), .A2(n21374), .ZN(n14918) );
  OAI21_X1 U16942 ( .B1(n17161), .B2(n14918), .A(n16379), .ZN(n14919) );
  AOI21_X1 U16943 ( .B1(n17161), .B2(n14922), .A(n14919), .ZN(n14920) );
  INV_X1 U16944 ( .A(n14920), .ZN(n14921) );
  OAI21_X1 U16945 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n17169) );
  NOR3_X1 U16946 ( .A1(n15036), .A2(n17169), .A3(P1_FLUSH_REG_SCAN_IN), .ZN(
        n14925) );
  INV_X1 U16947 ( .A(n21582), .ZN(n21578) );
  NAND2_X1 U16948 ( .A1(n21896), .A2(n21900), .ZN(n21869) );
  OAI21_X1 U16949 ( .B1(n21759), .B2(n21923), .A(n21869), .ZN(n21858) );
  AOI21_X1 U16950 ( .B1(n21895), .B2(n21896), .A(n21858), .ZN(n21928) );
  NAND2_X1 U16951 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21881), .ZN(n14933) );
  AND2_X1 U16952 ( .A1(n21868), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14929) );
  NAND2_X1 U16953 ( .A1(n21759), .A2(n14929), .ZN(n14934) );
  NOR2_X1 U16954 ( .A1(n21810), .A2(n14934), .ZN(n21816) );
  AOI21_X1 U16955 ( .B1(n14933), .B2(n21823), .A(n21816), .ZN(n14930) );
  OAI21_X1 U16956 ( .B1(n21928), .B2(n21821), .A(n14930), .ZN(n14931) );
  NAND2_X1 U16957 ( .A1(n17190), .A2(n14931), .ZN(n14932) );
  OAI21_X1 U16958 ( .B1(n17190), .B2(n13778), .A(n14932), .ZN(P1_U3475) );
  INV_X1 U16959 ( .A(n14933), .ZN(n16373) );
  INV_X1 U16960 ( .A(n21858), .ZN(n14935) );
  MUX2_X1 U16961 ( .A(n14935), .B(n14934), .S(n14926), .Z(n14936) );
  OAI21_X1 U16962 ( .B1(n16373), .B2(n21872), .A(n14936), .ZN(n14937) );
  NAND2_X1 U16963 ( .A1(n17190), .A2(n14937), .ZN(n14938) );
  OAI21_X1 U16964 ( .B1(n17190), .B2(n21875), .A(n14938), .ZN(P1_U3476) );
  INV_X1 U16965 ( .A(n14970), .ZN(n14976) );
  NAND3_X1 U16966 ( .A1(n14962), .A2(n13081), .A3(n15013), .ZN(n14942) );
  INV_X1 U16967 ( .A(n14939), .ZN(n14940) );
  NAND2_X1 U16968 ( .A1(n14940), .A2(n17066), .ZN(n14958) );
  AOI22_X1 U16969 ( .A1(n14942), .A2(n14958), .B1(n14941), .B2(n14981), .ZN(
        n14946) );
  NOR2_X1 U16970 ( .A1(n12629), .A2(n12906), .ZN(n14959) );
  INV_X1 U16971 ( .A(n14941), .ZN(n14943) );
  NAND2_X1 U16972 ( .A1(n14981), .A2(n14943), .ZN(n17067) );
  OAI211_X1 U16973 ( .C1(n14959), .C2(n11975), .A(n17067), .B(n14958), .ZN(
        n14944) );
  INV_X1 U16974 ( .A(n14944), .ZN(n14945) );
  MUX2_X1 U16975 ( .A(n14946), .B(n14945), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14947) );
  INV_X1 U16976 ( .A(n14947), .ZN(n14948) );
  AOI21_X1 U16977 ( .B1(n14819), .B2(n14976), .A(n14948), .ZN(n17076) );
  INV_X1 U16978 ( .A(n14949), .ZN(n14951) );
  NOR2_X1 U16979 ( .A1(n12599), .A2(n15029), .ZN(n14950) );
  NAND2_X1 U16980 ( .A1(n14951), .A2(n14950), .ZN(n14957) );
  NAND2_X1 U16981 ( .A1(n15017), .A2(n15015), .ZN(n14952) );
  AND2_X1 U16982 ( .A1(n14953), .A2(n14952), .ZN(n14956) );
  NAND4_X1 U16983 ( .A1(n14957), .A2(n14956), .A3(n14955), .A4(n14954), .ZN(
        n15441) );
  MUX2_X1 U16984 ( .A(n11832), .B(n17076), .S(n15441), .Z(n14999) );
  NAND2_X1 U16985 ( .A1(n15331), .A2(n14976), .ZN(n14966) );
  NAND2_X1 U16986 ( .A1(n13081), .A2(n14958), .ZN(n14960) );
  OAI22_X1 U16987 ( .A1(n17067), .A2(n11139), .B1(n14959), .B2(n14960), .ZN(
        n14964) );
  INV_X1 U16988 ( .A(n14960), .ZN(n14961) );
  AOI21_X1 U16989 ( .B1(n14962), .B2(n15013), .A(n14961), .ZN(n14963) );
  NOR2_X1 U16990 ( .A1(n14964), .A2(n14963), .ZN(n14965) );
  NAND2_X1 U16991 ( .A1(n14966), .A2(n14965), .ZN(n17072) );
  NAND2_X1 U16992 ( .A1(n17072), .A2(n15441), .ZN(n14969) );
  NAND2_X1 U16993 ( .A1(n15441), .A2(n17067), .ZN(n14967) );
  NAND2_X1 U16994 ( .A1(n14967), .A2(n10990), .ZN(n14968) );
  NAND2_X1 U16995 ( .A1(n14969), .A2(n14968), .ZN(n14990) );
  INV_X1 U16996 ( .A(n14990), .ZN(n14997) );
  OR2_X1 U16997 ( .A1(n12950), .A2(n14970), .ZN(n14975) );
  INV_X1 U16998 ( .A(n14981), .ZN(n14973) );
  AND2_X1 U16999 ( .A1(n11120), .A2(n14971), .ZN(n14977) );
  MUX2_X1 U17000 ( .A(n14973), .B(n14977), .S(n14972), .Z(n14974) );
  NAND2_X1 U17001 ( .A1(n14975), .A2(n14974), .ZN(n15439) );
  NAND2_X1 U17002 ( .A1(n14681), .A2(n14976), .ZN(n14985) );
  INV_X1 U17003 ( .A(n14977), .ZN(n14983) );
  INV_X1 U17004 ( .A(n11969), .ZN(n14980) );
  INV_X1 U17005 ( .A(n14978), .ZN(n14979) );
  NAND2_X1 U17006 ( .A1(n14980), .A2(n14979), .ZN(n14982) );
  AOI22_X1 U17007 ( .A1(n14983), .A2(n14982), .B1(n14981), .B2(n11139), .ZN(
        n14984) );
  NAND2_X1 U17008 ( .A1(n14985), .A2(n14984), .ZN(n17061) );
  OAI21_X1 U17009 ( .B1(n15439), .B2(n19302), .A(n17061), .ZN(n14988) );
  OAI21_X1 U17010 ( .B1(n15439), .B2(n19353), .A(n14986), .ZN(n14987) );
  NAND2_X1 U17011 ( .A1(n14988), .A2(n14987), .ZN(n14989) );
  NAND2_X1 U17012 ( .A1(n14989), .A2(n15441), .ZN(n14992) );
  NOR2_X1 U17013 ( .A1(n14992), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14991) );
  OR2_X1 U17014 ( .A1(n14991), .A2(n14990), .ZN(n14994) );
  NAND2_X1 U17015 ( .A1(n14992), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14993) );
  NAND2_X1 U17016 ( .A1(n14994), .A2(n14993), .ZN(n14998) );
  OR2_X1 U17017 ( .A1(n14998), .A2(n14999), .ZN(n14995) );
  AND2_X1 U17018 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n14995), .ZN(
        n14996) );
  OAI22_X1 U17019 ( .A1(n14999), .A2(n14997), .B1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n14996), .ZN(n15028) );
  NAND2_X1 U17020 ( .A1(n14999), .A2(n14998), .ZN(n15027) );
  OR2_X1 U17021 ( .A1(n17134), .A2(n15000), .ZN(n15001) );
  OAI21_X1 U17022 ( .B1(n15003), .B2(n15002), .A(n15001), .ZN(n15009) );
  INV_X1 U17023 ( .A(n15004), .ZN(n15005) );
  AND2_X1 U17024 ( .A1(n15006), .A2(n15005), .ZN(n15007) );
  AOI21_X1 U17025 ( .B1(n15009), .B2(n15008), .A(n15007), .ZN(n15012) );
  NAND2_X1 U17026 ( .A1(n15010), .A2(n15128), .ZN(n15011) );
  OAI211_X1 U17027 ( .C1(n15128), .C2(n15013), .A(n15012), .B(n15011), .ZN(
        n18720) );
  NOR2_X1 U17028 ( .A1(n15015), .A2(n15014), .ZN(n15016) );
  AND2_X1 U17029 ( .A1(n15017), .A2(n15016), .ZN(n18719) );
  OAI21_X1 U17030 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18719), .ZN(n15023) );
  INV_X1 U17031 ( .A(n18655), .ZN(n15018) );
  NAND3_X1 U17032 ( .A1(n15020), .A2(n15019), .A3(n15018), .ZN(n15021) );
  NAND3_X1 U17033 ( .A1(n15023), .A2(n15022), .A3(n15021), .ZN(n15024) );
  NOR2_X1 U17034 ( .A1(n18720), .A2(n15024), .ZN(n15025) );
  OAI21_X1 U17035 ( .B1(n15441), .B2(n18660), .A(n15025), .ZN(n15026) );
  AOI21_X1 U17036 ( .B1(n15028), .B2(n15027), .A(n15026), .ZN(n18712) );
  NAND3_X1 U17037 ( .A1(n18712), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n17057), 
        .ZN(n15032) );
  NOR2_X1 U17038 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n15029), .ZN(n15295) );
  AND2_X1 U17039 ( .A1(n15030), .A2(n15295), .ZN(n15307) );
  AOI22_X1 U17040 ( .A1(n15032), .A2(n15129), .B1(n15031), .B2(n15307), .ZN(
        n18704) );
  INV_X1 U17041 ( .A(n18704), .ZN(n15034) );
  NOR2_X1 U17042 ( .A1(n18711), .A2(n17419), .ZN(n17136) );
  AOI21_X1 U17043 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n18711), .A(n17136), 
        .ZN(n15033) );
  OAI21_X1 U17044 ( .B1(n15034), .B2(n12654), .A(n15033), .ZN(P2_U3593) );
  NOR3_X1 U17045 ( .A1(n15036), .A2(n17169), .A3(n15035), .ZN(n21590) );
  INV_X1 U17046 ( .A(n21772), .ZN(n15685) );
  OAI22_X1 U17047 ( .A1(n14035), .A2(n21923), .B1(n15685), .B2(n16373), .ZN(
        n15037) );
  OAI21_X1 U17048 ( .B1(n21590), .B2(n15037), .A(n17190), .ZN(n15038) );
  OAI21_X1 U17049 ( .B1(n17190), .B2(n21885), .A(n15038), .ZN(P1_U3478) );
  NOR2_X1 U17050 ( .A1(n15050), .A2(n17095), .ZN(n15087) );
  NAND2_X1 U17051 ( .A1(n15087), .A2(n15086), .ZN(n15085) );
  XNOR2_X1 U17052 ( .A(n15085), .B(n15054), .ZN(n15044) );
  NAND2_X1 U17053 ( .A1(n15040), .A2(n15041), .ZN(n15042) );
  NAND2_X1 U17054 ( .A1(n15039), .A2(n15042), .ZN(n16986) );
  INV_X1 U17055 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n15435) );
  MUX2_X1 U17056 ( .A(n16986), .B(n15435), .S(n16513), .Z(n15043) );
  OAI21_X1 U17057 ( .B1(n15044), .B2(n16524), .A(n15043), .ZN(P2_U2878) );
  NAND2_X1 U17058 ( .A1(n15046), .A2(n15045), .ZN(n15048) );
  INV_X1 U17059 ( .A(n14896), .ZN(n15047) );
  NAND2_X1 U17060 ( .A1(n15048), .A2(n15047), .ZN(n17037) );
  NOR2_X1 U17061 ( .A1(n15049), .A2(n19479), .ZN(n15051) );
  OAI211_X1 U17062 ( .C1(n15051), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15147), .B(n15050), .ZN(n15053) );
  NAND2_X1 U17063 ( .A1(n16513), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n15052) );
  OAI211_X1 U17064 ( .C1(n17037), .C2(n16513), .A(n15053), .B(n15052), .ZN(
        P2_U2881) );
  INV_X1 U17065 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n15305) );
  NOR2_X1 U17066 ( .A1(n15085), .A2(n15054), .ZN(n15057) );
  NAND2_X1 U17067 ( .A1(n15087), .A2(n15055), .ZN(n15111) );
  OAI211_X1 U17068 ( .C1(n15057), .C2(n15056), .A(n15147), .B(n15111), .ZN(
        n15064) );
  INV_X1 U17069 ( .A(n15058), .ZN(n15061) );
  NAND2_X1 U17070 ( .A1(n15039), .A2(n15059), .ZN(n15060) );
  NAND2_X1 U17071 ( .A1(n15061), .A2(n15060), .ZN(n16972) );
  INV_X1 U17072 ( .A(n16972), .ZN(n15062) );
  NAND2_X1 U17073 ( .A1(n15062), .A2(n16473), .ZN(n15063) );
  OAI211_X1 U17074 ( .C1(n16473), .C2(n15305), .A(n15064), .B(n15063), .ZN(
        P2_U2877) );
  XOR2_X1 U17075 ( .A(n15065), .B(n15066), .Z(n15249) );
  INV_X1 U17076 ( .A(n15249), .ZN(n15099) );
  INV_X1 U17077 ( .A(n17194), .ZN(n15067) );
  AOI21_X1 U17078 ( .B1(n15069), .B2(n15068), .A(n15067), .ZN(n21314) );
  AOI22_X1 U17079 ( .A1(n21314), .A2(n19985), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n17196), .ZN(n15070) );
  OAI21_X1 U17080 ( .B1(n15099), .B2(n15965), .A(n15070), .ZN(P1_U2869) );
  NAND2_X1 U17081 ( .A1(n15072), .A2(n15073), .ZN(n15074) );
  NAND2_X1 U17082 ( .A1(n15071), .A2(n15074), .ZN(n18452) );
  AND2_X1 U17083 ( .A1(n14822), .A2(n15075), .ZN(n15077) );
  AND2_X1 U17084 ( .A1(n15077), .A2(n15076), .ZN(n15110) );
  OAI211_X1 U17085 ( .C1(n15110), .C2(n15079), .A(n15078), .B(n15147), .ZN(
        n15081) );
  NAND2_X1 U17086 ( .A1(n16513), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15080) );
  OAI211_X1 U17087 ( .C1(n18452), .C2(n16513), .A(n15081), .B(n15080), .ZN(
        P2_U2875) );
  INV_X1 U17088 ( .A(n15082), .ZN(n15084) );
  OAI21_X1 U17089 ( .B1(n15084), .B2(n15083), .A(n15040), .ZN(n18427) );
  OAI211_X1 U17090 ( .C1(n15087), .C2(n15086), .A(n15085), .B(n15147), .ZN(
        n15089) );
  NAND2_X1 U17091 ( .A1(n16513), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n15088) );
  OAI211_X1 U17092 ( .C1(n18427), .C2(n16513), .A(n15089), .B(n15088), .ZN(
        P2_U2879) );
  OAI21_X1 U17093 ( .B1(n15091), .B2(n15093), .A(n15092), .ZN(n21312) );
  AOI22_X1 U17094 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n21348), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n15094) );
  OAI21_X1 U17095 ( .B1(n20043), .B2(n15259), .A(n15094), .ZN(n15095) );
  AOI21_X1 U17096 ( .B1(n15249), .B2(n21732), .A(n15095), .ZN(n15096) );
  OAI21_X1 U17097 ( .B1(n21312), .B2(n21574), .A(n15096), .ZN(P1_U2996) );
  INV_X1 U17098 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19890) );
  OR2_X1 U17099 ( .A1(n21731), .A2(BUF1_REG_3__SCAN_IN), .ZN(n15098) );
  INV_X1 U17100 ( .A(DATAI_3_), .ZN(n17337) );
  NAND2_X1 U17101 ( .A1(n21731), .A2(n17337), .ZN(n15097) );
  NAND2_X1 U17102 ( .A1(n15098), .A2(n15097), .ZN(n22022) );
  OAI222_X1 U17103 ( .A1(n15099), .A2(n16033), .B1(n16039), .B2(n19890), .C1(
        n22022), .C2(n16040), .ZN(P1_U2901) );
  NAND2_X1 U17104 ( .A1(n15103), .A2(n15102), .ZN(n15104) );
  AND2_X1 U17105 ( .A1(n15101), .A2(n15104), .ZN(n21379) );
  INV_X1 U17106 ( .A(n21379), .ZN(n15107) );
  INV_X1 U17107 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19892) );
  OR2_X1 U17108 ( .A1(n21731), .A2(BUF1_REG_4__SCAN_IN), .ZN(n15106) );
  INV_X1 U17109 ( .A(DATAI_4_), .ZN(n17292) );
  NAND2_X1 U17110 ( .A1(n21731), .A2(n17292), .ZN(n15105) );
  NAND2_X1 U17111 ( .A1(n15106), .A2(n15105), .ZN(n22068) );
  OAI222_X1 U17112 ( .A1(n15107), .A2(n16033), .B1(n19892), .B2(n16039), .C1(
        n22068), .C2(n16040), .ZN(P1_U2900) );
  OR2_X1 U17113 ( .A1(n15058), .A2(n15108), .ZN(n15109) );
  NAND2_X1 U17114 ( .A1(n15072), .A2(n15109), .ZN(n18442) );
  INV_X1 U17115 ( .A(n18442), .ZN(n16968) );
  INV_X1 U17116 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n18434) );
  NOR2_X1 U17117 ( .A1(n16473), .A2(n18434), .ZN(n15114) );
  AOI211_X1 U17118 ( .C1(n15112), .C2(n15111), .A(n16524), .B(n15110), .ZN(
        n15113) );
  AOI211_X1 U17119 ( .C1(n16968), .C2(n16473), .A(n15114), .B(n15113), .ZN(
        n15115) );
  INV_X1 U17120 ( .A(n15115), .ZN(P2_U2876) );
  INV_X1 U17121 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n18460) );
  INV_X1 U17122 ( .A(n15078), .ZN(n15117) );
  OAI211_X1 U17123 ( .C1(n15117), .C2(n15116), .A(n15147), .B(n15188), .ZN(
        n15122) );
  AND2_X1 U17124 ( .A1(n15071), .A2(n15119), .ZN(n15120) );
  NOR2_X1 U17125 ( .A1(n15118), .A2(n15120), .ZN(n18466) );
  NAND2_X1 U17126 ( .A1(n18466), .A2(n16473), .ZN(n15121) );
  OAI211_X1 U17127 ( .C1(n16473), .C2(n18460), .A(n15122), .B(n15121), .ZN(
        P2_U2874) );
  AOI21_X1 U17128 ( .B1(n15124), .B2(n15101), .A(n15123), .ZN(n21393) );
  INV_X1 U17129 ( .A(n21393), .ZN(n15153) );
  OR2_X1 U17130 ( .A1(n21731), .A2(BUF1_REG_5__SCAN_IN), .ZN(n15126) );
  INV_X1 U17131 ( .A(DATAI_5_), .ZN(n17293) );
  NAND2_X1 U17132 ( .A1(n21731), .A2(n17293), .ZN(n15125) );
  NAND2_X1 U17133 ( .A1(n15126), .A2(n15125), .ZN(n22114) );
  OAI222_X1 U17134 ( .A1(n16033), .A2(n15153), .B1(n16039), .B2(n14070), .C1(
        n22114), .C2(n16040), .ZN(P1_U2899) );
  INV_X1 U17135 ( .A(n17097), .ZN(n15127) );
  INV_X1 U17136 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n22214) );
  NAND2_X1 U17137 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n18711), .ZN(n18374) );
  NAND2_X1 U17138 ( .A1(n15129), .A2(n18374), .ZN(n18705) );
  INV_X1 U17139 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n20705) );
  OAI22_X2 U17140 ( .A1(n22214), .A2(n19707), .B1(n20705), .B2(n19706), .ZN(
        n19369) );
  INV_X1 U17141 ( .A(n19369), .ZN(n19282) );
  INV_X1 U17142 ( .A(n15140), .ZN(n15133) );
  NOR2_X1 U17143 ( .A1(n15132), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19235) );
  INV_X1 U17144 ( .A(n19235), .ZN(n19364) );
  NOR2_X1 U17145 ( .A1(n15133), .A2(n19364), .ZN(n15136) );
  NAND3_X1 U17146 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19257), .A3(
        n14986), .ZN(n19280) );
  NOR2_X1 U17147 ( .A1(n19353), .A2(n19280), .ZN(n19656) );
  INV_X1 U17148 ( .A(n19656), .ZN(n19745) );
  AOI21_X1 U17149 ( .B1(n19745), .B2(n19355), .A(n19700), .ZN(n15135) );
  AND2_X1 U17150 ( .A1(n19424), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n15226) );
  NAND2_X1 U17151 ( .A1(n19579), .A2(n15226), .ZN(n19358) );
  OR2_X1 U17152 ( .A1(n19431), .A2(n19358), .ZN(n15139) );
  NAND2_X1 U17153 ( .A1(n19280), .A2(n15139), .ZN(n15134) );
  OAI21_X1 U17154 ( .B1(n15136), .B2(n15135), .A(n15134), .ZN(n19749) );
  AOI22_X2 U17155 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19699), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19698), .ZN(n19372) );
  NAND2_X1 U17156 ( .A1(n19424), .A2(n19694), .ZN(n19341) );
  NAND2_X1 U17157 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19362), .ZN(n19641) );
  NAND2_X1 U17158 ( .A1(n12635), .A2(n19702), .ZN(n19281) );
  OAI22_X1 U17159 ( .A1(n19372), .A2(n19746), .B1(n19281), .B2(n19745), .ZN(
        n15137) );
  AOI21_X1 U17160 ( .B1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n19749), .A(
        n15137), .ZN(n15145) );
  NOR2_X1 U17161 ( .A1(n19355), .A2(n19280), .ZN(n15138) );
  NAND2_X1 U17162 ( .A1(n15139), .A2(n15138), .ZN(n15142) );
  OAI21_X1 U17163 ( .B1(n15140), .B2(n19656), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15141) );
  NAND2_X1 U17164 ( .A1(n15142), .A2(n15141), .ZN(n19748) );
  NAND2_X1 U17165 ( .A1(n19748), .A2(n15143), .ZN(n15144) );
  OAI211_X1 U17166 ( .C1(n19754), .C2(n19282), .A(n15145), .B(n15144), .ZN(
        P2_U3127) );
  OAI211_X1 U17167 ( .C1(n15187), .C2(n15148), .A(n15146), .B(n15147), .ZN(
        n15150) );
  NAND2_X1 U17168 ( .A1(n15717), .A2(n16473), .ZN(n15149) );
  OAI211_X1 U17169 ( .C1(n16473), .C2(n12442), .A(n15150), .B(n15149), .ZN(
        P2_U2872) );
  OR2_X1 U17170 ( .A1(n11086), .A2(n15151), .ZN(n15152) );
  NAND2_X1 U17171 ( .A1(n19973), .A2(n15152), .ZN(n21383) );
  INV_X1 U17172 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n15154) );
  OAI222_X1 U17173 ( .A1(n21383), .A2(n19979), .B1(n15154), .B2(n19989), .C1(
        n15153), .C2(n15965), .ZN(P1_U2867) );
  XNOR2_X1 U17174 ( .A(n15155), .B(n15156), .ZN(n15177) );
  AOI21_X1 U17175 ( .B1(n15339), .B2(n15285), .A(n15219), .ZN(n15336) );
  INV_X1 U17176 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n17482) );
  OAI22_X1 U17177 ( .A1(n15339), .A2(n17417), .B1(n17482), .B2(n18680), .ZN(
        n15159) );
  NOR2_X1 U17178 ( .A1(n15157), .A2(n17410), .ZN(n15158) );
  AOI211_X1 U17179 ( .C1(n17407), .C2(n15336), .A(n15159), .B(n15158), .ZN(
        n15163) );
  NAND3_X1 U17180 ( .A1(n15174), .A2(n16766), .A3(n15161), .ZN(n15162) );
  OAI211_X1 U17181 ( .C1(n15177), .C2(n17411), .A(n15163), .B(n15162), .ZN(
        P2_U3011) );
  XNOR2_X1 U17182 ( .A(n15165), .B(n15164), .ZN(n19430) );
  OAI22_X1 U17183 ( .A1(n18662), .A2(n19430), .B1(n17482), .B2(n18680), .ZN(
        n15173) );
  INV_X1 U17184 ( .A(n15660), .ZN(n15166) );
  NOR2_X1 U17185 ( .A1(n17005), .A2(n15166), .ZN(n15168) );
  NOR2_X1 U17186 ( .A1(n17002), .A2(n15659), .ZN(n15167) );
  OR2_X1 U17187 ( .A1(n15168), .A2(n15167), .ZN(n16997) );
  INV_X1 U17188 ( .A(n17052), .ZN(n15169) );
  NOR2_X1 U17189 ( .A1(n17002), .A2(n15169), .ZN(n15170) );
  NOR2_X1 U17190 ( .A1(n15170), .A2(n18665), .ZN(n15671) );
  INV_X1 U17191 ( .A(n17002), .ZN(n15171) );
  NAND2_X1 U17192 ( .A1(n15171), .A2(n15670), .ZN(n15668) );
  OAI211_X1 U17193 ( .C1(n15660), .C2(n17005), .A(n15671), .B(n15668), .ZN(
        n15211) );
  MUX2_X1 U17194 ( .A(n16997), .B(n15211), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n15172) );
  AOI211_X1 U17195 ( .C1(n18685), .C2(n14819), .A(n15173), .B(n15172), .ZN(
        n15176) );
  NAND3_X1 U17196 ( .A1(n15174), .A2(n15725), .A3(n15161), .ZN(n15175) );
  OAI211_X1 U17197 ( .C1(n15177), .C2(n18664), .A(n15176), .B(n15175), .ZN(
        P2_U3043) );
  OR2_X1 U17198 ( .A1(n15123), .A2(n15178), .ZN(n15180) );
  AND2_X1 U17199 ( .A1(n15180), .A2(n15179), .ZN(n21405) );
  INV_X1 U17200 ( .A(n21405), .ZN(n15183) );
  OR2_X1 U17201 ( .A1(n21731), .A2(BUF1_REG_6__SCAN_IN), .ZN(n15182) );
  INV_X1 U17202 ( .A(n21730), .ZN(n16036) );
  INV_X1 U17203 ( .A(DATAI_6_), .ZN(n17334) );
  NAND2_X1 U17204 ( .A1(n16036), .A2(n17334), .ZN(n15181) );
  NAND2_X1 U17205 ( .A1(n15182), .A2(n15181), .ZN(n22164) );
  OAI222_X1 U17206 ( .A1(n15183), .A2(n16033), .B1(n16039), .B2(n14080), .C1(
        n22164), .C2(n16040), .ZN(P1_U2898) );
  OR2_X1 U17207 ( .A1(n15118), .A2(n15184), .ZN(n15185) );
  NAND2_X1 U17208 ( .A1(n15186), .A2(n15185), .ZN(n18476) );
  NOR2_X1 U17209 ( .A1(n18476), .A2(n16513), .ZN(n15191) );
  AOI211_X1 U17210 ( .C1(n15189), .C2(n15188), .A(n16524), .B(n15187), .ZN(
        n15190) );
  AOI211_X1 U17211 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n16513), .A(n15191), .B(
        n15190), .ZN(n15192) );
  INV_X1 U17212 ( .A(n15192), .ZN(P2_U2873) );
  AOI21_X1 U17213 ( .B1(n15195), .B2(n15193), .A(n15194), .ZN(n15196) );
  INV_X1 U17214 ( .A(n15196), .ZN(n15401) );
  XNOR2_X1 U17215 ( .A(n15197), .B(n15198), .ZN(n16900) );
  INV_X1 U17216 ( .A(n16900), .ZN(n18505) );
  OAI22_X1 U17217 ( .A1(n19189), .A2(n19640), .B1(n15199), .B2(n19686), .ZN(
        n15200) );
  AOI21_X1 U17218 ( .B1(n18505), .B2(n19633), .A(n15200), .ZN(n15202) );
  AOI22_X1 U17219 ( .A1(n19185), .A2(BUF2_REG_17__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n15201) );
  OAI211_X1 U17220 ( .C1(n15401), .C2(n19636), .A(n15202), .B(n15201), .ZN(
        P2_U2902) );
  NAND2_X1 U17221 ( .A1(n15179), .A2(n15204), .ZN(n15205) );
  AND2_X1 U17222 ( .A1(n15347), .A2(n15205), .ZN(n20011) );
  INV_X1 U17223 ( .A(n20011), .ZN(n21414) );
  AOI21_X1 U17224 ( .B1(n15206), .B2(n19975), .A(n15376), .ZN(n21411) );
  AOI22_X1 U17225 ( .A1(n21411), .A2(n19985), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n17196), .ZN(n15207) );
  OAI21_X1 U17226 ( .B1(n21414), .B2(n15965), .A(n15207), .ZN(P1_U2865) );
  XNOR2_X1 U17227 ( .A(n15208), .B(n15209), .ZN(n15225) );
  XNOR2_X1 U17228 ( .A(n15210), .B(n18678), .ZN(n15223) );
  NAND2_X1 U17229 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16997), .ZN(
        n18676) );
  AOI21_X1 U17230 ( .B1(n15212), .B2(n18671), .A(n15211), .ZN(n18694) );
  NAND2_X1 U17231 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n18532), .ZN(n15213) );
  OAI221_X1 U17232 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18676), .C1(
        n18678), .C2(n18694), .A(n15213), .ZN(n15217) );
  XNOR2_X1 U17233 ( .A(n15214), .B(n15215), .ZN(n19481) );
  OAI22_X1 U17234 ( .A1(n19481), .A2(n18662), .B1(n18666), .B2(n18399), .ZN(
        n15216) );
  AOI211_X1 U17235 ( .C1(n15223), .C2(n15725), .A(n15217), .B(n15216), .ZN(
        n15218) );
  OAI21_X1 U17236 ( .B1(n15225), .B2(n18664), .A(n15218), .ZN(P2_U3042) );
  OAI21_X1 U17237 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n15219), .A(
        n15282), .ZN(n18402) );
  OAI22_X1 U17238 ( .A1(n12266), .A2(n18680), .B1(n16782), .B2(n18402), .ZN(
        n15220) );
  AOI21_X1 U17239 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16750), .A(
        n15220), .ZN(n15221) );
  OAI21_X1 U17240 ( .B1(n17410), .B2(n18399), .A(n15221), .ZN(n15222) );
  AOI21_X1 U17241 ( .B1(n15223), .B2(n16766), .A(n15222), .ZN(n15224) );
  OAI21_X1 U17242 ( .B1(n15225), .B2(n17411), .A(n15224), .ZN(P2_U3010) );
  INV_X1 U17243 ( .A(n15226), .ZN(n19313) );
  NAND3_X1 U17244 ( .A1(n14986), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19245) );
  OAI21_X1 U17245 ( .B1(n19225), .B2(n19313), .A(n19245), .ZN(n15230) );
  NAND2_X1 U17246 ( .A1(n15231), .A2(n19235), .ZN(n15228) );
  NOR2_X1 U17247 ( .A1(n19353), .A2(n19245), .ZN(n19719) );
  OAI21_X1 U17248 ( .B1(n19346), .B2(n19719), .A(n19362), .ZN(n15227) );
  NAND2_X1 U17249 ( .A1(n15228), .A2(n15227), .ZN(n15229) );
  NAND2_X1 U17250 ( .A1(n15230), .A2(n15229), .ZN(n19721) );
  INV_X1 U17251 ( .A(n19721), .ZN(n19594) );
  OAI21_X1 U17252 ( .B1(n15231), .B2(n19719), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15232) );
  OAI21_X1 U17253 ( .B1(n19245), .B2(n19355), .A(n15232), .ZN(n19720) );
  INV_X1 U17254 ( .A(n19719), .ZN(n19237) );
  INV_X1 U17255 ( .A(n19372), .ZN(n17109) );
  AOI22_X1 U17256 ( .A1(n19728), .A2(n19369), .B1(n19590), .B2(n17109), .ZN(
        n15234) );
  OAI21_X1 U17257 ( .B1(n19281), .B2(n19237), .A(n15234), .ZN(n15235) );
  AOI21_X1 U17258 ( .B1(n19720), .B2(n15143), .A(n15235), .ZN(n15236) );
  OAI21_X1 U17259 ( .B1(n19594), .B2(n15237), .A(n15236), .ZN(P2_U3159) );
  INV_X1 U17260 ( .A(n15146), .ZN(n15238) );
  OAI21_X1 U17261 ( .B1(n15238), .B2(n11413), .A(n15193), .ZN(n15320) );
  INV_X1 U17262 ( .A(n19701), .ZN(n15242) );
  OAI21_X1 U17263 ( .B1(n11060), .B2(n15239), .A(n15197), .ZN(n18495) );
  OAI22_X1 U17264 ( .A1(n18495), .A2(n19688), .B1(n15240), .B2(n19686), .ZN(
        n15241) );
  AOI21_X1 U17265 ( .B1(n16574), .B2(n15242), .A(n15241), .ZN(n15244) );
  AOI22_X1 U17266 ( .A1(n19185), .A2(BUF2_REG_16__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n15243) );
  OAI211_X1 U17267 ( .C1(n15320), .C2(n19636), .A(n15244), .B(n15243), .ZN(
        P2_U2903) );
  OR2_X1 U17268 ( .A1(n21731), .A2(BUF1_REG_7__SCAN_IN), .ZN(n15246) );
  INV_X1 U17269 ( .A(DATAI_7_), .ZN(n17231) );
  NAND2_X1 U17270 ( .A1(n16036), .A2(n17231), .ZN(n15245) );
  NAND2_X1 U17271 ( .A1(n15246), .A2(n15245), .ZN(n22211) );
  OAI222_X1 U17272 ( .A1(n21414), .A2(n16033), .B1(n16039), .B2(n14018), .C1(
        n22211), .C2(n16040), .ZN(P1_U2897) );
  INV_X1 U17273 ( .A(n15248), .ZN(n15247) );
  NAND2_X1 U17274 ( .A1(n15247), .A2(n11044), .ZN(n21373) );
  OAI21_X1 U17275 ( .B1(n15248), .B2(n15814), .A(n21553), .ZN(n21392) );
  NAND2_X1 U17276 ( .A1(n15249), .A2(n21392), .ZN(n15262) );
  NAND2_X1 U17277 ( .A1(n21551), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n15258) );
  OAI221_X1 U17278 ( .B1(n21403), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n21403), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n14514), .ZN(n15252) );
  NAND2_X1 U17279 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n15252), .ZN(n15255) );
  INV_X1 U17280 ( .A(n21403), .ZN(n21528) );
  INV_X1 U17281 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n15253) );
  NAND4_X1 U17282 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(n21528), .A4(n15253), .ZN(n15254) );
  NAND2_X1 U17283 ( .A1(n15255), .A2(n15254), .ZN(n15256) );
  AOI21_X1 U17284 ( .B1(n21564), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15256), .ZN(n15257) );
  OAI211_X1 U17285 ( .C1(n21560), .C2(n15259), .A(n15258), .B(n15257), .ZN(
        n15260) );
  AOI21_X1 U17286 ( .B1(n21519), .B2(n21314), .A(n15260), .ZN(n15261) );
  OAI211_X1 U17287 ( .C1(n15263), .C2(n21373), .A(n15262), .B(n15261), .ZN(
        P1_U2837) );
  INV_X1 U17288 ( .A(n21392), .ZN(n15274) );
  AOI22_X1 U17289 ( .A1(n21528), .A2(n15268), .B1(n21519), .B2(n14720), .ZN(
        n15271) );
  INV_X1 U17290 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15265) );
  NAND2_X1 U17291 ( .A1(n21521), .A2(n15265), .ZN(n15267) );
  NAND2_X1 U17292 ( .A1(n21564), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15266) );
  OAI211_X1 U17293 ( .C1(n15268), .C2(n14514), .A(n15267), .B(n15266), .ZN(
        n15269) );
  AOI21_X1 U17294 ( .B1(n21551), .B2(P1_EBX_REG_1__SCAN_IN), .A(n15269), .ZN(
        n15270) );
  OAI211_X1 U17295 ( .C1(n15264), .C2(n21373), .A(n15271), .B(n15270), .ZN(
        n15272) );
  INV_X1 U17296 ( .A(n15272), .ZN(n15273) );
  OAI21_X1 U17297 ( .B1(n15275), .B2(n15274), .A(n15273), .ZN(P1_U2839) );
  INV_X1 U17298 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15278) );
  AOI22_X2 U17299 ( .A1(n15761), .A2(n18711), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n15280), .ZN(n15429) );
  AOI21_X1 U17300 ( .B1(n15281), .B2(n16768), .A(n15288), .ZN(n16771) );
  AOI21_X1 U17301 ( .B1(n17418), .B2(n15286), .A(n15287), .ZN(n18412) );
  AOI21_X1 U17302 ( .B1(n17406), .B2(n15282), .A(n11015), .ZN(n17396) );
  OAI22_X1 U17303 ( .A1(n18711), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n15283) );
  INV_X1 U17304 ( .A(n15283), .ZN(n18384) );
  AOI22_X1 U17305 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15284), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18711), .ZN(n16456) );
  NOR2_X1 U17306 ( .A1(n18384), .A2(n16456), .ZN(n16455) );
  OAI21_X1 U17307 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n15285), .ZN(n15680) );
  NAND2_X1 U17308 ( .A1(n16455), .A2(n15680), .ZN(n15334) );
  NOR2_X1 U17309 ( .A1(n15336), .A2(n15334), .ZN(n18403) );
  NAND2_X1 U17310 ( .A1(n18403), .A2(n18402), .ZN(n15415) );
  NOR2_X1 U17311 ( .A1(n17396), .A2(n15415), .ZN(n15356) );
  OAI21_X1 U17312 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11015), .A(
        n15286), .ZN(n15568) );
  NAND2_X1 U17313 ( .A1(n15356), .A2(n15568), .ZN(n18411) );
  NOR2_X1 U17314 ( .A1(n18412), .A2(n18411), .ZN(n18424) );
  OAI21_X1 U17315 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n15287), .A(
        n15281), .ZN(n18425) );
  NAND2_X1 U17316 ( .A1(n18424), .A2(n18425), .ZN(n15430) );
  NOR2_X1 U17317 ( .A1(n16771), .A2(n15430), .ZN(n15472) );
  NOR2_X1 U17318 ( .A1(n18517), .A2(n15472), .ZN(n15290) );
  OR2_X1 U17319 ( .A1(n15288), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15289) );
  NAND2_X1 U17320 ( .A1(n15470), .A2(n15289), .ZN(n16748) );
  XNOR2_X1 U17321 ( .A(n15290), .B(n16748), .ZN(n15313) );
  AND2_X1 U17322 ( .A1(n18716), .A2(n21597), .ZN(n15293) );
  NAND2_X1 U17323 ( .A1(n19293), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18717) );
  OR3_X1 U17324 ( .A1(n12654), .A2(n18717), .A3(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n18714) );
  NAND3_X1 U17325 ( .A1(n18714), .A2(n18701), .A3(n18680), .ZN(n15292) );
  INV_X1 U17326 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15294) );
  INV_X1 U17327 ( .A(n15293), .ZN(n15300) );
  NAND2_X1 U17328 ( .A1(n15294), .A2(n15300), .ZN(n15296) );
  AOI21_X1 U17329 ( .B1(n12651), .B2(n15296), .A(n15295), .ZN(n15297) );
  INV_X1 U17330 ( .A(n15299), .ZN(n15302) );
  NAND2_X1 U17331 ( .A1(n15300), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15301) );
  AOI22_X1 U17332 ( .A1(n15303), .A2(n18642), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18641), .ZN(n15304) );
  OAI211_X1 U17333 ( .C1(n15305), .C2(n18598), .A(n15304), .B(n18680), .ZN(
        n15306) );
  AOI21_X1 U17334 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n18639), .A(n15306), 
        .ZN(n15311) );
  INV_X1 U17335 ( .A(n15308), .ZN(n15309) );
  XNOR2_X1 U17336 ( .A(n15426), .B(n15309), .ZN(n19207) );
  NAND2_X1 U17337 ( .A1(n18644), .A2(n19207), .ZN(n15310) );
  OAI211_X1 U17338 ( .C1(n18601), .C2(n16972), .A(n15311), .B(n15310), .ZN(
        n15312) );
  AOI21_X1 U17339 ( .B1(n15313), .B2(n18617), .A(n15312), .ZN(n15314) );
  INV_X1 U17340 ( .A(n15314), .ZN(P2_U2845) );
  AND2_X1 U17341 ( .A1(n15316), .A2(n15315), .ZN(n15318) );
  OR2_X1 U17342 ( .A1(n15318), .A2(n15317), .ZN(n18490) );
  INV_X1 U17343 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n18481) );
  MUX2_X1 U17344 ( .A(n18490), .B(n18481), .S(n16513), .Z(n15319) );
  OAI21_X1 U17345 ( .B1(n15320), .B2(n16524), .A(n15319), .ZN(P2_U2871) );
  NOR2_X1 U17346 ( .A1(n18517), .A2(n16455), .ZN(n15321) );
  XNOR2_X1 U17347 ( .A(n15321), .B(n15680), .ZN(n15322) );
  NAND2_X1 U17348 ( .A1(n15322), .A2(n18617), .ZN(n15333) );
  OAI21_X1 U17349 ( .B1(n15325), .B2(n15324), .A(n15323), .ZN(n19578) );
  NAND2_X1 U17350 ( .A1(n19578), .A2(n18644), .ZN(n15328) );
  INV_X1 U17351 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n17480) );
  OAI22_X1 U17352 ( .A1(n11919), .A2(n18598), .B1(n17480), .B2(n18627), .ZN(
        n15326) );
  AOI21_X1 U17353 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18641), .A(
        n15326), .ZN(n15327) );
  OAI211_X1 U17354 ( .C1(n18529), .C2(n15329), .A(n15328), .B(n15327), .ZN(
        n15330) );
  AOI21_X1 U17355 ( .B1(n15331), .B2(n18645), .A(n15330), .ZN(n15332) );
  OAI211_X1 U17356 ( .C1(n18400), .C2(n19579), .A(n15333), .B(n15332), .ZN(
        P2_U2853) );
  NAND2_X1 U17357 ( .A1(n18606), .A2(n15334), .ZN(n15335) );
  XNOR2_X1 U17358 ( .A(n15336), .B(n15335), .ZN(n15337) );
  NAND2_X1 U17359 ( .A1(n15337), .A2(n18617), .ZN(n15346) );
  INV_X1 U17360 ( .A(n19430), .ZN(n19531) );
  OAI22_X1 U17361 ( .A1(n15338), .A2(n18598), .B1(n17482), .B2(n18627), .ZN(
        n15341) );
  NOR2_X1 U17362 ( .A1(n18596), .A2(n15339), .ZN(n15340) );
  AOI211_X1 U17363 ( .C1(n18644), .C2(n19531), .A(n15341), .B(n15340), .ZN(
        n15342) );
  OAI21_X1 U17364 ( .B1(n15343), .B2(n18529), .A(n15342), .ZN(n15344) );
  AOI21_X1 U17365 ( .B1(n14819), .B2(n18645), .A(n15344), .ZN(n15345) );
  OAI211_X1 U17366 ( .C1(n19431), .C2(n18400), .A(n15346), .B(n15345), .ZN(
        P2_U2852) );
  XOR2_X1 U17367 ( .A(n15348), .B(n15347), .Z(n21426) );
  INV_X1 U17368 ( .A(n21426), .ZN(n15378) );
  OR2_X1 U17369 ( .A1(n21731), .A2(BUF1_REG_8__SCAN_IN), .ZN(n15350) );
  INV_X1 U17370 ( .A(DATAI_8_), .ZN(n17325) );
  NAND2_X1 U17371 ( .A1(n16036), .A2(n17325), .ZN(n15349) );
  NAND2_X1 U17372 ( .A1(n15350), .A2(n15349), .ZN(n21684) );
  INV_X1 U17373 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n15351) );
  OAI222_X1 U17374 ( .A1(n16033), .A2(n15378), .B1(n21684), .B2(n16040), .C1(
        n15351), .C2(n16039), .ZN(P1_U2896) );
  NOR2_X1 U17375 ( .A1(n15353), .A2(n15352), .ZN(n15354) );
  NOR2_X1 U17376 ( .A1(n18517), .A2(n15356), .ZN(n15357) );
  XNOR2_X1 U17377 ( .A(n15357), .B(n15568), .ZN(n15358) );
  AOI22_X1 U17378 ( .A1(n18644), .A2(n11076), .B1(n18617), .B2(n15358), .ZN(
        n15365) );
  INV_X1 U17379 ( .A(n17037), .ZN(n15363) );
  INV_X1 U17380 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n15359) );
  OAI21_X1 U17381 ( .B1(n15359), .B2(n18598), .A(n18680), .ZN(n15360) );
  AOI21_X1 U17382 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18641), .A(
        n15360), .ZN(n15361) );
  OAI21_X1 U17383 ( .B1(n18627), .B2(n12688), .A(n15361), .ZN(n15362) );
  AOI21_X1 U17384 ( .B1(n15363), .B2(n18645), .A(n15362), .ZN(n15364) );
  OAI211_X1 U17385 ( .C1(n15366), .C2(n18529), .A(n15365), .B(n15364), .ZN(
        P2_U2849) );
  INV_X1 U17386 ( .A(n15367), .ZN(n15368) );
  OAI21_X1 U17387 ( .B1(n15194), .B2(n15369), .A(n15368), .ZN(n15409) );
  OR2_X1 U17388 ( .A1(n15398), .A2(n15371), .ZN(n15372) );
  NOR2_X1 U17389 ( .A1(n16473), .A2(n12443), .ZN(n15373) );
  AOI21_X1 U17390 ( .B1(n18520), .B2(n16473), .A(n15373), .ZN(n15374) );
  OAI21_X1 U17391 ( .B1(n15409), .B2(n16524), .A(n15374), .ZN(P2_U2869) );
  NOR2_X1 U17392 ( .A1(n15376), .A2(n15375), .ZN(n15377) );
  OR2_X1 U17393 ( .A1(n15386), .A2(n15377), .ZN(n21423) );
  INV_X1 U17394 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21422) );
  OAI222_X1 U17395 ( .A1(n21423), .A2(n19979), .B1(n19989), .B2(n21422), .C1(
        n15965), .C2(n15378), .ZN(P1_U2864) );
  INV_X1 U17396 ( .A(n15381), .ZN(n15382) );
  OAI21_X1 U17397 ( .B1(n15380), .B2(n15383), .A(n15381), .ZN(n15582) );
  OR2_X1 U17398 ( .A1(n15386), .A2(n15385), .ZN(n15387) );
  NAND2_X1 U17399 ( .A1(n15384), .A2(n15387), .ZN(n15559) );
  OAI22_X1 U17400 ( .A1(n15559), .A2(n19979), .B1(n15388), .B2(n19989), .ZN(
        n15389) );
  INV_X1 U17401 ( .A(n15389), .ZN(n15390) );
  OAI21_X1 U17402 ( .B1(n15582), .B2(n15965), .A(n15390), .ZN(P1_U2863) );
  OAI22_X1 U17403 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n11170), .B1(n15559), 
        .B2(n21572), .ZN(n15394) );
  INV_X1 U17404 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21431) );
  INV_X1 U17405 ( .A(n14514), .ZN(n21359) );
  AOI21_X1 U17406 ( .B1(n21528), .B2(n15742), .A(n21359), .ZN(n21429) );
  AOI22_X1 U17407 ( .A1(n21551), .A2(P1_EBX_REG_9__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n21564), .ZN(n15392) );
  NAND2_X1 U17408 ( .A1(n15391), .A2(n14514), .ZN(n21476) );
  OAI211_X1 U17409 ( .C1(n21431), .C2(n21429), .A(n15392), .B(n21476), .ZN(
        n15393) );
  AOI211_X1 U17410 ( .C1(n15579), .C2(n21521), .A(n15394), .B(n15393), .ZN(
        n15395) );
  OAI21_X1 U17411 ( .B1(n15582), .B2(n21553), .A(n15395), .ZN(P1_U2831) );
  NOR2_X1 U17412 ( .A1(n15317), .A2(n15396), .ZN(n15397) );
  OR2_X1 U17413 ( .A1(n15398), .A2(n15397), .ZN(n16898) );
  NOR2_X1 U17414 ( .A1(n16898), .A2(n16513), .ZN(n15399) );
  AOI21_X1 U17415 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n16513), .A(n15399), .ZN(
        n15400) );
  OAI21_X1 U17416 ( .B1(n15401), .B2(n16524), .A(n15400), .ZN(P2_U2870) );
  INV_X1 U17417 ( .A(n19584), .ZN(n15406) );
  OAI21_X1 U17418 ( .B1(n15403), .B2(n15402), .A(n15451), .ZN(n18524) );
  OAI22_X1 U17419 ( .A1(n19688), .A2(n18524), .B1(n15404), .B2(n19686), .ZN(
        n15405) );
  AOI21_X1 U17420 ( .B1(n16574), .B2(n15406), .A(n15405), .ZN(n15408) );
  AOI22_X1 U17421 ( .A1(n19185), .A2(BUF2_REG_18__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15407) );
  OAI211_X1 U17422 ( .C1(n15409), .C2(n19636), .A(n15408), .B(n15407), .ZN(
        P2_U2901) );
  INV_X1 U17423 ( .A(n15410), .ZN(n15411) );
  NAND2_X1 U17424 ( .A1(n15412), .A2(n15411), .ZN(n15413) );
  AND2_X1 U17425 ( .A1(n15414), .A2(n15413), .ZN(n19420) );
  NAND2_X1 U17426 ( .A1(n18606), .A2(n15415), .ZN(n15416) );
  XNOR2_X1 U17427 ( .A(n17396), .B(n15416), .ZN(n15417) );
  AOI22_X1 U17428 ( .A1(n18644), .A2(n19420), .B1(n18617), .B2(n15417), .ZN(
        n15423) );
  INV_X1 U17429 ( .A(n17402), .ZN(n18684) );
  OAI21_X1 U17430 ( .B1(n15418), .B2(n18598), .A(n18680), .ZN(n15419) );
  AOI21_X1 U17431 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18641), .A(
        n15419), .ZN(n15420) );
  OAI21_X1 U17432 ( .B1(n18627), .B2(n12270), .A(n15420), .ZN(n15421) );
  AOI21_X1 U17433 ( .B1(n18684), .B2(n18645), .A(n15421), .ZN(n15422) );
  OAI211_X1 U17434 ( .C1(n15424), .C2(n18529), .A(n15423), .B(n15422), .ZN(
        P2_U2850) );
  OAI21_X1 U17435 ( .B1(n15425), .B2(n15427), .A(n15426), .ZN(n15428) );
  INV_X1 U17436 ( .A(n15428), .ZN(n19212) );
  NAND2_X1 U17437 ( .A1(n15429), .A2(n15430), .ZN(n15431) );
  XNOR2_X1 U17438 ( .A(n16771), .B(n15431), .ZN(n15432) );
  AOI22_X1 U17439 ( .A1(n19212), .A2(n18644), .B1(n18617), .B2(n15432), .ZN(
        n15438) );
  AOI22_X1 U17440 ( .A1(n15433), .A2(n18642), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18641), .ZN(n15434) );
  OAI211_X1 U17441 ( .C1(n15435), .C2(n18598), .A(n15434), .B(n18680), .ZN(
        n15436) );
  AOI21_X1 U17442 ( .B1(P2_REIP_REG_9__SCAN_IN), .B2(n18639), .A(n15436), .ZN(
        n15437) );
  OAI211_X1 U17443 ( .C1(n16986), .C2(n18601), .A(n15438), .B(n15437), .ZN(
        P2_U2846) );
  NOR2_X1 U17444 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17071) );
  INV_X1 U17445 ( .A(n18706), .ZN(n17060) );
  AOI22_X1 U17446 ( .A1(n18517), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18384), .B2(n15429), .ZN(n17058) );
  AOI222_X1 U17447 ( .A1(n15439), .A2(n17071), .B1(n17060), .B2(n19694), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n17058), .ZN(n15446) );
  NAND2_X1 U17448 ( .A1(n15441), .A2(n15440), .ZN(n15444) );
  NOR2_X1 U17449 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12654), .ZN(n15442) );
  AOI21_X1 U17450 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17136), .A(n15442), .ZN(
        n15443) );
  NAND2_X1 U17451 ( .A1(n15444), .A2(n15443), .ZN(n18661) );
  INV_X1 U17452 ( .A(n18661), .ZN(n17063) );
  NAND2_X1 U17453 ( .A1(n17063), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15445) );
  OAI21_X1 U17454 ( .B1(n15446), .B2(n17063), .A(n15445), .ZN(P2_U3601) );
  OR2_X1 U17455 ( .A1(n21731), .A2(BUF1_REG_9__SCAN_IN), .ZN(n15448) );
  INV_X1 U17456 ( .A(DATAI_9_), .ZN(n17326) );
  NAND2_X1 U17457 ( .A1(n16036), .A2(n17326), .ZN(n15447) );
  NAND2_X1 U17458 ( .A1(n15448), .A2(n15447), .ZN(n21689) );
  INV_X1 U17459 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n15449) );
  OAI222_X1 U17460 ( .A1(n16033), .A2(n15582), .B1(n21689), .B2(n16040), .C1(
        n15449), .C2(n16039), .ZN(P1_U2895) );
  OAI21_X1 U17461 ( .B1(n15367), .B2(n15450), .A(n15493), .ZN(n15492) );
  INV_X1 U17462 ( .A(n19538), .ZN(n15454) );
  XNOR2_X1 U17463 ( .A(n11405), .B(n15451), .ZN(n16878) );
  INV_X1 U17464 ( .A(n16878), .ZN(n18533) );
  OAI22_X1 U17465 ( .A1(n19688), .A2(n18533), .B1(n15452), .B2(n19686), .ZN(
        n15453) );
  AOI21_X1 U17466 ( .B1(n16574), .B2(n15454), .A(n15453), .ZN(n15456) );
  AOI22_X1 U17467 ( .A1(n19185), .A2(BUF2_REG_19__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n15455) );
  OAI211_X1 U17468 ( .C1(n15492), .C2(n19636), .A(n15456), .B(n15455), .ZN(
        P2_U2900) );
  NOR2_X1 U17469 ( .A1(n15382), .A2(n15458), .ZN(n15459) );
  INV_X1 U17470 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n15462) );
  OR2_X1 U17471 ( .A1(n21731), .A2(BUF1_REG_10__SCAN_IN), .ZN(n15461) );
  INV_X1 U17472 ( .A(DATAI_10_), .ZN(n17328) );
  NAND2_X1 U17473 ( .A1(n16036), .A2(n17328), .ZN(n15460) );
  NAND2_X1 U17474 ( .A1(n15461), .A2(n15460), .ZN(n21694) );
  OAI222_X1 U17475 ( .A1(n21440), .A2(n16033), .B1(n15462), .B2(n16039), .C1(
        n21694), .C2(n16040), .ZN(P1_U2894) );
  INV_X1 U17476 ( .A(n15463), .ZN(n15487) );
  AOI21_X1 U17477 ( .B1(n15465), .B2(n15464), .A(n11060), .ZN(n19191) );
  INV_X1 U17478 ( .A(n19191), .ZN(n15484) );
  NOR2_X1 U17479 ( .A1(n18701), .A2(n15429), .ZN(n16457) );
  INV_X1 U17480 ( .A(n15466), .ZN(n15482) );
  INV_X1 U17481 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15468) );
  AOI22_X1 U17482 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n18640), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n18639), .ZN(n15467) );
  OAI211_X1 U17483 ( .C1(n15468), .C2(n18596), .A(n18680), .B(n15467), .ZN(
        n15481) );
  NOR2_X1 U17484 ( .A1(n15475), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15469) );
  OR2_X1 U17485 ( .A1(n15477), .A2(n15469), .ZN(n16709) );
  INV_X1 U17486 ( .A(n16709), .ZN(n18459) );
  NAND2_X1 U17487 ( .A1(n15470), .A2(n16735), .ZN(n15471) );
  AND2_X1 U17488 ( .A1(n15474), .A2(n15471), .ZN(n18440) );
  NAND2_X1 U17489 ( .A1(n15472), .A2(n16748), .ZN(n18432) );
  NOR2_X1 U17490 ( .A1(n18440), .A2(n18432), .ZN(n18449) );
  AND2_X1 U17491 ( .A1(n15474), .A2(n15473), .ZN(n15476) );
  OR2_X1 U17492 ( .A1(n15476), .A2(n15475), .ZN(n18450) );
  NAND2_X1 U17493 ( .A1(n18449), .A2(n18450), .ZN(n18457) );
  NOR2_X1 U17494 ( .A1(n18459), .A2(n18457), .ZN(n18473) );
  NOR2_X1 U17495 ( .A1(n15477), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15478) );
  OR2_X1 U17496 ( .A1(n12561), .A2(n15478), .ZN(n18474) );
  NAND2_X1 U17497 ( .A1(n18473), .A2(n18474), .ZN(n15479) );
  NOR2_X1 U17498 ( .A1(n15482), .A2(n15479), .ZN(n18487) );
  NAND2_X1 U17499 ( .A1(n18606), .A2(n18617), .ZN(n18647) );
  AOI211_X1 U17500 ( .C1(n15482), .C2(n15479), .A(n18487), .B(n18647), .ZN(
        n15480) );
  AOI211_X1 U17501 ( .C1(n16457), .C2(n15482), .A(n15481), .B(n15480), .ZN(
        n15483) );
  OAI21_X1 U17502 ( .B1(n15484), .B2(n18638), .A(n15483), .ZN(n15485) );
  AOI21_X1 U17503 ( .B1(n15717), .B2(n18645), .A(n15485), .ZN(n15486) );
  OAI21_X1 U17504 ( .B1(n15487), .B2(n18529), .A(n15486), .ZN(P2_U2840) );
  NAND2_X1 U17505 ( .A1(n15370), .A2(n15488), .ZN(n15489) );
  NAND2_X1 U17506 ( .A1(n15503), .A2(n15489), .ZN(n18534) );
  NOR2_X1 U17507 ( .A1(n18534), .A2(n16513), .ZN(n15490) );
  AOI21_X1 U17508 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n16513), .A(n15490), .ZN(
        n15491) );
  OAI21_X1 U17509 ( .B1(n15492), .B2(n16524), .A(n15491), .ZN(P2_U2868) );
  OAI21_X1 U17510 ( .B1(n13053), .B2(n11412), .A(n15517), .ZN(n15507) );
  AND2_X1 U17511 ( .A1(n15495), .A2(n15494), .ZN(n15496) );
  OR2_X1 U17512 ( .A1(n15496), .A2(n13335), .ZN(n18550) );
  OAI22_X1 U17513 ( .A1(n19688), .A2(n18550), .B1(n19686), .B2(n15497), .ZN(
        n15498) );
  AOI21_X1 U17514 ( .B1(n16574), .B2(n15499), .A(n15498), .ZN(n15501) );
  AOI22_X1 U17515 ( .A1(n19185), .A2(BUF2_REG_20__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n15500) );
  OAI211_X1 U17516 ( .C1(n15507), .C2(n19636), .A(n15501), .B(n15500), .ZN(
        P2_U2899) );
  NAND2_X1 U17517 ( .A1(n15503), .A2(n15502), .ZN(n15504) );
  NAND2_X1 U17518 ( .A1(n15505), .A2(n15504), .ZN(n18542) );
  INV_X1 U17519 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n18539) );
  MUX2_X1 U17520 ( .A(n18542), .B(n18539), .S(n16513), .Z(n15506) );
  OAI21_X1 U17521 ( .B1(n15507), .B2(n16524), .A(n15506), .ZN(P2_U2867) );
  OR2_X1 U17522 ( .A1(n15457), .A2(n15509), .ZN(n15510) );
  NAND2_X1 U17523 ( .A1(n10984), .A2(n15510), .ZN(n15584) );
  INV_X1 U17524 ( .A(n15511), .ZN(n15583) );
  XNOR2_X1 U17525 ( .A(n15584), .B(n15583), .ZN(n21447) );
  NAND2_X1 U17526 ( .A1(n16353), .A2(n15512), .ZN(n15513) );
  NAND2_X1 U17527 ( .A1(n16331), .A2(n15513), .ZN(n21446) );
  OAI22_X1 U17528 ( .A1(n21446), .A2(n19979), .B1(n15514), .B2(n19989), .ZN(
        n15515) );
  INV_X1 U17529 ( .A(n15515), .ZN(n15516) );
  OAI21_X1 U17530 ( .B1(n21447), .B2(n15965), .A(n15516), .ZN(P1_U2861) );
  INV_X1 U17531 ( .A(n15517), .ZN(n15521) );
  INV_X1 U17532 ( .A(n15518), .ZN(n15520) );
  INV_X1 U17533 ( .A(n15519), .ZN(n16516) );
  OAI21_X1 U17534 ( .B1(n15521), .B2(n15520), .A(n16516), .ZN(n15575) );
  INV_X1 U17535 ( .A(n16448), .ZN(n15524) );
  OAI22_X1 U17536 ( .A1(n19189), .A2(n19436), .B1(n15522), .B2(n19686), .ZN(
        n15523) );
  AOI21_X1 U17537 ( .B1(n19633), .B2(n15524), .A(n15523), .ZN(n15526) );
  AOI22_X1 U17538 ( .A1(n19185), .A2(BUF2_REG_21__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n15525) );
  OAI211_X1 U17539 ( .C1(n15575), .C2(n19636), .A(n15526), .B(n15525), .ZN(
        P2_U2898) );
  INV_X1 U17540 ( .A(n15528), .ZN(n15529) );
  AOI21_X1 U17541 ( .B1(n15530), .B2(n15527), .A(n15529), .ZN(n15547) );
  NAND2_X1 U17542 ( .A1(n20033), .A2(n21425), .ZN(n15531) );
  NAND2_X1 U17543 ( .A1(n21348), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n15541) );
  OAI211_X1 U17544 ( .C1(n16164), .C2(n15532), .A(n15531), .B(n15541), .ZN(
        n15533) );
  AOI21_X1 U17545 ( .B1(n21426), .B2(n21732), .A(n15533), .ZN(n15534) );
  OAI21_X1 U17546 ( .B1(n15547), .B2(n21574), .A(n15534), .ZN(P1_U2991) );
  NAND2_X1 U17547 ( .A1(n21302), .A2(n15535), .ZN(n15537) );
  INV_X1 U17548 ( .A(n15538), .ZN(n15556) );
  NAND3_X1 U17549 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21337), .A3(
        n21319), .ZN(n21334) );
  INV_X1 U17550 ( .A(n21284), .ZN(n16284) );
  AOI21_X1 U17551 ( .B1(n21299), .B2(n15555), .A(n16284), .ZN(n15557) );
  NAND3_X1 U17552 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15557), .A3(
        n15538), .ZN(n15539) );
  NAND2_X1 U17553 ( .A1(n16328), .A2(n21284), .ZN(n16240) );
  NAND2_X1 U17554 ( .A1(n15539), .A2(n16240), .ZN(n21336) );
  INV_X1 U17555 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15540) );
  AOI21_X1 U17556 ( .B1(n21334), .B2(n21336), .A(n15540), .ZN(n15545) );
  INV_X1 U17557 ( .A(n15541), .ZN(n15544) );
  NOR2_X1 U17558 ( .A1(n21423), .A2(n21338), .ZN(n15543) );
  INV_X1 U17559 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21323) );
  NOR4_X1 U17560 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16358), .A3(
        n21337), .A4(n21323), .ZN(n15542) );
  NOR4_X1 U17561 ( .A1(n15545), .A2(n15544), .A3(n15543), .A4(n15542), .ZN(
        n15546) );
  OAI21_X1 U17562 ( .B1(n15547), .B2(n21339), .A(n15546), .ZN(P1_U3023) );
  OR2_X1 U17563 ( .A1(n16036), .A2(n20071), .ZN(n15549) );
  NAND2_X1 U17564 ( .A1(n16036), .A2(DATAI_11_), .ZN(n15548) );
  AND2_X1 U17565 ( .A1(n15549), .A2(n15548), .ZN(n21699) );
  INV_X1 U17566 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15550) );
  OAI222_X1 U17567 ( .A1(n21447), .A2(n16033), .B1(n21699), .B2(n16040), .C1(
        n15550), .C2(n16039), .ZN(P1_U2893) );
  OAI21_X1 U17568 ( .B1(n15551), .B2(n15553), .A(n10998), .ZN(n15576) );
  INV_X1 U17569 ( .A(n15576), .ZN(n15563) );
  INV_X1 U17570 ( .A(n21302), .ZN(n15554) );
  NOR3_X1 U17571 ( .A1(n15555), .A2(n15554), .A3(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21330) );
  NAND2_X1 U17572 ( .A1(n21305), .A2(n15556), .ZN(n21328) );
  NAND2_X1 U17573 ( .A1(n15557), .A2(n21328), .ZN(n21325) );
  NOR2_X1 U17574 ( .A1(n21330), .A2(n21325), .ZN(n21324) );
  OAI21_X1 U17575 ( .B1(n16328), .B2(n15558), .A(n21324), .ZN(n16354) );
  OAI22_X1 U17576 ( .A1(n15559), .A2(n21338), .B1(n21431), .B2(n21288), .ZN(
        n15561) );
  NOR3_X1 U17577 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16358), .A3(
        n15560), .ZN(n16355) );
  AOI211_X1 U17578 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n16354), .A(
        n15561), .B(n16355), .ZN(n15562) );
  OAI21_X1 U17579 ( .B1(n15563), .B2(n21339), .A(n15562), .ZN(P1_U3022) );
  XNOR2_X1 U17580 ( .A(n11002), .B(n15565), .ZN(n17039) );
  OR2_X1 U17581 ( .A1(n15566), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17036) );
  NAND3_X1 U17582 ( .A1(n17036), .A2(n16766), .A3(n15567), .ZN(n15572) );
  NOR2_X1 U17583 ( .A1(n17410), .A2(n17037), .ZN(n15570) );
  OAI22_X1 U17584 ( .A1(n12688), .A2(n18680), .B1(n16782), .B2(n15568), .ZN(
        n15569) );
  AOI211_X1 U17585 ( .C1(n16750), .C2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n15570), .B(n15569), .ZN(n15571) );
  OAI211_X1 U17586 ( .C1(n17411), .C2(n17039), .A(n15572), .B(n15571), .ZN(
        P2_U3008) );
  NAND2_X1 U17587 ( .A1(n16513), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15574) );
  NAND2_X1 U17588 ( .A1(n16451), .A2(n16473), .ZN(n15573) );
  OAI211_X1 U17589 ( .C1(n15575), .C2(n16524), .A(n15574), .B(n15573), .ZN(
        P2_U2866) );
  NAND2_X1 U17590 ( .A1(n15576), .A2(n20039), .ZN(n15581) );
  INV_X1 U17591 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15577) );
  OAI22_X1 U17592 ( .A1(n16164), .A2(n15577), .B1(n21288), .B2(n21431), .ZN(
        n15578) );
  AOI21_X1 U17593 ( .B1(n20033), .B2(n15579), .A(n15578), .ZN(n15580) );
  OAI211_X1 U17594 ( .C1(n20022), .C2(n15582), .A(n15581), .B(n15580), .ZN(
        P1_U2990) );
  OAI21_X1 U17595 ( .B1(n15584), .B2(n15583), .A(n10984), .ZN(n15592) );
  AND2_X1 U17596 ( .A1(n15592), .A2(n15591), .ZN(n15594) );
  NAND2_X1 U17597 ( .A1(n15586), .A2(n15585), .ZN(n15599) );
  OAI21_X1 U17598 ( .B1(n15594), .B2(n15587), .A(n15599), .ZN(n16165) );
  OR2_X1 U17599 ( .A1(n16036), .A2(n20075), .ZN(n15589) );
  NAND2_X1 U17600 ( .A1(n21731), .A2(DATAI_13_), .ZN(n15588) );
  AND2_X1 U17601 ( .A1(n15589), .A2(n15588), .ZN(n21709) );
  INV_X1 U17602 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n15590) );
  OAI222_X1 U17603 ( .A1(n16033), .A2(n16165), .B1(n21709), .B2(n16040), .C1(
        n15590), .C2(n16039), .ZN(P1_U2891) );
  NOR2_X1 U17604 ( .A1(n15592), .A2(n15591), .ZN(n15593) );
  INV_X1 U17605 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15597) );
  OR2_X1 U17606 ( .A1(n16036), .A2(BUF1_REG_12__SCAN_IN), .ZN(n15596) );
  INV_X1 U17607 ( .A(DATAI_12_), .ZN(n17322) );
  NAND2_X1 U17608 ( .A1(n16036), .A2(n17322), .ZN(n15595) );
  NAND2_X1 U17609 ( .A1(n15596), .A2(n15595), .ZN(n21704) );
  OAI222_X1 U17610 ( .A1(n21464), .A2(n16033), .B1(n15597), .B2(n16039), .C1(
        n21704), .C2(n16040), .ZN(P1_U2892) );
  INV_X1 U17611 ( .A(n15970), .ZN(n15598) );
  AOI21_X1 U17612 ( .B1(n15600), .B2(n15599), .A(n15598), .ZN(n16155) );
  INV_X1 U17613 ( .A(n16155), .ZN(n15622) );
  NAND2_X1 U17614 ( .A1(n15738), .A2(n15601), .ZN(n15602) );
  AND2_X1 U17615 ( .A1(n15974), .A2(n15602), .ZN(n21273) );
  AOI22_X1 U17616 ( .A1(n21273), .A2(n19985), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n17196), .ZN(n15603) );
  OAI21_X1 U17617 ( .B1(n15622), .B2(n15965), .A(n15603), .ZN(P1_U2858) );
  NAND2_X1 U17618 ( .A1(n21475), .A2(n21567), .ZN(n21473) );
  INV_X1 U17619 ( .A(n21473), .ZN(n15604) );
  OAI21_X1 U17620 ( .B1(n15605), .B2(P1_REIP_REG_14__SCAN_IN), .A(n15604), 
        .ZN(n15611) );
  INV_X1 U17621 ( .A(n16153), .ZN(n15609) );
  AOI22_X1 U17622 ( .A1(n21273), .A2(n21519), .B1(n21551), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n15606) );
  OAI211_X1 U17623 ( .C1(n21546), .C2(n15607), .A(n15606), .B(n21476), .ZN(
        n15608) );
  AOI21_X1 U17624 ( .B1(n21521), .B2(n15609), .A(n15608), .ZN(n15610) );
  OAI211_X1 U17625 ( .C1(n15622), .C2(n21553), .A(n15611), .B(n15610), .ZN(
        P1_U2826) );
  INV_X1 U17626 ( .A(n15957), .ZN(n15613) );
  OAI21_X1 U17627 ( .B1(n15614), .B2(n15612), .A(n15613), .ZN(n21479) );
  NAND2_X1 U17628 ( .A1(n15616), .A2(n21731), .ZN(n15658) );
  OAI22_X1 U17629 ( .A1(n16027), .A2(n21976), .B1(n16039), .B2(n14801), .ZN(
        n15615) );
  AOI21_X1 U17630 ( .B1(n16029), .B2(DATAI_18_), .A(n15615), .ZN(n15618) );
  NAND2_X1 U17631 ( .A1(n16030), .A2(BUF1_REG_18__SCAN_IN), .ZN(n15617) );
  OAI211_X1 U17632 ( .C1(n21479), .C2(n16033), .A(n15618), .B(n15617), .ZN(
        P1_U2886) );
  INV_X1 U17633 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20077) );
  OR2_X1 U17634 ( .A1(n16036), .A2(n20077), .ZN(n15620) );
  NAND2_X1 U17635 ( .A1(n21731), .A2(DATAI_14_), .ZN(n15619) );
  AND2_X1 U17636 ( .A1(n15620), .A2(n15619), .ZN(n21714) );
  INV_X1 U17637 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n15621) );
  OAI222_X1 U17638 ( .A1(n16033), .A2(n15622), .B1(n21714), .B2(n16040), .C1(
        n15621), .C2(n16039), .ZN(P1_U2890) );
  INV_X1 U17639 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17532) );
  NAND2_X1 U17640 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .ZN(n17534) );
  AND3_X1 U17641 ( .A1(n20768), .A2(n18916), .A3(n15624), .ZN(n15625) );
  INV_X1 U17642 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n20207) );
  NAND3_X1 U17643 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n17501) );
  NOR3_X1 U17644 ( .A1(n20207), .A2(n20189), .A3(n17501), .ZN(n17635) );
  NAND3_X1 U17645 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17874), .A3(n17635), .ZN(
        n17524) );
  NOR2_X1 U17646 ( .A1(n17534), .A2(n17524), .ZN(n17633) );
  NAND3_X1 U17647 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n17633), .ZN(n17632) );
  NOR2_X1 U17648 ( .A1(n17532), .A2(n17632), .ZN(n17619) );
  INV_X1 U17649 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17531) );
  NOR2_X1 U17650 ( .A1(n20274), .A2(n17531), .ZN(n15626) );
  NOR2_X1 U17651 ( .A1(n20622), .A2(n17524), .ZN(n17536) );
  INV_X1 U17652 ( .A(n17536), .ZN(n17527) );
  NOR2_X1 U17653 ( .A1(n17534), .A2(n17527), .ZN(n17519) );
  AOI21_X1 U17654 ( .B1(n15626), .B2(n17519), .A(P3_EBX_REG_10__SCAN_IN), .ZN(
        n15627) );
  NOR2_X1 U17655 ( .A1(n17619), .A2(n15627), .ZN(n15639) );
  AOI22_X1 U17656 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15631) );
  AOI22_X1 U17657 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15630) );
  AOI22_X1 U17658 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15629) );
  AOI22_X1 U17659 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15628) );
  NAND4_X1 U17660 ( .A1(n15631), .A2(n15630), .A3(n15629), .A4(n15628), .ZN(
        n15637) );
  AOI22_X1 U17661 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15635) );
  AOI22_X1 U17662 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15634) );
  AOI22_X1 U17663 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15633) );
  BUF_X1 U17664 ( .A(n17838), .Z(n17860) );
  AOI22_X1 U17665 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15632) );
  NAND4_X1 U17666 ( .A1(n15635), .A2(n15634), .A3(n15633), .A4(n15632), .ZN(
        n15636) );
  NOR2_X1 U17667 ( .A1(n15637), .A2(n15636), .ZN(n20613) );
  INV_X1 U17668 ( .A(n20613), .ZN(n15638) );
  INV_X1 U17669 ( .A(n17874), .ZN(n17877) );
  MUX2_X1 U17670 ( .A(n15639), .B(n15638), .S(n17878), .Z(P3_U2693) );
  INV_X1 U17671 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n20198) );
  OAI21_X1 U17672 ( .B1(n15640), .B2(n11420), .A(n20198), .ZN(n17115) );
  NAND2_X1 U17673 ( .A1(n15641), .A2(n17115), .ZN(n21230) );
  INV_X1 U17674 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20789) );
  NAND2_X1 U17675 ( .A1(n20789), .A2(n21246), .ZN(n20808) );
  NOR2_X1 U17676 ( .A1(n21230), .A2(n20808), .ZN(n15647) );
  OAI21_X1 U17677 ( .B1(n17125), .B2(n20105), .A(n20598), .ZN(n15644) );
  INV_X1 U17678 ( .A(n21234), .ZN(n21217) );
  NOR2_X1 U17679 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21246), .ZN(n18752) );
  INV_X1 U17680 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21260) );
  NOR2_X1 U17681 ( .A1(n20789), .A2(n17117), .ZN(n17885) );
  NAND2_X1 U17682 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n17885), .ZN(n21244) );
  NOR2_X1 U17683 ( .A1(n21260), .A2(n21244), .ZN(n15646) );
  MUX2_X1 U17684 ( .A(n15647), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n20833), .Z(P3_U3284) );
  AOI21_X1 U17685 ( .B1(n15648), .B2(n15832), .A(n15729), .ZN(n15822) );
  AOI21_X1 U17686 ( .B1(n20038), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15649), .ZN(n15650) );
  OAI21_X1 U17687 ( .B1(n20043), .B2(n15823), .A(n15650), .ZN(n15651) );
  AOI21_X1 U17688 ( .B1(n15822), .B2(n21732), .A(n15651), .ZN(n15652) );
  OAI21_X1 U17689 ( .B1(n15653), .B2(n21574), .A(n15652), .ZN(P1_U2970) );
  INV_X1 U17690 ( .A(DATAI_31_), .ZN(n22213) );
  NAND3_X1 U17691 ( .A1(n15654), .A2(n13429), .A3(n16039), .ZN(n15657) );
  AOI22_X1 U17692 ( .A1(n16030), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n15655), .ZN(n15656) );
  OAI211_X1 U17693 ( .C1(n15658), .C2(n22213), .A(n15657), .B(n15656), .ZN(
        P1_U2873) );
  AOI21_X1 U17694 ( .B1(n15660), .B2(n15659), .A(n17005), .ZN(n15661) );
  INV_X1 U17695 ( .A(n15661), .ZN(n15675) );
  XOR2_X1 U17696 ( .A(n15663), .B(n15662), .Z(n15683) );
  INV_X1 U17697 ( .A(n15664), .ZN(n15665) );
  NAND2_X1 U17698 ( .A1(n15666), .A2(n15665), .ZN(n15676) );
  NAND3_X1 U17699 ( .A1(n15725), .A2(n15677), .A3(n15676), .ZN(n15667) );
  NAND2_X1 U17700 ( .A1(n18500), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n15679) );
  OAI211_X1 U17701 ( .C1(n15668), .C2(n17052), .A(n15667), .B(n15679), .ZN(
        n15673) );
  INV_X1 U17702 ( .A(n19578), .ZN(n15669) );
  OAI22_X1 U17703 ( .A1(n15671), .A2(n15670), .B1(n15669), .B2(n18662), .ZN(
        n15672) );
  AOI211_X1 U17704 ( .C1(n15683), .C2(n13329), .A(n15673), .B(n15672), .ZN(
        n15674) );
  OAI211_X1 U17705 ( .C1(n18666), .C2(n11943), .A(n15675), .B(n15674), .ZN(
        P2_U3044) );
  AND3_X1 U17706 ( .A1(n15677), .A2(n16766), .A3(n15676), .ZN(n15682) );
  NAND2_X1 U17707 ( .A1(n16750), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15678) );
  OAI211_X1 U17708 ( .C1(n16782), .C2(n15680), .A(n15679), .B(n15678), .ZN(
        n15681) );
  AOI211_X1 U17709 ( .C1(n15683), .C2(n12546), .A(n15682), .B(n15681), .ZN(
        n15684) );
  OAI21_X1 U17710 ( .B1(n11943), .B2(n17410), .A(n15684), .ZN(P2_U3012) );
  AOI21_X1 U17711 ( .B1(n17152), .B2(n16385), .A(n16393), .ZN(n15688) );
  OAI22_X1 U17712 ( .A1(n15685), .A2(n16375), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13490), .ZN(n17153) );
  OAI22_X1 U17713 ( .A1(n16379), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16380), .ZN(n15686) );
  AOI21_X1 U17714 ( .B1(n17153), .B2(n16385), .A(n15686), .ZN(n15687) );
  OAI22_X1 U17715 ( .A1(n15688), .A2(n13797), .B1(n16393), .B2(n15687), .ZN(
        P1_U3474) );
  NAND2_X1 U17716 ( .A1(n18688), .A2(n17005), .ZN(n16906) );
  AND3_X1 U17717 ( .A1(n15689), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n16856), .ZN(n15692) );
  NOR2_X1 U17718 ( .A1(n17005), .A2(n15689), .ZN(n15690) );
  NOR2_X1 U17719 ( .A1(n15691), .A2(n15690), .ZN(n16862) );
  OAI21_X1 U17720 ( .B1(n15692), .B2(n17002), .A(n16862), .ZN(n15722) );
  AOI21_X2 U17721 ( .B1(n16676), .B2(n16906), .A(n15722), .ZN(n16909) );
  INV_X1 U17722 ( .A(n16684), .ZN(n15694) );
  OAI22_X2 U17723 ( .A1(n15694), .A2(n18688), .B1(n15693), .B2(n16855), .ZN(
        n16897) );
  NAND2_X1 U17724 ( .A1(n16897), .A2(n16905), .ZN(n15701) );
  INV_X1 U17725 ( .A(n16673), .ZN(n15695) );
  AOI21_X1 U17726 ( .B1(n15697), .B2(n15696), .A(n15695), .ZN(n16689) );
  NOR2_X1 U17727 ( .A1(n18490), .A2(n18666), .ZN(n15699) );
  NAND2_X1 U17728 ( .A1(n18500), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16686) );
  OAI21_X1 U17729 ( .B1(n18495), .B2(n18662), .A(n16686), .ZN(n15698) );
  AOI211_X1 U17730 ( .C1(n16689), .C2(n13329), .A(n15699), .B(n15698), .ZN(
        n15700) );
  OAI211_X1 U17731 ( .C1(n16909), .C2(n16905), .A(n15701), .B(n15700), .ZN(
        P2_U3030) );
  INV_X1 U17732 ( .A(n18624), .ZN(n15711) );
  NAND3_X1 U17733 ( .A1(n15705), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15704), .ZN(n15708) );
  INV_X1 U17734 ( .A(n15706), .ZN(n15707) );
  OAI21_X1 U17735 ( .B1(n15711), .B2(n18666), .A(n15710), .ZN(n15712) );
  AOI21_X1 U17736 ( .B1(n15713), .B2(n15725), .A(n15712), .ZN(n15714) );
  OAI21_X1 U17737 ( .B1(n15715), .B2(n18664), .A(n15714), .ZN(P2_U3016) );
  INV_X1 U17738 ( .A(n15716), .ZN(n15726) );
  NAND2_X1 U17739 ( .A1(n15717), .A2(n18685), .ZN(n15721) );
  INV_X1 U17740 ( .A(n15718), .ZN(n15719) );
  AOI21_X1 U17741 ( .B1(n19191), .B2(n12928), .A(n15719), .ZN(n15720) );
  OAI211_X1 U17742 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16855), .A(
        n15721), .B(n15720), .ZN(n15723) );
  OR2_X1 U17743 ( .A1(n15723), .A2(n11396), .ZN(n15724) );
  AOI21_X1 U17744 ( .B1(n15726), .B2(n15725), .A(n15724), .ZN(n15727) );
  OAI21_X1 U17745 ( .B1(n18664), .B2(n15728), .A(n15727), .ZN(P2_U3031) );
  INV_X1 U17746 ( .A(n16055), .ZN(n15983) );
  INV_X1 U17747 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n15737) );
  INV_X1 U17748 ( .A(n15731), .ZN(n15732) );
  AOI22_X1 U17749 ( .A1(n15734), .A2(n15733), .B1(n15732), .B2(n15836), .ZN(
        n15736) );
  OAI222_X1 U17750 ( .A1(n15983), .A2(n15965), .B1(n15737), .B2(n19989), .C1(
        n19979), .C2(n16170), .ZN(P1_U2842) );
  OAI21_X1 U17751 ( .B1(n16333), .B2(n15739), .A(n15738), .ZN(n16315) );
  INV_X1 U17752 ( .A(n16315), .ZN(n15740) );
  AOI22_X1 U17753 ( .A1(n15740), .A2(n19985), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n17196), .ZN(n15741) );
  OAI21_X1 U17754 ( .B1(n16165), .B2(n15965), .A(n15741), .ZN(P1_U2859) );
  INV_X1 U17755 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21435) );
  NOR4_X1 U17756 ( .A1(n21359), .A2(n21435), .A3(n21431), .A4(n15742), .ZN(
        n21434) );
  NAND3_X1 U17757 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(n21434), .ZN(n15743) );
  NAND2_X1 U17758 ( .A1(n21567), .A2(n15743), .ZN(n21457) );
  INV_X1 U17759 ( .A(n21551), .ZN(n21562) );
  OAI22_X1 U17760 ( .A1(n16315), .A2(n21572), .B1(n15744), .B2(n21562), .ZN(
        n15745) );
  AOI211_X1 U17761 ( .C1(n21564), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n21492), .B(n15745), .ZN(n15746) );
  OAI221_X1 U17762 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15747), .C1(n19922), 
        .C2(n21457), .A(n15746), .ZN(n15748) );
  AOI21_X1 U17763 ( .B1(n21521), .B2(n16168), .A(n15748), .ZN(n15749) );
  OAI21_X1 U17764 ( .B1(n16165), .B2(n21553), .A(n15749), .ZN(P1_U2827) );
  AND2_X1 U17765 ( .A1(n16416), .A2(n15750), .ZN(n15751) );
  OR2_X1 U17766 ( .A1(n15751), .A2(n11016), .ZN(n18608) );
  NOR2_X1 U17767 ( .A1(n16782), .A2(n18608), .ZN(n15752) );
  AOI211_X1 U17768 ( .C1(n16750), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15753), .B(n15752), .ZN(n15754) );
  OAI21_X1 U17769 ( .B1(n18602), .B2(n17410), .A(n15754), .ZN(n15755) );
  AOI21_X1 U17770 ( .B1(n15756), .B2(n16766), .A(n15755), .ZN(n15757) );
  OAI21_X1 U17771 ( .B1(n15758), .B2(n17411), .A(n15757), .ZN(P2_U2986) );
  NAND2_X1 U17772 ( .A1(n16750), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15759) );
  OAI211_X1 U17773 ( .C1(n16782), .C2(n15761), .A(n15760), .B(n15759), .ZN(
        n15762) );
  INV_X1 U17774 ( .A(n15762), .ZN(n15763) );
  OAI21_X1 U17775 ( .B1(n16472), .B2(n17410), .A(n15763), .ZN(n15764) );
  AOI21_X1 U17776 ( .B1(n15765), .B2(n16766), .A(n15764), .ZN(n15766) );
  OAI21_X1 U17777 ( .B1(n15767), .B2(n17411), .A(n15766), .ZN(P2_U2983) );
  NOR2_X1 U17778 ( .A1(n18613), .A2(n16513), .ZN(n15768) );
  AOI21_X1 U17779 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n16513), .A(n15768), .ZN(
        n15769) );
  OAI21_X1 U17780 ( .B1(n15770), .B2(n16524), .A(n15769), .ZN(P2_U2858) );
  NAND2_X1 U17781 ( .A1(n15772), .A2(n15771), .ZN(n15775) );
  INV_X1 U17782 ( .A(n15773), .ZN(n15774) );
  NAND2_X1 U17783 ( .A1(n15775), .A2(n15774), .ZN(n15802) );
  AOI22_X1 U17784 ( .A1(n10966), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11975), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15779) );
  AOI22_X1 U17785 ( .A1(n15777), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10964), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15778) );
  NAND2_X1 U17786 ( .A1(n15779), .A2(n15778), .ZN(n15799) );
  AOI22_X1 U17787 ( .A1(n15780), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11842), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15782) );
  AOI21_X1 U17788 ( .B1(n15792), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n15784), .ZN(n15781) );
  OAI211_X1 U17789 ( .C1(n15787), .C2(n15783), .A(n15782), .B(n15781), .ZN(
        n15798) );
  INV_X1 U17790 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17112) );
  OAI21_X1 U17791 ( .B1(n10968), .B2(n17112), .A(n15784), .ZN(n15790) );
  OAI22_X1 U17792 ( .A1(n11793), .A2(n15788), .B1(n15787), .B2(n15786), .ZN(
        n15789) );
  AOI211_X1 U17793 ( .C1(n11975), .C2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n15790), .B(n15789), .ZN(n15796) );
  AOI22_X1 U17794 ( .A1(n15792), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10965), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15795) );
  AOI22_X1 U17795 ( .A1(n11842), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n15776), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15794) );
  NAND3_X1 U17796 ( .A1(n15796), .A2(n15795), .A3(n15794), .ZN(n15797) );
  OAI21_X1 U17797 ( .B1(n15799), .B2(n15798), .A(n15797), .ZN(n15800) );
  INV_X1 U17798 ( .A(n15800), .ZN(n15801) );
  XNOR2_X1 U17799 ( .A(n15802), .B(n15801), .ZN(n15812) );
  OAI22_X1 U17800 ( .A1(n19189), .A2(n19194), .B1(n19686), .B2(n15804), .ZN(
        n15805) );
  AOI21_X1 U17801 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n19184), .A(n15805), .ZN(
        n15807) );
  NAND2_X1 U17802 ( .A1(n19185), .A2(BUF2_REG_30__SCAN_IN), .ZN(n15806) );
  OAI211_X1 U17803 ( .C1(n15803), .C2(n19688), .A(n15807), .B(n15806), .ZN(
        n15808) );
  INV_X1 U17804 ( .A(n15808), .ZN(n15809) );
  OAI21_X1 U17805 ( .B1(n15812), .B2(n19636), .A(n15809), .ZN(P2_U2889) );
  NAND2_X1 U17806 ( .A1(n18624), .A2(n16473), .ZN(n15811) );
  NAND2_X1 U17807 ( .A1(n16513), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15810) );
  OAI211_X1 U17808 ( .C1(n15812), .C2(n16524), .A(n15811), .B(n15810), .ZN(
        P2_U2857) );
  INV_X1 U17809 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n17288) );
  NAND2_X1 U17810 ( .A1(n15813), .A2(n17288), .ZN(n15816) );
  NAND2_X1 U17811 ( .A1(n15814), .A2(n10981), .ZN(n15815) );
  MUX2_X1 U17812 ( .A(n15816), .B(n15815), .S(n21262), .Z(P1_U3487) );
  XNOR2_X1 U17813 ( .A(n15827), .B(P1_REIP_REG_30__SCAN_IN), .ZN(n15820) );
  AOI22_X1 U17814 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n21564), .B1(
        n21521), .B2(n16051), .ZN(n15818) );
  NAND2_X1 U17815 ( .A1(n21551), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n15817) );
  NAND2_X1 U17816 ( .A1(n15818), .A2(n15817), .ZN(n15819) );
  INV_X1 U17817 ( .A(n15822), .ZN(n15987) );
  OAI22_X1 U17818 ( .A1(n15824), .A2(n21546), .B1(n21560), .B2(n15823), .ZN(
        n15826) );
  NOR2_X1 U17819 ( .A1(n15903), .A2(n21572), .ZN(n15825) );
  INV_X1 U17820 ( .A(n21567), .ZN(n21534) );
  NOR2_X1 U17821 ( .A1(n21534), .A2(n19943), .ZN(n15828) );
  OAI21_X1 U17822 ( .B1(n15839), .B2(n15828), .A(n15827), .ZN(n15829) );
  OAI211_X1 U17823 ( .C1(n15987), .C2(n21553), .A(n15830), .B(n15829), .ZN(
        P1_U2811) );
  INV_X1 U17824 ( .A(n15862), .ZN(n15835) );
  AOI21_X1 U17825 ( .B1(n15835), .B2(n15848), .A(n15834), .ZN(n15837) );
  NOR2_X1 U17826 ( .A1(n15837), .A2(n15836), .ZN(n16186) );
  INV_X1 U17827 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n15906) );
  AOI22_X1 U17828 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n21564), .B1(
        n21521), .B2(n16069), .ZN(n15838) );
  OAI21_X1 U17829 ( .B1(n21562), .B2(n15906), .A(n15838), .ZN(n15842) );
  AOI21_X1 U17830 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n21567), .A(n15855), 
        .ZN(n15840) );
  NOR2_X1 U17831 ( .A1(n15840), .A2(n15839), .ZN(n15841) );
  AOI211_X1 U17832 ( .C1(n21519), .C2(n16186), .A(n15842), .B(n15841), .ZN(
        n15843) );
  OAI21_X1 U17833 ( .B1(n16066), .B2(n21553), .A(n15843), .ZN(P1_U2812) );
  AOI21_X1 U17834 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n21567), .A(n15857), 
        .ZN(n15854) );
  AOI21_X1 U17836 ( .B1(n15846), .B2(n15845), .A(n15831), .ZN(n16075) );
  NAND2_X1 U17837 ( .A1(n16075), .A2(n21568), .ZN(n15853) );
  OAI22_X1 U17838 ( .A1(n15847), .A2(n21546), .B1(n21560), .B2(n16073), .ZN(
        n15851) );
  XNOR2_X1 U17839 ( .A(n15862), .B(n15848), .ZN(n16196) );
  INV_X1 U17840 ( .A(n16196), .ZN(n15849) );
  NOR2_X1 U17841 ( .A1(n15849), .A2(n21572), .ZN(n15850) );
  AOI211_X1 U17842 ( .C1(n21551), .C2(P1_EBX_REG_27__SCAN_IN), .A(n15851), .B(
        n15850), .ZN(n15852) );
  OAI211_X1 U17843 ( .C1(n15855), .C2(n15854), .A(n15853), .B(n15852), .ZN(
        P1_U2813) );
  OAI21_X1 U17844 ( .B1(n15909), .B2(n15856), .A(n15845), .ZN(n16084) );
  INV_X1 U17845 ( .A(n15857), .ZN(n15867) );
  INV_X1 U17846 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15859) );
  INV_X1 U17847 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15858) );
  OAI22_X1 U17848 ( .A1(n21565), .A2(n15859), .B1(n21534), .B2(n15858), .ZN(
        n15866) );
  NAND2_X1 U17849 ( .A1(n15913), .A2(n15860), .ZN(n15861) );
  NAND2_X1 U17850 ( .A1(n15862), .A2(n15861), .ZN(n16209) );
  AOI22_X1 U17851 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n21564), .B1(
        n21521), .B2(n16079), .ZN(n15864) );
  NAND2_X1 U17852 ( .A1(n21551), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n15863) );
  OAI211_X1 U17853 ( .C1(n16209), .C2(n21572), .A(n15864), .B(n15863), .ZN(
        n15865) );
  AOI21_X1 U17854 ( .B1(n15867), .B2(n15866), .A(n15865), .ZN(n15868) );
  OAI21_X1 U17855 ( .B1(n16084), .B2(n21553), .A(n15868), .ZN(P1_U2814) );
  NOR2_X1 U17856 ( .A1(n15970), .A2(n15869), .ZN(n15881) );
  INV_X1 U17857 ( .A(n15881), .ZN(n15870) );
  AOI21_X1 U17858 ( .B1(n15871), .B2(n15870), .A(n15612), .ZN(n20034) );
  INV_X1 U17859 ( .A(n20034), .ZN(n16026) );
  XOR2_X1 U17860 ( .A(n15873), .B(n15872), .Z(n19984) );
  AOI22_X1 U17861 ( .A1(n21551), .A2(P1_EBX_REG_17__SCAN_IN), .B1(n21521), 
        .B2(n20032), .ZN(n15874) );
  OAI211_X1 U17862 ( .C1(n21546), .C2(n15875), .A(n15874), .B(n21476), .ZN(
        n15877) );
  AOI211_X1 U17863 ( .C1(n15880), .C2(n19927), .A(n21534), .B(n21483), .ZN(
        n15876) );
  AOI211_X1 U17864 ( .C1(n21519), .C2(n19984), .A(n15877), .B(n15876), .ZN(
        n15878) );
  OAI21_X1 U17865 ( .B1(n16026), .B2(n21553), .A(n15878), .ZN(P1_U2823) );
  AOI21_X1 U17866 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n21567), .A(n15879), 
        .ZN(n15891) );
  INV_X1 U17867 ( .A(n15880), .ZN(n15890) );
  AOI21_X1 U17868 ( .B1(n15968), .B2(n15882), .A(n15881), .ZN(n16144) );
  NAND2_X1 U17869 ( .A1(n16144), .A2(n21568), .ZN(n15889) );
  NOR2_X1 U17870 ( .A1(n15972), .A2(n15883), .ZN(n15884) );
  OR2_X1 U17871 ( .A1(n15872), .A2(n15884), .ZN(n15966) );
  INV_X1 U17872 ( .A(n15966), .ZN(n21344) );
  AOI22_X1 U17873 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n21551), .B1(n21521), 
        .B2(n16140), .ZN(n15885) );
  OAI211_X1 U17874 ( .C1(n21546), .C2(n15886), .A(n15885), .B(n21476), .ZN(
        n15887) );
  AOI21_X1 U17875 ( .B1(n21344), .B2(n21519), .A(n15887), .ZN(n15888) );
  OAI211_X1 U17876 ( .C1(n15891), .C2(n15890), .A(n15889), .B(n15888), .ZN(
        P1_U2824) );
  INV_X1 U17877 ( .A(n15892), .ZN(n15893) );
  NAND2_X1 U17878 ( .A1(n15893), .A2(n21392), .ZN(n15900) );
  NAND2_X1 U17879 ( .A1(n21546), .A2(n21560), .ZN(n15894) );
  AOI22_X1 U17880 ( .A1(n21551), .A2(P1_EBX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n15894), .ZN(n15899) );
  INV_X1 U17881 ( .A(n15895), .ZN(n16364) );
  INV_X1 U17882 ( .A(n21373), .ZN(n15896) );
  AOI22_X1 U17883 ( .A1(n21519), .A2(n16364), .B1(n15896), .B2(n21772), .ZN(
        n15898) );
  NAND2_X1 U17884 ( .A1(n21567), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n15897) );
  NAND4_X1 U17885 ( .A1(n15900), .A2(n15899), .A3(n15898), .A4(n15897), .ZN(
        P1_U2840) );
  INV_X1 U17886 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15901) );
  OAI22_X1 U17887 ( .A1(n15902), .A2(n19979), .B1(n19989), .B2(n15901), .ZN(
        P1_U2841) );
  OAI222_X1 U17888 ( .A1(n15965), .A2(n15987), .B1(n15904), .B2(n19989), .C1(
        n15903), .C2(n19979), .ZN(P1_U2843) );
  INV_X1 U17889 ( .A(n16186), .ZN(n15905) );
  OAI222_X1 U17890 ( .A1(n15965), .A2(n16066), .B1(n15906), .B2(n19989), .C1(
        n15905), .C2(n19979), .ZN(P1_U2844) );
  INV_X1 U17891 ( .A(n16075), .ZN(n15994) );
  AOI22_X1 U17892 ( .A1(n16196), .A2(n19985), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n17196), .ZN(n15907) );
  OAI21_X1 U17893 ( .B1(n15994), .B2(n15965), .A(n15907), .ZN(P1_U2845) );
  INV_X1 U17894 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15908) );
  OAI222_X1 U17895 ( .A1(n15965), .A2(n16084), .B1(n15908), .B2(n19989), .C1(
        n16209), .C2(n19979), .ZN(P1_U2846) );
  AOI21_X1 U17896 ( .B1(n15910), .B2(n15919), .A(n15909), .ZN(n21569) );
  INV_X1 U17897 ( .A(n15965), .ZN(n19986) );
  OR2_X1 U17898 ( .A1(n15920), .A2(n15911), .ZN(n15912) );
  NAND2_X1 U17899 ( .A1(n15913), .A2(n15912), .ZN(n21573) );
  OAI22_X1 U17900 ( .A1(n21573), .A2(n19979), .B1(n21561), .B2(n19989), .ZN(
        n15914) );
  AOI21_X1 U17901 ( .B1(n21569), .B2(n19986), .A(n15914), .ZN(n15915) );
  INV_X1 U17902 ( .A(n15915), .ZN(P1_U2847) );
  NAND2_X1 U17903 ( .A1(n15916), .A2(n15917), .ZN(n15918) );
  NAND2_X1 U17904 ( .A1(n15919), .A2(n15918), .ZN(n21554) );
  INV_X1 U17905 ( .A(n15920), .ZN(n15921) );
  OAI21_X1 U17906 ( .B1(n15922), .B2(n15929), .A(n15921), .ZN(n21548) );
  INV_X1 U17907 ( .A(n21548), .ZN(n15923) );
  AOI22_X1 U17908 ( .A1(n15923), .A2(n19985), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n17196), .ZN(n15924) );
  OAI21_X1 U17909 ( .B1(n21554), .B2(n15965), .A(n15924), .ZN(P1_U2848) );
  OR2_X1 U17910 ( .A1(n15925), .A2(n15926), .ZN(n15927) );
  NAND2_X1 U17911 ( .A1(n15916), .A2(n15927), .ZN(n21538) );
  AND2_X1 U17912 ( .A1(n15937), .A2(n15928), .ZN(n15930) );
  OR2_X1 U17913 ( .A1(n15930), .A2(n15929), .ZN(n21537) );
  INV_X1 U17914 ( .A(n21537), .ZN(n15931) );
  AOI22_X1 U17915 ( .A1(n15931), .A2(n19985), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n17196), .ZN(n15932) );
  OAI21_X1 U17916 ( .B1(n21538), .B2(n15965), .A(n15932), .ZN(P1_U2849) );
  INV_X1 U17918 ( .A(n15925), .ZN(n15935) );
  OAI21_X1 U17919 ( .B1(n15936), .B2(n15934), .A(n15935), .ZN(n21523) );
  INV_X1 U17920 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15940) );
  INV_X1 U17921 ( .A(n15937), .ZN(n15938) );
  AOI21_X1 U17922 ( .B1(n15939), .B2(n15943), .A(n15938), .ZN(n21520) );
  INV_X1 U17923 ( .A(n21520), .ZN(n16248) );
  OAI222_X1 U17924 ( .A1(n15965), .A2(n21523), .B1(n15940), .B2(n19989), .C1(
        n16248), .C2(n19979), .ZN(P1_U2850) );
  AOI21_X1 U17925 ( .B1(n15942), .B2(n15941), .A(n15934), .ZN(n21515) );
  INV_X1 U17926 ( .A(n21515), .ZN(n16015) );
  OAI21_X1 U17927 ( .B1(n15951), .B2(n15944), .A(n15943), .ZN(n21513) );
  INV_X1 U17928 ( .A(n21513), .ZN(n16258) );
  AOI22_X1 U17929 ( .A1(n16258), .A2(n19985), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n17196), .ZN(n15945) );
  OAI21_X1 U17930 ( .B1(n16015), .B2(n15965), .A(n15945), .ZN(P1_U2851) );
  NAND2_X1 U17931 ( .A1(n15946), .A2(n15947), .ZN(n15948) );
  NAND2_X1 U17932 ( .A1(n15941), .A2(n15948), .ZN(n21504) );
  INV_X1 U17933 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15952) );
  NOR2_X1 U17934 ( .A1(n15954), .A2(n15949), .ZN(n15950) );
  OR2_X1 U17935 ( .A1(n15951), .A2(n15950), .ZN(n21503) );
  OAI222_X1 U17936 ( .A1(n15965), .A2(n21504), .B1(n15952), .B2(n19989), .C1(
        n21503), .C2(n19979), .ZN(P1_U2852) );
  AND2_X1 U17937 ( .A1(n15963), .A2(n15953), .ZN(n15955) );
  OR2_X1 U17938 ( .A1(n15955), .A2(n15954), .ZN(n21501) );
  OR2_X1 U17939 ( .A1(n15957), .A2(n15956), .ZN(n15958) );
  OAI222_X1 U17940 ( .A1(n19979), .A2(n21501), .B1(n15959), .B2(n19989), .C1(
        n16022), .C2(n15965), .ZN(P1_U2853) );
  INV_X1 U17941 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15964) );
  NAND2_X1 U17942 ( .A1(n15961), .A2(n15960), .ZN(n15962) );
  NAND2_X1 U17943 ( .A1(n15963), .A2(n15962), .ZN(n21486) );
  OAI222_X1 U17944 ( .A1(n15965), .A2(n21479), .B1(n19989), .B2(n15964), .C1(
        n21486), .C2(n19979), .ZN(P1_U2854) );
  INV_X1 U17945 ( .A(n16144), .ZN(n16034) );
  INV_X1 U17946 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15967) );
  OAI222_X1 U17947 ( .A1(n15965), .A2(n16034), .B1(n15967), .B2(n19989), .C1(
        n15966), .C2(n19979), .ZN(P1_U2856) );
  INV_X1 U17948 ( .A(n15968), .ZN(n15969) );
  AOI21_X1 U17949 ( .B1(n15971), .B2(n15970), .A(n15969), .ZN(n21471) );
  INV_X1 U17950 ( .A(n15972), .ZN(n15976) );
  NAND2_X1 U17951 ( .A1(n15974), .A2(n15973), .ZN(n15975) );
  NAND2_X1 U17952 ( .A1(n15976), .A2(n15975), .ZN(n21469) );
  OAI22_X1 U17953 ( .A1(n21469), .A2(n19979), .B1(n15977), .B2(n19989), .ZN(
        n15978) );
  AOI21_X1 U17954 ( .B1(n21471), .B2(n19986), .A(n15978), .ZN(n15979) );
  INV_X1 U17955 ( .A(n15979), .ZN(P1_U2857) );
  OAI22_X1 U17956 ( .A1(n16027), .A2(n21714), .B1(n16039), .B2(n21716), .ZN(
        n15980) );
  AOI21_X1 U17957 ( .B1(n16029), .B2(DATAI_30_), .A(n15980), .ZN(n15982) );
  NAND2_X1 U17958 ( .A1(n16030), .A2(BUF1_REG_30__SCAN_IN), .ZN(n15981) );
  OAI211_X1 U17959 ( .C1(n15983), .C2(n16033), .A(n15982), .B(n15981), .ZN(
        P1_U2874) );
  OAI22_X1 U17960 ( .A1(n16027), .A2(n21709), .B1(n16039), .B2(n21711), .ZN(
        n15984) );
  AOI21_X1 U17961 ( .B1(n16029), .B2(DATAI_29_), .A(n15984), .ZN(n15986) );
  NAND2_X1 U17962 ( .A1(n16030), .A2(BUF1_REG_29__SCAN_IN), .ZN(n15985) );
  OAI211_X1 U17963 ( .C1(n15987), .C2(n16033), .A(n15986), .B(n15985), .ZN(
        P1_U2875) );
  OAI22_X1 U17964 ( .A1(n16027), .A2(n21704), .B1(n16039), .B2(n21706), .ZN(
        n15988) );
  AOI21_X1 U17965 ( .B1(n16029), .B2(DATAI_28_), .A(n15988), .ZN(n15990) );
  NAND2_X1 U17966 ( .A1(n16030), .A2(BUF1_REG_28__SCAN_IN), .ZN(n15989) );
  OAI211_X1 U17967 ( .C1(n16066), .C2(n16033), .A(n15990), .B(n15989), .ZN(
        P1_U2876) );
  OAI22_X1 U17968 ( .A1(n16027), .A2(n21699), .B1(n16039), .B2(n21701), .ZN(
        n15991) );
  AOI21_X1 U17969 ( .B1(n16029), .B2(DATAI_27_), .A(n15991), .ZN(n15993) );
  NAND2_X1 U17970 ( .A1(n16030), .A2(BUF1_REG_27__SCAN_IN), .ZN(n15992) );
  OAI211_X1 U17971 ( .C1(n15994), .C2(n16033), .A(n15993), .B(n15992), .ZN(
        P1_U2877) );
  OAI22_X1 U17972 ( .A1(n16027), .A2(n21694), .B1(n16039), .B2(n21696), .ZN(
        n15995) );
  AOI21_X1 U17973 ( .B1(n16029), .B2(DATAI_26_), .A(n15995), .ZN(n15997) );
  NAND2_X1 U17974 ( .A1(n16030), .A2(BUF1_REG_26__SCAN_IN), .ZN(n15996) );
  OAI211_X1 U17975 ( .C1(n16084), .C2(n16033), .A(n15997), .B(n15996), .ZN(
        P1_U2878) );
  INV_X1 U17976 ( .A(n21569), .ZN(n16001) );
  OAI22_X1 U17977 ( .A1(n16027), .A2(n21689), .B1(n16039), .B2(n21691), .ZN(
        n15998) );
  AOI21_X1 U17978 ( .B1(n16029), .B2(DATAI_25_), .A(n15998), .ZN(n16000) );
  NAND2_X1 U17979 ( .A1(n16030), .A2(BUF1_REG_25__SCAN_IN), .ZN(n15999) );
  OAI211_X1 U17980 ( .C1(n16001), .C2(n16033), .A(n16000), .B(n15999), .ZN(
        P1_U2879) );
  OAI22_X1 U17981 ( .A1(n16027), .A2(n21684), .B1(n16039), .B2(n21686), .ZN(
        n16002) );
  AOI21_X1 U17982 ( .B1(n16029), .B2(DATAI_24_), .A(n16002), .ZN(n16004) );
  NAND2_X1 U17983 ( .A1(n16030), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16003) );
  OAI211_X1 U17984 ( .C1(n21554), .C2(n16033), .A(n16004), .B(n16003), .ZN(
        P1_U2880) );
  OAI22_X1 U17985 ( .A1(n16027), .A2(n22211), .B1(n16039), .B2(n14698), .ZN(
        n16005) );
  AOI21_X1 U17986 ( .B1(n16029), .B2(DATAI_23_), .A(n16005), .ZN(n16007) );
  NAND2_X1 U17987 ( .A1(n16030), .A2(BUF1_REG_23__SCAN_IN), .ZN(n16006) );
  OAI211_X1 U17988 ( .C1(n21538), .C2(n16033), .A(n16007), .B(n16006), .ZN(
        P1_U2881) );
  INV_X1 U17989 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n16008) );
  OAI22_X1 U17990 ( .A1(n16027), .A2(n22164), .B1(n16039), .B2(n16008), .ZN(
        n16009) );
  AOI21_X1 U17991 ( .B1(n16029), .B2(DATAI_22_), .A(n16009), .ZN(n16011) );
  NAND2_X1 U17992 ( .A1(n16030), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16010) );
  OAI211_X1 U17993 ( .C1(n21523), .C2(n16033), .A(n16011), .B(n16010), .ZN(
        P1_U2882) );
  OAI22_X1 U17994 ( .A1(n16027), .A2(n22114), .B1(n16039), .B2(n14701), .ZN(
        n16012) );
  AOI21_X1 U17995 ( .B1(n16029), .B2(DATAI_21_), .A(n16012), .ZN(n16014) );
  NAND2_X1 U17996 ( .A1(n16030), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16013) );
  OAI211_X1 U17997 ( .C1(n16015), .C2(n16033), .A(n16014), .B(n16013), .ZN(
        P1_U2883) );
  OAI22_X1 U17998 ( .A1(n16027), .A2(n22068), .B1(n16039), .B2(n14793), .ZN(
        n16016) );
  AOI21_X1 U17999 ( .B1(n16029), .B2(DATAI_20_), .A(n16016), .ZN(n16018) );
  NAND2_X1 U18000 ( .A1(n16030), .A2(BUF1_REG_20__SCAN_IN), .ZN(n16017) );
  OAI211_X1 U18001 ( .C1(n21504), .C2(n16033), .A(n16018), .B(n16017), .ZN(
        P1_U2884) );
  OAI22_X1 U18002 ( .A1(n16027), .A2(n22022), .B1(n16039), .B2(n14797), .ZN(
        n16019) );
  AOI21_X1 U18003 ( .B1(n16029), .B2(DATAI_19_), .A(n16019), .ZN(n16021) );
  NAND2_X1 U18004 ( .A1(n16030), .A2(BUF1_REG_19__SCAN_IN), .ZN(n16020) );
  OAI211_X1 U18005 ( .C1(n16022), .C2(n16033), .A(n16021), .B(n16020), .ZN(
        P1_U2885) );
  OAI22_X1 U18006 ( .A1(n16027), .A2(n21933), .B1(n16039), .B2(n14791), .ZN(
        n16023) );
  AOI21_X1 U18007 ( .B1(n16029), .B2(DATAI_17_), .A(n16023), .ZN(n16025) );
  NAND2_X1 U18008 ( .A1(n16030), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16024) );
  OAI211_X1 U18009 ( .C1(n16026), .C2(n16033), .A(n16025), .B(n16024), .ZN(
        P1_U2887) );
  OAI22_X1 U18010 ( .A1(n16027), .A2(n21729), .B1(n16039), .B2(n14789), .ZN(
        n16028) );
  AOI21_X1 U18011 ( .B1(n16029), .B2(DATAI_16_), .A(n16028), .ZN(n16032) );
  NAND2_X1 U18012 ( .A1(n16030), .A2(BUF1_REG_16__SCAN_IN), .ZN(n16031) );
  OAI211_X1 U18013 ( .C1(n16034), .C2(n16033), .A(n16032), .B(n16031), .ZN(
        P1_U2888) );
  INV_X1 U18014 ( .A(n21471), .ZN(n16041) );
  INV_X1 U18015 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16035) );
  OR2_X1 U18016 ( .A1(n16036), .A2(n16035), .ZN(n16038) );
  NAND2_X1 U18017 ( .A1(n21731), .A2(DATAI_15_), .ZN(n16037) );
  AND2_X1 U18018 ( .A1(n16038), .A2(n16037), .ZN(n21725) );
  INV_X1 U18019 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19908) );
  OAI222_X1 U18020 ( .A1(n16033), .A2(n16041), .B1(n16040), .B2(n21725), .C1(
        n16039), .C2(n19908), .ZN(P1_U2889) );
  NOR2_X1 U18021 ( .A1(n16336), .A2(n16180), .ZN(n16048) );
  INV_X1 U18022 ( .A(n16042), .ZN(n16047) );
  INV_X1 U18023 ( .A(n16043), .ZN(n16044) );
  NAND2_X1 U18024 ( .A1(n16045), .A2(n16044), .ZN(n16046) );
  XNOR2_X1 U18025 ( .A(n16050), .B(n16049), .ZN(n16179) );
  INV_X1 U18026 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16053) );
  NAND2_X1 U18027 ( .A1(n20033), .A2(n16051), .ZN(n16052) );
  NAND2_X1 U18028 ( .A1(n21348), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16173) );
  OAI211_X1 U18029 ( .C1(n16053), .C2(n16164), .A(n16052), .B(n16173), .ZN(
        n16054) );
  AOI21_X1 U18030 ( .B1(n16055), .B2(n21732), .A(n16054), .ZN(n16056) );
  OAI21_X1 U18031 ( .B1(n16179), .B2(n21574), .A(n16056), .ZN(P1_U2969) );
  NAND2_X1 U18032 ( .A1(n16102), .A2(n16057), .ZN(n16062) );
  NAND2_X1 U18033 ( .A1(n16062), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16061) );
  NOR2_X1 U18034 ( .A1(n16058), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16059) );
  MUX2_X1 U18035 ( .A(n16059), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n16336), .Z(n16060) );
  OAI211_X1 U18036 ( .C1(n16062), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16061), .B(n16060), .ZN(n16064) );
  XNOR2_X1 U18037 ( .A(n16064), .B(n16063), .ZN(n16188) );
  NAND2_X1 U18038 ( .A1(n21348), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16182) );
  OAI21_X1 U18039 ( .B1(n16164), .B2(n16065), .A(n16182), .ZN(n16068) );
  NOR2_X1 U18040 ( .A1(n16066), .A2(n20022), .ZN(n16067) );
  OAI21_X1 U18041 ( .B1(n21574), .B2(n16188), .A(n16070), .ZN(P1_U2971) );
  XNOR2_X1 U18042 ( .A(n13755), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16071) );
  XNOR2_X1 U18043 ( .A(n16045), .B(n16071), .ZN(n16199) );
  INV_X1 U18044 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n17284) );
  NOR2_X1 U18045 ( .A1(n21288), .A2(n17284), .ZN(n16193) );
  AOI21_X1 U18046 ( .B1(n20038), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16193), .ZN(n16072) );
  OAI21_X1 U18047 ( .B1(n20043), .B2(n16073), .A(n16072), .ZN(n16074) );
  AOI21_X1 U18048 ( .B1(n16075), .B2(n21732), .A(n16074), .ZN(n16076) );
  OAI21_X1 U18049 ( .B1(n16199), .B2(n21574), .A(n16076), .ZN(P1_U2972) );
  NAND2_X1 U18050 ( .A1(n21348), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n16203) );
  OAI21_X1 U18051 ( .B1(n16164), .B2(n16077), .A(n16203), .ZN(n16078) );
  AOI21_X1 U18052 ( .B1(n16079), .B2(n20033), .A(n16078), .ZN(n16083) );
  NAND2_X1 U18053 ( .A1(n16081), .A2(n16202), .ZN(n16200) );
  NAND3_X1 U18054 ( .A1(n16080), .A2(n16200), .A3(n20039), .ZN(n16082) );
  OAI211_X1 U18055 ( .C1(n16084), .C2(n20022), .A(n16083), .B(n16082), .ZN(
        P1_U2973) );
  OAI21_X1 U18056 ( .B1(n16102), .B2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16085), .ZN(n16088) );
  INV_X1 U18057 ( .A(n13759), .ZN(n16086) );
  MUX2_X1 U18058 ( .A(n16232), .B(n16086), .S(n16336), .Z(n16087) );
  NAND2_X1 U18059 ( .A1(n16088), .A2(n16087), .ZN(n16089) );
  XNOR2_X1 U18060 ( .A(n16089), .B(n16212), .ZN(n16217) );
  NAND2_X1 U18061 ( .A1(n21348), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n16211) );
  NAND2_X1 U18062 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16090) );
  OAI211_X1 U18063 ( .C1(n20043), .C2(n21559), .A(n16211), .B(n16090), .ZN(
        n16091) );
  AOI21_X1 U18064 ( .B1(n21569), .B2(n21732), .A(n16091), .ZN(n16092) );
  OAI21_X1 U18065 ( .B1(n21574), .B2(n16217), .A(n16092), .ZN(P1_U2974) );
  NAND2_X1 U18066 ( .A1(n16337), .A2(n16232), .ZN(n16094) );
  NAND3_X1 U18067 ( .A1(n16102), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n13755), .ZN(n16093) );
  OAI21_X1 U18068 ( .B1(n16102), .B2(n16094), .A(n16093), .ZN(n16095) );
  XOR2_X1 U18069 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n16095), .Z(
        n16218) );
  INV_X1 U18070 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n16096) );
  NOR2_X1 U18071 ( .A1(n21288), .A2(n16096), .ZN(n16223) );
  AOI21_X1 U18072 ( .B1(n20038), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16223), .ZN(n16098) );
  NAND2_X1 U18073 ( .A1(n20033), .A2(n21544), .ZN(n16097) );
  OAI211_X1 U18074 ( .C1(n21554), .C2(n20022), .A(n16098), .B(n16097), .ZN(
        n16099) );
  AOI21_X1 U18075 ( .B1(n16218), .B2(n20039), .A(n16099), .ZN(n16100) );
  INV_X1 U18076 ( .A(n16100), .ZN(P1_U2975) );
  XNOR2_X1 U18077 ( .A(n13755), .B(n16232), .ZN(n16101) );
  XNOR2_X1 U18078 ( .A(n16102), .B(n16101), .ZN(n16227) );
  NAND2_X1 U18079 ( .A1(n16227), .A2(n20039), .ZN(n16105) );
  NOR2_X1 U18080 ( .A1(n21288), .A2(n21535), .ZN(n16230) );
  NOR2_X1 U18081 ( .A1(n20043), .A2(n21543), .ZN(n16103) );
  AOI211_X1 U18082 ( .C1(n20038), .C2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16230), .B(n16103), .ZN(n16104) );
  OAI211_X1 U18083 ( .C1(n20022), .C2(n21538), .A(n16105), .B(n16104), .ZN(
        P1_U2976) );
  NAND2_X1 U18084 ( .A1(n16107), .A2(n16106), .ZN(n16108) );
  XOR2_X1 U18085 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n16108), .Z(
        n16252) );
  NAND2_X1 U18086 ( .A1(n21348), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n16247) );
  OAI21_X1 U18087 ( .B1(n16164), .B2(n16109), .A(n16247), .ZN(n16111) );
  NOR2_X1 U18088 ( .A1(n21523), .A2(n20022), .ZN(n16110) );
  AOI211_X1 U18089 ( .C1(n20033), .C2(n21522), .A(n16111), .B(n16110), .ZN(
        n16112) );
  OAI21_X1 U18090 ( .B1(n21574), .B2(n16252), .A(n16112), .ZN(P1_U2977) );
  MUX2_X1 U18091 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n13754), .S(
        n16337), .Z(n16121) );
  MUX2_X1 U18092 ( .A(n16114), .B(n16276), .S(n16122), .Z(n16115) );
  NAND2_X1 U18093 ( .A1(n16121), .A2(n16115), .ZN(n16116) );
  XNOR2_X1 U18094 ( .A(n16116), .B(n16253), .ZN(n16261) );
  NOR2_X1 U18095 ( .A1(n21288), .A2(n21527), .ZN(n16257) );
  NOR2_X1 U18096 ( .A1(n16164), .A2(n16117), .ZN(n16118) );
  AOI211_X1 U18097 ( .C1(n20033), .C2(n21510), .A(n16257), .B(n16118), .ZN(
        n16120) );
  NAND2_X1 U18098 ( .A1(n21515), .A2(n21732), .ZN(n16119) );
  OAI211_X1 U18099 ( .C1(n16261), .C2(n21574), .A(n16120), .B(n16119), .ZN(
        P1_U2978) );
  OAI21_X1 U18100 ( .B1(n16276), .B2(n16114), .A(n16121), .ZN(n16123) );
  XNOR2_X1 U18101 ( .A(n16123), .B(n16122), .ZN(n16270) );
  NAND2_X1 U18102 ( .A1(n21348), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16266) );
  OAI21_X1 U18103 ( .B1(n16164), .B2(n21509), .A(n16266), .ZN(n16125) );
  NOR2_X1 U18104 ( .A1(n21504), .A2(n20022), .ZN(n16124) );
  AOI211_X1 U18105 ( .C1(n20033), .C2(n21502), .A(n16125), .B(n16124), .ZN(
        n16126) );
  OAI21_X1 U18106 ( .B1(n16270), .B2(n21574), .A(n16126), .ZN(P1_U2979) );
  OR2_X1 U18107 ( .A1(n16128), .A2(n16127), .ZN(n16281) );
  NAND3_X1 U18108 ( .A1(n16281), .A2(n20039), .A3(n16129), .ZN(n16132) );
  NAND2_X1 U18109 ( .A1(n21348), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n16288) );
  OAI21_X1 U18110 ( .B1(n16164), .B2(n21478), .A(n16288), .ZN(n16130) );
  AOI21_X1 U18111 ( .B1(n21482), .B2(n20033), .A(n16130), .ZN(n16131) );
  OAI211_X1 U18112 ( .C1(n20022), .C2(n21479), .A(n16132), .B(n16131), .ZN(
        P1_U2981) );
  AND3_X1 U18113 ( .A1(n16149), .A2(n16134), .A3(n16133), .ZN(n16136) );
  OAI211_X1 U18114 ( .C1(n16136), .C2(n16336), .A(n16135), .B(n16157), .ZN(
        n20028) );
  MUX2_X1 U18115 ( .A(n16337), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .S(
        n20028), .Z(n16137) );
  OAI21_X1 U18116 ( .B1(n16138), .B2(n16336), .A(n16137), .ZN(n16139) );
  INV_X1 U18117 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21353) );
  XNOR2_X1 U18118 ( .A(n16139), .B(n21353), .ZN(n21343) );
  INV_X1 U18119 ( .A(n16140), .ZN(n16142) );
  AOI22_X1 U18120 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n21348), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16141) );
  OAI21_X1 U18121 ( .B1(n20043), .B2(n16142), .A(n16141), .ZN(n16143) );
  AOI21_X1 U18122 ( .B1(n16144), .B2(n21732), .A(n16143), .ZN(n16145) );
  OAI21_X1 U18123 ( .B1(n21343), .B2(n21574), .A(n16145), .ZN(P1_U2983) );
  AOI21_X1 U18124 ( .B1(n16146), .B2(n16293), .A(n16147), .ZN(n16148) );
  AOI21_X1 U18125 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16337), .A(
        n16148), .ZN(n16151) );
  MUX2_X1 U18126 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n16149), .S(
        n16336), .Z(n16150) );
  XNOR2_X1 U18127 ( .A(n16151), .B(n16150), .ZN(n21272) );
  AOI22_X1 U18128 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n21348), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16152) );
  OAI21_X1 U18129 ( .B1(n20043), .B2(n16153), .A(n16152), .ZN(n16154) );
  AOI21_X1 U18130 ( .B1(n16155), .B2(n21732), .A(n16154), .ZN(n16156) );
  OAI21_X1 U18131 ( .B1(n21272), .B2(n21574), .A(n16156), .ZN(P1_U2985) );
  OAI21_X1 U18132 ( .B1(n16146), .B2(n16158), .A(n16157), .ZN(n16325) );
  INV_X1 U18133 ( .A(n16159), .ZN(n16160) );
  NOR3_X1 U18134 ( .A1(n16325), .A2(n16321), .A3(n16160), .ZN(n16323) );
  NOR2_X1 U18135 ( .A1(n16323), .A2(n16321), .ZN(n16161) );
  XOR2_X1 U18136 ( .A(n16162), .B(n16161), .Z(n16320) );
  INV_X1 U18137 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16163) );
  NAND2_X1 U18138 ( .A1(n21348), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n16314) );
  OAI21_X1 U18139 ( .B1(n16164), .B2(n16163), .A(n16314), .ZN(n16167) );
  NOR2_X1 U18140 ( .A1(n16165), .A2(n20022), .ZN(n16166) );
  AOI211_X1 U18141 ( .C1(n20033), .C2(n16168), .A(n16167), .B(n16166), .ZN(
        n16169) );
  OAI21_X1 U18142 ( .B1(n16320), .B2(n21574), .A(n16169), .ZN(P1_U2986) );
  INV_X1 U18143 ( .A(n16170), .ZN(n16177) );
  OAI21_X1 U18144 ( .B1(n16172), .B2(n16171), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16174) );
  OAI211_X1 U18145 ( .C1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n16175), .A(
        n16174), .B(n16173), .ZN(n16176) );
  AOI21_X1 U18146 ( .B1(n16177), .B2(n21345), .A(n16176), .ZN(n16178) );
  OAI21_X1 U18147 ( .B1(n16179), .B2(n21339), .A(n16178), .ZN(P1_U3001) );
  NAND2_X1 U18148 ( .A1(n16189), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16184) );
  NAND3_X1 U18149 ( .A1(n16195), .A2(n16181), .A3(n16180), .ZN(n16183) );
  OAI211_X1 U18150 ( .C1(n16184), .C2(n16190), .A(n16183), .B(n16182), .ZN(
        n16185) );
  AOI21_X1 U18151 ( .B1(n16186), .B2(n21345), .A(n16185), .ZN(n16187) );
  OAI21_X1 U18152 ( .B1(n16188), .B2(n21339), .A(n16187), .ZN(P1_U3003) );
  INV_X1 U18153 ( .A(n16189), .ZN(n16191) );
  NOR3_X1 U18154 ( .A1(n16191), .A2(n16190), .A3(n16194), .ZN(n16192) );
  AOI211_X1 U18155 ( .C1(n16195), .C2(n16194), .A(n16193), .B(n16192), .ZN(
        n16198) );
  NAND2_X1 U18156 ( .A1(n16196), .A2(n21345), .ZN(n16197) );
  OAI211_X1 U18157 ( .C1(n16199), .C2(n21339), .A(n16198), .B(n16197), .ZN(
        P1_U3004) );
  NAND3_X1 U18158 ( .A1(n16080), .A2(n16200), .A3(n21346), .ZN(n16208) );
  NAND3_X1 U18159 ( .A1(n16231), .A2(n16201), .A3(n16212), .ZN(n16210) );
  AOI21_X1 U18160 ( .B1(n16213), .B2(n16210), .A(n16202), .ZN(n16206) );
  OAI21_X1 U18161 ( .B1(n16204), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16203), .ZN(n16205) );
  NOR2_X1 U18162 ( .A1(n16206), .A2(n16205), .ZN(n16207) );
  OAI211_X1 U18163 ( .C1(n21338), .C2(n16209), .A(n16208), .B(n16207), .ZN(
        P1_U3005) );
  INV_X1 U18164 ( .A(n21573), .ZN(n16215) );
  OAI211_X1 U18165 ( .C1(n16213), .C2(n16212), .A(n16211), .B(n16210), .ZN(
        n16214) );
  AOI21_X1 U18166 ( .B1(n16215), .B2(n21345), .A(n16214), .ZN(n16216) );
  OAI21_X1 U18167 ( .B1(n16217), .B2(n21339), .A(n16216), .ZN(P1_U3006) );
  NAND2_X1 U18168 ( .A1(n16218), .A2(n21346), .ZN(n16226) );
  INV_X1 U18169 ( .A(n16219), .ZN(n16228) );
  OAI21_X1 U18170 ( .B1(n16220), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16228), .ZN(n16224) );
  INV_X1 U18171 ( .A(n16231), .ZN(n16221) );
  NOR3_X1 U18172 ( .A1(n16221), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16232), .ZN(n16222) );
  AOI211_X1 U18173 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n16224), .A(
        n16223), .B(n16222), .ZN(n16225) );
  OAI211_X1 U18174 ( .C1(n21338), .C2(n21548), .A(n16226), .B(n16225), .ZN(
        P1_U3007) );
  NAND2_X1 U18175 ( .A1(n16227), .A2(n21346), .ZN(n16234) );
  NOR2_X1 U18176 ( .A1(n16228), .A2(n16232), .ZN(n16229) );
  AOI211_X1 U18177 ( .C1(n16232), .C2(n16231), .A(n16230), .B(n16229), .ZN(
        n16233) );
  OAI211_X1 U18178 ( .C1(n21338), .C2(n21537), .A(n16234), .B(n16233), .ZN(
        P1_U3008) );
  INV_X1 U18179 ( .A(n16235), .ZN(n16236) );
  OR2_X1 U18180 ( .A1(n21285), .A2(n16236), .ZN(n16239) );
  OR2_X1 U18181 ( .A1(n16237), .A2(n21289), .ZN(n16238) );
  NAND3_X1 U18182 ( .A1(n16239), .A2(n21284), .A3(n16238), .ZN(n16272) );
  NOR2_X1 U18183 ( .A1(n16272), .A2(n16242), .ZN(n16255) );
  INV_X1 U18184 ( .A(n16240), .ZN(n16254) );
  NOR2_X1 U18185 ( .A1(n16358), .A2(n16326), .ZN(n16329) );
  NAND3_X1 U18186 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16282), .A3(
        n16329), .ZN(n21352) );
  NOR2_X1 U18187 ( .A1(n21352), .A2(n16241), .ZN(n16280) );
  INV_X1 U18188 ( .A(n16242), .ZN(n16243) );
  NAND3_X1 U18189 ( .A1(n16277), .A2(n16243), .A3(n16253), .ZN(n16259) );
  OAI21_X1 U18190 ( .B1(n16255), .B2(n16254), .A(n16259), .ZN(n16250) );
  INV_X1 U18191 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16244) );
  NAND3_X1 U18192 ( .A1(n16277), .A2(n16245), .A3(n16244), .ZN(n16246) );
  OAI211_X1 U18193 ( .C1(n16248), .C2(n21338), .A(n16247), .B(n16246), .ZN(
        n16249) );
  AOI21_X1 U18194 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16250), .A(
        n16249), .ZN(n16251) );
  OAI21_X1 U18195 ( .B1(n16252), .B2(n21339), .A(n16251), .ZN(P1_U3009) );
  NOR3_X1 U18196 ( .A1(n16255), .A2(n16254), .A3(n16253), .ZN(n16256) );
  AOI211_X1 U18197 ( .C1(n16258), .C2(n21345), .A(n16257), .B(n16256), .ZN(
        n16260) );
  OAI211_X1 U18198 ( .C1(n16261), .C2(n21339), .A(n16260), .B(n16259), .ZN(
        P1_U3010) );
  NOR2_X1 U18199 ( .A1(n16276), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16268) );
  INV_X1 U18200 ( .A(n16262), .ZN(n16283) );
  INV_X1 U18201 ( .A(n16312), .ZN(n16263) );
  NOR2_X1 U18202 ( .A1(n21283), .A2(n16316), .ZN(n16313) );
  AOI22_X1 U18203 ( .A1(n21305), .A2(n16283), .B1(n16263), .B2(n16313), .ZN(
        n21276) );
  AOI21_X1 U18204 ( .B1(n21276), .B2(n16365), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16264) );
  OAI21_X1 U18205 ( .B1(n16264), .B2(n16272), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16265) );
  OAI211_X1 U18206 ( .C1(n21503), .C2(n21338), .A(n16266), .B(n16265), .ZN(
        n16267) );
  AOI21_X1 U18207 ( .B1(n16277), .B2(n16268), .A(n16267), .ZN(n16269) );
  OAI21_X1 U18208 ( .B1(n16270), .B2(n21339), .A(n16269), .ZN(P1_U3011) );
  XNOR2_X1 U18209 ( .A(n16336), .B(n16276), .ZN(n16271) );
  XNOR2_X1 U18210 ( .A(n16114), .B(n16271), .ZN(n20040) );
  INV_X1 U18211 ( .A(n20040), .ZN(n16279) );
  NAND2_X1 U18212 ( .A1(n21348), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n16274) );
  NAND2_X1 U18213 ( .A1(n16272), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16273) );
  OAI211_X1 U18214 ( .C1(n21501), .C2(n21338), .A(n16274), .B(n16273), .ZN(
        n16275) );
  AOI21_X1 U18215 ( .B1(n16277), .B2(n16276), .A(n16275), .ZN(n16278) );
  OAI21_X1 U18216 ( .B1(n16279), .B2(n21339), .A(n16278), .ZN(P1_U3012) );
  INV_X1 U18217 ( .A(n16280), .ZN(n16292) );
  NAND3_X1 U18218 ( .A1(n16281), .A2(n21346), .A3(n16129), .ZN(n16291) );
  INV_X1 U18219 ( .A(n16316), .ZN(n16308) );
  OAI21_X1 U18220 ( .B1(n21285), .B2(n16308), .A(n16282), .ZN(n16285) );
  NOR2_X1 U18221 ( .A1(n16283), .A2(n21289), .ZN(n16310) );
  AOI211_X1 U18222 ( .C1(n16286), .C2(n16285), .A(n16310), .B(n16284), .ZN(
        n21349) );
  OAI21_X1 U18223 ( .B1(n16328), .B2(n16287), .A(n21349), .ZN(n16304) );
  OAI21_X1 U18224 ( .B1(n21486), .B2(n21338), .A(n16288), .ZN(n16289) );
  AOI21_X1 U18225 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n16304), .A(
        n16289), .ZN(n16290) );
  OAI211_X1 U18226 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n16292), .A(
        n16291), .B(n16290), .ZN(P1_U3013) );
  INV_X1 U18227 ( .A(n16293), .ZN(n16295) );
  INV_X1 U18228 ( .A(n16135), .ZN(n16294) );
  AOI211_X1 U18229 ( .C1(n16337), .C2(n16296), .A(n16295), .B(n16294), .ZN(
        n16298) );
  INV_X1 U18230 ( .A(n16298), .ZN(n16297) );
  NAND2_X1 U18231 ( .A1(n16297), .A2(n16302), .ZN(n16300) );
  NAND2_X1 U18232 ( .A1(n16298), .A2(n21353), .ZN(n16299) );
  MUX2_X1 U18233 ( .A(n16300), .B(n16299), .S(n16337), .Z(n16301) );
  XNOR2_X1 U18234 ( .A(n16301), .B(n13917), .ZN(n20037) );
  AOI22_X1 U18235 ( .A1(n19984), .A2(n21345), .B1(n21348), .B2(
        P1_REIP_REG_17__SCAN_IN), .ZN(n16307) );
  INV_X1 U18236 ( .A(n16302), .ZN(n16303) );
  OAI21_X1 U18237 ( .B1(n21352), .B2(n16303), .A(n13917), .ZN(n16305) );
  NAND2_X1 U18238 ( .A1(n16305), .A2(n16304), .ZN(n16306) );
  OAI211_X1 U18239 ( .C1(n20037), .C2(n21339), .A(n16307), .B(n16306), .ZN(
        P1_U3014) );
  AOI21_X1 U18240 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16308), .A(
        n16365), .ZN(n16309) );
  NOR2_X1 U18241 ( .A1(n16310), .A2(n16309), .ZN(n16311) );
  OAI211_X1 U18242 ( .C1(n16313), .C2(n16312), .A(n16311), .B(n16366), .ZN(
        n21277) );
  OAI21_X1 U18243 ( .B1(n16315), .B2(n21338), .A(n16314), .ZN(n16318) );
  AOI221_X1 U18244 ( .B1(n16316), .B2(n21276), .C1(n16365), .C2(n21276), .A(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16317) );
  AOI211_X1 U18245 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n21277), .A(
        n16318), .B(n16317), .ZN(n16319) );
  OAI21_X1 U18246 ( .B1(n16320), .B2(n21339), .A(n16319), .ZN(P1_U3018) );
  INV_X1 U18247 ( .A(n16321), .ZN(n16322) );
  OAI21_X1 U18248 ( .B1(n16133), .B2(n16336), .A(n16322), .ZN(n16324) );
  AOI21_X1 U18249 ( .B1(n16325), .B2(n16324), .A(n16323), .ZN(n20026) );
  INV_X1 U18250 ( .A(n16326), .ZN(n16327) );
  OAI21_X1 U18251 ( .B1(n16328), .B2(n16327), .A(n21324), .ZN(n16347) );
  AOI22_X1 U18252 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16347), .B1(
        n16329), .B2(n16133), .ZN(n16335) );
  AND2_X1 U18253 ( .A1(n16331), .A2(n16330), .ZN(n16332) );
  NOR2_X1 U18254 ( .A1(n16333), .A2(n16332), .ZN(n21455) );
  AOI22_X1 U18255 ( .A1(n21455), .A2(n21345), .B1(n21348), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16334) );
  OAI211_X1 U18256 ( .C1(n20026), .C2(n21339), .A(n16335), .B(n16334), .ZN(
        P1_U3019) );
  NOR2_X1 U18257 ( .A1(n10998), .A2(n16336), .ZN(n16340) );
  INV_X1 U18258 ( .A(n16146), .ZN(n16339) );
  INV_X1 U18259 ( .A(n10998), .ZN(n16338) );
  MUX2_X1 U18260 ( .A(n16339), .B(n16338), .S(n16337), .Z(n16350) );
  MUX2_X1 U18261 ( .A(n13755), .B(n16340), .S(n16349), .Z(n16341) );
  NAND3_X1 U18262 ( .A1(n16343), .A2(n16342), .A3(n21319), .ZN(n16345) );
  NOR2_X1 U18263 ( .A1(n21288), .A2(n21453), .ZN(n20020) );
  INV_X1 U18264 ( .A(n20020), .ZN(n16344) );
  OAI211_X1 U18265 ( .C1(n21338), .C2(n21446), .A(n16345), .B(n16344), .ZN(
        n16346) );
  AOI21_X1 U18266 ( .B1(n16347), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16346), .ZN(n16348) );
  OAI21_X1 U18267 ( .B1(n20018), .B2(n21339), .A(n16348), .ZN(P1_U3020) );
  OAI21_X1 U18268 ( .B1(n16350), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16349), .ZN(n20017) );
  NAND2_X1 U18269 ( .A1(n15384), .A2(n16351), .ZN(n16352) );
  AND2_X1 U18270 ( .A1(n16353), .A2(n16352), .ZN(n21438) );
  OAI21_X1 U18271 ( .B1(n16355), .B2(n16354), .A(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16356) );
  OAI21_X1 U18272 ( .B1(n21288), .B2(n21435), .A(n16356), .ZN(n16360) );
  NOR3_X1 U18273 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16358), .A3(
        n16357), .ZN(n16359) );
  AOI211_X1 U18274 ( .C1(n21345), .C2(n21438), .A(n16360), .B(n16359), .ZN(
        n16361) );
  OAI21_X1 U18275 ( .B1(n20017), .B2(n21339), .A(n16361), .ZN(P1_U3021) );
  OR2_X1 U18276 ( .A1(n16362), .A2(n21339), .ZN(n16371) );
  AOI21_X1 U18277 ( .B1(n21345), .B2(n16364), .A(n16363), .ZN(n16370) );
  NAND2_X1 U18278 ( .A1(n16366), .A2(n16365), .ZN(n16367) );
  NAND2_X1 U18279 ( .A1(n16367), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16368) );
  NAND4_X1 U18280 ( .A1(n16371), .A2(n16370), .A3(n16369), .A4(n16368), .ZN(
        P1_U3031) );
  OAI21_X1 U18281 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n21759), .A(n21858), 
        .ZN(n16372) );
  OAI21_X1 U18282 ( .B1(n16373), .B2(n15264), .A(n16372), .ZN(n16374) );
  MUX2_X1 U18283 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n16374), .S(
        n17190), .Z(P1_U3477) );
  NOR3_X1 U18284 ( .A1(n13490), .A2(n14915), .A3(n14762), .ZN(n16377) );
  NOR2_X1 U18285 ( .A1(n15264), .A2(n16375), .ZN(n16376) );
  AOI211_X1 U18286 ( .C1(n17152), .C2(n13551), .A(n16377), .B(n16376), .ZN(
        n17156) );
  INV_X1 U18287 ( .A(n16385), .ZN(n16383) );
  OAI22_X1 U18288 ( .A1(n16378), .A2(n21300), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16387) );
  NOR2_X1 U18289 ( .A1(n16379), .A2(n21283), .ZN(n16389) );
  NOR3_X1 U18290 ( .A1(n14915), .A2(n14762), .A3(n16380), .ZN(n16381) );
  AOI21_X1 U18291 ( .B1(n16387), .B2(n16389), .A(n16381), .ZN(n16382) );
  OAI21_X1 U18292 ( .B1(n17156), .B2(n16383), .A(n16382), .ZN(n16384) );
  MUX2_X1 U18293 ( .A(n16384), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n16393), .Z(P1_U3473) );
  NAND2_X1 U18294 ( .A1(n16386), .A2(n16385), .ZN(n16392) );
  INV_X1 U18295 ( .A(n16387), .ZN(n16388) );
  AOI22_X1 U18296 ( .A1(n16390), .A2(n21587), .B1(n16389), .B2(n16388), .ZN(
        n16391) );
  NAND2_X1 U18297 ( .A1(n16392), .A2(n16391), .ZN(n16394) );
  MUX2_X1 U18298 ( .A(n16394), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n16393), .Z(P1_U3472) );
  NAND2_X1 U18299 ( .A1(n16679), .A2(n16397), .ZN(n16396) );
  INV_X1 U18300 ( .A(n16399), .ZN(n16395) );
  OAI21_X1 U18301 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16398), .A(
        n16397), .ZN(n18488) );
  NAND2_X1 U18302 ( .A1(n18487), .A2(n18488), .ZN(n18496) );
  NOR2_X1 U18303 ( .A1(n18497), .A2(n18496), .ZN(n18516) );
  OAI21_X1 U18304 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n16399), .A(
        n16401), .ZN(n18518) );
  NAND2_X1 U18305 ( .A1(n18516), .A2(n18518), .ZN(n18525) );
  INV_X1 U18306 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16400) );
  AOI21_X1 U18307 ( .B1(n16401), .B2(n16400), .A(n16403), .ZN(n18527) );
  OAI21_X1 U18308 ( .B1(n16403), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16402), .ZN(n18546) );
  NAND2_X1 U18309 ( .A1(n18606), .A2(n18545), .ZN(n16445) );
  OR2_X1 U18310 ( .A1(n11079), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16404) );
  NAND2_X1 U18311 ( .A1(n16406), .A2(n16404), .ZN(n18559) );
  NAND2_X1 U18312 ( .A1(n18606), .A2(n18557), .ZN(n18567) );
  INV_X1 U18313 ( .A(n16408), .ZN(n16405) );
  AOI21_X1 U18314 ( .B1(n16628), .B2(n16406), .A(n16405), .ZN(n16631) );
  INV_X1 U18315 ( .A(n16631), .ZN(n18568) );
  NAND2_X1 U18316 ( .A1(n18606), .A2(n18566), .ZN(n16431) );
  NAND2_X1 U18317 ( .A1(n16408), .A2(n16407), .ZN(n16409) );
  NAND2_X1 U18318 ( .A1(n16410), .A2(n16409), .ZN(n16619) );
  AOI21_X1 U18319 ( .B1(n16605), .B2(n16410), .A(n16411), .ZN(n16608) );
  INV_X1 U18320 ( .A(n16608), .ZN(n18579) );
  OR2_X1 U18321 ( .A1(n16411), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16412) );
  NAND2_X1 U18322 ( .A1(n16414), .A2(n16412), .ZN(n18590) );
  NAND2_X1 U18323 ( .A1(n18606), .A2(n18588), .ZN(n16417) );
  NAND2_X1 U18324 ( .A1(n16414), .A2(n16413), .ZN(n16415) );
  NAND2_X1 U18325 ( .A1(n16416), .A2(n16415), .ZN(n16580) );
  OAI211_X1 U18326 ( .C1(n16417), .C2(n16580), .A(n18617), .B(n18605), .ZN(
        n16428) );
  OR2_X1 U18327 ( .A1(n16418), .A2(n16419), .ZN(n16420) );
  NAND2_X1 U18328 ( .A1(n13358), .A2(n16420), .ZN(n16583) );
  INV_X1 U18329 ( .A(n16583), .ZN(n16794) );
  AND2_X1 U18330 ( .A1(n16538), .A2(n16421), .ZN(n16423) );
  OR2_X1 U18331 ( .A1(n16423), .A2(n16422), .ZN(n16791) );
  AOI22_X1 U18332 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n18640), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n18639), .ZN(n16425) );
  NAND2_X1 U18333 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18641), .ZN(
        n16424) );
  OAI211_X1 U18334 ( .C1(n16791), .C2(n18638), .A(n16425), .B(n16424), .ZN(
        n16426) );
  AOI21_X1 U18335 ( .B1(n16794), .B2(n18645), .A(n16426), .ZN(n16427) );
  OAI211_X1 U18336 ( .C1(n16429), .C2(n18529), .A(n16428), .B(n16427), .ZN(
        P2_U2828) );
  OAI211_X1 U18337 ( .C1(n16431), .C2(n16619), .A(n18617), .B(n16430), .ZN(
        n16441) );
  INV_X1 U18338 ( .A(n16432), .ZN(n16511) );
  AND2_X1 U18339 ( .A1(n16511), .A2(n16433), .ZN(n16434) );
  NOR2_X1 U18340 ( .A1(n11414), .A2(n16434), .ZN(n16616) );
  XOR2_X1 U18341 ( .A(n16436), .B(n16435), .Z(n16822) );
  NAND2_X1 U18342 ( .A1(n16822), .A2(n18644), .ZN(n16438) );
  AOI22_X1 U18343 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n18640), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18639), .ZN(n16437) );
  OAI211_X1 U18344 ( .C1(n16407), .C2(n18596), .A(n16438), .B(n16437), .ZN(
        n16439) );
  AOI21_X1 U18345 ( .B1(n16616), .B2(n18645), .A(n16439), .ZN(n16440) );
  OAI211_X1 U18346 ( .C1(n18529), .C2(n16442), .A(n16441), .B(n16440), .ZN(
        P2_U2831) );
  OAI211_X1 U18347 ( .C1(n16445), .C2(n16444), .A(n18617), .B(n16443), .ZN(
        n16453) );
  INV_X1 U18348 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n16446) );
  OAI22_X1 U18349 ( .A1(n16446), .A2(n18598), .B1(n13296), .B2(n18627), .ZN(
        n16450) );
  OAI22_X1 U18350 ( .A1(n18638), .A2(n16448), .B1(n16447), .B2(n18596), .ZN(
        n16449) );
  AOI211_X1 U18351 ( .C1(n16451), .C2(n18645), .A(n16450), .B(n16449), .ZN(
        n16452) );
  OAI211_X1 U18352 ( .C1(n18529), .C2(n16454), .A(n16453), .B(n16452), .ZN(
        P2_U2834) );
  AOI211_X1 U18353 ( .C1(n18384), .C2(n16456), .A(n18517), .B(n16455), .ZN(
        n17059) );
  NAND2_X1 U18354 ( .A1(n17059), .A2(n18617), .ZN(n16471) );
  INV_X1 U18355 ( .A(n16457), .ZN(n18509) );
  AOI22_X1 U18356 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18641), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n18639), .ZN(n16458) );
  OAI21_X1 U18357 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18509), .A(
        n16458), .ZN(n16459) );
  AOI21_X1 U18358 ( .B1(n18640), .B2(P2_EBX_REG_1__SCAN_IN), .A(n16459), .ZN(
        n16467) );
  INV_X1 U18359 ( .A(n16460), .ZN(n16463) );
  INV_X1 U18360 ( .A(n16461), .ZN(n16462) );
  NAND2_X1 U18361 ( .A1(n16463), .A2(n16462), .ZN(n16464) );
  NAND2_X1 U18362 ( .A1(n16465), .A2(n16464), .ZN(n19632) );
  NAND2_X1 U18363 ( .A1(n19632), .A2(n18644), .ZN(n16466) );
  OAI211_X1 U18364 ( .C1(n18529), .C2(n16468), .A(n16467), .B(n16466), .ZN(
        n16469) );
  AOI21_X1 U18365 ( .B1(n14681), .B2(n18645), .A(n16469), .ZN(n16470) );
  OAI211_X1 U18366 ( .C1(n19424), .C2(n18400), .A(n16471), .B(n16470), .ZN(
        P2_U2854) );
  INV_X1 U18367 ( .A(n16472), .ZN(n18646) );
  MUX2_X1 U18368 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n18646), .S(n16473), .Z(
        P2_U2856) );
  INV_X1 U18369 ( .A(n16475), .ZN(n16476) );
  NOR2_X1 U18370 ( .A1(n10994), .A2(n16476), .ZN(n16478) );
  XNOR2_X1 U18371 ( .A(n16478), .B(n16477), .ZN(n16530) );
  NOR2_X1 U18372 ( .A1(n18602), .A2(n16513), .ZN(n16479) );
  AOI21_X1 U18373 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16513), .A(n16479), .ZN(
        n16480) );
  OAI21_X1 U18374 ( .B1(n16530), .B2(n16524), .A(n16480), .ZN(P2_U2859) );
  INV_X1 U18375 ( .A(n10994), .ZN(n16482) );
  NAND2_X1 U18376 ( .A1(n16482), .A2(n16481), .ZN(n16483) );
  XOR2_X1 U18377 ( .A(n16484), .B(n16483), .Z(n16535) );
  NOR2_X1 U18378 ( .A1(n16583), .A2(n16513), .ZN(n16485) );
  AOI21_X1 U18379 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16513), .A(n16485), .ZN(
        n16486) );
  OAI21_X1 U18380 ( .B1(n16535), .B2(n16524), .A(n16486), .ZN(P2_U2860) );
  AOI21_X1 U18381 ( .B1(n16489), .B2(n16488), .A(n10993), .ZN(n16490) );
  INV_X1 U18382 ( .A(n16490), .ZN(n16544) );
  NOR2_X1 U18383 ( .A1(n16500), .A2(n16491), .ZN(n16492) );
  OR2_X1 U18384 ( .A1(n16418), .A2(n16492), .ZN(n18586) );
  NOR2_X1 U18385 ( .A1(n18586), .A2(n16513), .ZN(n16493) );
  AOI21_X1 U18386 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n16513), .A(n16493), .ZN(
        n16494) );
  OAI21_X1 U18387 ( .B1(n16544), .B2(n16524), .A(n16494), .ZN(P2_U2861) );
  OAI21_X1 U18388 ( .B1(n16495), .B2(n16497), .A(n16496), .ZN(n16556) );
  NOR2_X1 U18389 ( .A1(n11414), .A2(n16498), .ZN(n16499) );
  OR2_X1 U18390 ( .A1(n16500), .A2(n16499), .ZN(n18575) );
  NOR2_X1 U18391 ( .A1(n18575), .A2(n16513), .ZN(n16501) );
  AOI21_X1 U18392 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n16513), .A(n16501), .ZN(
        n16502) );
  OAI21_X1 U18393 ( .B1(n16556), .B2(n16524), .A(n16502), .ZN(P2_U2862) );
  AOI21_X1 U18394 ( .B1(n11075), .B2(n16504), .A(n16503), .ZN(n16505) );
  INV_X1 U18395 ( .A(n16505), .ZN(n16561) );
  INV_X1 U18396 ( .A(n16616), .ZN(n16826) );
  NOR2_X1 U18397 ( .A1(n16826), .A2(n16513), .ZN(n16506) );
  AOI21_X1 U18398 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16513), .A(n16506), .ZN(
        n16507) );
  OAI21_X1 U18399 ( .B1(n16561), .B2(n16524), .A(n16507), .ZN(P2_U2863) );
  XNOR2_X1 U18400 ( .A(n16515), .B(n16508), .ZN(n16568) );
  NAND2_X1 U18401 ( .A1(n16522), .A2(n16509), .ZN(n16510) );
  NAND2_X1 U18402 ( .A1(n16511), .A2(n16510), .ZN(n16832) );
  NOR2_X1 U18403 ( .A1(n16832), .A2(n16513), .ZN(n16512) );
  AOI21_X1 U18404 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16513), .A(n16512), .ZN(
        n16514) );
  OAI21_X1 U18405 ( .B1(n16568), .B2(n16524), .A(n16514), .ZN(P2_U2864) );
  AOI21_X1 U18406 ( .B1(n16517), .B2(n16516), .A(n16515), .ZN(n16518) );
  INV_X1 U18407 ( .A(n16518), .ZN(n16577) );
  OR2_X1 U18408 ( .A1(n16520), .A2(n16519), .ZN(n16521) );
  NAND2_X1 U18409 ( .A1(n16522), .A2(n16521), .ZN(n18554) );
  MUX2_X1 U18410 ( .A(n18554), .B(n12495), .S(n16513), .Z(n16523) );
  OAI21_X1 U18411 ( .B1(n16577), .B2(n16524), .A(n16523), .ZN(P2_U2865) );
  OAI22_X1 U18412 ( .A1(n18611), .A2(n19688), .B1(n19686), .B2(n16525), .ZN(
        n16526) );
  AOI21_X1 U18413 ( .B1(n16574), .B2(n16527), .A(n16526), .ZN(n16529) );
  AOI22_X1 U18414 ( .A1(n19185), .A2(BUF2_REG_28__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n16528) );
  OAI211_X1 U18415 ( .C1(n16530), .C2(n19636), .A(n16529), .B(n16528), .ZN(
        P2_U2891) );
  AOI22_X1 U18416 ( .A1(n16574), .A2(n19203), .B1(n19631), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16532) );
  AOI22_X1 U18417 ( .A1(n19185), .A2(BUF2_REG_27__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n16531) );
  OAI211_X1 U18418 ( .C1(n16791), .C2(n19688), .A(n16532), .B(n16531), .ZN(
        n16533) );
  INV_X1 U18419 ( .A(n16533), .ZN(n16534) );
  OAI21_X1 U18420 ( .B1(n16535), .B2(n19636), .A(n16534), .ZN(P2_U2892) );
  NAND2_X1 U18421 ( .A1(n16548), .A2(n16536), .ZN(n16537) );
  NAND2_X1 U18422 ( .A1(n16538), .A2(n16537), .ZN(n18585) );
  OAI22_X1 U18423 ( .A1(n18585), .A2(n19688), .B1(n19686), .B2(n16539), .ZN(
        n16540) );
  AOI21_X1 U18424 ( .B1(n16574), .B2(n16541), .A(n16540), .ZN(n16543) );
  AOI22_X1 U18425 ( .A1(n19185), .A2(BUF2_REG_26__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n16542) );
  OAI211_X1 U18426 ( .C1(n16544), .C2(n19636), .A(n16543), .B(n16542), .ZN(
        P2_U2893) );
  OR2_X1 U18427 ( .A1(n16546), .A2(n16545), .ZN(n16547) );
  NAND2_X1 U18428 ( .A1(n16548), .A2(n16547), .ZN(n18574) );
  OAI22_X1 U18429 ( .A1(n18574), .A2(n19688), .B1(n19686), .B2(n14852), .ZN(
        n16554) );
  INV_X1 U18430 ( .A(n19185), .ZN(n16552) );
  INV_X1 U18431 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n16551) );
  INV_X1 U18432 ( .A(n19184), .ZN(n16550) );
  INV_X1 U18433 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16549) );
  OAI22_X1 U18434 ( .A1(n16552), .A2(n16551), .B1(n16550), .B2(n16549), .ZN(
        n16553) );
  AOI211_X1 U18435 ( .C1(n16574), .C2(n19211), .A(n16554), .B(n16553), .ZN(
        n16555) );
  OAI21_X1 U18436 ( .B1(n16556), .B2(n19636), .A(n16555), .ZN(P2_U2894) );
  OAI22_X1 U18437 ( .A1(n19189), .A2(n19215), .B1(n19686), .B2(n16557), .ZN(
        n16558) );
  AOI21_X1 U18438 ( .B1(n16822), .B2(n19633), .A(n16558), .ZN(n16560) );
  AOI22_X1 U18439 ( .A1(n19185), .A2(BUF2_REG_24__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n16559) );
  OAI211_X1 U18440 ( .C1(n16561), .C2(n19636), .A(n16560), .B(n16559), .ZN(
        P2_U2895) );
  AOI22_X1 U18441 ( .A1(n19185), .A2(BUF2_REG_23__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16565) );
  AND2_X1 U18442 ( .A1(n11063), .A2(n16562), .ZN(n16563) );
  NOR2_X1 U18443 ( .A1(n16435), .A2(n16563), .ZN(n18564) );
  AOI22_X1 U18444 ( .A1(n19633), .A2(n18564), .B1(n19631), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16564) );
  OAI211_X1 U18445 ( .C1(n19218), .C2(n19189), .A(n16565), .B(n16564), .ZN(
        n16566) );
  INV_X1 U18446 ( .A(n16566), .ZN(n16567) );
  OAI21_X1 U18447 ( .B1(n16568), .B2(n19636), .A(n16567), .ZN(P2_U2896) );
  INV_X1 U18448 ( .A(n13334), .ZN(n16570) );
  OAI21_X1 U18449 ( .B1(n16570), .B2(n11226), .A(n11063), .ZN(n18562) );
  OAI22_X1 U18450 ( .A1(n19688), .A2(n18562), .B1(n19686), .B2(n16571), .ZN(
        n16572) );
  AOI21_X1 U18451 ( .B1(n16574), .B2(n16573), .A(n16572), .ZN(n16576) );
  AOI22_X1 U18452 ( .A1(n19185), .A2(BUF2_REG_22__SCAN_IN), .B1(n19184), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16575) );
  OAI211_X1 U18453 ( .C1(n16577), .C2(n19636), .A(n16576), .B(n16575), .ZN(
        P2_U2897) );
  XNOR2_X1 U18454 ( .A(n16578), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16798) );
  INV_X1 U18455 ( .A(n16591), .ZN(n16579) );
  AOI21_X1 U18456 ( .B1(n12524), .B2(n16579), .A(n11144), .ZN(n16795) );
  NOR2_X1 U18457 ( .A1(n18680), .A2(n17492), .ZN(n16788) );
  NOR2_X1 U18458 ( .A1(n16782), .A2(n16580), .ZN(n16581) );
  AOI211_X1 U18459 ( .C1(n16750), .C2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16788), .B(n16581), .ZN(n16582) );
  OAI21_X1 U18460 ( .B1(n16583), .B2(n17410), .A(n16582), .ZN(n16584) );
  AOI21_X1 U18461 ( .B1(n16795), .B2(n16766), .A(n16584), .ZN(n16585) );
  OAI21_X1 U18462 ( .B1(n16798), .B2(n17411), .A(n16585), .ZN(P2_U2987) );
  AOI21_X1 U18463 ( .B1(n16586), .B2(n16599), .A(n16601), .ZN(n16588) );
  MUX2_X1 U18464 ( .A(n16599), .B(n16588), .S(n16587), .Z(n16589) );
  NAND2_X1 U18465 ( .A1(n16590), .A2(n16589), .ZN(n16808) );
  AOI21_X1 U18466 ( .B1(n16799), .B2(n11037), .A(n16591), .ZN(n16806) );
  NOR2_X1 U18467 ( .A1(n18680), .A2(n17491), .ZN(n16800) );
  NOR2_X1 U18468 ( .A1(n16782), .A2(n18590), .ZN(n16592) );
  AOI211_X1 U18469 ( .C1(n16750), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16800), .B(n16592), .ZN(n16593) );
  OAI21_X1 U18470 ( .B1(n18586), .B2(n17410), .A(n16593), .ZN(n16594) );
  AOI21_X1 U18471 ( .B1(n16806), .B2(n16766), .A(n16594), .ZN(n16595) );
  OAI21_X1 U18472 ( .B1(n16808), .B2(n17411), .A(n16595), .ZN(P2_U2988) );
  OAI21_X1 U18473 ( .B1(n16596), .B2(n16597), .A(n16812), .ZN(n16598) );
  NAND2_X1 U18474 ( .A1(n16598), .A2(n11037), .ZN(n16819) );
  INV_X1 U18475 ( .A(n16599), .ZN(n16600) );
  NOR2_X1 U18476 ( .A1(n16601), .A2(n16600), .ZN(n16602) );
  XNOR2_X1 U18477 ( .A(n16586), .B(n16602), .ZN(n16809) );
  NAND2_X1 U18478 ( .A1(n16809), .A2(n12546), .ZN(n16610) );
  NOR2_X1 U18479 ( .A1(n18680), .A2(n16603), .ZN(n16810) );
  INV_X1 U18480 ( .A(n16810), .ZN(n16604) );
  OAI21_X1 U18481 ( .B1(n17417), .B2(n16605), .A(n16604), .ZN(n16607) );
  NOR2_X1 U18482 ( .A1(n18575), .A2(n17410), .ZN(n16606) );
  AOI211_X1 U18483 ( .C1(n17407), .C2(n16608), .A(n16607), .B(n16606), .ZN(
        n16609) );
  OAI211_X1 U18484 ( .C1(n16819), .C2(n17408), .A(n16610), .B(n16609), .ZN(
        P2_U2989) );
  INV_X1 U18485 ( .A(n16612), .ZN(n16613) );
  NOR2_X1 U18486 ( .A1(n16614), .A2(n16613), .ZN(n16615) );
  XNOR2_X1 U18487 ( .A(n16611), .B(n16615), .ZN(n16830) );
  XNOR2_X1 U18488 ( .A(n16596), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16828) );
  NAND2_X1 U18489 ( .A1(n16616), .A2(n16711), .ZN(n16618) );
  NOR2_X1 U18490 ( .A1(n18680), .A2(n17490), .ZN(n16821) );
  AOI21_X1 U18491 ( .B1(n16750), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16821), .ZN(n16617) );
  OAI211_X1 U18492 ( .C1(n16782), .C2(n16619), .A(n16618), .B(n16617), .ZN(
        n16620) );
  AOI21_X1 U18493 ( .B1(n16828), .B2(n16766), .A(n16620), .ZN(n16621) );
  OAI21_X1 U18494 ( .B1(n16830), .B2(n17411), .A(n16621), .ZN(P2_U2990) );
  OAI21_X1 U18495 ( .B1(n16622), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16596), .ZN(n16842) );
  INV_X1 U18496 ( .A(n16624), .ZN(n16626) );
  NOR2_X1 U18497 ( .A1(n16626), .A2(n16625), .ZN(n16627) );
  XNOR2_X1 U18498 ( .A(n11001), .B(n16627), .ZN(n16831) );
  NAND2_X1 U18499 ( .A1(n16831), .A2(n12546), .ZN(n16633) );
  NAND2_X1 U18500 ( .A1(n18500), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16835) );
  OAI21_X1 U18501 ( .B1(n17417), .B2(n16628), .A(n16835), .ZN(n16630) );
  NOR2_X1 U18502 ( .A1(n16832), .A2(n17410), .ZN(n16629) );
  AOI211_X1 U18503 ( .C1(n17407), .C2(n16631), .A(n16630), .B(n16629), .ZN(
        n16632) );
  OAI211_X1 U18504 ( .C1(n17408), .C2(n16842), .A(n16633), .B(n16632), .ZN(
        P2_U2991) );
  INV_X1 U18505 ( .A(n16635), .ZN(n16636) );
  NOR2_X1 U18506 ( .A1(n16637), .A2(n16636), .ZN(n16638) );
  XNOR2_X1 U18507 ( .A(n16634), .B(n16638), .ZN(n16853) );
  AOI21_X1 U18508 ( .B1(n16847), .B2(n13292), .A(n16622), .ZN(n16851) );
  NOR2_X1 U18509 ( .A1(n18680), .A2(n17489), .ZN(n16843) );
  NOR2_X1 U18510 ( .A1(n16782), .A2(n18559), .ZN(n16639) );
  AOI211_X1 U18511 ( .C1(n16750), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16843), .B(n16639), .ZN(n16640) );
  OAI21_X1 U18512 ( .B1(n18554), .B2(n17410), .A(n16640), .ZN(n16641) );
  AOI21_X1 U18513 ( .B1(n16851), .B2(n16766), .A(n16641), .ZN(n16642) );
  OAI21_X1 U18514 ( .B1(n16853), .B2(n17411), .A(n16642), .ZN(P2_U2992) );
  XNOR2_X1 U18515 ( .A(n16643), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16874) );
  XNOR2_X1 U18516 ( .A(n16650), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16872) );
  INV_X1 U18517 ( .A(n18546), .ZN(n16645) );
  NAND2_X1 U18518 ( .A1(n18532), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n16867) );
  OAI21_X1 U18519 ( .B1(n17417), .B2(n11299), .A(n16867), .ZN(n16644) );
  AOI21_X1 U18520 ( .B1(n17407), .B2(n16645), .A(n16644), .ZN(n16646) );
  OAI21_X1 U18521 ( .B1(n18542), .B2(n17410), .A(n16646), .ZN(n16647) );
  AOI21_X1 U18522 ( .B1(n16872), .B2(n16766), .A(n16647), .ZN(n16648) );
  OAI21_X1 U18523 ( .B1(n16874), .B2(n17411), .A(n16648), .ZN(P2_U2994) );
  OAI21_X1 U18524 ( .B1(n16665), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n16650), .ZN(n16885) );
  INV_X1 U18525 ( .A(n16663), .ZN(n16651) );
  NOR2_X1 U18526 ( .A1(n11050), .A2(n16651), .ZN(n16655) );
  NAND2_X1 U18527 ( .A1(n16653), .A2(n16652), .ZN(n16654) );
  XNOR2_X1 U18528 ( .A(n16655), .B(n16654), .ZN(n16883) );
  NOR2_X1 U18529 ( .A1(n18680), .A2(n17487), .ZN(n16877) );
  AOI21_X1 U18530 ( .B1(n16750), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16877), .ZN(n16657) );
  NAND2_X1 U18531 ( .A1(n17407), .A2(n18527), .ZN(n16656) );
  OAI211_X1 U18532 ( .C1(n18534), .C2(n17410), .A(n16657), .B(n16656), .ZN(
        n16658) );
  AOI21_X1 U18533 ( .B1(n16883), .B2(n12546), .A(n16658), .ZN(n16659) );
  OAI21_X1 U18534 ( .B1(n16885), .B2(n17408), .A(n16659), .ZN(P2_U2995) );
  AOI21_X1 U18535 ( .B1(n16663), .B2(n16661), .A(n16660), .ZN(n16662) );
  AOI21_X1 U18536 ( .B1(n11050), .B2(n16663), .A(n16662), .ZN(n16896) );
  NAND2_X1 U18537 ( .A1(n16684), .A2(n16664), .ZN(n16677) );
  AOI21_X1 U18538 ( .B1(n16891), .B2(n16677), .A(n16665), .ZN(n16886) );
  NAND2_X1 U18539 ( .A1(n16886), .A2(n16766), .ZN(n16669) );
  NOR2_X1 U18540 ( .A1(n18680), .A2(n18512), .ZN(n16887) );
  AOI21_X1 U18541 ( .B1(n16750), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16887), .ZN(n16666) );
  OAI21_X1 U18542 ( .B1(n16782), .B2(n18518), .A(n16666), .ZN(n16667) );
  AOI21_X1 U18543 ( .B1(n18520), .B2(n16711), .A(n16667), .ZN(n16668) );
  OAI211_X1 U18544 ( .C1(n16896), .C2(n17411), .A(n16669), .B(n16668), .ZN(
        P2_U2996) );
  NAND2_X1 U18545 ( .A1(n16671), .A2(n16670), .ZN(n16675) );
  NAND2_X1 U18546 ( .A1(n16673), .A2(n16672), .ZN(n16674) );
  XOR2_X1 U18547 ( .A(n16675), .B(n16674), .Z(n16904) );
  OAI21_X1 U18548 ( .B1(n16676), .B2(n16905), .A(n16907), .ZN(n16678) );
  NAND3_X1 U18549 ( .A1(n16678), .A2(n16766), .A3(n16677), .ZN(n16683) );
  NAND2_X1 U18550 ( .A1(n18500), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16899) );
  OAI21_X1 U18551 ( .B1(n17417), .B2(n16679), .A(n16899), .ZN(n16681) );
  NOR2_X1 U18552 ( .A1(n16898), .A2(n17410), .ZN(n16680) );
  AOI211_X1 U18553 ( .C1(n17407), .C2(n18497), .A(n16681), .B(n16680), .ZN(
        n16682) );
  OAI211_X1 U18554 ( .C1(n16904), .C2(n17411), .A(n16683), .B(n16682), .ZN(
        P2_U2997) );
  XNOR2_X1 U18555 ( .A(n16684), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16691) );
  NOR2_X1 U18556 ( .A1(n18490), .A2(n17410), .ZN(n16688) );
  NAND2_X1 U18557 ( .A1(n16750), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16685) );
  OAI211_X1 U18558 ( .C1(n16782), .C2(n18488), .A(n16686), .B(n16685), .ZN(
        n16687) );
  AOI211_X1 U18559 ( .C1(n16689), .C2(n12546), .A(n16688), .B(n16687), .ZN(
        n16690) );
  OAI21_X1 U18560 ( .B1(n16691), .B2(n17408), .A(n16690), .ZN(P2_U2998) );
  INV_X1 U18561 ( .A(n12549), .ZN(n16693) );
  OAI21_X1 U18562 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16692), .A(
        n16693), .ZN(n16929) );
  OAI21_X1 U18563 ( .B1(n16696), .B2(n16695), .A(n16694), .ZN(n16927) );
  NOR2_X1 U18564 ( .A1(n18680), .A2(n16697), .ZN(n16917) );
  NOR2_X1 U18565 ( .A1(n16782), .A2(n18474), .ZN(n16698) );
  AOI211_X1 U18566 ( .C1(n16750), .C2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16917), .B(n16698), .ZN(n16699) );
  OAI21_X1 U18567 ( .B1(n18476), .B2(n17410), .A(n16699), .ZN(n16700) );
  AOI21_X1 U18568 ( .B1(n16927), .B2(n12546), .A(n16700), .ZN(n16701) );
  OAI21_X1 U18569 ( .B1(n17408), .B2(n16929), .A(n16701), .ZN(P2_U3000) );
  NAND2_X1 U18570 ( .A1(n16703), .A2(n16702), .ZN(n16704) );
  XNOR2_X1 U18571 ( .A(n12550), .B(n16704), .ZN(n16944) );
  INV_X1 U18572 ( .A(n16727), .ZN(n16706) );
  AOI21_X1 U18573 ( .B1(n16706), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16707) );
  NOR2_X1 U18574 ( .A1(n16707), .A2(n16692), .ZN(n16930) );
  NAND2_X1 U18575 ( .A1(n16930), .A2(n16766), .ZN(n16713) );
  NOR2_X1 U18576 ( .A1(n18680), .A2(n17485), .ZN(n16935) );
  AOI21_X1 U18577 ( .B1(n16750), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16935), .ZN(n16708) );
  OAI21_X1 U18578 ( .B1(n16782), .B2(n16709), .A(n16708), .ZN(n16710) );
  AOI21_X1 U18579 ( .B1(n18466), .B2(n16711), .A(n16710), .ZN(n16712) );
  OAI211_X1 U18580 ( .C1(n17411), .C2(n16944), .A(n16713), .B(n16712), .ZN(
        P2_U3001) );
  XNOR2_X1 U18581 ( .A(n16727), .B(n16714), .ZN(n16955) );
  INV_X1 U18582 ( .A(n16715), .ZN(n16717) );
  NAND2_X1 U18583 ( .A1(n16717), .A2(n16716), .ZN(n16721) );
  NAND2_X1 U18584 ( .A1(n16719), .A2(n16718), .ZN(n16720) );
  XNOR2_X1 U18585 ( .A(n16721), .B(n16720), .ZN(n16952) );
  NOR2_X1 U18586 ( .A1(n18680), .A2(n17484), .ZN(n16946) );
  NOR2_X1 U18587 ( .A1(n16782), .A2(n18450), .ZN(n16722) );
  AOI211_X1 U18588 ( .C1(n16750), .C2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16946), .B(n16722), .ZN(n16723) );
  OAI21_X1 U18589 ( .B1(n17410), .B2(n18452), .A(n16723), .ZN(n16724) );
  AOI21_X1 U18590 ( .B1(n16952), .B2(n12546), .A(n16724), .ZN(n16725) );
  OAI21_X1 U18591 ( .B1(n16955), .B2(n17408), .A(n16725), .ZN(P2_U3002) );
  OAI21_X1 U18592 ( .B1(n16726), .B2(n16977), .A(n16965), .ZN(n16728) );
  NAND2_X1 U18593 ( .A1(n16728), .A2(n16727), .ZN(n16971) );
  NAND2_X1 U18594 ( .A1(n16730), .A2(n16729), .ZN(n16734) );
  NOR2_X1 U18595 ( .A1(n16732), .A2(n16731), .ZN(n16733) );
  XOR2_X1 U18596 ( .A(n16734), .B(n16733), .Z(n16956) );
  NAND2_X1 U18597 ( .A1(n18500), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n16960) );
  OAI21_X1 U18598 ( .B1(n17417), .B2(n16735), .A(n16960), .ZN(n16736) );
  AOI21_X1 U18599 ( .B1(n17407), .B2(n18440), .A(n16736), .ZN(n16737) );
  OAI21_X1 U18600 ( .B1(n18442), .B2(n17410), .A(n16737), .ZN(n16738) );
  AOI21_X1 U18601 ( .B1(n16956), .B2(n12546), .A(n16738), .ZN(n16739) );
  OAI21_X1 U18602 ( .B1(n17408), .B2(n16971), .A(n16739), .ZN(P2_U3003) );
  XNOR2_X1 U18603 ( .A(n16726), .B(n16977), .ZN(n16982) );
  OR2_X1 U18604 ( .A1(n11058), .A2(n16740), .ZN(n16741) );
  NAND2_X1 U18605 ( .A1(n16741), .A2(n16754), .ZN(n16746) );
  INV_X1 U18606 ( .A(n16742), .ZN(n16744) );
  NAND2_X1 U18607 ( .A1(n16744), .A2(n16743), .ZN(n16745) );
  XNOR2_X1 U18608 ( .A(n16746), .B(n16745), .ZN(n16980) );
  NOR2_X1 U18609 ( .A1(n18680), .A2(n16747), .ZN(n16974) );
  NOR2_X1 U18610 ( .A1(n16782), .A2(n16748), .ZN(n16749) );
  AOI211_X1 U18611 ( .C1(n16750), .C2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16974), .B(n16749), .ZN(n16751) );
  OAI21_X1 U18612 ( .B1(n17410), .B2(n16972), .A(n16751), .ZN(n16752) );
  AOI21_X1 U18613 ( .B1(n16980), .B2(n12546), .A(n16752), .ZN(n16753) );
  OAI21_X1 U18614 ( .B1(n16982), .B2(n17408), .A(n16753), .ZN(P2_U3004) );
  INV_X1 U18615 ( .A(n16754), .ZN(n16755) );
  NOR2_X1 U18616 ( .A1(n16756), .A2(n16755), .ZN(n16763) );
  NAND2_X1 U18617 ( .A1(n16758), .A2(n16757), .ZN(n17020) );
  OR2_X1 U18618 ( .A1(n17020), .A2(n16759), .ZN(n16761) );
  NAND2_X1 U18619 ( .A1(n16761), .A2(n16760), .ZN(n16762) );
  XOR2_X1 U18620 ( .A(n16763), .B(n16762), .Z(n16994) );
  INV_X1 U18621 ( .A(n16764), .ZN(n16765) );
  NAND2_X1 U18622 ( .A1(n16765), .A2(n16991), .ZN(n16983) );
  NAND3_X1 U18623 ( .A1(n16983), .A2(n16766), .A3(n16726), .ZN(n16773) );
  OAI22_X1 U18624 ( .A1(n17417), .A2(n16768), .B1(n16767), .B2(n18680), .ZN(
        n16770) );
  NOR2_X1 U18625 ( .A1(n16986), .A2(n17410), .ZN(n16769) );
  AOI211_X1 U18626 ( .C1(n17407), .C2(n16771), .A(n16770), .B(n16769), .ZN(
        n16772) );
  OAI211_X1 U18627 ( .C1(n16994), .C2(n17411), .A(n16773), .B(n16772), .ZN(
        P2_U3005) );
  OAI21_X1 U18628 ( .B1(n16776), .B2(n16775), .A(n16774), .ZN(n17015) );
  NAND2_X1 U18629 ( .A1(n16778), .A2(n16777), .ZN(n16781) );
  OR2_X1 U18630 ( .A1(n17020), .A2(n17017), .ZN(n16779) );
  NAND2_X1 U18631 ( .A1(n16779), .A2(n17016), .ZN(n16780) );
  XOR2_X1 U18632 ( .A(n16781), .B(n16780), .Z(n17013) );
  OAI22_X1 U18633 ( .A1(n12710), .A2(n18680), .B1(n16782), .B2(n18425), .ZN(
        n16785) );
  INV_X1 U18634 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16783) );
  OAI22_X1 U18635 ( .A1(n18427), .A2(n17410), .B1(n16783), .B2(n17417), .ZN(
        n16784) );
  AOI211_X1 U18636 ( .C1(n17013), .C2(n12546), .A(n16785), .B(n16784), .ZN(
        n16786) );
  OAI21_X1 U18637 ( .B1(n17015), .B2(n17408), .A(n16786), .ZN(P2_U3006) );
  NOR2_X1 U18638 ( .A1(n16787), .A2(n12524), .ZN(n16793) );
  INV_X1 U18639 ( .A(n16788), .ZN(n16789) );
  OAI211_X1 U18640 ( .C1(n16791), .C2(n18662), .A(n16790), .B(n16789), .ZN(
        n16792) );
  AOI211_X1 U18641 ( .C1(n16794), .C2(n18685), .A(n16793), .B(n16792), .ZN(
        n16797) );
  NAND2_X1 U18642 ( .A1(n16795), .A2(n15725), .ZN(n16796) );
  OAI211_X1 U18643 ( .C1(n16798), .C2(n18664), .A(n16797), .B(n16796), .ZN(
        P2_U3019) );
  XNOR2_X1 U18644 ( .A(n16799), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16801) );
  AOI21_X1 U18645 ( .B1(n16801), .B2(n16811), .A(n16800), .ZN(n16802) );
  OAI21_X1 U18646 ( .B1(n18585), .B2(n18662), .A(n16802), .ZN(n16803) );
  AOI21_X1 U18647 ( .B1(n16816), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16803), .ZN(n16804) );
  OAI21_X1 U18648 ( .B1(n18586), .B2(n18666), .A(n16804), .ZN(n16805) );
  AOI21_X1 U18649 ( .B1(n16806), .B2(n15725), .A(n16805), .ZN(n16807) );
  OAI21_X1 U18650 ( .B1(n16808), .B2(n18664), .A(n16807), .ZN(P2_U3020) );
  NAND2_X1 U18651 ( .A1(n16809), .A2(n13329), .ZN(n16818) );
  AOI21_X1 U18652 ( .B1(n16812), .B2(n16811), .A(n16810), .ZN(n16813) );
  OAI21_X1 U18653 ( .B1(n18574), .B2(n18662), .A(n16813), .ZN(n16815) );
  NOR2_X1 U18654 ( .A1(n18575), .A2(n18666), .ZN(n16814) );
  AOI211_X1 U18655 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n16816), .A(
        n16815), .B(n16814), .ZN(n16817) );
  OAI211_X1 U18656 ( .C1(n18688), .C2(n16819), .A(n16818), .B(n16817), .ZN(
        P2_U3021) );
  AOI211_X1 U18657 ( .C1(n12928), .C2(n16822), .A(n16821), .B(n16820), .ZN(
        n16825) );
  NAND2_X1 U18658 ( .A1(n16823), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16824) );
  OAI211_X1 U18659 ( .C1(n16826), .C2(n18666), .A(n16825), .B(n16824), .ZN(
        n16827) );
  AOI21_X1 U18660 ( .B1(n16828), .B2(n15725), .A(n16827), .ZN(n16829) );
  OAI21_X1 U18661 ( .B1(n16830), .B2(n18664), .A(n16829), .ZN(P2_U3022) );
  NAND2_X1 U18662 ( .A1(n16831), .A2(n13329), .ZN(n16841) );
  INV_X1 U18663 ( .A(n16832), .ZN(n18565) );
  NAND3_X1 U18664 ( .A1(n16990), .A2(n16833), .A3(n16847), .ZN(n16845) );
  AOI21_X1 U18665 ( .B1(n16848), .B2(n16845), .A(n16834), .ZN(n16839) );
  NAND2_X1 U18666 ( .A1(n12928), .A2(n18564), .ZN(n16836) );
  OAI211_X1 U18667 ( .C1(n16837), .C2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16836), .B(n16835), .ZN(n16838) );
  AOI211_X1 U18668 ( .C1(n18565), .C2(n18685), .A(n16839), .B(n16838), .ZN(
        n16840) );
  OAI211_X1 U18669 ( .C1(n16842), .C2(n18688), .A(n16841), .B(n16840), .ZN(
        P2_U3023) );
  NOR2_X1 U18670 ( .A1(n18554), .A2(n18666), .ZN(n16850) );
  INV_X1 U18671 ( .A(n18562), .ZN(n16844) );
  AOI21_X1 U18672 ( .B1(n12928), .B2(n16844), .A(n16843), .ZN(n16846) );
  OAI211_X1 U18673 ( .C1(n16848), .C2(n16847), .A(n16846), .B(n16845), .ZN(
        n16849) );
  AOI211_X1 U18674 ( .C1(n16851), .C2(n15725), .A(n16850), .B(n16849), .ZN(
        n16852) );
  OAI21_X1 U18675 ( .B1(n16853), .B2(n18664), .A(n16852), .ZN(P2_U3024) );
  INV_X1 U18676 ( .A(n16858), .ZN(n16854) );
  NOR2_X1 U18677 ( .A1(n16855), .A2(n16854), .ZN(n16863) );
  NAND2_X1 U18678 ( .A1(n16863), .A2(n16891), .ZN(n16890) );
  NOR2_X1 U18679 ( .A1(n16857), .A2(n12915), .ZN(n16859) );
  OAI21_X1 U18680 ( .B1(n17002), .B2(n16859), .A(n16858), .ZN(n16860) );
  NAND2_X1 U18681 ( .A1(n16860), .A2(n18671), .ZN(n16861) );
  AND2_X1 U18682 ( .A1(n16862), .A2(n16861), .ZN(n16892) );
  NAND2_X1 U18683 ( .A1(n16890), .A2(n16892), .ZN(n16879) );
  INV_X1 U18684 ( .A(n16863), .ZN(n16875) );
  OAI21_X1 U18685 ( .B1(n16891), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16864) );
  OAI21_X1 U18686 ( .B1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n16864), .ZN(n16868) );
  INV_X1 U18687 ( .A(n18550), .ZN(n16865) );
  NAND2_X1 U18688 ( .A1(n12928), .A2(n16865), .ZN(n16866) );
  OAI211_X1 U18689 ( .C1(n16875), .C2(n16868), .A(n16867), .B(n16866), .ZN(
        n16869) );
  AOI21_X1 U18690 ( .B1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n16879), .A(
        n16869), .ZN(n16870) );
  OAI21_X1 U18691 ( .B1(n18542), .B2(n18666), .A(n16870), .ZN(n16871) );
  AOI21_X1 U18692 ( .B1(n16872), .B2(n15725), .A(n16871), .ZN(n16873) );
  OAI21_X1 U18693 ( .B1(n16874), .B2(n18664), .A(n16873), .ZN(P2_U3026) );
  NOR3_X1 U18694 ( .A1(n16875), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16891), .ZN(n16876) );
  AOI211_X1 U18695 ( .C1(n12928), .C2(n16878), .A(n16877), .B(n16876), .ZN(
        n16881) );
  NAND2_X1 U18696 ( .A1(n16879), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16880) );
  OAI211_X1 U18697 ( .C1(n18534), .C2(n18666), .A(n16881), .B(n16880), .ZN(
        n16882) );
  AOI21_X1 U18698 ( .B1(n16883), .B2(n13329), .A(n16882), .ZN(n16884) );
  OAI21_X1 U18699 ( .B1(n16885), .B2(n18688), .A(n16884), .ZN(P2_U3027) );
  NAND2_X1 U18700 ( .A1(n16886), .A2(n15725), .ZN(n16895) );
  INV_X1 U18701 ( .A(n18524), .ZN(n16888) );
  AOI21_X1 U18702 ( .B1(n12928), .B2(n16888), .A(n16887), .ZN(n16889) );
  OAI211_X1 U18703 ( .C1(n16892), .C2(n16891), .A(n16890), .B(n16889), .ZN(
        n16893) );
  AOI21_X1 U18704 ( .B1(n18520), .B2(n18685), .A(n16893), .ZN(n16894) );
  OAI211_X1 U18705 ( .C1(n16896), .C2(n18664), .A(n16895), .B(n16894), .ZN(
        P2_U3028) );
  NAND3_X1 U18706 ( .A1(n16897), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16907), .ZN(n16903) );
  INV_X1 U18707 ( .A(n16898), .ZN(n18506) );
  OAI21_X1 U18708 ( .B1(n16900), .B2(n18662), .A(n16899), .ZN(n16901) );
  AOI21_X1 U18709 ( .B1(n18506), .B2(n18685), .A(n16901), .ZN(n16902) );
  OAI211_X1 U18710 ( .C1(n16904), .C2(n18664), .A(n16903), .B(n16902), .ZN(
        n16911) );
  OAI21_X1 U18711 ( .B1(n18671), .B2(n16906), .A(n16905), .ZN(n16908) );
  AOI21_X1 U18712 ( .B1(n16909), .B2(n16908), .A(n16907), .ZN(n16910) );
  OR2_X1 U18713 ( .A1(n16911), .A2(n16910), .ZN(P2_U3029) );
  AND2_X1 U18714 ( .A1(n16990), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16964) );
  NAND2_X1 U18715 ( .A1(n16964), .A2(n16912), .ZN(n16919) );
  NOR2_X1 U18716 ( .A1(n16919), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16949) );
  NAND2_X1 U18717 ( .A1(n18671), .A2(n16991), .ZN(n16913) );
  NAND2_X1 U18718 ( .A1(n16987), .A2(n16913), .ZN(n16963) );
  AND2_X1 U18719 ( .A1(n18671), .A2(n16914), .ZN(n16915) );
  OR2_X1 U18720 ( .A1(n16963), .A2(n16915), .ZN(n16951) );
  NOR2_X1 U18721 ( .A1(n16949), .A2(n16951), .ZN(n16939) );
  OR2_X1 U18722 ( .A1(n16919), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16934) );
  AOI21_X1 U18723 ( .B1(n16939), .B2(n16934), .A(n16920), .ZN(n16926) );
  OAI21_X1 U18724 ( .B1(n11062), .B2(n16916), .A(n15464), .ZN(n19196) );
  INV_X1 U18725 ( .A(n19196), .ZN(n16918) );
  AOI21_X1 U18726 ( .B1(n16918), .B2(n12928), .A(n16917), .ZN(n16924) );
  INV_X1 U18727 ( .A(n16919), .ZN(n16922) );
  NAND3_X1 U18728 ( .A1(n16922), .A2(n16921), .A3(n16920), .ZN(n16923) );
  OAI211_X1 U18729 ( .C1(n18476), .C2(n18666), .A(n16924), .B(n16923), .ZN(
        n16925) );
  AOI211_X1 U18730 ( .C1(n16927), .C2(n13329), .A(n16926), .B(n16925), .ZN(
        n16928) );
  OAI21_X1 U18731 ( .B1(n18688), .B2(n16929), .A(n16928), .ZN(P2_U3032) );
  NAND2_X1 U18732 ( .A1(n16930), .A2(n15725), .ZN(n16943) );
  AND2_X1 U18733 ( .A1(n16931), .A2(n16932), .ZN(n16933) );
  OR2_X1 U18734 ( .A1(n11062), .A2(n16933), .ZN(n18465) );
  INV_X1 U18735 ( .A(n16934), .ZN(n16936) );
  AOI21_X1 U18736 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16936), .A(
        n16935), .ZN(n16937) );
  OAI21_X1 U18737 ( .B1(n18662), .B2(n18465), .A(n16937), .ZN(n16941) );
  NOR2_X1 U18738 ( .A1(n16939), .A2(n16938), .ZN(n16940) );
  AOI211_X1 U18739 ( .C1(n18466), .C2(n18685), .A(n16941), .B(n16940), .ZN(
        n16942) );
  OAI211_X1 U18740 ( .C1(n16944), .C2(n18664), .A(n16943), .B(n16942), .ZN(
        P2_U3033) );
  OAI21_X1 U18741 ( .B1(n12789), .B2(n11411), .A(n16931), .ZN(n19202) );
  INV_X1 U18742 ( .A(n19202), .ZN(n16947) );
  AOI21_X1 U18743 ( .B1(n12928), .B2(n16947), .A(n16946), .ZN(n16948) );
  OAI21_X1 U18744 ( .B1(n18452), .B2(n18666), .A(n16948), .ZN(n16950) );
  AOI211_X1 U18745 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16951), .A(
        n16950), .B(n16949), .ZN(n16954) );
  NAND2_X1 U18746 ( .A1(n16952), .A2(n13329), .ZN(n16953) );
  OAI211_X1 U18747 ( .C1(n16955), .C2(n18688), .A(n16954), .B(n16953), .ZN(
        P2_U3034) );
  NAND2_X1 U18748 ( .A1(n16956), .A2(n13329), .ZN(n16970) );
  OR2_X1 U18749 ( .A1(n16958), .A2(n16957), .ZN(n16959) );
  AND2_X1 U18750 ( .A1(n16945), .A2(n16959), .ZN(n19204) );
  INV_X1 U18751 ( .A(n19204), .ZN(n16962) );
  NAND3_X1 U18752 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16964), .A3(
        n16965), .ZN(n16961) );
  OAI211_X1 U18753 ( .C1(n18662), .C2(n16962), .A(n16961), .B(n16960), .ZN(
        n16967) );
  INV_X1 U18754 ( .A(n16963), .ZN(n16978) );
  NAND2_X1 U18755 ( .A1(n16964), .A2(n16977), .ZN(n16975) );
  AOI21_X1 U18756 ( .B1(n16978), .B2(n16975), .A(n16965), .ZN(n16966) );
  AOI211_X1 U18757 ( .C1(n16968), .C2(n18685), .A(n16967), .B(n16966), .ZN(
        n16969) );
  OAI211_X1 U18758 ( .C1(n16971), .C2(n18688), .A(n16970), .B(n16969), .ZN(
        P2_U3035) );
  NOR2_X1 U18759 ( .A1(n16972), .A2(n18666), .ZN(n16973) );
  AOI211_X1 U18760 ( .C1(n12928), .C2(n19207), .A(n16974), .B(n16973), .ZN(
        n16976) );
  OAI211_X1 U18761 ( .C1(n16978), .C2(n16977), .A(n16976), .B(n16975), .ZN(
        n16979) );
  AOI21_X1 U18762 ( .B1(n16980), .B2(n13329), .A(n16979), .ZN(n16981) );
  OAI21_X1 U18763 ( .B1(n16982), .B2(n18688), .A(n16981), .ZN(P2_U3036) );
  NAND3_X1 U18764 ( .A1(n16983), .A2(n15725), .A3(n16726), .ZN(n16993) );
  NAND2_X1 U18765 ( .A1(n12928), .A2(n19212), .ZN(n16985) );
  NAND2_X1 U18766 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18500), .ZN(n16984) );
  OAI211_X1 U18767 ( .C1(n16986), .C2(n18666), .A(n16985), .B(n16984), .ZN(
        n16989) );
  NOR2_X1 U18768 ( .A1(n16987), .A2(n16991), .ZN(n16988) );
  AOI211_X1 U18769 ( .C1(n16991), .C2(n16990), .A(n16989), .B(n16988), .ZN(
        n16992) );
  OAI211_X1 U18770 ( .C1(n18664), .C2(n16994), .A(n16993), .B(n16992), .ZN(
        P2_U3037) );
  INV_X1 U18771 ( .A(n16995), .ZN(n16996) );
  NAND2_X1 U18772 ( .A1(n16997), .A2(n16996), .ZN(n17028) );
  AOI211_X1 U18773 ( .C1(n17000), .C2(n16999), .A(n16998), .B(n17028), .ZN(
        n17012) );
  OAI22_X1 U18774 ( .A1(n17003), .A2(n17005), .B1(n17002), .B2(n17001), .ZN(
        n17004) );
  NOR2_X1 U18775 ( .A1(n18665), .A2(n17004), .ZN(n17040) );
  OAI21_X1 U18776 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17005), .A(
        n17040), .ZN(n17033) );
  NAND2_X1 U18777 ( .A1(n17033), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17010) );
  OAI21_X1 U18778 ( .B1(n17007), .B2(n17006), .A(n11235), .ZN(n19217) );
  INV_X1 U18779 ( .A(n19217), .ZN(n17008) );
  AOI22_X1 U18780 ( .A1(n12928), .A2(n17008), .B1(n18532), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n17009) );
  OAI211_X1 U18781 ( .C1(n18427), .C2(n18666), .A(n17010), .B(n17009), .ZN(
        n17011) );
  AOI211_X1 U18782 ( .C1(n17013), .C2(n13329), .A(n17012), .B(n17011), .ZN(
        n17014) );
  OAI21_X1 U18783 ( .B1(n17015), .B2(n18688), .A(n17014), .ZN(P2_U3038) );
  INV_X1 U18784 ( .A(n17016), .ZN(n17018) );
  NOR2_X1 U18785 ( .A1(n17018), .A2(n17017), .ZN(n17019) );
  XNOR2_X1 U18786 ( .A(n17020), .B(n17019), .ZN(n17412) );
  NOR2_X1 U18787 ( .A1(n17022), .A2(n17021), .ZN(n17409) );
  INV_X1 U18788 ( .A(n17409), .ZN(n17024) );
  NAND3_X1 U18789 ( .A1(n17024), .A2(n15725), .A3(n17023), .ZN(n17035) );
  INV_X1 U18790 ( .A(n18416), .ZN(n17026) );
  NOR2_X1 U18791 ( .A1(n12281), .A2(n18680), .ZN(n17025) );
  AOI21_X1 U18792 ( .B1(n18685), .B2(n17026), .A(n17025), .ZN(n17027) );
  OAI21_X1 U18793 ( .B1(n17028), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17027), .ZN(n17032) );
  XNOR2_X1 U18794 ( .A(n17030), .B(n17029), .ZN(n19221) );
  NOR2_X1 U18795 ( .A1(n19221), .A2(n18662), .ZN(n17031) );
  AOI211_X1 U18796 ( .C1(n17033), .C2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n17032), .B(n17031), .ZN(n17034) );
  OAI211_X1 U18797 ( .C1(n17412), .C2(n18664), .A(n17035), .B(n17034), .ZN(
        P2_U3039) );
  NAND3_X1 U18798 ( .A1(n17036), .A2(n15725), .A3(n15567), .ZN(n17047) );
  OAI22_X1 U18799 ( .A1(n18666), .A2(n17037), .B1(n12688), .B2(n18680), .ZN(
        n17038) );
  AOI21_X1 U18800 ( .B1(n11076), .B2(n12928), .A(n17038), .ZN(n17046) );
  OR2_X1 U18801 ( .A1(n17039), .A2(n18664), .ZN(n17045) );
  NOR2_X1 U18802 ( .A1(n18675), .A2(n18676), .ZN(n17042) );
  INV_X1 U18803 ( .A(n17040), .ZN(n17041) );
  MUX2_X1 U18804 ( .A(n17042), .B(n17041), .S(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n17043) );
  INV_X1 U18805 ( .A(n17043), .ZN(n17044) );
  NAND4_X1 U18806 ( .A1(n17047), .A2(n17046), .A3(n17045), .A4(n17044), .ZN(
        P2_U3040) );
  INV_X1 U18807 ( .A(n19632), .ZN(n19423) );
  OAI21_X1 U18808 ( .B1(n18662), .B2(n19423), .A(n17048), .ZN(n17049) );
  AOI21_X1 U18809 ( .B1(n17050), .B2(n13329), .A(n17049), .ZN(n17056) );
  AOI22_X1 U18810 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18665), .B1(
        n15725), .B2(n17051), .ZN(n17055) );
  NAND2_X1 U18811 ( .A1(n14681), .A2(n18685), .ZN(n17054) );
  OAI211_X1 U18812 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n18671), .B(n17052), .ZN(n17053) );
  NAND4_X1 U18813 ( .A1(n17056), .A2(n17055), .A3(n17054), .A4(n17053), .ZN(
        P2_U3045) );
  NOR2_X1 U18814 ( .A1(n17058), .A2(n17057), .ZN(n17069) );
  AOI21_X1 U18815 ( .B1(n18517), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n17059), .ZN(n17065) );
  INV_X1 U18816 ( .A(n19424), .ZN(n19421) );
  AOI222_X1 U18817 ( .A1(n17071), .A2(n17061), .B1(n17069), .B2(n17065), .C1(
        n19421), .C2(n17060), .ZN(n17064) );
  NAND2_X1 U18818 ( .A1(n17063), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17062) );
  OAI21_X1 U18819 ( .B1(n17064), .B2(n17063), .A(n17062), .ZN(P2_U3600) );
  INV_X1 U18820 ( .A(n17065), .ZN(n17070) );
  INV_X1 U18821 ( .A(n17071), .ZN(n18696) );
  NOR3_X1 U18822 ( .A1(n17067), .A2(n18696), .A3(n17066), .ZN(n17068) );
  AOI21_X1 U18823 ( .B1(n17070), .B2(n17069), .A(n17068), .ZN(n17074) );
  NAND2_X1 U18824 ( .A1(n17072), .A2(n17071), .ZN(n17073) );
  OAI211_X1 U18825 ( .C1(n19579), .C2(n18706), .A(n17074), .B(n17073), .ZN(
        n17075) );
  MUX2_X1 U18826 ( .A(n10990), .B(n17075), .S(n18661), .Z(P2_U3599) );
  OAI22_X1 U18827 ( .A1(n19431), .A2(n18706), .B1(n17076), .B2(n18696), .ZN(
        n17077) );
  MUX2_X1 U18828 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17077), .S(
        n18661), .Z(P2_U3596) );
  OAI21_X1 U18829 ( .B1(n19709), .B2(n19811), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n17078) );
  NAND2_X1 U18830 ( .A1(n17078), .A2(n19346), .ZN(n17087) );
  INV_X1 U18831 ( .A(n17079), .ZN(n19704) );
  INV_X1 U18832 ( .A(n12097), .ZN(n17080) );
  NOR2_X1 U18833 ( .A1(n17080), .A2(n19364), .ZN(n17081) );
  OAI22_X1 U18834 ( .A1(n17087), .A2(n19704), .B1(n19361), .B2(n17081), .ZN(
        n17082) );
  NAND2_X1 U18835 ( .A1(n19257), .A2(n17436), .ZN(n19352) );
  INV_X1 U18836 ( .A(n19352), .ZN(n19326) );
  NAND2_X1 U18837 ( .A1(n17101), .A2(n19326), .ZN(n17091) );
  NAND2_X1 U18838 ( .A1(n17083), .A2(n19702), .ZN(n19585) );
  OAI22_X1 U18839 ( .A1(n19630), .A2(n19817), .B1(n17091), .B2(n19585), .ZN(
        n17084) );
  AOI21_X1 U18840 ( .B1(n19811), .B2(n19627), .A(n17084), .ZN(n17089) );
  INV_X1 U18841 ( .A(n17091), .ZN(n19809) );
  NOR2_X1 U18842 ( .A1(n19704), .A2(n19809), .ZN(n17086) );
  OAI21_X1 U18843 ( .B1(n12097), .B2(n19809), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17085) );
  NOR2_X2 U18844 ( .A1(n19584), .A2(n19700), .ZN(n19626) );
  NAND2_X1 U18845 ( .A1(n19813), .A2(n19626), .ZN(n17088) );
  OAI211_X1 U18846 ( .C1(n19680), .C2(n17090), .A(n17089), .B(n17088), .ZN(
        P2_U3050) );
  OAI22_X1 U18847 ( .A1(n19817), .A2(n19282), .B1(n17091), .B2(n19281), .ZN(
        n17092) );
  AOI21_X1 U18848 ( .B1(n19811), .B2(n17109), .A(n17092), .ZN(n17094) );
  NAND2_X1 U18849 ( .A1(n19813), .A2(n15143), .ZN(n17093) );
  OAI211_X1 U18850 ( .C1(n19680), .C2(n17095), .A(n17094), .B(n17093), .ZN(
        P2_U3055) );
  INV_X1 U18851 ( .A(n17096), .ZN(n19247) );
  OAI21_X1 U18852 ( .B1(n19788), .B2(n19781), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n17098) );
  NAND2_X1 U18853 ( .A1(n17098), .A2(n19346), .ZN(n17103) );
  NOR2_X1 U18854 ( .A1(n19327), .A2(n17101), .ZN(n17099) );
  NOR2_X1 U18855 ( .A1(n17100), .A2(n17099), .ZN(n19244) );
  NAND2_X1 U18856 ( .A1(n19244), .A2(n17436), .ZN(n17107) );
  NOR2_X1 U18857 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19257), .ZN(
        n19312) );
  NAND2_X1 U18858 ( .A1(n17101), .A2(n19312), .ZN(n17104) );
  INV_X1 U18859 ( .A(n17104), .ZN(n19780) );
  OAI21_X1 U18860 ( .B1(n12105), .B2(n19780), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17102) );
  INV_X1 U18861 ( .A(n17103), .ZN(n17108) );
  NOR2_X1 U18862 ( .A1(n19700), .A2(n17104), .ZN(n17105) );
  AOI211_X1 U18863 ( .C1(n12105), .C2(n19235), .A(n19361), .B(n17105), .ZN(
        n17106) );
  AOI22_X1 U18864 ( .A1(n17109), .A2(n19781), .B1(n19357), .B2(n19780), .ZN(
        n17111) );
  NAND2_X1 U18865 ( .A1(n19788), .A2(n19369), .ZN(n17110) );
  OAI211_X1 U18866 ( .C1(n19786), .C2(n17112), .A(n17111), .B(n17110), .ZN(
        n17113) );
  AOI21_X1 U18867 ( .B1(n15143), .B2(n19782), .A(n17113), .ZN(n17114) );
  INV_X1 U18868 ( .A(n17114), .ZN(P2_U3087) );
  NAND2_X1 U18869 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18773) );
  NAND2_X1 U18870 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18240) );
  INV_X1 U18871 ( .A(n18240), .ZN(n18182) );
  NOR2_X1 U18872 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17885), .ZN(n20104) );
  INV_X1 U18873 ( .A(n20104), .ZN(n17890) );
  NOR2_X1 U18874 ( .A1(n18182), .A2(n17890), .ZN(n17118) );
  NAND2_X1 U18875 ( .A1(n18802), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18769) );
  OR2_X1 U18876 ( .A1(n17115), .A2(n17861), .ZN(n17887) );
  NOR2_X1 U18877 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n17887), .ZN(n17116) );
  NAND2_X1 U18878 ( .A1(n20198), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20787) );
  OAI21_X1 U18879 ( .B1(n17116), .B2(n21244), .A(n18956), .ZN(n18290) );
  NAND2_X1 U18880 ( .A1(n18769), .A2(n18290), .ZN(n18291) );
  AOI221_X1 U18881 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18773), .C1(n17118), 
        .C2(n18773), .A(n18291), .ZN(n18288) );
  NAND3_X1 U18882 ( .A1(n17117), .A2(n21246), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18798) );
  INV_X1 U18883 ( .A(n18798), .ZN(n18774) );
  INV_X1 U18884 ( .A(n17118), .ZN(n17119) );
  OAI21_X1 U18885 ( .B1(n18802), .B2(n21246), .A(n17119), .ZN(n18289) );
  OAI221_X1 U18886 ( .B1(n18774), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18774), .C2(n18289), .A(n18290), .ZN(n18286) );
  AOI22_X1 U18887 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18288), .B1(
        n18286), .B2(n18795), .ZN(P3_U2865) );
  INV_X1 U18888 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17120) );
  INV_X1 U18889 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21649) );
  AOI221_X1 U18890 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n21649), .C1(
        P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18364), 
        .ZN(n21605) );
  INV_X1 U18891 ( .A(BS16), .ZN(n17347) );
  NAND2_X1 U18892 ( .A1(n21654), .A2(n21649), .ZN(n21606) );
  AOI21_X1 U18893 ( .B1(n17347), .B2(n21606), .A(n17121), .ZN(n21601) );
  AOI21_X1 U18894 ( .B1(n17120), .B2(n17121), .A(n21601), .ZN(P3_U3280) );
  AND2_X1 U18895 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n17121), .ZN(P3_U3028) );
  AND2_X1 U18896 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17121), .ZN(P3_U3027) );
  AND2_X1 U18897 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17121), .ZN(P3_U3026) );
  AND2_X1 U18898 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17121), .ZN(P3_U3025) );
  AND2_X1 U18899 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17121), .ZN(P3_U3024) );
  AND2_X1 U18900 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n17121), .ZN(P3_U3023) );
  AND2_X1 U18901 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17121), .ZN(P3_U3022) );
  AND2_X1 U18902 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17121), .ZN(P3_U3021) );
  AND2_X1 U18903 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17121), .ZN(
        P3_U3020) );
  AND2_X1 U18904 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17121), .ZN(
        P3_U3019) );
  AND2_X1 U18905 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17121), .ZN(
        P3_U3018) );
  AND2_X1 U18906 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17121), .ZN(
        P3_U3017) );
  AND2_X1 U18907 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17121), .ZN(
        P3_U3016) );
  AND2_X1 U18908 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17121), .ZN(
        P3_U3015) );
  AND2_X1 U18909 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17121), .ZN(
        P3_U3014) );
  AND2_X1 U18910 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17121), .ZN(
        P3_U3013) );
  AND2_X1 U18911 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17121), .ZN(
        P3_U3012) );
  AND2_X1 U18912 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17121), .ZN(
        P3_U3011) );
  AND2_X1 U18913 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17121), .ZN(
        P3_U3010) );
  AND2_X1 U18914 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17121), .ZN(
        P3_U3009) );
  AND2_X1 U18915 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n17121), .ZN(
        P3_U3008) );
  AND2_X1 U18916 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n17121), .ZN(
        P3_U3007) );
  AND2_X1 U18917 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17121), .ZN(
        P3_U3006) );
  AND2_X1 U18918 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17121), .ZN(
        P3_U3005) );
  AND2_X1 U18919 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n17121), .ZN(
        P3_U3004) );
  AND2_X1 U18920 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n17121), .ZN(
        P3_U3003) );
  AND2_X1 U18921 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n17121), .ZN(
        P3_U3002) );
  AND2_X1 U18922 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n17121), .ZN(
        P3_U3001) );
  AND2_X1 U18923 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n17121), .ZN(
        P3_U3000) );
  AND2_X1 U18924 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n17121), .ZN(
        P3_U2999) );
  AOI21_X1 U18925 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17123)
         );
  INV_X1 U18926 ( .A(n21244), .ZN(n17122) );
  NOR4_X1 U18927 ( .A1(n20789), .A2(n17883), .A3(n21652), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n21201) );
  AOI211_X1 U18928 ( .C1(n18240), .C2(n17123), .A(n17122), .B(n21201), .ZN(
        P3_U2998) );
  NOR2_X1 U18929 ( .A1(n17124), .A2(n18290), .ZN(P3_U2867) );
  NAND2_X1 U18930 ( .A1(n17883), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18281) );
  INV_X1 U18931 ( .A(n18281), .ZN(n18076) );
  NAND2_X1 U18932 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18076), .ZN(n20102) );
  INV_X2 U18933 ( .A(n20102), .ZN(n18353) );
  NOR2_X4 U18934 ( .A1(n18353), .A2(n18337), .ZN(n18348) );
  AND2_X1 U18935 ( .A1(n18348), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U18936 ( .A1(n17884), .A2(n20101), .ZN(n17127) );
  OAI22_X1 U18937 ( .A1(P3_READREQUEST_REG_SCAN_IN), .A2(n17127), .B1(n20108), 
        .B2(n20101), .ZN(n17126) );
  INV_X1 U18938 ( .A(n17126), .ZN(P3_U3298) );
  NOR2_X1 U18939 ( .A1(P3_MEMORYFETCH_REG_SCAN_IN), .A2(n17127), .ZN(n17128)
         );
  NOR2_X1 U18940 ( .A1(n20584), .A2(n17128), .ZN(P3_U3299) );
  AND2_X1 U18941 ( .A1(n21640), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21631) );
  AOI21_X1 U18942 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21631), .A(n17129), 
        .ZN(n17131) );
  INV_X1 U18943 ( .A(n17131), .ZN(n21600) );
  NOR2_X1 U18944 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n21629) );
  OAI21_X1 U18945 ( .B1(BS16), .B2(n21629), .A(n21600), .ZN(n21598) );
  OAI21_X1 U18946 ( .B1(n21600), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n21598), 
        .ZN(n17130) );
  INV_X1 U18947 ( .A(n17130), .ZN(P2_U3591) );
  AND2_X1 U18948 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17131), .ZN(P2_U3208) );
  AND2_X1 U18949 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17131), .ZN(P2_U3207) );
  AND2_X1 U18950 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17132), .ZN(P2_U3206) );
  AND2_X1 U18951 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17131), .ZN(P2_U3205) );
  AND2_X1 U18952 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17132), .ZN(P2_U3204) );
  AND2_X1 U18953 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17131), .ZN(P2_U3203) );
  AND2_X1 U18954 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17132), .ZN(P2_U3202) );
  AND2_X1 U18955 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17132), .ZN(P2_U3201) );
  AND2_X1 U18956 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n17132), .ZN(
        P2_U3200) );
  AND2_X1 U18957 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n17132), .ZN(
        P2_U3199) );
  AND2_X1 U18958 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n17132), .ZN(
        P2_U3198) );
  AND2_X1 U18959 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n17132), .ZN(
        P2_U3197) );
  AND2_X1 U18960 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n17131), .ZN(
        P2_U3196) );
  AND2_X1 U18961 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n17131), .ZN(
        P2_U3195) );
  AND2_X1 U18962 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n17131), .ZN(
        P2_U3194) );
  AND2_X1 U18963 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17131), .ZN(
        P2_U3193) );
  AND2_X1 U18964 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17131), .ZN(
        P2_U3192) );
  AND2_X1 U18965 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17131), .ZN(
        P2_U3191) );
  AND2_X1 U18966 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17131), .ZN(
        P2_U3190) );
  AND2_X1 U18967 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17131), .ZN(
        P2_U3189) );
  AND2_X1 U18968 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17131), .ZN(
        P2_U3188) );
  AND2_X1 U18969 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17131), .ZN(
        P2_U3187) );
  AND2_X1 U18970 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17132), .ZN(
        P2_U3186) );
  AND2_X1 U18971 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17132), .ZN(
        P2_U3185) );
  AND2_X1 U18972 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17132), .ZN(
        P2_U3184) );
  AND2_X1 U18973 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17132), .ZN(
        P2_U3183) );
  AND2_X1 U18974 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17132), .ZN(
        P2_U3182) );
  AND2_X1 U18975 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17132), .ZN(
        P2_U3181) );
  AND2_X1 U18976 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17132), .ZN(
        P2_U3180) );
  AND2_X1 U18977 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17132), .ZN(
        P2_U3179) );
  OAI221_X1 U18978 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(
        P2_STATEBS16_REG_SCAN_IN), .C1(n18711), .C2(n18716), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n17133) );
  AOI21_X1 U18979 ( .B1(n17133), .B2(n19293), .A(n17136), .ZN(P2_U3178) );
  INV_X1 U18980 ( .A(n17134), .ZN(n17135) );
  INV_X1 U18981 ( .A(n17435), .ZN(n17429) );
  NOR2_X1 U18982 ( .A1(n17137), .A2(n17429), .ZN(P2_U3047) );
  AND2_X1 U18983 ( .A1(n17464), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U18984 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17141) );
  NOR4_X1 U18985 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17140) );
  NOR4_X1 U18986 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17139) );
  NOR4_X1 U18987 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17138) );
  NAND4_X1 U18988 ( .A1(n17141), .A2(n17140), .A3(n17139), .A4(n17138), .ZN(
        n17147) );
  NOR4_X1 U18989 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17145) );
  AOI211_X1 U18990 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17144) );
  NOR4_X1 U18991 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17143) );
  NOR4_X1 U18992 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17142) );
  NAND4_X1 U18993 ( .A1(n17145), .A2(n17144), .A3(n17143), .A4(n17142), .ZN(
        n17146) );
  NOR2_X1 U18994 ( .A1(n17147), .A2(n17146), .ZN(n17444) );
  INV_X1 U18995 ( .A(n17444), .ZN(n17442) );
  NOR2_X1 U18996 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17442), .ZN(n17437) );
  OR3_X1 U18997 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17441) );
  INV_X1 U18998 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U18999 ( .A1(n17437), .A2(n17441), .B1(n17442), .B2(n17148), .ZN(
        P2_U2821) );
  INV_X1 U19000 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U19001 ( .A1(n17437), .A2(n12645), .B1(n17442), .B2(n17149), .ZN(
        P2_U2820) );
  INV_X1 U19002 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17150) );
  INV_X1 U19003 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21614) );
  INV_X1 U19004 ( .A(n22329), .ZN(n22328) );
  AND2_X1 U19005 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21619), .ZN(n17192) );
  AOI221_X1 U19006 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n17347), .C1(
        P1_STATE_REG_2__SCAN_IN), .C2(n17347), .A(n17151), .ZN(n21595) );
  AOI21_X1 U19007 ( .B1(n17150), .B2(n17151), .A(n21595), .ZN(P1_U3464) );
  AND2_X1 U19008 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n17151), .ZN(P1_U3193) );
  AND2_X1 U19009 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n17151), .ZN(P1_U3192) );
  AND2_X1 U19010 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n17151), .ZN(P1_U3191) );
  AND2_X1 U19011 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n17151), .ZN(P1_U3190) );
  AND2_X1 U19012 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n17151), .ZN(P1_U3189) );
  AND2_X1 U19013 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n17151), .ZN(P1_U3188) );
  AND2_X1 U19014 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n17151), .ZN(P1_U3187) );
  AND2_X1 U19015 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n17151), .ZN(P1_U3186) );
  AND2_X1 U19016 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n17151), .ZN(
        P1_U3185) );
  AND2_X1 U19017 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n17151), .ZN(
        P1_U3184) );
  AND2_X1 U19018 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n17151), .ZN(
        P1_U3183) );
  AND2_X1 U19019 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n17151), .ZN(
        P1_U3182) );
  AND2_X1 U19020 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n17151), .ZN(
        P1_U3181) );
  AND2_X1 U19021 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n17151), .ZN(
        P1_U3180) );
  AND2_X1 U19022 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n17151), .ZN(
        P1_U3179) );
  AND2_X1 U19023 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n17151), .ZN(
        P1_U3178) );
  AND2_X1 U19024 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n17151), .ZN(
        P1_U3177) );
  AND2_X1 U19025 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n17151), .ZN(
        P1_U3176) );
  AND2_X1 U19026 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n17151), .ZN(
        P1_U3175) );
  AND2_X1 U19027 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n17151), .ZN(
        P1_U3174) );
  AND2_X1 U19028 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n17151), .ZN(
        P1_U3173) );
  AND2_X1 U19029 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n17151), .ZN(
        P1_U3172) );
  AND2_X1 U19030 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n17151), .ZN(
        P1_U3171) );
  AND2_X1 U19031 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n17151), .ZN(
        P1_U3170) );
  AND2_X1 U19032 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n17151), .ZN(
        P1_U3169) );
  AND2_X1 U19033 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n17151), .ZN(
        P1_U3168) );
  AND2_X1 U19034 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n17151), .ZN(
        P1_U3167) );
  AND2_X1 U19035 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n17151), .ZN(
        P1_U3166) );
  AND2_X1 U19036 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n17151), .ZN(
        P1_U3165) );
  AND2_X1 U19037 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n17151), .ZN(
        P1_U3164) );
  AOI21_X1 U19038 ( .B1(n21616), .B2(n21917), .A(n17186), .ZN(n17184) );
  INV_X1 U19039 ( .A(n17152), .ZN(n17155) );
  INV_X1 U19040 ( .A(n17153), .ZN(n17154) );
  OAI211_X1 U19041 ( .C1(n13797), .C2(n17155), .A(n17154), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17158) );
  INV_X1 U19042 ( .A(n17156), .ZN(n17157) );
  OAI21_X1 U19043 ( .B1(n21763), .B2(n17158), .A(n17157), .ZN(n17160) );
  NAND2_X1 U19044 ( .A1(n17158), .A2(n21763), .ZN(n17159) );
  OAI21_X1 U19045 ( .B1(n17161), .B2(n17160), .A(n17159), .ZN(n17162) );
  AOI222_X1 U19046 ( .A1(n21875), .A2(n17163), .B1(n21875), .B2(n17162), .C1(
        n17163), .C2(n17162), .ZN(n17166) );
  INV_X1 U19047 ( .A(n17164), .ZN(n17165) );
  AOI222_X1 U19048 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17166), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17165), .C1(n17166), 
        .C2(n17165), .ZN(n17176) );
  OAI21_X1 U19049 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n17167), .ZN(n17173) );
  INV_X1 U19050 ( .A(n17168), .ZN(n17172) );
  INV_X1 U19051 ( .A(n17169), .ZN(n17170) );
  NAND4_X1 U19052 ( .A1(n17173), .A2(n17172), .A3(n17171), .A4(n17170), .ZN(
        n17174) );
  AOI211_X1 U19053 ( .C1(n17176), .C2(n17191), .A(n17175), .B(n17174), .ZN(
        n21593) );
  NOR2_X1 U19054 ( .A1(n17177), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21265) );
  NAND3_X1 U19055 ( .A1(n10996), .A2(n21265), .A3(n17178), .ZN(n17182) );
  OAI21_X1 U19056 ( .B1(n21667), .B2(n17180), .A(n17179), .ZN(n17181) );
  AND2_X1 U19057 ( .A1(n17182), .A2(n17181), .ZN(n17188) );
  OAI221_X1 U19058 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n21593), 
        .A(n17188), .ZN(n21584) );
  NAND3_X1 U19059 ( .A1(n17184), .A2(n17183), .A3(n21584), .ZN(n21589) );
  AOI21_X1 U19060 ( .B1(n17186), .B2(n17185), .A(n17184), .ZN(n17187) );
  OAI21_X1 U19061 ( .B1(n17188), .B2(n17187), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n17189) );
  OAI21_X1 U19062 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n21589), .A(n17189), 
        .ZN(P1_U3162) );
  NOR2_X1 U19063 ( .A1(n17191), .A2(n17190), .ZN(P1_U3032) );
  AND2_X1 U19064 ( .A1(n19894), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U19065 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17287) );
  AOI21_X1 U19066 ( .B1(n17192), .B2(n17287), .A(n22328), .ZN(P1_U2802) );
  AND2_X1 U19067 ( .A1(n17194), .A2(n17193), .ZN(n17195) );
  NOR2_X1 U19068 ( .A1(n11086), .A2(n17195), .ZN(n21371) );
  AOI222_X1 U19069 ( .A1(n17196), .A2(P1_EBX_REG_4__SCAN_IN), .B1(n19985), 
        .B2(n21371), .C1(n21379), .C2(n19986), .ZN(n17393) );
  OAI22_X1 U19070 ( .A1(n21527), .A2(keyinput_126), .B1(keyinput_127), .B2(
        P1_REIP_REG_20__SCAN_IN), .ZN(n17197) );
  AOI221_X1 U19071 ( .B1(n21527), .B2(keyinput_126), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_127), .A(n17197), .ZN(n17391)
         );
  INV_X1 U19072 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21524) );
  INV_X1 U19073 ( .A(keyinput_125), .ZN(n17282) );
  INV_X1 U19074 ( .A(keyinput_124), .ZN(n17280) );
  INV_X1 U19075 ( .A(keyinput_123), .ZN(n17278) );
  INV_X1 U19076 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n17376) );
  INV_X1 U19077 ( .A(keyinput_119), .ZN(n17272) );
  INV_X1 U19078 ( .A(keyinput_118), .ZN(n17270) );
  INV_X1 U19079 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19963) );
  OAI22_X1 U19080 ( .A1(n19963), .A2(keyinput_114), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_115), .ZN(n17198) );
  AOI221_X1 U19081 ( .B1(n19963), .B2(keyinput_114), .C1(keyinput_115), .C2(
        P1_BYTEENABLE_REG_3__SCAN_IN), .A(n17198), .ZN(n17268) );
  INV_X1 U19082 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n17357) );
  AOI22_X1 U19083 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(keyinput_103), .B1(n17288), 
        .B2(keyinput_102), .ZN(n17199) );
  OAI221_X1 U19084 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_103), .C1(n17288), 
        .C2(keyinput_102), .A(n17199), .ZN(n17252) );
  OAI22_X1 U19085 ( .A1(READY1), .A2(keyinput_100), .B1(READY2), .B2(
        keyinput_101), .ZN(n17200) );
  AOI221_X1 U19086 ( .B1(READY1), .B2(keyinput_100), .C1(keyinput_101), .C2(
        READY2), .A(n17200), .ZN(n17249) );
  INV_X1 U19087 ( .A(NA), .ZN(n21655) );
  INV_X1 U19088 ( .A(keyinput_98), .ZN(n17247) );
  INV_X1 U19089 ( .A(HOLD), .ZN(n21653) );
  OAI22_X1 U19090 ( .A1(DATAI_1_), .A2(keyinput_95), .B1(keyinput_96), .B2(
        DATAI_0_), .ZN(n17201) );
  AOI221_X1 U19091 ( .B1(DATAI_1_), .B2(keyinput_95), .C1(DATAI_0_), .C2(
        keyinput_96), .A(n17201), .ZN(n17244) );
  INV_X1 U19092 ( .A(keyinput_90), .ZN(n17237) );
  INV_X1 U19093 ( .A(DATAI_11_), .ZN(n17323) );
  OAI22_X1 U19094 ( .A1(n17323), .A2(keyinput_85), .B1(keyinput_84), .B2(
        DATAI_12_), .ZN(n17202) );
  AOI221_X1 U19095 ( .B1(n17323), .B2(keyinput_85), .C1(DATAI_12_), .C2(
        keyinput_84), .A(n17202), .ZN(n17235) );
  INV_X1 U19096 ( .A(DATAI_28_), .ZN(n22069) );
  OAI22_X1 U19097 ( .A1(n22069), .A2(keyinput_68), .B1(DATAI_27_), .B2(
        keyinput_69), .ZN(n17203) );
  AOI221_X1 U19098 ( .B1(n22069), .B2(keyinput_68), .C1(keyinput_69), .C2(
        DATAI_27_), .A(n17203), .ZN(n17212) );
  INV_X1 U19099 ( .A(DATAI_29_), .ZN(n22115) );
  INV_X1 U19100 ( .A(keyinput_67), .ZN(n17208) );
  INV_X1 U19101 ( .A(keyinput_66), .ZN(n17206) );
  INV_X1 U19102 ( .A(DATAI_30_), .ZN(n22165) );
  AOI22_X1 U19103 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_64), .B1(
        DATAI_31_), .B2(keyinput_65), .ZN(n17204) );
  OAI221_X1 U19104 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_64), .C1(
        DATAI_31_), .C2(keyinput_65), .A(n17204), .ZN(n17205) );
  OAI221_X1 U19105 ( .B1(DATAI_30_), .B2(n17206), .C1(n22165), .C2(keyinput_66), .A(n17205), .ZN(n17207) );
  OAI221_X1 U19106 ( .B1(DATAI_29_), .B2(keyinput_67), .C1(n22115), .C2(n17208), .A(n17207), .ZN(n17211) );
  INV_X1 U19107 ( .A(DATAI_26_), .ZN(n21977) );
  AOI22_X1 U19108 ( .A1(DATAI_25_), .A2(keyinput_71), .B1(n21977), .B2(
        keyinput_70), .ZN(n17209) );
  OAI221_X1 U19109 ( .B1(DATAI_25_), .B2(keyinput_71), .C1(n21977), .C2(
        keyinput_70), .A(n17209), .ZN(n17210) );
  AOI21_X1 U19110 ( .B1(n17212), .B2(n17211), .A(n17210), .ZN(n17228) );
  INV_X1 U19111 ( .A(DATAI_21_), .ZN(n22118) );
  AOI22_X1 U19112 ( .A1(DATAI_24_), .A2(keyinput_72), .B1(n22118), .B2(
        keyinput_75), .ZN(n17213) );
  OAI221_X1 U19113 ( .B1(DATAI_24_), .B2(keyinput_72), .C1(n22118), .C2(
        keyinput_75), .A(n17213), .ZN(n17216) );
  INV_X1 U19114 ( .A(DATAI_22_), .ZN(n22168) );
  AOI22_X1 U19115 ( .A1(DATAI_23_), .A2(keyinput_73), .B1(n22168), .B2(
        keyinput_74), .ZN(n17214) );
  OAI221_X1 U19116 ( .B1(DATAI_23_), .B2(keyinput_73), .C1(n22168), .C2(
        keyinput_74), .A(n17214), .ZN(n17215) );
  AOI211_X1 U19117 ( .C1(keyinput_76), .C2(DATAI_20_), .A(n17216), .B(n17215), 
        .ZN(n17217) );
  OAI21_X1 U19118 ( .B1(keyinput_76), .B2(DATAI_20_), .A(n17217), .ZN(n17227)
         );
  INV_X1 U19119 ( .A(DATAI_14_), .ZN(n17316) );
  OAI22_X1 U19120 ( .A1(n17316), .A2(keyinput_82), .B1(keyinput_78), .B2(
        DATAI_18_), .ZN(n17218) );
  AOI221_X1 U19121 ( .B1(n17316), .B2(keyinput_82), .C1(DATAI_18_), .C2(
        keyinput_78), .A(n17218), .ZN(n17226) );
  INV_X1 U19122 ( .A(DATAI_15_), .ZN(n17310) );
  OAI22_X1 U19123 ( .A1(n17310), .A2(keyinput_81), .B1(keyinput_80), .B2(
        DATAI_16_), .ZN(n17219) );
  AOI221_X1 U19124 ( .B1(n17310), .B2(keyinput_81), .C1(DATAI_16_), .C2(
        keyinput_80), .A(n17219), .ZN(n17223) );
  INV_X1 U19125 ( .A(DATAI_13_), .ZN(n17221) );
  INV_X1 U19126 ( .A(DATAI_17_), .ZN(n21936) );
  OAI22_X1 U19127 ( .A1(n17221), .A2(keyinput_83), .B1(n21936), .B2(
        keyinput_79), .ZN(n17220) );
  AOI221_X1 U19128 ( .B1(n17221), .B2(keyinput_83), .C1(keyinput_79), .C2(
        n21936), .A(n17220), .ZN(n17222) );
  OAI211_X1 U19129 ( .C1(DATAI_19_), .C2(keyinput_77), .A(n17223), .B(n17222), 
        .ZN(n17224) );
  AOI21_X1 U19130 ( .B1(DATAI_19_), .B2(keyinput_77), .A(n17224), .ZN(n17225)
         );
  OAI211_X1 U19131 ( .C1(n17228), .C2(n17227), .A(n17226), .B(n17225), .ZN(
        n17234) );
  AOI22_X1 U19132 ( .A1(n17325), .A2(keyinput_88), .B1(n17326), .B2(
        keyinput_87), .ZN(n17229) );
  OAI221_X1 U19133 ( .B1(n17325), .B2(keyinput_88), .C1(n17326), .C2(
        keyinput_87), .A(n17229), .ZN(n17233) );
  AOI22_X1 U19134 ( .A1(DATAI_10_), .A2(keyinput_86), .B1(n17231), .B2(
        keyinput_89), .ZN(n17230) );
  OAI221_X1 U19135 ( .B1(DATAI_10_), .B2(keyinput_86), .C1(n17231), .C2(
        keyinput_89), .A(n17230), .ZN(n17232) );
  AOI211_X1 U19136 ( .C1(n17235), .C2(n17234), .A(n17233), .B(n17232), .ZN(
        n17236) );
  AOI221_X1 U19137 ( .B1(DATAI_6_), .B2(keyinput_90), .C1(n17334), .C2(n17237), 
        .A(n17236), .ZN(n17242) );
  AOI22_X1 U19138 ( .A1(n17292), .A2(keyinput_92), .B1(n17293), .B2(
        keyinput_91), .ZN(n17238) );
  OAI221_X1 U19139 ( .B1(n17292), .B2(keyinput_92), .C1(n17293), .C2(
        keyinput_91), .A(n17238), .ZN(n17241) );
  OAI22_X1 U19140 ( .A1(n17337), .A2(keyinput_93), .B1(DATAI_2_), .B2(
        keyinput_94), .ZN(n17239) );
  AOI221_X1 U19141 ( .B1(n17337), .B2(keyinput_93), .C1(keyinput_94), .C2(
        DATAI_2_), .A(n17239), .ZN(n17240) );
  OAI21_X1 U19142 ( .B1(n17242), .B2(n17241), .A(n17240), .ZN(n17243) );
  AOI22_X1 U19143 ( .A1(keyinput_97), .A2(n21653), .B1(n17244), .B2(n17243), 
        .ZN(n17245) );
  OAI21_X1 U19144 ( .B1(n21653), .B2(keyinput_97), .A(n17245), .ZN(n17246) );
  OAI221_X1 U19145 ( .B1(NA), .B2(keyinput_98), .C1(n21655), .C2(n17247), .A(
        n17246), .ZN(n17248) );
  OAI211_X1 U19146 ( .C1(BS16), .C2(keyinput_99), .A(n17249), .B(n17248), .ZN(
        n17250) );
  AOI21_X1 U19147 ( .B1(BS16), .B2(keyinput_99), .A(n17250), .ZN(n17251) );
  OAI22_X1 U19148 ( .A1(n17252), .A2(n17251), .B1(n17357), .B2(keyinput_104), 
        .ZN(n17253) );
  AOI21_X1 U19149 ( .B1(n17357), .B2(keyinput_104), .A(n17253), .ZN(n17260) );
  INV_X1 U19150 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20048) );
  OAI22_X1 U19151 ( .A1(n20048), .A2(keyinput_106), .B1(keyinput_105), .B2(
        P1_M_IO_N_REG_SCAN_IN), .ZN(n17254) );
  AOI221_X1 U19152 ( .B1(n20048), .B2(keyinput_106), .C1(P1_M_IO_N_REG_SCAN_IN), .C2(keyinput_105), .A(n17254), .ZN(n17259) );
  INV_X1 U19153 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21615) );
  AOI22_X1 U19154 ( .A1(n21575), .A2(keyinput_110), .B1(n21615), .B2(
        keyinput_107), .ZN(n17255) );
  OAI221_X1 U19155 ( .B1(n21575), .B2(keyinput_110), .C1(n21615), .C2(
        keyinput_107), .A(n17255), .ZN(n17258) );
  AOI22_X1 U19156 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_109), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_108), .ZN(n17256) );
  OAI221_X1 U19157 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_109), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_108), .A(n17256), .ZN(n17257)
         );
  AOI211_X1 U19158 ( .C1(n17260), .C2(n17259), .A(n17258), .B(n17257), .ZN(
        n17263) );
  AOI22_X1 U19159 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput_111), .B1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_113), .ZN(n17261) );
  OAI221_X1 U19160 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_111), .C1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_113), .A(n17261), .ZN(
        n17262) );
  AOI211_X1 U19161 ( .C1(P1_BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_112), .A(
        n17263), .B(n17262), .ZN(n17264) );
  OAI21_X1 U19162 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_112), .A(
        n17264), .ZN(n17267) );
  AOI22_X1 U19163 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_117), .B1(
        n19947), .B2(keyinput_116), .ZN(n17265) );
  OAI221_X1 U19164 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_117), .C1(
        n19947), .C2(keyinput_116), .A(n17265), .ZN(n17266) );
  AOI21_X1 U19165 ( .B1(n17268), .B2(n17267), .A(n17266), .ZN(n17269) );
  AOI221_X1 U19166 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_118), .C1(
        n19943), .C2(n17270), .A(n17269), .ZN(n17271) );
  AOI221_X1 U19167 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_119), .C1(
        n17376), .C2(n17272), .A(n17271), .ZN(n17275) );
  AOI22_X1 U19168 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(keyinput_122), .B1(
        n17284), .B2(keyinput_120), .ZN(n17273) );
  OAI221_X1 U19169 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_122), .C1(
        n17284), .C2(keyinput_120), .A(n17273), .ZN(n17274) );
  AOI211_X1 U19170 ( .C1(P1_REIP_REG_26__SCAN_IN), .C2(keyinput_121), .A(
        n17275), .B(n17274), .ZN(n17276) );
  OAI21_X1 U19171 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_121), .A(n17276), .ZN(n17277) );
  OAI221_X1 U19172 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_123), .C1(
        n16096), .C2(n17278), .A(n17277), .ZN(n17279) );
  OAI221_X1 U19173 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_124), .C1(
        n21535), .C2(n17280), .A(n17279), .ZN(n17281) );
  OAI221_X1 U19174 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_125), .C1(
        n21524), .C2(n17282), .A(n17281), .ZN(n17390) );
  INV_X1 U19175 ( .A(keyinput_61), .ZN(n17385) );
  INV_X1 U19176 ( .A(keyinput_60), .ZN(n17383) );
  INV_X1 U19177 ( .A(keyinput_59), .ZN(n17381) );
  OAI22_X1 U19178 ( .A1(n17284), .A2(keyinput_56), .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_58), .ZN(n17283) );
  AOI221_X1 U19179 ( .B1(n17284), .B2(keyinput_56), .C1(keyinput_58), .C2(
        P1_REIP_REG_25__SCAN_IN), .A(n17283), .ZN(n17378) );
  INV_X1 U19180 ( .A(keyinput_55), .ZN(n17375) );
  INV_X1 U19181 ( .A(keyinput_54), .ZN(n17373) );
  INV_X1 U19182 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19970) );
  OAI22_X1 U19183 ( .A1(n19970), .A2(keyinput_48), .B1(n20100), .B2(
        keyinput_47), .ZN(n17285) );
  AOI221_X1 U19184 ( .B1(n19970), .B2(keyinput_48), .C1(keyinput_47), .C2(
        n20100), .A(n17285), .ZN(n17365) );
  OAI22_X1 U19185 ( .A1(n17288), .A2(keyinput_38), .B1(n17287), .B2(
        keyinput_39), .ZN(n17286) );
  AOI221_X1 U19186 ( .B1(n17288), .B2(keyinput_38), .C1(keyinput_39), .C2(
        n17287), .A(n17286), .ZN(n17353) );
  INV_X1 U19187 ( .A(READY2), .ZN(n17351) );
  INV_X1 U19188 ( .A(keyinput_34), .ZN(n17345) );
  AOI22_X1 U19189 ( .A1(DATAI_0_), .A2(keyinput_32), .B1(n17290), .B2(
        keyinput_31), .ZN(n17289) );
  OAI221_X1 U19190 ( .B1(DATAI_0_), .B2(keyinput_32), .C1(n17290), .C2(
        keyinput_31), .A(n17289), .ZN(n17342) );
  OAI22_X1 U19191 ( .A1(n17293), .A2(keyinput_27), .B1(n17292), .B2(
        keyinput_28), .ZN(n17291) );
  AOI221_X1 U19192 ( .B1(n17293), .B2(keyinput_27), .C1(keyinput_28), .C2(
        n17292), .A(n17291), .ZN(n17340) );
  INV_X1 U19193 ( .A(keyinput_26), .ZN(n17335) );
  INV_X1 U19194 ( .A(DATAI_20_), .ZN(n22071) );
  INV_X1 U19195 ( .A(DATAI_23_), .ZN(n22218) );
  AOI22_X1 U19196 ( .A1(n22071), .A2(keyinput_12), .B1(n22218), .B2(keyinput_9), .ZN(n17294) );
  OAI221_X1 U19197 ( .B1(n22071), .B2(keyinput_12), .C1(n22218), .C2(
        keyinput_9), .A(n17294), .ZN(n17298) );
  OAI22_X1 U19198 ( .A1(n22168), .A2(keyinput_10), .B1(DATAI_24_), .B2(
        keyinput_8), .ZN(n17295) );
  AOI221_X1 U19199 ( .B1(n22168), .B2(keyinput_10), .C1(keyinput_8), .C2(
        DATAI_24_), .A(n17295), .ZN(n17296) );
  OAI21_X1 U19200 ( .B1(keyinput_11), .B2(DATAI_21_), .A(n17296), .ZN(n17297)
         );
  AOI211_X1 U19201 ( .C1(keyinput_11), .C2(DATAI_21_), .A(n17298), .B(n17297), 
        .ZN(n17320) );
  INV_X1 U19202 ( .A(keyinput_3), .ZN(n17303) );
  INV_X1 U19203 ( .A(keyinput_2), .ZN(n17301) );
  OAI22_X1 U19204 ( .A1(DATAI_31_), .A2(keyinput_1), .B1(
        P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_0), .ZN(n17299) );
  AOI221_X1 U19205 ( .B1(DATAI_31_), .B2(keyinput_1), .C1(keyinput_0), .C2(
        P1_MEMORYFETCH_REG_SCAN_IN), .A(n17299), .ZN(n17300) );
  AOI221_X1 U19206 ( .B1(DATAI_30_), .B2(n17301), .C1(n22165), .C2(keyinput_2), 
        .A(n17300), .ZN(n17302) );
  AOI221_X1 U19207 ( .B1(DATAI_29_), .B2(keyinput_3), .C1(n22115), .C2(n17303), 
        .A(n17302), .ZN(n17308) );
  INV_X1 U19208 ( .A(DATAI_27_), .ZN(n22023) );
  AOI22_X1 U19209 ( .A1(n22023), .A2(keyinput_5), .B1(n22069), .B2(keyinput_4), 
        .ZN(n17304) );
  OAI221_X1 U19210 ( .B1(n22023), .B2(keyinput_5), .C1(n22069), .C2(keyinput_4), .A(n17304), .ZN(n17307) );
  OAI22_X1 U19211 ( .A1(n21977), .A2(keyinput_6), .B1(DATAI_25_), .B2(
        keyinput_7), .ZN(n17305) );
  AOI221_X1 U19212 ( .B1(n21977), .B2(keyinput_6), .C1(keyinput_7), .C2(
        DATAI_25_), .A(n17305), .ZN(n17306) );
  OAI21_X1 U19213 ( .B1(n17308), .B2(n17307), .A(n17306), .ZN(n17319) );
  AOI22_X1 U19214 ( .A1(DATAI_13_), .A2(keyinput_19), .B1(n17310), .B2(
        keyinput_17), .ZN(n17309) );
  OAI221_X1 U19215 ( .B1(DATAI_13_), .B2(keyinput_19), .C1(n17310), .C2(
        keyinput_17), .A(n17309), .ZN(n17318) );
  INV_X1 U19216 ( .A(DATAI_18_), .ZN(n21980) );
  OAI22_X1 U19217 ( .A1(n21980), .A2(keyinput_14), .B1(keyinput_15), .B2(
        DATAI_17_), .ZN(n17311) );
  AOI221_X1 U19218 ( .B1(n21980), .B2(keyinput_14), .C1(DATAI_17_), .C2(
        keyinput_15), .A(n17311), .ZN(n17315) );
  INV_X1 U19219 ( .A(DATAI_16_), .ZN(n21746) );
  INV_X1 U19220 ( .A(DATAI_19_), .ZN(n22026) );
  AOI22_X1 U19221 ( .A1(n21746), .A2(keyinput_16), .B1(n22026), .B2(
        keyinput_13), .ZN(n17312) );
  OAI221_X1 U19222 ( .B1(n21746), .B2(keyinput_16), .C1(n22026), .C2(
        keyinput_13), .A(n17312), .ZN(n17313) );
  AOI21_X1 U19223 ( .B1(keyinput_18), .B2(n17316), .A(n17313), .ZN(n17314) );
  OAI211_X1 U19224 ( .C1(keyinput_18), .C2(n17316), .A(n17315), .B(n17314), 
        .ZN(n17317) );
  AOI211_X1 U19225 ( .C1(n17320), .C2(n17319), .A(n17318), .B(n17317), .ZN(
        n17332) );
  AOI22_X1 U19226 ( .A1(n17323), .A2(keyinput_21), .B1(n17322), .B2(
        keyinput_20), .ZN(n17321) );
  OAI221_X1 U19227 ( .B1(n17323), .B2(keyinput_21), .C1(n17322), .C2(
        keyinput_20), .A(n17321), .ZN(n17331) );
  OAI22_X1 U19228 ( .A1(n17326), .A2(keyinput_23), .B1(n17325), .B2(
        keyinput_24), .ZN(n17324) );
  AOI221_X1 U19229 ( .B1(n17326), .B2(keyinput_23), .C1(keyinput_24), .C2(
        n17325), .A(n17324), .ZN(n17330) );
  OAI22_X1 U19230 ( .A1(n17328), .A2(keyinput_22), .B1(DATAI_7_), .B2(
        keyinput_25), .ZN(n17327) );
  AOI221_X1 U19231 ( .B1(n17328), .B2(keyinput_22), .C1(keyinput_25), .C2(
        DATAI_7_), .A(n17327), .ZN(n17329) );
  OAI211_X1 U19232 ( .C1(n17332), .C2(n17331), .A(n17330), .B(n17329), .ZN(
        n17333) );
  OAI221_X1 U19233 ( .B1(DATAI_6_), .B2(n17335), .C1(n17334), .C2(keyinput_26), 
        .A(n17333), .ZN(n17339) );
  AOI22_X1 U19234 ( .A1(DATAI_2_), .A2(keyinput_30), .B1(n17337), .B2(
        keyinput_29), .ZN(n17336) );
  OAI221_X1 U19235 ( .B1(DATAI_2_), .B2(keyinput_30), .C1(n17337), .C2(
        keyinput_29), .A(n17336), .ZN(n17338) );
  AOI21_X1 U19236 ( .B1(n17340), .B2(n17339), .A(n17338), .ZN(n17341) );
  OAI22_X1 U19237 ( .A1(keyinput_33), .A2(n21653), .B1(n17342), .B2(n17341), 
        .ZN(n17343) );
  AOI21_X1 U19238 ( .B1(keyinput_33), .B2(n21653), .A(n17343), .ZN(n17344) );
  AOI221_X1 U19239 ( .B1(NA), .B2(keyinput_34), .C1(n21655), .C2(n17345), .A(
        n17344), .ZN(n17349) );
  AOI22_X1 U19240 ( .A1(READY1), .A2(keyinput_36), .B1(n17347), .B2(
        keyinput_35), .ZN(n17346) );
  OAI221_X1 U19241 ( .B1(READY1), .B2(keyinput_36), .C1(n17347), .C2(
        keyinput_35), .A(n17346), .ZN(n17348) );
  AOI211_X1 U19242 ( .C1(n17351), .C2(keyinput_37), .A(n17349), .B(n17348), 
        .ZN(n17350) );
  OAI21_X1 U19243 ( .B1(n17351), .B2(keyinput_37), .A(n17350), .ZN(n17352) );
  AOI22_X1 U19244 ( .A1(n17353), .A2(n17352), .B1(P1_D_C_N_REG_SCAN_IN), .B2(
        keyinput_42), .ZN(n17354) );
  OAI21_X1 U19245 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_42), .A(n17354), 
        .ZN(n17363) );
  AOI22_X1 U19246 ( .A1(n17357), .A2(keyinput_40), .B1(keyinput_41), .B2(
        n17356), .ZN(n17355) );
  OAI221_X1 U19247 ( .B1(n17357), .B2(keyinput_40), .C1(n17356), .C2(
        keyinput_41), .A(n17355), .ZN(n17362) );
  OAI22_X1 U19248 ( .A1(n21575), .A2(keyinput_46), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_44), .ZN(n17358) );
  AOI221_X1 U19249 ( .B1(n21575), .B2(keyinput_46), .C1(keyinput_44), .C2(
        P1_STATEBS16_REG_SCAN_IN), .A(n17358), .ZN(n17361) );
  OAI22_X1 U19250 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_43), .B1(
        P1_MORE_REG_SCAN_IN), .B2(keyinput_45), .ZN(n17359) );
  AOI221_X1 U19251 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_43), 
        .C1(keyinput_45), .C2(P1_MORE_REG_SCAN_IN), .A(n17359), .ZN(n17360) );
  OAI211_X1 U19252 ( .C1(n17363), .C2(n17362), .A(n17361), .B(n17360), .ZN(
        n17364) );
  OAI211_X1 U19253 ( .C1(P1_BYTEENABLE_REG_1__SCAN_IN), .C2(keyinput_49), .A(
        n17365), .B(n17364), .ZN(n17366) );
  AOI21_X1 U19254 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_49), .A(
        n17366), .ZN(n17371) );
  AOI22_X1 U19255 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_50), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_51), .ZN(n17367) );
  OAI221_X1 U19256 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_50), .C1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_51), .A(n17367), .ZN(
        n17370) );
  OAI22_X1 U19257 ( .A1(n19947), .A2(keyinput_52), .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_53), .ZN(n17368) );
  AOI221_X1 U19258 ( .B1(n19947), .B2(keyinput_52), .C1(keyinput_53), .C2(
        P1_REIP_REG_30__SCAN_IN), .A(n17368), .ZN(n17369) );
  OAI21_X1 U19259 ( .B1(n17371), .B2(n17370), .A(n17369), .ZN(n17372) );
  OAI221_X1 U19260 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n17373), .C1(n19943), 
        .C2(keyinput_54), .A(n17372), .ZN(n17374) );
  OAI221_X1 U19261 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_55), .C1(
        n17376), .C2(n17375), .A(n17374), .ZN(n17377) );
  OAI211_X1 U19262 ( .C1(P1_REIP_REG_26__SCAN_IN), .C2(keyinput_57), .A(n17378), .B(n17377), .ZN(n17379) );
  AOI21_X1 U19263 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_57), .A(n17379), 
        .ZN(n17380) );
  AOI221_X1 U19264 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(keyinput_59), .C1(
        n16096), .C2(n17381), .A(n17380), .ZN(n17382) );
  AOI221_X1 U19265 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_60), .C1(
        n21535), .C2(n17383), .A(n17382), .ZN(n17384) );
  AOI221_X1 U19266 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_61), .C1(
        n21524), .C2(n17385), .A(n17384), .ZN(n17389) );
  INV_X1 U19267 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U19268 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_62), .B1(n17387), .B2(keyinput_63), .ZN(n17386) );
  OAI221_X1 U19269 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_62), .C1(
        n17387), .C2(keyinput_63), .A(n17386), .ZN(n17388) );
  AOI211_X1 U19270 ( .C1(n17391), .C2(n17390), .A(n17389), .B(n17388), .ZN(
        n17392) );
  XNOR2_X1 U19271 ( .A(n17393), .B(n17392), .ZN(P1_U2868) );
  INV_X1 U19272 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17395) );
  OAI22_X1 U19273 ( .A1(n18371), .A2(n17395), .B1(n18711), .B2(n17394), .ZN(
        P2_U2816) );
  AOI22_X1 U19274 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n18532), .B1(n17407), 
        .B2(n17396), .ZN(n17405) );
  INV_X1 U19275 ( .A(n17397), .ZN(n17399) );
  XNOR2_X1 U19276 ( .A(n17398), .B(n17399), .ZN(n18683) );
  OAI21_X1 U19277 ( .B1(n17401), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n17400), .ZN(n18689) );
  OAI22_X1 U19278 ( .A1(n18689), .A2(n17408), .B1(n17410), .B2(n17402), .ZN(
        n17403) );
  AOI21_X1 U19279 ( .B1(n12546), .B2(n18683), .A(n17403), .ZN(n17404) );
  OAI211_X1 U19280 ( .C1(n17406), .C2(n17417), .A(n17405), .B(n17404), .ZN(
        P2_U3009) );
  AOI22_X1 U19281 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n18532), .B1(n17407), 
        .B2(n18412), .ZN(n17416) );
  NOR2_X1 U19282 ( .A1(n17409), .A2(n17408), .ZN(n17414) );
  OAI22_X1 U19283 ( .A1(n17412), .A2(n17411), .B1(n17410), .B2(n18416), .ZN(
        n17413) );
  AOI21_X1 U19284 ( .B1(n17414), .B2(n17023), .A(n17413), .ZN(n17415) );
  OAI211_X1 U19285 ( .C1(n17418), .C2(n17417), .A(n17416), .B(n17415), .ZN(
        P2_U3007) );
  NOR2_X1 U19286 ( .A1(n17420), .A2(n17419), .ZN(n18703) );
  NOR2_X1 U19287 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12654), .ZN(
        n17421) );
  AOI211_X1 U19288 ( .C1(n19694), .C2(n18372), .A(n18703), .B(n17421), .ZN(
        n17422) );
  AOI22_X1 U19289 ( .A1(n17435), .A2(n19353), .B1(n17422), .B2(n17429), .ZN(
        P2_U3605) );
  NAND2_X1 U19290 ( .A1(n19421), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19224) );
  INV_X1 U19291 ( .A(n19224), .ZN(n17424) );
  INV_X1 U19292 ( .A(n18372), .ZN(n17423) );
  AOI21_X1 U19293 ( .B1(n17424), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n17423), 
        .ZN(n17431) );
  NAND2_X1 U19294 ( .A1(n17424), .A2(n19579), .ZN(n19328) );
  INV_X1 U19295 ( .A(n19328), .ZN(n17425) );
  AOI222_X1 U19296 ( .A1(n19578), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n17426), 
        .B2(n17431), .C1(n19346), .C2(n17425), .ZN(n17427) );
  AOI22_X1 U19297 ( .A1(n17435), .A2(n19257), .B1(n17427), .B2(n17429), .ZN(
        P2_U3603) );
  OR2_X1 U19298 ( .A1(n19355), .A2(n21597), .ZN(n19343) );
  NAND2_X1 U19299 ( .A1(n19424), .A2(n19343), .ZN(n17428) );
  AOI22_X1 U19300 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19632), .B1(n17431), 
        .B2(n17428), .ZN(n17430) );
  AOI22_X1 U19301 ( .A1(n17435), .A2(n14986), .B1(n17430), .B2(n17429), .ZN(
        P2_U3604) );
  INV_X1 U19302 ( .A(n19431), .ZN(n19359) );
  AOI22_X1 U19303 ( .A1(n19359), .A2(n17431), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19531), .ZN(n17434) );
  AOI21_X1 U19304 ( .B1(n19248), .B2(n19298), .A(n19343), .ZN(n17432) );
  NOR2_X1 U19305 ( .A1(n17435), .A2(n17432), .ZN(n17433) );
  AOI22_X1 U19306 ( .A1(n17436), .A2(n17435), .B1(n17434), .B2(n17433), .ZN(
        P2_U3602) );
  INV_X1 U19307 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21599) );
  NAND2_X1 U19308 ( .A1(n17437), .A2(n21599), .ZN(n17440) );
  OAI21_X1 U19309 ( .B1(n12645), .B2(n12646), .A(n17444), .ZN(n17438) );
  OAI21_X1 U19310 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17444), .A(n17438), 
        .ZN(n17439) );
  OAI221_X1 U19311 ( .B1(n17440), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17440), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17439), .ZN(P2_U2822) );
  INV_X1 U19312 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17443) );
  OAI221_X1 U19313 ( .B1(n17444), .B2(n17443), .C1(n17442), .C2(n17441), .A(
        n17440), .ZN(P2_U2823) );
  OAI22_X1 U19314 ( .A1(n17499), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n17495), .ZN(n17445) );
  INV_X1 U19315 ( .A(n17445), .ZN(P2_U3611) );
  INV_X1 U19316 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17446) );
  AOI22_X1 U19317 ( .A1(n17495), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17446), 
        .B2(n17499), .ZN(P2_U3608) );
  AOI21_X1 U19318 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n21600), .ZN(n17447) );
  INV_X1 U19319 ( .A(n17447), .ZN(P2_U2815) );
  AOI22_X1 U19320 ( .A1(n17473), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17449) );
  OAI21_X1 U19321 ( .B1(n19685), .B2(n17475), .A(n17449), .ZN(P2_U2951) );
  INV_X1 U19322 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U19323 ( .A1(n17473), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17450) );
  OAI21_X1 U19324 ( .B1(n17451), .B2(n17475), .A(n17450), .ZN(P2_U2950) );
  INV_X1 U19325 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U19326 ( .A1(n17473), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17452) );
  OAI21_X1 U19327 ( .B1(n17453), .B2(n17475), .A(n17452), .ZN(P2_U2949) );
  INV_X1 U19328 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U19329 ( .A1(n17465), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17454) );
  OAI21_X1 U19330 ( .B1(n17455), .B2(n17475), .A(n17454), .ZN(P2_U2948) );
  AOI22_X1 U19331 ( .A1(n17473), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17456) );
  OAI21_X1 U19332 ( .B1(n19480), .B2(n17475), .A(n17456), .ZN(P2_U2947) );
  INV_X1 U19333 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U19334 ( .A1(n17465), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17457) );
  OAI21_X1 U19335 ( .B1(n17458), .B2(n17475), .A(n17457), .ZN(P2_U2946) );
  INV_X1 U19336 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U19337 ( .A1(n17465), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17459) );
  OAI21_X1 U19338 ( .B1(n17460), .B2(n17475), .A(n17459), .ZN(P2_U2945) );
  INV_X1 U19339 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19219) );
  AOI22_X1 U19340 ( .A1(n17465), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17461) );
  OAI21_X1 U19341 ( .B1(n19219), .B2(n17475), .A(n17461), .ZN(P2_U2944) );
  INV_X1 U19342 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19216) );
  AOI22_X1 U19343 ( .A1(n17465), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17462) );
  OAI21_X1 U19344 ( .B1(n19216), .B2(n17475), .A(n17462), .ZN(P2_U2943) );
  AOI22_X1 U19345 ( .A1(n17473), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17463) );
  OAI21_X1 U19346 ( .B1(n19214), .B2(n17475), .A(n17463), .ZN(P2_U2942) );
  INV_X1 U19347 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17467) );
  AOI22_X1 U19348 ( .A1(n17465), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17466) );
  OAI21_X1 U19349 ( .B1(n17467), .B2(n17475), .A(n17466), .ZN(P2_U2941) );
  AOI22_X1 U19350 ( .A1(n17473), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17468) );
  OAI21_X1 U19351 ( .B1(n19206), .B2(n17475), .A(n17468), .ZN(P2_U2940) );
  INV_X1 U19352 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19201) );
  AOI22_X1 U19353 ( .A1(n17473), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17469) );
  OAI21_X1 U19354 ( .B1(n19201), .B2(n17475), .A(n17469), .ZN(P2_U2939) );
  INV_X1 U19355 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n17471) );
  AOI22_X1 U19356 ( .A1(n17473), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17470) );
  OAI21_X1 U19357 ( .B1(n17471), .B2(n17475), .A(n17470), .ZN(P2_U2938) );
  INV_X1 U19358 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19195) );
  AOI22_X1 U19359 ( .A1(n17473), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17472) );
  OAI21_X1 U19360 ( .B1(n19195), .B2(n17475), .A(n17472), .ZN(P2_U2937) );
  AOI22_X1 U19361 ( .A1(n17473), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17464), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17474) );
  OAI21_X1 U19362 ( .B1(n17476), .B2(n17475), .A(n17474), .ZN(P2_U2936) );
  AOI21_X1 U19363 ( .B1(n17478), .B2(n17477), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n17479) );
  AOI21_X1 U19364 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n17495), .A(n17479), 
        .ZN(P2_U2817) );
  NOR2_X1 U19365 ( .A1(n21640), .A2(n17499), .ZN(n21627) );
  INV_X2 U19366 ( .A(n21627), .ZN(n21638) );
  OAI222_X1 U19367 ( .A1(n21638), .A2(n12646), .B1(n19821), .B2(n17495), .C1(
        n17480), .C2(n17496), .ZN(P2_U3212) );
  INV_X1 U19368 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n17481) );
  OAI222_X1 U19369 ( .A1(n17496), .A2(n17482), .B1(n17481), .B2(n17495), .C1(
        n17480), .C2(n21638), .ZN(P2_U3213) );
  INV_X1 U19370 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n17483) );
  OAI222_X1 U19371 ( .A1(n17496), .A2(n12266), .B1(n17483), .B2(n17495), .C1(
        n17482), .C2(n21638), .ZN(P2_U3214) );
  INV_X1 U19372 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19825) );
  OAI222_X1 U19373 ( .A1(n17496), .A2(n12270), .B1(n19825), .B2(n17495), .C1(
        n12266), .C2(n21638), .ZN(P2_U3215) );
  INV_X1 U19374 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19827) );
  OAI222_X1 U19375 ( .A1(n17496), .A2(n12688), .B1(n19827), .B2(n17495), .C1(
        n12270), .C2(n21638), .ZN(P2_U3216) );
  INV_X1 U19376 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19829) );
  OAI222_X1 U19377 ( .A1(n17496), .A2(n12281), .B1(n19829), .B2(n17495), .C1(
        n12688), .C2(n21638), .ZN(P2_U3217) );
  INV_X1 U19378 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19831) );
  OAI222_X1 U19379 ( .A1(n17496), .A2(n12710), .B1(n19831), .B2(n17495), .C1(
        n12281), .C2(n21638), .ZN(P2_U3218) );
  INV_X1 U19380 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19834) );
  OAI222_X1 U19381 ( .A1(n17496), .A2(n16767), .B1(n19834), .B2(n17495), .C1(
        n12710), .C2(n21638), .ZN(P2_U3219) );
  INV_X1 U19382 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19836) );
  OAI222_X1 U19383 ( .A1(n21638), .A2(n16767), .B1(n19836), .B2(n17495), .C1(
        n16747), .C2(n17496), .ZN(P2_U3220) );
  INV_X1 U19384 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19838) );
  OAI222_X1 U19385 ( .A1(n21638), .A2(n16747), .B1(n19838), .B2(n17495), .C1(
        n18433), .C2(n17496), .ZN(P2_U3221) );
  INV_X1 U19386 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19840) );
  OAI222_X1 U19387 ( .A1(n21638), .A2(n18433), .B1(n19840), .B2(n17495), .C1(
        n17484), .C2(n17496), .ZN(P2_U3222) );
  INV_X1 U19388 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19842) );
  OAI222_X1 U19389 ( .A1(n21638), .A2(n17484), .B1(n19842), .B2(n17495), .C1(
        n17485), .C2(n17496), .ZN(P2_U3223) );
  INV_X1 U19390 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19844) );
  OAI222_X1 U19391 ( .A1(n21638), .A2(n17485), .B1(n19844), .B2(n17495), .C1(
        n16697), .C2(n17496), .ZN(P2_U3224) );
  INV_X1 U19392 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19846) );
  OAI222_X1 U19393 ( .A1(n21638), .A2(n16697), .B1(n19846), .B2(n17495), .C1(
        n12844), .C2(n17496), .ZN(P2_U3225) );
  INV_X1 U19394 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19848) );
  OAI222_X1 U19395 ( .A1(n21638), .A2(n12844), .B1(n19848), .B2(n17495), .C1(
        n17486), .C2(n17496), .ZN(P2_U3226) );
  INV_X1 U19396 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19850) );
  OAI222_X1 U19397 ( .A1(n21638), .A2(n17486), .B1(n19850), .B2(n17495), .C1(
        n18498), .C2(n17496), .ZN(P2_U3227) );
  INV_X1 U19398 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19852) );
  OAI222_X1 U19399 ( .A1(n21638), .A2(n18498), .B1(n19852), .B2(n17495), .C1(
        n18512), .C2(n17496), .ZN(P2_U3228) );
  INV_X1 U19400 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19854) );
  OAI222_X1 U19401 ( .A1(n17496), .A2(n17487), .B1(n19854), .B2(n17495), .C1(
        n18512), .C2(n21638), .ZN(P2_U3229) );
  INV_X1 U19402 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19856) );
  OAI222_X1 U19403 ( .A1(n21638), .A2(n17487), .B1(n19856), .B2(n17495), .C1(
        n17488), .C2(n17496), .ZN(P2_U3230) );
  INV_X1 U19404 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19858) );
  OAI222_X1 U19405 ( .A1(n17496), .A2(n13296), .B1(n19858), .B2(n17495), .C1(
        n17488), .C2(n21638), .ZN(P2_U3231) );
  INV_X1 U19406 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19860) );
  OAI222_X1 U19407 ( .A1(n17496), .A2(n17489), .B1(n19860), .B2(n17495), .C1(
        n13296), .C2(n21638), .ZN(P2_U3232) );
  INV_X1 U19408 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19862) );
  OAI222_X1 U19409 ( .A1(n17496), .A2(n12331), .B1(n19862), .B2(n17495), .C1(
        n17489), .C2(n21638), .ZN(P2_U3233) );
  INV_X1 U19410 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19864) );
  OAI222_X1 U19411 ( .A1(n17496), .A2(n17490), .B1(n19864), .B2(n17495), .C1(
        n12331), .C2(n21638), .ZN(P2_U3234) );
  INV_X1 U19412 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19866) );
  OAI222_X1 U19413 ( .A1(n17496), .A2(n16603), .B1(n19866), .B2(n17495), .C1(
        n17490), .C2(n21638), .ZN(P2_U3235) );
  INV_X1 U19414 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19868) );
  OAI222_X1 U19415 ( .A1(n21638), .A2(n16603), .B1(n19868), .B2(n17495), .C1(
        n17491), .C2(n17496), .ZN(P2_U3236) );
  INV_X1 U19416 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19870) );
  OAI222_X1 U19417 ( .A1(n17496), .A2(n17492), .B1(n19870), .B2(n17495), .C1(
        n17491), .C2(n21638), .ZN(P2_U3237) );
  INV_X1 U19418 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19872) );
  OAI222_X1 U19419 ( .A1(n21638), .A2(n17492), .B1(n19872), .B2(n17495), .C1(
        n17493), .C2(n17496), .ZN(P2_U3238) );
  INV_X1 U19420 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19874) );
  OAI222_X1 U19421 ( .A1(n17496), .A2(n17494), .B1(n19874), .B2(n17495), .C1(
        n17493), .C2(n21638), .ZN(P2_U3239) );
  INV_X1 U19422 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19876) );
  OAI222_X1 U19423 ( .A1(n21638), .A2(n17494), .B1(n19876), .B2(n17495), .C1(
        n18626), .C2(n17496), .ZN(P2_U3240) );
  INV_X1 U19424 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19879) );
  OAI222_X1 U19425 ( .A1(n17496), .A2(n12877), .B1(n19879), .B2(n17495), .C1(
        n18626), .C2(n21638), .ZN(P2_U3241) );
  OAI22_X1 U19426 ( .A1(n17499), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n17495), .ZN(n17497) );
  INV_X1 U19427 ( .A(n17497), .ZN(P2_U3588) );
  OAI22_X1 U19428 ( .A1(n17499), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n17495), .ZN(n17498) );
  INV_X1 U19429 ( .A(n17498), .ZN(P2_U3587) );
  MUX2_X1 U19430 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n17499), .Z(P2_U3586) );
  OAI22_X1 U19431 ( .A1(n17499), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n17495), .ZN(n17500) );
  INV_X1 U19432 ( .A(n17500), .ZN(P2_U3585) );
  AND2_X1 U19433 ( .A1(n17874), .A2(n17635), .ZN(n17528) );
  NAND2_X1 U19434 ( .A1(n20768), .A2(n17874), .ZN(n17880) );
  NOR2_X1 U19435 ( .A1(n17501), .A2(n17880), .ZN(n17507) );
  AOI22_X1 U19436 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17872), .B1(
        P3_EBX_REG_3__SCAN_IN), .B2(n17507), .ZN(n17502) );
  OAI22_X1 U19437 ( .A1(n17528), .A2(n17502), .B1(n17717), .B2(n17872), .ZN(
        P3_U2699) );
  INV_X1 U19438 ( .A(n17507), .ZN(n17504) );
  INV_X1 U19439 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17608) );
  NAND3_X1 U19440 ( .A1(n17504), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17872), .ZN(
        n17503) );
  OAI221_X1 U19441 ( .B1(n17504), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17872), 
        .C2(n17608), .A(n17503), .ZN(P3_U2700) );
  NOR2_X1 U19442 ( .A1(n17505), .A2(n17875), .ZN(n17506) );
  AOI21_X1 U19443 ( .B1(n17874), .B2(n17506), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17508) );
  AOI221_X1 U19444 ( .B1(n17508), .B2(n17872), .C1(n17706), .C2(n17878), .A(
        n17507), .ZN(P3_U2701) );
  OR2_X1 U19445 ( .A1(n17878), .A2(n17633), .ZN(n17523) );
  AOI22_X1 U19446 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17518) );
  AOI22_X1 U19447 ( .A1(n17861), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17517) );
  AOI22_X1 U19448 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17849), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17509) );
  OAI21_X1 U19449 ( .B1(n11093), .B2(n17684), .A(n17509), .ZN(n17515) );
  AOI22_X1 U19450 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U19451 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17512) );
  AOI22_X1 U19452 ( .A1(n17832), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17511) );
  AOI22_X1 U19453 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17833), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17510) );
  NAND4_X1 U19454 ( .A1(n17513), .A2(n17512), .A3(n17511), .A4(n17510), .ZN(
        n17514) );
  AOI211_X1 U19455 ( .C1(n17725), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n17515), .B(n17514), .ZN(n17516) );
  NAND3_X1 U19456 ( .A1(n17518), .A2(n17517), .A3(n17516), .ZN(n20769) );
  AOI22_X1 U19457 ( .A1(n17878), .A2(n20769), .B1(n17519), .B2(n17531), .ZN(
        n17520) );
  OAI21_X1 U19458 ( .B1(n17531), .B2(n17523), .A(n17520), .ZN(P3_U2695) );
  NOR2_X1 U19459 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17527), .ZN(n17521) );
  AOI22_X1 U19460 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17878), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n17521), .ZN(n17522) );
  OAI21_X1 U19461 ( .B1(n20251), .B2(n17523), .A(n17522), .ZN(P3_U2696) );
  INV_X1 U19462 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17526) );
  NAND2_X1 U19463 ( .A1(n17872), .A2(n17524), .ZN(n17529) );
  NAND2_X1 U19464 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17878), .ZN(
        n17525) );
  OAI221_X1 U19465 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17527), .C1(n17526), 
        .C2(n17529), .A(n17525), .ZN(P3_U2697) );
  NOR2_X1 U19466 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17528), .ZN(n17530) );
  INV_X1 U19467 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17746) );
  OAI22_X1 U19468 ( .A1(n17530), .A2(n17529), .B1(n17746), .B2(n17872), .ZN(
        P3_U2698) );
  NOR4_X1 U19469 ( .A1(n20305), .A2(n17532), .A3(n20274), .A4(n17531), .ZN(
        n17560) );
  INV_X1 U19470 ( .A(n17560), .ZN(n17535) );
  NAND4_X1 U19471 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .A4(P3_EBX_REG_12__SCAN_IN), .ZN(n17533)
         );
  NOR3_X1 U19472 ( .A1(n17535), .A2(n17534), .A3(n17533), .ZN(n17636) );
  NAND2_X1 U19473 ( .A1(n17636), .A2(n17536), .ZN(n17549) );
  INV_X1 U19474 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17548) );
  NAND2_X1 U19475 ( .A1(n17872), .A2(n17549), .ZN(n17562) );
  AOI22_X1 U19476 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17546) );
  AOI22_X1 U19477 ( .A1(n17848), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17545) );
  AOI22_X1 U19478 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17537) );
  OAI21_X1 U19479 ( .B1(n17747), .B2(n17684), .A(n17537), .ZN(n17543) );
  AOI22_X1 U19480 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17849), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17541) );
  AOI22_X1 U19481 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17540) );
  AOI22_X1 U19482 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17833), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U19483 ( .A1(n17832), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17538) );
  NAND4_X1 U19484 ( .A1(n17541), .A2(n17540), .A3(n17539), .A4(n17538), .ZN(
        n17542) );
  AOI211_X1 U19485 ( .C1(n17725), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n17543), .B(n17542), .ZN(n17544) );
  NAND3_X1 U19486 ( .A1(n17546), .A2(n17545), .A3(n17544), .ZN(n20746) );
  NAND2_X1 U19487 ( .A1(n17878), .A2(n20746), .ZN(n17547) );
  OAI221_X1 U19488 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17549), .C1(n17548), 
        .C2(n17562), .A(n17547), .ZN(P3_U2687) );
  AOI22_X1 U19489 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17559) );
  AOI22_X1 U19490 ( .A1(n11561), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17558) );
  AOI22_X1 U19491 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17550) );
  OAI21_X1 U19492 ( .B1(n11093), .B2(n17695), .A(n17550), .ZN(n17556) );
  AOI22_X1 U19493 ( .A1(n17718), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17554) );
  AOI22_X1 U19494 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17553) );
  AOI22_X1 U19495 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17552) );
  AOI22_X1 U19496 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17551) );
  NAND4_X1 U19497 ( .A1(n17554), .A2(n17553), .A3(n17552), .A4(n17551), .ZN(
        n17555) );
  AOI211_X1 U19498 ( .C1(n17851), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n17556), .B(n17555), .ZN(n17557) );
  NAND3_X1 U19499 ( .A1(n17559), .A2(n17558), .A3(n17557), .ZN(n20762) );
  INV_X1 U19500 ( .A(n20762), .ZN(n17564) );
  INV_X1 U19501 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20346) );
  INV_X1 U19502 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20335) );
  NOR2_X1 U19503 ( .A1(n20346), .A2(n20335), .ZN(n17561) );
  INV_X1 U19504 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17575) );
  NAND2_X1 U19505 ( .A1(n17560), .A2(n17633), .ZN(n17618) );
  NOR2_X1 U19506 ( .A1(n17575), .A2(n17618), .ZN(n17603) );
  AOI21_X1 U19507 ( .B1(n17561), .B2(n17603), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n17563) );
  OAI22_X1 U19508 ( .A1(n17564), .A2(n17872), .B1(n17563), .B2(n17562), .ZN(
        P3_U2688) );
  AOI22_X1 U19509 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17574) );
  AOI22_X1 U19510 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17573) );
  AOI22_X1 U19511 ( .A1(n17838), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17565) );
  OAI21_X1 U19512 ( .B1(n11093), .B2(n17746), .A(n17565), .ZN(n17571) );
  AOI22_X1 U19513 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17569) );
  AOI22_X1 U19514 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17568) );
  AOI22_X1 U19515 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17567) );
  AOI22_X1 U19516 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17566) );
  NAND4_X1 U19517 ( .A1(n17569), .A2(n17568), .A3(n17567), .A4(n17566), .ZN(
        n17570) );
  AOI211_X1 U19518 ( .C1(n17858), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n17571), .B(n17570), .ZN(n17572) );
  NAND3_X1 U19519 ( .A1(n17574), .A2(n17573), .A3(n17572), .ZN(n20601) );
  INV_X1 U19520 ( .A(n20601), .ZN(n17577) );
  NOR3_X1 U19521 ( .A1(n20622), .A2(n17575), .A3(n17618), .ZN(n17589) );
  OAI21_X1 U19522 ( .B1(n17878), .B2(n17603), .A(P3_EBX_REG_13__SCAN_IN), .ZN(
        n17578) );
  OAI21_X1 U19523 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17589), .A(n17578), .ZN(
        n17576) );
  OAI21_X1 U19524 ( .B1(n17577), .B2(n17872), .A(n17576), .ZN(P3_U2690) );
  NAND2_X1 U19525 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17578), .ZN(n17592) );
  AOI22_X1 U19526 ( .A1(n17861), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17588) );
  AOI22_X1 U19527 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17587) );
  AOI22_X1 U19528 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17579) );
  OAI21_X1 U19529 ( .B1(n11093), .B2(n17730), .A(n17579), .ZN(n17585) );
  AOI22_X1 U19530 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17583) );
  AOI22_X1 U19531 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17582) );
  AOI22_X1 U19532 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17581) );
  AOI22_X1 U19533 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17580) );
  NAND4_X1 U19534 ( .A1(n17583), .A2(n17582), .A3(n17581), .A4(n17580), .ZN(
        n17584) );
  AOI211_X1 U19535 ( .C1(n17851), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17585), .B(n17584), .ZN(n17586) );
  NAND3_X1 U19536 ( .A1(n17588), .A2(n17587), .A3(n17586), .ZN(n20756) );
  INV_X1 U19537 ( .A(n20756), .ZN(n17591) );
  NAND3_X1 U19538 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17589), .A3(n20346), 
        .ZN(n17590) );
  OAI221_X1 U19539 ( .B1(n17878), .B2(n17592), .C1(n17872), .C2(n17591), .A(
        n17590), .ZN(P3_U2689) );
  AOI22_X1 U19540 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17596) );
  AOI22_X1 U19541 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17595) );
  AOI22_X1 U19542 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17594) );
  AOI22_X1 U19543 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17593) );
  NAND4_X1 U19544 ( .A1(n17596), .A2(n17595), .A3(n17594), .A4(n17593), .ZN(
        n17602) );
  AOI22_X1 U19545 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17600) );
  AOI22_X1 U19546 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17599) );
  AOI22_X1 U19547 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17598) );
  AOI22_X1 U19548 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17597) );
  NAND4_X1 U19549 ( .A1(n17600), .A2(n17599), .A3(n17598), .A4(n17597), .ZN(
        n17601) );
  NOR2_X1 U19550 ( .A1(n17602), .A2(n17601), .ZN(n20606) );
  INV_X1 U19551 ( .A(n17618), .ZN(n17605) );
  NOR2_X1 U19552 ( .A1(n17878), .A2(n17603), .ZN(n17604) );
  OAI21_X1 U19553 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17605), .A(n17604), .ZN(
        n17606) );
  OAI21_X1 U19554 ( .B1(n20606), .B2(n17872), .A(n17606), .ZN(P3_U2691) );
  AOI22_X1 U19555 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17617) );
  AOI22_X1 U19556 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17616) );
  AOI22_X1 U19557 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17607) );
  OAI21_X1 U19558 ( .B1(n11093), .B2(n17608), .A(n17607), .ZN(n17614) );
  AOI22_X1 U19559 ( .A1(n17838), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17612) );
  AOI22_X1 U19560 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17611) );
  AOI22_X1 U19561 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17610) );
  AOI22_X1 U19562 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17609) );
  NAND4_X1 U19563 ( .A1(n17612), .A2(n17611), .A3(n17610), .A4(n17609), .ZN(
        n17613) );
  AOI211_X1 U19564 ( .C1(n17791), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17614), .B(n17613), .ZN(n17615) );
  NAND3_X1 U19565 ( .A1(n17617), .A2(n17616), .A3(n17615), .ZN(n20609) );
  INV_X1 U19566 ( .A(n20609), .ZN(n17621) );
  OAI21_X1 U19567 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17619), .A(n17618), .ZN(
        n17620) );
  AOI22_X1 U19568 ( .A1(n17878), .A2(n17621), .B1(n17620), .B2(n17872), .ZN(
        P3_U2692) );
  AOI22_X1 U19569 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17718), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17824), .ZN(n17625) );
  AOI22_X1 U19570 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17838), .ZN(n17624) );
  AOI22_X1 U19571 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17832), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17852), .ZN(n17623) );
  AOI22_X1 U19572 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17853), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n10977), .ZN(n17622) );
  NAND4_X1 U19573 ( .A1(n17625), .A2(n17624), .A3(n17623), .A4(n17622), .ZN(
        n17631) );
  AOI22_X1 U19574 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17858), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17629) );
  AOI22_X1 U19575 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17849), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17628) );
  AOI22_X1 U19576 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17627) );
  AOI22_X1 U19577 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17626) );
  NAND4_X1 U19578 ( .A1(n17629), .A2(n17628), .A3(n17627), .A4(n17626), .ZN(
        n17630) );
  NOR2_X1 U19579 ( .A1(n17631), .A2(n17630), .ZN(n20617) );
  OAI221_X1 U19580 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(P3_EBX_REG_8__SCAN_IN), 
        .C1(P3_EBX_REG_9__SCAN_IN), .C2(n17633), .A(n17632), .ZN(n17634) );
  AOI22_X1 U19581 ( .A1(n17878), .A2(n20617), .B1(n17634), .B2(n17872), .ZN(
        P3_U2694) );
  INV_X1 U19582 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n20579) );
  INV_X1 U19583 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n20435) );
  INV_X1 U19584 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n20400) );
  INV_X1 U19585 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20384) );
  NAND4_X1 U19586 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17636), .A4(n17635), .ZN(n17869) );
  NOR2_X1 U19587 ( .A1(n20384), .A2(n17869), .ZN(n17868) );
  NAND2_X1 U19588 ( .A1(n17874), .A2(n17868), .ZN(n17817) );
  NAND2_X1 U19589 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17846), .ZN(n17845) );
  NOR2_X1 U19590 ( .A1(n20435), .A2(n17845), .ZN(n17744) );
  INV_X1 U19591 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n20491) );
  INV_X1 U19592 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n20476) );
  INV_X1 U19593 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20448) );
  NAND4_X1 U19594 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_28__SCAN_IN), 
        .A3(P3_EBX_REG_27__SCAN_IN), .A4(P3_EBX_REG_26__SCAN_IN), .ZN(n17637)
         );
  NOR4_X1 U19595 ( .A1(n20491), .A2(n20476), .A3(n20448), .A4(n17637), .ZN(
        n17638) );
  NAND4_X1 U19596 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n17744), .A4(n17638), .ZN(n17641) );
  NOR2_X1 U19597 ( .A1(n20579), .A2(n17641), .ZN(n17743) );
  NAND2_X1 U19598 ( .A1(n17872), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17640) );
  NAND2_X1 U19599 ( .A1(n17743), .A2(n20768), .ZN(n17639) );
  OAI22_X1 U19600 ( .A1(n17743), .A2(n17640), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17639), .ZN(P3_U2672) );
  NAND2_X1 U19601 ( .A1(n20579), .A2(n17641), .ZN(n17642) );
  NAND2_X1 U19602 ( .A1(n17642), .A2(n17872), .ZN(n17742) );
  AOI22_X1 U19603 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17849), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17646) );
  AOI22_X1 U19604 ( .A1(n17861), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17645) );
  AOI22_X1 U19605 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17644) );
  AOI22_X1 U19606 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17643) );
  NAND4_X1 U19607 ( .A1(n17646), .A2(n17645), .A3(n17644), .A4(n17643), .ZN(
        n17652) );
  AOI22_X1 U19608 ( .A1(n17838), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17650) );
  AOI22_X1 U19609 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17649) );
  AOI22_X1 U19610 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17648) );
  AOI22_X1 U19611 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17647) );
  NAND4_X1 U19612 ( .A1(n17650), .A2(n17649), .A3(n17648), .A4(n17647), .ZN(
        n17651) );
  NOR2_X1 U19613 ( .A1(n17652), .A2(n17651), .ZN(n17741) );
  AOI22_X1 U19614 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17656) );
  AOI22_X1 U19615 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17655) );
  AOI22_X1 U19616 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17654) );
  AOI22_X1 U19617 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17653) );
  NAND4_X1 U19618 ( .A1(n17656), .A2(n17655), .A3(n17654), .A4(n17653), .ZN(
        n17662) );
  AOI22_X1 U19619 ( .A1(n17718), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17660) );
  AOI22_X1 U19620 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17659) );
  AOI22_X1 U19621 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17850), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17658) );
  AOI22_X1 U19622 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17657) );
  NAND4_X1 U19623 ( .A1(n17660), .A2(n17659), .A3(n17658), .A4(n17657), .ZN(
        n17661) );
  NOR2_X1 U19624 ( .A1(n17662), .A2(n17661), .ZN(n17767) );
  AOI22_X1 U19625 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17718), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17666) );
  AOI22_X1 U19626 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17665) );
  AOI22_X1 U19627 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17664) );
  AOI22_X1 U19628 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17663) );
  NAND4_X1 U19629 ( .A1(n17666), .A2(n17665), .A3(n17664), .A4(n17663), .ZN(
        n17672) );
  AOI22_X1 U19630 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17670) );
  AOI22_X1 U19631 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17669) );
  AOI22_X1 U19632 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17668) );
  AOI22_X1 U19633 ( .A1(n17861), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17667) );
  NAND4_X1 U19634 ( .A1(n17670), .A2(n17669), .A3(n17668), .A4(n17667), .ZN(
        n17671) );
  NOR2_X1 U19635 ( .A1(n17672), .A2(n17671), .ZN(n17772) );
  AOI22_X1 U19636 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17823), .ZN(n17676) );
  AOI22_X1 U19637 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17718), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17675) );
  AOI22_X1 U19638 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17852), .B1(
        n17833), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17674) );
  AOI22_X1 U19639 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17832), .ZN(n17673) );
  NAND4_X1 U19640 ( .A1(n17676), .A2(n17675), .A3(n17674), .A4(n17673), .ZN(
        n17682) );
  AOI22_X1 U19641 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17824), .ZN(n17680) );
  AOI22_X1 U19642 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17849), .ZN(n17679) );
  AOI22_X1 U19643 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17861), .ZN(n17678) );
  AOI22_X1 U19644 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17848), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17838), .ZN(n17677) );
  NAND4_X1 U19645 ( .A1(n17680), .A2(n17679), .A3(n17678), .A4(n17677), .ZN(
        n17681) );
  NOR2_X1 U19646 ( .A1(n17682), .A2(n17681), .ZN(n17781) );
  AOI22_X1 U19647 ( .A1(n17861), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17693) );
  AOI22_X1 U19648 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17692) );
  AOI22_X1 U19649 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17683) );
  OAI21_X1 U19650 ( .B1(n17731), .B2(n17684), .A(n17683), .ZN(n17690) );
  AOI22_X1 U19651 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17688) );
  AOI22_X1 U19652 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17687) );
  AOI22_X1 U19653 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17686) );
  AOI22_X1 U19654 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17685) );
  NAND4_X1 U19655 ( .A1(n17688), .A2(n17687), .A3(n17686), .A4(n17685), .ZN(
        n17689) );
  AOI211_X1 U19656 ( .C1(n17791), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n17690), .B(n17689), .ZN(n17691) );
  NAND3_X1 U19657 ( .A1(n17693), .A2(n17692), .A3(n17691), .ZN(n17786) );
  AOI22_X1 U19658 ( .A1(n17838), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17704) );
  AOI22_X1 U19659 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17703) );
  AOI22_X1 U19660 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17694) );
  OAI21_X1 U19661 ( .B1(n17747), .B2(n17695), .A(n17694), .ZN(n17701) );
  AOI22_X1 U19662 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17699) );
  AOI22_X1 U19663 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17849), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17698) );
  AOI22_X1 U19664 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17833), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17697) );
  AOI22_X1 U19665 ( .A1(n17832), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17696) );
  NAND4_X1 U19666 ( .A1(n17699), .A2(n17698), .A3(n17697), .A4(n17696), .ZN(
        n17700) );
  AOI211_X1 U19667 ( .C1(n17725), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n17701), .B(n17700), .ZN(n17702) );
  NAND3_X1 U19668 ( .A1(n17704), .A2(n17703), .A3(n17702), .ZN(n17787) );
  NAND2_X1 U19669 ( .A1(n17786), .A2(n17787), .ZN(n17785) );
  NOR2_X1 U19670 ( .A1(n17781), .A2(n17785), .ZN(n17780) );
  AOI22_X1 U19671 ( .A1(n17718), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17715) );
  AOI22_X1 U19672 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17714) );
  AOI22_X1 U19673 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17705) );
  OAI21_X1 U19674 ( .B1(n17731), .B2(n17706), .A(n17705), .ZN(n17712) );
  AOI22_X1 U19675 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17710) );
  AOI22_X1 U19676 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17709) );
  AOI22_X1 U19677 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17708) );
  AOI22_X1 U19678 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17707) );
  NAND4_X1 U19679 ( .A1(n17710), .A2(n17709), .A3(n17708), .A4(n17707), .ZN(
        n17711) );
  AOI211_X1 U19680 ( .C1(n17791), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n17712), .B(n17711), .ZN(n17713) );
  NAND3_X1 U19681 ( .A1(n17715), .A2(n17714), .A3(n17713), .ZN(n17777) );
  NAND2_X1 U19682 ( .A1(n17780), .A2(n17777), .ZN(n17776) );
  NOR2_X1 U19683 ( .A1(n17772), .A2(n17776), .ZN(n17771) );
  AOI22_X1 U19684 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17860), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17728) );
  AOI22_X1 U19685 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17727) );
  AOI22_X1 U19686 ( .A1(n10971), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17849), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17716) );
  OAI21_X1 U19687 ( .B1(n17731), .B2(n17717), .A(n17716), .ZN(n17724) );
  AOI22_X1 U19688 ( .A1(n17718), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17722) );
  AOI22_X1 U19689 ( .A1(n17861), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17721) );
  AOI22_X1 U19690 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17720) );
  AOI22_X1 U19691 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17719) );
  NAND4_X1 U19692 ( .A1(n17722), .A2(n17721), .A3(n17720), .A4(n17719), .ZN(
        n17723) );
  AOI211_X1 U19693 ( .C1(n17725), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n17724), .B(n17723), .ZN(n17726) );
  NAND3_X1 U19694 ( .A1(n17728), .A2(n17727), .A3(n17726), .ZN(n17758) );
  NAND2_X1 U19695 ( .A1(n17771), .A2(n17758), .ZN(n17766) );
  NOR2_X1 U19696 ( .A1(n17767), .A2(n17766), .ZN(n17765) );
  AOI22_X1 U19697 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17740) );
  AOI22_X1 U19698 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17739) );
  AOI22_X1 U19699 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17729) );
  OAI21_X1 U19700 ( .B1(n17731), .B2(n17730), .A(n17729), .ZN(n17737) );
  AOI22_X1 U19701 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17735) );
  AOI22_X1 U19702 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17838), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17734) );
  AOI22_X1 U19703 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17733) );
  AOI22_X1 U19704 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17732) );
  NAND4_X1 U19705 ( .A1(n17735), .A2(n17734), .A3(n17733), .A4(n17732), .ZN(
        n17736) );
  AOI211_X1 U19706 ( .C1(n17849), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n17737), .B(n17736), .ZN(n17738) );
  NAND3_X1 U19707 ( .A1(n17740), .A2(n17739), .A3(n17738), .ZN(n17762) );
  NAND2_X1 U19708 ( .A1(n17765), .A2(n17762), .ZN(n17761) );
  XNOR2_X1 U19709 ( .A(n17741), .B(n17761), .ZN(n20707) );
  OAI22_X1 U19710 ( .A1(n17743), .A2(n17742), .B1(n20707), .B2(n17872), .ZN(
        P3_U2673) );
  NOR2_X1 U19711 ( .A1(n20622), .A2(n17845), .ZN(n17815) );
  NAND2_X1 U19712 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17815), .ZN(n17759) );
  NOR2_X1 U19713 ( .A1(n17878), .A2(n17744), .ZN(n17814) );
  AOI22_X1 U19714 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17756) );
  AOI22_X1 U19715 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17838), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17755) );
  AOI22_X1 U19716 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17745) );
  OAI21_X1 U19717 ( .B1(n17747), .B2(n17746), .A(n17745), .ZN(n17753) );
  AOI22_X1 U19718 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U19719 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17750) );
  AOI22_X1 U19720 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U19721 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17748) );
  NAND4_X1 U19722 ( .A1(n17751), .A2(n17750), .A3(n17749), .A4(n17748), .ZN(
        n17752) );
  AOI211_X1 U19723 ( .C1(n17791), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n17753), .B(n17752), .ZN(n17754) );
  NAND3_X1 U19724 ( .A1(n17756), .A2(n17755), .A3(n17754), .ZN(n20654) );
  AOI22_X1 U19725 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17814), .B1(n17878), 
        .B2(n20654), .ZN(n17757) );
  OAI21_X1 U19726 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17759), .A(n17757), .ZN(
        P3_U2682) );
  OAI21_X1 U19727 ( .B1(n17771), .B2(n17758), .A(n17766), .ZN(n20727) );
  NAND2_X1 U19728 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17775), .ZN(n17770) );
  OAI211_X1 U19729 ( .C1(n17775), .C2(P3_EBX_REG_27__SCAN_IN), .A(n17872), .B(
        n17770), .ZN(n17760) );
  OAI21_X1 U19730 ( .B1(n17872), .B2(n20727), .A(n17760), .ZN(P3_U2676) );
  NAND3_X1 U19731 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n17775), .ZN(n17764) );
  OAI21_X1 U19732 ( .B1(n17765), .B2(n17762), .A(n17761), .ZN(n20715) );
  NAND3_X1 U19733 ( .A1(n17764), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17872), 
        .ZN(n17763) );
  OAI221_X1 U19734 ( .B1(n17764), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17872), 
        .C2(n20715), .A(n17763), .ZN(P3_U2674) );
  AND2_X1 U19735 ( .A1(n17872), .A2(n17764), .ZN(n17768) );
  AOI21_X1 U19736 ( .B1(n17767), .B2(n17766), .A(n17765), .ZN(n20720) );
  AOI22_X1 U19737 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17768), .B1(n20720), 
        .B2(n17878), .ZN(n17769) );
  OAI21_X1 U19738 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17770), .A(n17769), .ZN(
        P3_U2675) );
  AOI21_X1 U19739 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17872), .A(n17779), .ZN(
        n17774) );
  AOI21_X1 U19740 ( .B1(n17772), .B2(n17776), .A(n17771), .ZN(n20696) );
  INV_X1 U19741 ( .A(n20696), .ZN(n17773) );
  OAI22_X1 U19742 ( .A1(n17775), .A2(n17774), .B1(n17773), .B2(n17872), .ZN(
        P3_U2677) );
  INV_X1 U19743 ( .A(n17784), .ZN(n17789) );
  AOI22_X1 U19744 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17872), .B1(
        P3_EBX_REG_24__SCAN_IN), .B2(n17789), .ZN(n17778) );
  OAI21_X1 U19745 ( .B1(n17780), .B2(n17777), .A(n17776), .ZN(n20695) );
  OAI22_X1 U19746 ( .A1(n17779), .A2(n17778), .B1(n20695), .B2(n17872), .ZN(
        P3_U2678) );
  AOI21_X1 U19747 ( .B1(n17781), .B2(n17785), .A(n17780), .ZN(n20732) );
  INV_X1 U19748 ( .A(n20732), .ZN(n17783) );
  NAND3_X1 U19749 ( .A1(n17784), .A2(P3_EBX_REG_24__SCAN_IN), .A3(n17872), 
        .ZN(n17782) );
  OAI221_X1 U19750 ( .B1(n17784), .B2(P3_EBX_REG_24__SCAN_IN), .C1(n17872), 
        .C2(n17783), .A(n17782), .ZN(P3_U2679) );
  AOI21_X1 U19751 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17872), .A(n17803), .ZN(
        n17788) );
  OAI21_X1 U19752 ( .B1(n17787), .B2(n17786), .A(n17785), .ZN(n20738) );
  OAI22_X1 U19753 ( .A1(n17789), .A2(n17788), .B1(n17872), .B2(n20738), .ZN(
        P3_U2680) );
  AOI21_X1 U19754 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17872), .A(n17790), .ZN(
        n17802) );
  AOI22_X1 U19755 ( .A1(n17791), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17795) );
  AOI22_X1 U19756 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17794) );
  AOI22_X1 U19757 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17793) );
  AOI22_X1 U19758 ( .A1(n11437), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17792) );
  NAND4_X1 U19759 ( .A1(n17795), .A2(n17794), .A3(n17793), .A4(n17792), .ZN(
        n17801) );
  AOI22_X1 U19760 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17799) );
  AOI22_X1 U19761 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17798) );
  AOI22_X1 U19762 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17797) );
  AOI22_X1 U19763 ( .A1(n17838), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17796) );
  NAND4_X1 U19764 ( .A1(n17799), .A2(n17798), .A3(n17797), .A4(n17796), .ZN(
        n17800) );
  NOR2_X1 U19765 ( .A1(n17801), .A2(n17800), .ZN(n20666) );
  OAI22_X1 U19766 ( .A1(n17803), .A2(n17802), .B1(n20666), .B2(n17872), .ZN(
        P3_U2681) );
  AOI22_X1 U19767 ( .A1(n17848), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17807) );
  AOI22_X1 U19768 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17806) );
  AOI22_X1 U19769 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17805) );
  AOI22_X1 U19770 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17804) );
  NAND4_X1 U19771 ( .A1(n17807), .A2(n17806), .A3(n17805), .A4(n17804), .ZN(
        n17813) );
  AOI22_X1 U19772 ( .A1(n10972), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17838), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17811) );
  AOI22_X1 U19773 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17810) );
  AOI22_X1 U19774 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17849), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17809) );
  AOI22_X1 U19775 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17808) );
  NAND4_X1 U19776 ( .A1(n17811), .A2(n17810), .A3(n17809), .A4(n17808), .ZN(
        n17812) );
  NOR2_X1 U19777 ( .A1(n17813), .A2(n17812), .ZN(n20664) );
  OAI21_X1 U19778 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17815), .A(n17814), .ZN(
        n17816) );
  OAI21_X1 U19779 ( .B1(n20664), .B2(n17872), .A(n17816), .ZN(P3_U2683) );
  AOI21_X1 U19780 ( .B1(n20400), .B2(n17817), .A(n17878), .ZN(n17818) );
  INV_X1 U19781 ( .A(n17818), .ZN(n17831) );
  AOI22_X1 U19782 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17838), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17822) );
  AOI22_X1 U19783 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17821) );
  AOI22_X1 U19784 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17820) );
  AOI22_X1 U19785 ( .A1(n17833), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17819) );
  NAND4_X1 U19786 ( .A1(n17822), .A2(n17821), .A3(n17820), .A4(n17819), .ZN(
        n17830) );
  AOI22_X1 U19787 ( .A1(n17823), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17828) );
  AOI22_X1 U19788 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17827) );
  AOI22_X1 U19789 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17826) );
  AOI22_X1 U19790 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10972), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17825) );
  NAND4_X1 U19791 ( .A1(n17828), .A2(n17827), .A3(n17826), .A4(n17825), .ZN(
        n17829) );
  NOR2_X1 U19792 ( .A1(n17830), .A2(n17829), .ZN(n20685) );
  OAI22_X1 U19793 ( .A1(n17846), .A2(n17831), .B1(n20685), .B2(n17872), .ZN(
        P3_U2685) );
  AOI22_X1 U19794 ( .A1(n17850), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17837) );
  AOI22_X1 U19795 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17836) );
  AOI22_X1 U19796 ( .A1(n10977), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17832), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17835) );
  AOI22_X1 U19797 ( .A1(n17853), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17852), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17834) );
  NAND4_X1 U19798 ( .A1(n17837), .A2(n17836), .A3(n17835), .A4(n17834), .ZN(
        n17844) );
  AOI22_X1 U19799 ( .A1(n17838), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17842) );
  AOI22_X1 U19800 ( .A1(n17849), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17841) );
  AOI22_X1 U19801 ( .A1(n17858), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17823), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17840) );
  AOI22_X1 U19802 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10971), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17839) );
  NAND4_X1 U19803 ( .A1(n17842), .A2(n17841), .A3(n17840), .A4(n17839), .ZN(
        n17843) );
  NOR2_X1 U19804 ( .A1(n17844), .A2(n17843), .ZN(n20680) );
  OAI21_X1 U19805 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17846), .A(n17845), .ZN(
        n17847) );
  AOI22_X1 U19806 ( .A1(n17878), .A2(n20680), .B1(n17847), .B2(n17872), .ZN(
        P3_U2684) );
  AOI22_X1 U19807 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17849), .B1(
        n17848), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17857) );
  AOI22_X1 U19808 ( .A1(n17851), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17850), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17856) );
  AOI22_X1 U19809 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17852), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17832), .ZN(n17855) );
  AOI22_X1 U19810 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17833), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17853), .ZN(n17854) );
  NAND4_X1 U19811 ( .A1(n17857), .A2(n17856), .A3(n17855), .A4(n17854), .ZN(
        n17867) );
  AOI22_X1 U19812 ( .A1(n17725), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17858), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17865) );
  AOI22_X1 U19813 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17823), .B1(
        n17859), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17864) );
  AOI22_X1 U19814 ( .A1(n17860), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17863) );
  AOI22_X1 U19815 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10972), .B1(
        n17861), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17862) );
  NAND4_X1 U19816 ( .A1(n17865), .A2(n17864), .A3(n17863), .A4(n17862), .ZN(
        n17866) );
  NOR2_X1 U19817 ( .A1(n17867), .A2(n17866), .ZN(n20689) );
  AOI211_X1 U19818 ( .C1(n20384), .C2(n17869), .A(n17868), .B(n17880), .ZN(
        n17870) );
  AOI21_X1 U19819 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17877), .A(n17870), .ZN(
        n17871) );
  OAI21_X1 U19820 ( .B1(n20689), .B2(n17872), .A(n17871), .ZN(P3_U2686) );
  OAI222_X1 U19821 ( .A1(n17880), .A2(n17876), .B1(n17875), .B2(n17874), .C1(
        n17873), .C2(n17872), .ZN(P3_U2702) );
  AOI22_X1 U19822 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17878), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17877), .ZN(n17879) );
  OAI21_X1 U19823 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17880), .A(n17879), .ZN(
        P3_U2703) );
  INV_X1 U19824 ( .A(n17881), .ZN(n21227) );
  OAI21_X1 U19825 ( .B1(n21227), .B2(n20113), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17882) );
  OAI21_X1 U19826 ( .B1(n17884), .B2(n17883), .A(n17882), .ZN(P3_U2634) );
  INV_X1 U19827 ( .A(n17885), .ZN(n17886) );
  AOI21_X1 U19828 ( .B1(n21260), .B2(n17887), .A(n17886), .ZN(n21251) );
  INV_X1 U19829 ( .A(n18769), .ZN(n18750) );
  OAI21_X1 U19830 ( .B1(n21251), .B2(n18750), .A(n18290), .ZN(n17888) );
  OAI221_X1 U19831 ( .B1(n18802), .B2(n17890), .C1(n18802), .C2(n18290), .A(
        n17888), .ZN(P3_U2863) );
  NOR2_X2 U19832 ( .A1(n21259), .A2(n20106), .ZN(n18279) );
  NAND2_X1 U19833 ( .A1(n20625), .A2(n18279), .ZN(n18195) );
  INV_X1 U19834 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n20985) );
  NOR3_X1 U19835 ( .A1(n10978), .A2(n20985), .A3(n20982), .ZN(n18124) );
  INV_X1 U19836 ( .A(n17889), .ZN(n21136) );
  INV_X1 U19837 ( .A(n20984), .ZN(n20973) );
  OAI22_X1 U19838 ( .A1(n21136), .A2(n18285), .B1(n20973), .B2(n18195), .ZN(
        n17927) );
  AOI21_X1 U19839 ( .B1(n18124), .B2(n21135), .A(n17927), .ZN(n18127) );
  NOR2_X1 U19840 ( .A1(n17891), .A2(n20169), .ZN(n18114) );
  AOI21_X1 U19841 ( .B1(n18182), .B2(n17891), .A(n18251), .ZN(n18119) );
  OAI21_X1 U19842 ( .B1(n18114), .B2(n18281), .A(n18119), .ZN(n17905) );
  INV_X1 U19843 ( .A(n18074), .ZN(n18035) );
  NOR3_X1 U19844 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18035), .A3(
        n17891), .ZN(n17906) );
  INV_X1 U19845 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21152) );
  NAND2_X1 U19846 ( .A1(n17907), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20413) );
  OAI21_X1 U19847 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18114), .A(
        n20413), .ZN(n20398) );
  OAI22_X1 U19848 ( .A1(n11764), .A2(n21152), .B1(n18116), .B2(n20398), .ZN(
        n17892) );
  AOI211_X1 U19849 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17905), .A(
        n17906), .B(n17892), .ZN(n17896) );
  AOI21_X1 U19850 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18189), .A(
        n17987), .ZN(n17894) );
  XNOR2_X1 U19851 ( .A(n17894), .B(n17899), .ZN(n21150) );
  NOR2_X1 U19852 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21135), .ZN(
        n21149) );
  AOI22_X1 U19853 ( .A1(n18197), .A2(n21150), .B1(n21149), .B2(n18124), .ZN(
        n17895) );
  OAI211_X1 U19854 ( .C1(n18127), .C2(n17902), .A(n17896), .B(n17895), .ZN(
        P3_U2812) );
  INV_X1 U19855 ( .A(n10978), .ZN(n18161) );
  NAND2_X1 U19856 ( .A1(n18161), .A2(n17897), .ZN(n18089) );
  INV_X1 U19857 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21123) );
  NOR2_X1 U19858 ( .A1(n17898), .A2(n21123), .ZN(n20834) );
  NAND2_X1 U19859 ( .A1(n21136), .A2(n20834), .ZN(n21112) );
  NAND2_X1 U19860 ( .A1(n20973), .A2(n20834), .ZN(n21113) );
  AOI22_X1 U19861 ( .A1(n18225), .A2(n21112), .B1(n18141), .B2(n21113), .ZN(
        n17993) );
  NOR2_X1 U19862 ( .A1(n17900), .A2(n17899), .ZN(n17971) );
  NOR3_X1 U19863 ( .A1(n18190), .A2(n17902), .A3(n17901), .ZN(n17986) );
  NOR2_X1 U19864 ( .A1(n17971), .A2(n17986), .ZN(n17903) );
  XOR2_X1 U19865 ( .A(n17903), .B(n21123), .Z(n21120) );
  INV_X1 U19866 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n20408) );
  NOR2_X1 U19867 ( .A1(n11764), .A2(n20408), .ZN(n21119) );
  INV_X1 U19868 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n20409) );
  AOI21_X1 U19869 ( .B1(n20409), .B2(n20413), .A(n17978), .ZN(n17904) );
  INV_X1 U19870 ( .A(n17904), .ZN(n20416) );
  OAI21_X1 U19871 ( .B1(n17906), .B2(n17905), .A(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17909) );
  NAND3_X1 U19872 ( .A1(n17907), .A2(n20409), .A3(n18074), .ZN(n17908) );
  OAI211_X1 U19873 ( .C1(n20416), .C2(n18116), .A(n17909), .B(n17908), .ZN(
        n17910) );
  AOI211_X1 U19874 ( .C1(n18197), .C2(n21120), .A(n21119), .B(n17910), .ZN(
        n17911) );
  OAI221_X1 U19875 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18089), 
        .C1(n21123), .C2(n17993), .A(n17911), .ZN(P3_U2811) );
  NAND3_X1 U19876 ( .A1(n17930), .A2(n20348), .A3(n18074), .ZN(n17925) );
  NOR2_X1 U19877 ( .A1(n17912), .A2(n20169), .ZN(n18132) );
  AOI21_X1 U19878 ( .B1(n18182), .B2(n17912), .A(n18251), .ZN(n18134) );
  OAI21_X1 U19879 ( .B1(n18132), .B2(n18281), .A(n18134), .ZN(n17922) );
  INV_X1 U19880 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20371) );
  NOR2_X1 U19881 ( .A1(n11764), .A2(n20371), .ZN(n20987) );
  NAND2_X1 U19882 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18132), .ZN(
        n20347) );
  OAI21_X1 U19883 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18132), .A(
        n20347), .ZN(n20353) );
  NOR2_X1 U19884 ( .A1(n18116), .A2(n20353), .ZN(n17913) );
  AOI211_X1 U19885 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17922), .A(
        n20987), .B(n17913), .ZN(n17918) );
  NOR3_X1 U19886 ( .A1(n11539), .A2(n18190), .A3(n20928), .ZN(n18158) );
  NAND2_X1 U19887 ( .A1(n20958), .A2(n18158), .ZN(n18128) );
  NAND2_X1 U19888 ( .A1(n17935), .A2(n17914), .ZN(n18129) );
  AOI22_X1 U19889 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18128), .B1(
        n18129), .B2(n18140), .ZN(n17915) );
  XOR2_X1 U19890 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17915), .Z(
        n20988) );
  OAI21_X1 U19891 ( .B1(n10978), .B2(n20982), .A(n20985), .ZN(n17916) );
  AOI22_X1 U19892 ( .A1(n18197), .A2(n20988), .B1(n17927), .B2(n17916), .ZN(
        n17917) );
  OAI211_X1 U19893 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17925), .A(
        n17918), .B(n17917), .ZN(P3_U2815) );
  AOI22_X1 U19894 ( .A1(n18189), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n11551), .B2(n18190), .ZN(n17919) );
  XNOR2_X1 U19895 ( .A(n17920), .B(n17919), .ZN(n21167) );
  OAI21_X1 U19896 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n20378), .ZN(n17924) );
  INV_X1 U19897 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17921) );
  AOI22_X1 U19898 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18118), .B1(
        n17921), .B2(n20347), .ZN(n20362) );
  AOI22_X1 U19899 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17922), .B1(
        n18110), .B2(n20362), .ZN(n17923) );
  NAND2_X1 U19900 ( .A1(n10979), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n21165) );
  OAI211_X1 U19901 ( .C1(n17925), .C2(n17924), .A(n17923), .B(n21165), .ZN(
        n17926) );
  AOI221_X1 U19902 ( .B1(n18124), .B2(n11551), .C1(n17927), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n17926), .ZN(n17928) );
  OAI21_X1 U19903 ( .B1(n18144), .B2(n21167), .A(n17928), .ZN(P3_U2814) );
  NAND3_X1 U19904 ( .A1(n20934), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n20952), .ZN(n20957) );
  NAND2_X1 U19905 ( .A1(n17930), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17931) );
  AOI21_X1 U19906 ( .B1(n18076), .B2(n17931), .A(n18251), .ZN(n17929) );
  OAI21_X1 U19907 ( .B1(n17930), .B2(n18240), .A(n17929), .ZN(n17947) );
  INV_X1 U19908 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20321) );
  NOR2_X1 U19909 ( .A1(n11764), .A2(n20321), .ZN(n17933) );
  NAND2_X1 U19910 ( .A1(n17930), .A2(n18074), .ZN(n17944) );
  INV_X1 U19911 ( .A(n17931), .ZN(n18146) );
  NAND2_X1 U19912 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18146), .ZN(
        n17942) );
  OAI21_X1 U19913 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18146), .A(
        n17942), .ZN(n20311) );
  OAI22_X1 U19914 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17944), .B1(
        n20311), .B2(n18116), .ZN(n17932) );
  AOI211_X1 U19915 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17947), .A(
        n17933), .B(n17932), .ZN(n17940) );
  NOR2_X1 U19916 ( .A1(n20936), .A2(n17941), .ZN(n20948) );
  NAND2_X1 U19917 ( .A1(n21138), .A2(n20959), .ZN(n20951) );
  INV_X1 U19918 ( .A(n20951), .ZN(n17934) );
  OAI22_X1 U19919 ( .A1(n20948), .A2(n18285), .B1(n17934), .B2(n18195), .ZN(
        n17951) );
  INV_X1 U19920 ( .A(n20934), .ZN(n20938) );
  INV_X1 U19921 ( .A(n18158), .ZN(n18169) );
  NOR2_X1 U19922 ( .A1(n20938), .A2(n18169), .ZN(n17937) );
  NAND2_X1 U19923 ( .A1(n17935), .A2(n11543), .ZN(n18170) );
  INV_X1 U19924 ( .A(n18170), .ZN(n18157) );
  AOI22_X1 U19925 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17937), .B1(
        n17936), .B2(n18157), .ZN(n17938) );
  XOR2_X1 U19926 ( .A(n20952), .B(n17938), .Z(n20954) );
  AOI22_X1 U19927 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17951), .B1(
        n18197), .B2(n20954), .ZN(n17939) );
  OAI211_X1 U19928 ( .C1(n10978), .C2(n20957), .A(n17940), .B(n17939), .ZN(
        P3_U2818) );
  OR2_X1 U19929 ( .A1(n17941), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n21176) );
  INV_X1 U19930 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20331) );
  NOR2_X1 U19931 ( .A1(n11764), .A2(n20331), .ZN(n17946) );
  INV_X1 U19932 ( .A(n17942), .ZN(n18131) );
  XNOR2_X1 U19933 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n18131), .ZN(
        n20323) );
  OAI21_X1 U19934 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n20322), .ZN(n17943) );
  OAI22_X1 U19935 ( .A1(n18116), .A2(n20323), .B1(n17944), .B2(n17943), .ZN(
        n17945) );
  AOI211_X1 U19936 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17947), .A(
        n17946), .B(n17945), .ZN(n17953) );
  NAND3_X1 U19937 ( .A1(n18189), .A2(n11074), .A3(n20959), .ZN(n17948) );
  OAI21_X1 U19938 ( .B1(n18189), .B2(n17949), .A(n17948), .ZN(n17950) );
  XOR2_X1 U19939 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17950), .Z(
        n21169) );
  AOI22_X1 U19940 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17951), .B1(
        n18197), .B2(n21169), .ZN(n17952) );
  OAI211_X1 U19941 ( .C1(n10978), .C2(n21176), .A(n17953), .B(n17952), .ZN(
        P3_U2817) );
  INV_X1 U19942 ( .A(n17985), .ZN(n17954) );
  AOI21_X1 U19943 ( .B1(n17956), .B2(n17955), .A(n17954), .ZN(n18006) );
  XOR2_X1 U19944 ( .A(n21087), .B(n18006), .Z(n21005) );
  INV_X1 U19945 ( .A(n20430), .ZN(n17979) );
  NAND2_X1 U19946 ( .A1(n17979), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17996) );
  OAI21_X1 U19947 ( .B1(n17978), .B2(n18281), .A(n18280), .ZN(n17957) );
  AOI21_X1 U19948 ( .B1(n18182), .B2(n17996), .A(n17957), .ZN(n17981) );
  OAI21_X1 U19949 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18117), .A(
        n17981), .ZN(n17969) );
  INV_X1 U19950 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20442) );
  NOR2_X1 U19951 ( .A1(n20442), .A2(n17977), .ZN(n17958) );
  INV_X1 U19952 ( .A(n17995), .ZN(n17999) );
  OAI21_X1 U19953 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17958), .A(
        n17999), .ZN(n20456) );
  NOR2_X1 U19954 ( .A1(n18035), .A2(n17996), .ZN(n17970) );
  OAI211_X1 U19955 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17970), .B(n17997), .ZN(n17959) );
  NAND2_X1 U19956 ( .A1(n10979), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n21003) );
  OAI211_X1 U19957 ( .C1(n18116), .C2(n20456), .A(n17959), .B(n21003), .ZN(
        n17965) );
  INV_X1 U19958 ( .A(n17960), .ZN(n21088) );
  NOR2_X1 U19959 ( .A1(n21088), .A2(n18089), .ZN(n17963) );
  INV_X1 U19960 ( .A(n17961), .ZN(n21091) );
  INV_X1 U19961 ( .A(n20839), .ZN(n21092) );
  AOI22_X1 U19962 ( .A1(n18225), .A2(n21091), .B1(n18141), .B2(n21092), .ZN(
        n17976) );
  INV_X1 U19963 ( .A(n17976), .ZN(n17962) );
  MUX2_X1 U19964 ( .A(n17963), .B(n17962), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17964) );
  AOI211_X1 U19965 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n17969), .A(
        n17965), .B(n17964), .ZN(n17966) );
  OAI21_X1 U19966 ( .B1(n18144), .B2(n21005), .A(n17966), .ZN(P3_U2808) );
  INV_X1 U19967 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20846) );
  INV_X1 U19968 ( .A(n17977), .ZN(n17967) );
  AOI22_X1 U19969 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17977), .B1(
        n17967), .B2(n20442), .ZN(n20438) );
  OAI22_X1 U19970 ( .A1(n11764), .A2(n20846), .B1(n18116), .B2(n20438), .ZN(
        n17968) );
  AOI221_X1 U19971 ( .B1(n17970), .B2(n20442), .C1(n17969), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17968), .ZN(n17975) );
  INV_X1 U19972 ( .A(n20837), .ZN(n20841) );
  AOI22_X1 U19973 ( .A1(n20841), .A2(n17986), .B1(n17972), .B2(n17971), .ZN(
        n17973) );
  XOR2_X1 U19974 ( .A(n20999), .B(n17973), .Z(n20844) );
  INV_X1 U19975 ( .A(n18089), .ZN(n18043) );
  NOR2_X1 U19976 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n20837), .ZN(
        n20843) );
  AOI22_X1 U19977 ( .A1(n18197), .A2(n20844), .B1(n18043), .B2(n20843), .ZN(
        n17974) );
  OAI211_X1 U19978 ( .C1(n17976), .C2(n20999), .A(n17975), .B(n17974), .ZN(
        P3_U2809) );
  INV_X1 U19979 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17992) );
  OAI21_X1 U19980 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17978), .A(
        n17977), .ZN(n20432) );
  INV_X1 U19981 ( .A(n20432), .ZN(n17984) );
  INV_X1 U19982 ( .A(n18117), .ZN(n17983) );
  AOI21_X1 U19983 ( .B1(n17979), .B2(n19082), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17980) );
  NAND2_X1 U19984 ( .A1(n10979), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n21130) );
  OAI21_X1 U19985 ( .B1(n17981), .B2(n17980), .A(n21130), .ZN(n17982) );
  AOI221_X1 U19986 ( .B1(n18110), .B2(n17984), .C1(n17983), .C2(n17984), .A(
        n17982), .ZN(n17991) );
  OAI221_X1 U19987 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17987), 
        .C1(n21123), .C2(n17986), .A(n17985), .ZN(n17988) );
  XOR2_X1 U19988 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17988), .Z(
        n21132) );
  INV_X1 U19989 ( .A(n21132), .ZN(n17989) );
  NOR2_X1 U19990 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21123), .ZN(
        n21127) );
  AOI22_X1 U19991 ( .A1(n18197), .A2(n17989), .B1(n18043), .B2(n21127), .ZN(
        n17990) );
  OAI211_X1 U19992 ( .C1(n17993), .C2(n17992), .A(n17991), .B(n17990), .ZN(
        P3_U2810) );
  OAI21_X1 U19993 ( .B1(n21093), .B2(n21092), .A(n18141), .ZN(n18005) );
  OAI21_X1 U19994 ( .B1(n21093), .B2(n21091), .A(n18225), .ZN(n18004) );
  OAI22_X1 U19995 ( .A1(n21092), .A2(n18005), .B1(n21091), .B2(n18004), .ZN(
        n17994) );
  INV_X1 U19996 ( .A(n17994), .ZN(n18011) );
  OAI21_X1 U19997 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17995), .A(
        n18026), .ZN(n20466) );
  INV_X1 U19998 ( .A(n20466), .ZN(n18003) );
  NOR2_X1 U19999 ( .A1(n17997), .A2(n17996), .ZN(n18000) );
  NAND2_X1 U20000 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18000), .ZN(
        n18033) );
  AND2_X1 U20001 ( .A1(n18033), .A2(n19082), .ZN(n17998) );
  AOI211_X1 U20002 ( .C1(n18076), .C2(n17999), .A(n18251), .B(n17998), .ZN(
        n18013) );
  AOI21_X1 U20003 ( .B1(n18000), .B2(n19082), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18001) );
  INV_X1 U20004 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20474) );
  OAI22_X1 U20005 ( .A1(n18013), .A2(n18001), .B1(n11764), .B2(n20474), .ZN(
        n18002) );
  AOI221_X1 U20006 ( .B1(n18110), .B2(n18003), .C1(n17983), .C2(n18003), .A(
        n18002), .ZN(n18010) );
  NAND2_X1 U20007 ( .A1(n18005), .A2(n18004), .ZN(n18030) );
  OAI221_X1 U20008 ( .B1(n18007), .B2(n18189), .C1(n18007), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18006), .ZN(n18008) );
  XNOR2_X1 U20009 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n18008), .ZN(
        n21101) );
  AOI22_X1 U20010 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18030), .B1(
        n18197), .B2(n21101), .ZN(n18009) );
  OAI211_X1 U20011 ( .C1(n18011), .C2(n21087), .A(n18010), .B(n18009), .ZN(
        P3_U2807) );
  XOR2_X1 U20012 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18012), .Z(
        n21014) );
  OAI21_X1 U20013 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18117), .A(
        n18013), .ZN(n18028) );
  INV_X1 U20014 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20477) );
  NOR2_X1 U20015 ( .A1(n20477), .A2(n18026), .ZN(n18015) );
  INV_X1 U20016 ( .A(n18063), .ZN(n18014) );
  OAI21_X1 U20017 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18015), .A(
        n18014), .ZN(n20496) );
  NOR2_X1 U20018 ( .A1(n18035), .A2(n18033), .ZN(n18029) );
  OAI211_X1 U20019 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18029), .B(n18034), .ZN(n18016) );
  NAND2_X1 U20020 ( .A1(n10979), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21019) );
  OAI211_X1 U20021 ( .C1(n18116), .C2(n20496), .A(n18016), .B(n21019), .ZN(
        n18021) );
  XOR2_X1 U20022 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18017), .Z(
        n21013) );
  OAI21_X1 U20023 ( .B1(n18190), .B2(n18018), .A(n11019), .ZN(n18019) );
  XOR2_X1 U20024 ( .A(n18019), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n21016) );
  OAI22_X1 U20025 ( .A1(n18195), .A2(n21013), .B1(n18144), .B2(n21016), .ZN(
        n18020) );
  AOI211_X1 U20026 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18028), .A(
        n18021), .B(n18020), .ZN(n18022) );
  OAI21_X1 U20027 ( .B1(n18285), .B2(n21014), .A(n18022), .ZN(P3_U2805) );
  AOI21_X1 U20028 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18024), .A(
        n18023), .ZN(n21111) );
  INV_X1 U20029 ( .A(n18026), .ZN(n18025) );
  AOI22_X1 U20030 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18026), .B1(
        n18025), .B2(n20477), .ZN(n20482) );
  NAND2_X1 U20031 ( .A1(n10979), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n21109) );
  OAI21_X1 U20032 ( .B1(n18116), .B2(n20482), .A(n21109), .ZN(n18027) );
  AOI221_X1 U20033 ( .B1(n18029), .B2(n20477), .C1(n18028), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18027), .ZN(n18032) );
  NOR3_X1 U20034 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21088), .A3(
        n21093), .ZN(n21108) );
  AOI22_X1 U20035 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18030), .B1(
        n18043), .B2(n21108), .ZN(n18031) );
  OAI211_X1 U20036 ( .C1(n21111), .C2(n18144), .A(n18032), .B(n18031), .ZN(
        P3_U2806) );
  NOR2_X1 U20037 ( .A1(n18034), .A2(n18033), .ZN(n18061) );
  NAND2_X1 U20038 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18061), .ZN(
        n18038) );
  NOR3_X1 U20039 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18035), .A3(
        n18038), .ZN(n18051) );
  OAI21_X1 U20040 ( .B1(n18063), .B2(n18281), .A(n18280), .ZN(n18036) );
  AOI21_X1 U20041 ( .B1(n18182), .B2(n18038), .A(n18036), .ZN(n18066) );
  OAI21_X1 U20042 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18117), .A(
        n18066), .ZN(n18054) );
  OAI21_X1 U20043 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11061), .A(
        n18109), .ZN(n20544) );
  INV_X1 U20044 ( .A(n18037), .ZN(n18040) );
  NOR2_X1 U20045 ( .A1(n20517), .A2(n18038), .ZN(n18073) );
  NAND3_X1 U20046 ( .A1(n18073), .A2(n11288), .A3(n18074), .ZN(n18039) );
  OAI211_X1 U20047 ( .C1(n18116), .C2(n20544), .A(n18040), .B(n18039), .ZN(
        n18041) );
  AOI221_X1 U20048 ( .B1(n18051), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(
        n18054), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n18041), .ZN(
        n18050) );
  INV_X1 U20049 ( .A(n21022), .ZN(n21037) );
  AOI22_X1 U20050 ( .A1(n18225), .A2(n21040), .B1(n18141), .B2(n21037), .ZN(
        n18071) );
  NAND2_X1 U20051 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18071), .ZN(
        n18055) );
  OAI211_X1 U20052 ( .C1(n18225), .C2(n18141), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18055), .ZN(n18049) );
  NAND3_X1 U20053 ( .A1(n21054), .A2(n18043), .A3(n18042), .ZN(n18048) );
  OAI211_X1 U20054 ( .C1(n18046), .C2(n18045), .A(n18197), .B(n18044), .ZN(
        n18047) );
  NAND4_X1 U20055 ( .A1(n18050), .A2(n18049), .A3(n18048), .A4(n18047), .ZN(
        P3_U2802) );
  AOI21_X1 U20056 ( .B1(n20517), .B2(n18062), .A(n11061), .ZN(n20521) );
  AOI21_X1 U20057 ( .B1(n18110), .B2(n20521), .A(n18051), .ZN(n18059) );
  OAI21_X1 U20058 ( .B1(n18189), .B2(n18053), .A(n18052), .ZN(n21042) );
  AOI22_X1 U20059 ( .A1(n18197), .A2(n21042), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18054), .ZN(n18058) );
  NOR2_X1 U20060 ( .A1(n18090), .A2(n18089), .ZN(n18056) );
  OAI21_X1 U20061 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18056), .A(
        n18055), .ZN(n18057) );
  NAND2_X1 U20062 ( .A1(n10979), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21043) );
  NAND4_X1 U20063 ( .A1(n18059), .A2(n18058), .A3(n18057), .A4(n21043), .ZN(
        P3_U2803) );
  OAI221_X1 U20064 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18190), 
        .C1(n21025), .C2(n18018), .A(n11019), .ZN(n18060) );
  XOR2_X1 U20065 ( .A(n18070), .B(n18060), .Z(n21021) );
  NOR4_X1 U20066 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21010), .A3(
        n21025), .A4(n18089), .ZN(n18068) );
  AOI21_X1 U20067 ( .B1(n18061), .B2(n19082), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18065) );
  OAI21_X1 U20068 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18063), .A(
        n18062), .ZN(n20509) );
  OAI21_X1 U20069 ( .B1(n18110), .B2(n17983), .A(n11285), .ZN(n18064) );
  NAND2_X1 U20070 ( .A1(n10979), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n21032) );
  OAI211_X1 U20071 ( .C1(n18066), .C2(n18065), .A(n18064), .B(n21032), .ZN(
        n18067) );
  AOI211_X1 U20072 ( .C1(n18197), .C2(n21021), .A(n18068), .B(n18067), .ZN(
        n18069) );
  OAI21_X1 U20073 ( .B1(n18071), .B2(n18070), .A(n18069), .ZN(P3_U2804) );
  INV_X1 U20074 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21071) );
  INV_X1 U20075 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21075) );
  NAND2_X1 U20076 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n21051), .ZN(
        n18072) );
  XOR2_X1 U20077 ( .A(n21071), .B(n18072), .Z(n21082) );
  INV_X1 U20078 ( .A(n21082), .ZN(n18085) );
  INV_X1 U20079 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n20575) );
  NOR2_X1 U20080 ( .A1(n11764), .A2(n20575), .ZN(n21079) );
  NAND2_X1 U20081 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18073), .ZN(
        n18103) );
  NOR2_X1 U20082 ( .A1(n20549), .A2(n18103), .ZN(n18075) );
  NAND2_X1 U20083 ( .A1(n18075), .A2(n18074), .ZN(n18093) );
  XNOR2_X1 U20084 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18078) );
  NOR2_X1 U20085 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18117), .ZN(
        n18111) );
  NOR2_X1 U20086 ( .A1(n19083), .A2(n18075), .ZN(n18101) );
  AOI211_X1 U20087 ( .C1(n18109), .C2(n18076), .A(n18101), .B(n18251), .ZN(
        n18104) );
  INV_X1 U20088 ( .A(n18104), .ZN(n18077) );
  NOR2_X1 U20089 ( .A1(n18111), .A2(n18077), .ZN(n18092) );
  OAI22_X1 U20090 ( .A1(n18093), .A2(n18078), .B1(n18092), .B2(n20583), .ZN(
        n18079) );
  AOI211_X1 U20091 ( .C1(n11013), .C2(n18110), .A(n21079), .B(n18079), .ZN(
        n18084) );
  NAND3_X1 U20092 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21062) );
  NOR2_X1 U20093 ( .A1(n21037), .A2(n21062), .ZN(n21049) );
  NAND2_X1 U20094 ( .A1(n21049), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18080) );
  XOR2_X1 U20095 ( .A(n18080), .B(n21071), .Z(n21078) );
  NAND2_X1 U20096 ( .A1(n18097), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n18086) );
  NAND3_X1 U20097 ( .A1(n18098), .A2(n18081), .A3(n21075), .ZN(n18087) );
  INV_X1 U20098 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21074) );
  AOI22_X1 U20099 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18086), .B1(
        n18087), .B2(n21074), .ZN(n18082) );
  XNOR2_X1 U20100 ( .A(n21071), .B(n18082), .ZN(n21083) );
  AOI22_X1 U20101 ( .A1(n21078), .A2(n18141), .B1(n18197), .B2(n21083), .ZN(
        n18083) );
  OAI211_X1 U20102 ( .C1(n18085), .C2(n18285), .A(n18084), .B(n18083), .ZN(
        P3_U2799) );
  NAND2_X1 U20103 ( .A1(n18087), .A2(n18086), .ZN(n18088) );
  XOR2_X1 U20104 ( .A(n18088), .B(n21074), .Z(n21070) );
  NOR3_X1 U20105 ( .A1(n18090), .A2(n21062), .A3(n18089), .ZN(n18095) );
  OAI22_X1 U20106 ( .A1(n21049), .A2(n18195), .B1(n21051), .B2(n18285), .ZN(
        n18107) );
  INV_X1 U20107 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n20559) );
  XNOR2_X1 U20108 ( .A(n20559), .B(n18108), .ZN(n20573) );
  AOI22_X1 U20109 ( .A1(n10979), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n18110), 
        .B2(n20573), .ZN(n18091) );
  OAI221_X1 U20110 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18093), .C1(
        n20559), .C2(n18092), .A(n18091), .ZN(n18094) );
  AOI221_X1 U20111 ( .B1(n18095), .B2(n21074), .C1(n18107), .C2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(n18094), .ZN(n18096) );
  OAI21_X1 U20112 ( .B1(n21070), .B2(n18144), .A(n18096), .ZN(P3_U2800) );
  AOI21_X1 U20113 ( .B1(n18098), .B2(n18081), .A(n18097), .ZN(n18099) );
  XOR2_X1 U20114 ( .A(n18099), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n21060) );
  OAI211_X1 U20115 ( .C1(n18100), .C2(n18285), .A(n21055), .B(n21075), .ZN(
        n18106) );
  INV_X1 U20116 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20552) );
  NOR2_X1 U20117 ( .A1(n11764), .A2(n20552), .ZN(n21058) );
  INV_X1 U20118 ( .A(n18101), .ZN(n18102) );
  OAI22_X1 U20119 ( .A1(n18104), .A2(n20549), .B1(n18103), .B2(n18102), .ZN(
        n18105) );
  AOI211_X1 U20120 ( .C1(n18107), .C2(n18106), .A(n21058), .B(n18105), .ZN(
        n18113) );
  AOI21_X1 U20121 ( .B1(n20549), .B2(n18109), .A(n18108), .ZN(n20546) );
  OAI21_X1 U20122 ( .B1(n18111), .B2(n18110), .A(n20546), .ZN(n18112) );
  OAI211_X1 U20123 ( .C1(n21060), .C2(n18144), .A(n18113), .B(n18112), .ZN(
        P3_U2801) );
  INV_X1 U20124 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n20395) );
  NAND2_X1 U20125 ( .A1(n18118), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18115) );
  AOI21_X1 U20126 ( .B1(n20395), .B2(n18115), .A(n18114), .ZN(n20379) );
  AOI21_X1 U20127 ( .B1(n18118), .B2(n19082), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18120) );
  INV_X1 U20128 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n21158) );
  OAI22_X1 U20129 ( .A1(n18120), .A2(n18119), .B1(n11764), .B2(n21158), .ZN(
        n18121) );
  AOI21_X1 U20130 ( .B1(n20379), .B2(n18253), .A(n18121), .ZN(n18126) );
  OAI21_X1 U20131 ( .B1(n18123), .B2(n21147), .A(n18122), .ZN(n21156) );
  NOR2_X1 U20132 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n11551), .ZN(
        n21155) );
  AOI22_X1 U20133 ( .A1(n18197), .A2(n21156), .B1(n18124), .B2(n21155), .ZN(
        n18125) );
  OAI211_X1 U20134 ( .C1(n18127), .C2(n21147), .A(n18126), .B(n18125), .ZN(
        P3_U2813) );
  NAND2_X1 U20135 ( .A1(n18129), .A2(n18128), .ZN(n18130) );
  XOR2_X1 U20136 ( .A(n18130), .B(n18140), .Z(n20972) );
  NAND2_X1 U20137 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18131), .ZN(
        n18133) );
  AOI21_X1 U20138 ( .B1(n18135), .B2(n18133), .A(n18132), .ZN(n20340) );
  NOR3_X1 U20139 ( .A1(n18181), .A2(n20269), .A3(n19083), .ZN(n18175) );
  NAND2_X1 U20140 ( .A1(n20298), .A2(n18175), .ZN(n18148) );
  AOI221_X1 U20141 ( .B1(n20322), .B2(n18135), .C1(n18148), .C2(n18135), .A(
        n18134), .ZN(n18137) );
  INV_X1 U20142 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18362) );
  NOR2_X1 U20143 ( .A1(n11764), .A2(n18362), .ZN(n18136) );
  AOI211_X1 U20144 ( .C1(n20340), .C2(n18253), .A(n18137), .B(n18136), .ZN(
        n18143) );
  AOI21_X1 U20145 ( .B1(n18140), .B2(n18138), .A(n20974), .ZN(n20968) );
  AOI21_X1 U20146 ( .B1(n18140), .B2(n18139), .A(n20976), .ZN(n20965) );
  AOI22_X1 U20147 ( .A1(n18225), .A2(n20968), .B1(n18141), .B2(n20965), .ZN(
        n18142) );
  OAI211_X1 U20148 ( .C1(n20972), .C2(n18144), .A(n18143), .B(n18142), .ZN(
        P3_U2816) );
  NOR2_X1 U20149 ( .A1(n18181), .A2(n20169), .ZN(n20227) );
  INV_X1 U20150 ( .A(n20227), .ZN(n18145) );
  OR2_X1 U20151 ( .A1(n20269), .A2(n18145), .ZN(n18173) );
  NOR2_X1 U20152 ( .A1(n18156), .A2(n18173), .ZN(n18155) );
  INV_X1 U20153 ( .A(n18155), .ZN(n20299) );
  AOI21_X1 U20154 ( .B1(n20309), .B2(n20299), .A(n18146), .ZN(n20302) );
  NAND2_X1 U20155 ( .A1(n18280), .A2(n18240), .ZN(n18172) );
  NAND2_X1 U20156 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18175), .ZN(
        n18163) );
  OAI21_X1 U20157 ( .B1(n18275), .B2(n20309), .A(n18163), .ZN(n18147) );
  AOI22_X1 U20158 ( .A1(n20302), .A2(n18253), .B1(n18148), .B2(n18147), .ZN(
        n18154) );
  OAI22_X1 U20159 ( .A1(n21138), .A2(n18195), .B1(n18285), .B2(n18149), .ZN(
        n18168) );
  OAI22_X1 U20160 ( .A1(n20938), .A2(n18169), .B1(n18162), .B2(n18170), .ZN(
        n18150) );
  XOR2_X1 U20161 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18150), .Z(
        n20930) );
  AOI22_X1 U20162 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18168), .B1(
        n18197), .B2(n20930), .ZN(n18153) );
  NAND2_X1 U20163 ( .A1(n10979), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18152) );
  INV_X1 U20164 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20931) );
  OAI221_X1 U20165 ( .B1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n20934), 
        .C1(n20931), .C2(n20938), .A(n18161), .ZN(n18151) );
  NAND4_X1 U20166 ( .A1(n18154), .A2(n18153), .A3(n18152), .A4(n18151), .ZN(
        P3_U2819) );
  AOI21_X1 U20167 ( .B1(n18156), .B2(n18173), .A(n18155), .ZN(n20281) );
  AOI22_X1 U20168 ( .A1(n10979), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n20281), 
        .B2(n18253), .ZN(n18167) );
  AOI221_X1 U20169 ( .B1(n18189), .B2(n18169), .C1(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18169), .A(n21177), .ZN(
        n18160) );
  AOI221_X1 U20170 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18158), .C1(
        n21199), .C2(n18157), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18159) );
  AOI221_X1 U20171 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18160), .C1(
        n11547), .C2(n18160), .A(n18159), .ZN(n21178) );
  AOI22_X1 U20172 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18168), .B1(
        n18197), .B2(n21178), .ZN(n18166) );
  NAND3_X1 U20173 ( .A1(n20938), .A2(n18162), .A3(n18161), .ZN(n18165) );
  OAI211_X1 U20174 ( .C1(n18175), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18172), .B(n18163), .ZN(n18164) );
  NAND4_X1 U20175 ( .A1(n18167), .A2(n18166), .A3(n18165), .A4(n18164), .ZN(
        P3_U2820) );
  INV_X1 U20176 ( .A(n18168), .ZN(n18179) );
  NAND2_X1 U20177 ( .A1(n18170), .A2(n18169), .ZN(n18171) );
  XOR2_X1 U20178 ( .A(n18171), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n21195) );
  INV_X1 U20179 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20289) );
  NOR2_X1 U20180 ( .A1(n11764), .A2(n20289), .ZN(n18177) );
  INV_X1 U20181 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20262) );
  INV_X1 U20182 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18208) );
  NOR2_X1 U20183 ( .A1(n20262), .A2(n18208), .ZN(n18185) );
  NOR2_X1 U20184 ( .A1(n18181), .A2(n19083), .ZN(n18200) );
  AOI22_X1 U20185 ( .A1(n18185), .A2(n18200), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18172), .ZN(n18174) );
  INV_X1 U20186 ( .A(n18181), .ZN(n18184) );
  NAND3_X1 U20187 ( .A1(n18184), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20255) );
  NOR2_X1 U20188 ( .A1(n20262), .A2(n20255), .ZN(n18183) );
  OAI21_X1 U20189 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18183), .A(
        n18173), .ZN(n20272) );
  OAI22_X1 U20190 ( .A1(n18175), .A2(n18174), .B1(n18276), .B2(n20272), .ZN(
        n18176) );
  AOI211_X1 U20191 ( .C1(n18197), .C2(n21195), .A(n18177), .B(n18176), .ZN(
        n18178) );
  OAI221_X1 U20192 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n10978), .C1(
        n21199), .C2(n18179), .A(n18178), .ZN(P3_U2821) );
  AOI21_X1 U20193 ( .B1(n18182), .B2(n18181), .A(n18251), .ZN(n18207) );
  AOI21_X1 U20194 ( .B1(n20262), .B2(n20255), .A(n18183), .ZN(n20257) );
  NAND2_X1 U20195 ( .A1(n18184), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18186) );
  AOI211_X1 U20196 ( .C1(n20262), .C2(n18186), .A(n18185), .B(n19083), .ZN(
        n18188) );
  INV_X1 U20197 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20266) );
  NOR2_X1 U20198 ( .A1(n11764), .A2(n20266), .ZN(n18187) );
  AOI211_X1 U20199 ( .C1(n20257), .C2(n18253), .A(n18188), .B(n18187), .ZN(
        n18199) );
  AOI22_X1 U20200 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18190), .B1(
        n18189), .B2(n11543), .ZN(n18191) );
  XNOR2_X1 U20201 ( .A(n18192), .B(n18191), .ZN(n20922) );
  OAI21_X1 U20202 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18194), .A(
        n18193), .ZN(n20926) );
  OAI22_X1 U20203 ( .A1(n18285), .A2(n20926), .B1(n18195), .B2(n20922), .ZN(
        n18196) );
  AOI21_X1 U20204 ( .B1(n18197), .B2(n20922), .A(n18196), .ZN(n18198) );
  OAI211_X1 U20205 ( .C1(n20262), .C2(n18207), .A(n18199), .B(n18198), .ZN(
        P3_U2822) );
  OAI21_X1 U20206 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20227), .A(
        n20255), .ZN(n20242) );
  AOI22_X1 U20207 ( .A1(n10979), .A2(P3_REIP_REG_7__SCAN_IN), .B1(n18200), 
        .B2(n18208), .ZN(n18211) );
  AOI21_X1 U20208 ( .B1(n20918), .B2(n18202), .A(n18201), .ZN(n20913) );
  OAI21_X1 U20209 ( .B1(n18205), .B2(n18204), .A(n18203), .ZN(n18206) );
  XOR2_X1 U20210 ( .A(n18206), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n20917) );
  OAI22_X1 U20211 ( .A1(n18285), .A2(n20917), .B1(n18208), .B2(n18207), .ZN(
        n18209) );
  AOI21_X1 U20212 ( .B1(n18279), .B2(n20913), .A(n18209), .ZN(n18210) );
  OAI211_X1 U20213 ( .C1(n18276), .C2(n20242), .A(n18211), .B(n18210), .ZN(
        P3_U2823) );
  NAND2_X1 U20214 ( .A1(n18214), .A2(n19082), .ZN(n18221) );
  AOI21_X1 U20215 ( .B1(n11082), .B2(n18213), .A(n18212), .ZN(n20903) );
  AOI22_X1 U20216 ( .A1(n10979), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18279), 
        .B2(n20903), .ZN(n18220) );
  AOI21_X1 U20217 ( .B1(n19082), .B2(n18214), .A(n18275), .ZN(n18229) );
  INV_X1 U20218 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18215) );
  NAND2_X1 U20219 ( .A1(n18214), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18222) );
  AOI21_X1 U20220 ( .B1(n18215), .B2(n18222), .A(n20227), .ZN(n20231) );
  INV_X1 U20221 ( .A(n20231), .ZN(n20228) );
  OAI21_X1 U20222 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18217), .A(
        n18216), .ZN(n20906) );
  OAI22_X1 U20223 ( .A1(n18276), .A2(n20228), .B1(n18285), .B2(n20906), .ZN(
        n18218) );
  AOI21_X1 U20224 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18229), .A(
        n18218), .ZN(n18219) );
  OAI211_X1 U20225 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18221), .A(
        n18220), .B(n18219), .ZN(P3_U2824) );
  NOR2_X1 U20226 ( .A1(n20196), .A2(n20169), .ZN(n18242) );
  OAI21_X1 U20227 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18242), .A(
        n18222), .ZN(n20214) );
  XOR2_X1 U20228 ( .A(n18224), .B(n18223), .Z(n20892) );
  AOI22_X1 U20229 ( .A1(n10979), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18225), 
        .B2(n20892), .ZN(n18231) );
  AOI21_X1 U20230 ( .B1(n20891), .B2(n18227), .A(n18226), .ZN(n20895) );
  OAI21_X1 U20231 ( .B1(n18251), .B2(n20196), .A(n20225), .ZN(n18228) );
  AOI22_X1 U20232 ( .A1(n18279), .A2(n20895), .B1(n18229), .B2(n18228), .ZN(
        n18230) );
  OAI211_X1 U20233 ( .C1(n18276), .C2(n20214), .A(n18231), .B(n18230), .ZN(
        P3_U2825) );
  AOI21_X1 U20234 ( .B1(n20883), .B2(n18232), .A(n21050), .ZN(n18238) );
  AOI211_X1 U20235 ( .C1(n18235), .C2(n18234), .A(n18233), .B(n21210), .ZN(
        n18236) );
  AOI21_X1 U20236 ( .B1(n18238), .B2(n18237), .A(n18236), .ZN(n20885) );
  NOR2_X1 U20237 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19083), .ZN(
        n18239) );
  AOI22_X1 U20238 ( .A1(n10979), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18241), 
        .B2(n18239), .ZN(n18244) );
  OAI21_X1 U20239 ( .B1(n18241), .B2(n18240), .A(n18280), .ZN(n18256) );
  INV_X1 U20240 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20200) );
  NAND2_X1 U20241 ( .A1(n18241), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18252) );
  AOI21_X1 U20242 ( .B1(n20200), .B2(n18252), .A(n18242), .ZN(n20199) );
  AOI22_X1 U20243 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18256), .B1(
        n20199), .B2(n18253), .ZN(n18243) );
  OAI211_X1 U20244 ( .C1(n20885), .C2(n21259), .A(n18244), .B(n18243), .ZN(
        P3_U2826) );
  OAI21_X1 U20245 ( .B1(n18247), .B2(n18246), .A(n18245), .ZN(n20882) );
  AOI21_X1 U20246 ( .B1(n18250), .B2(n18249), .A(n18248), .ZN(n20879) );
  AOI22_X1 U20247 ( .A1(n10979), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18279), 
        .B2(n20879), .ZN(n18258) );
  OAI21_X1 U20248 ( .B1(n18251), .B2(n20180), .A(n20181), .ZN(n18255) );
  NOR2_X1 U20249 ( .A1(n20180), .A2(n20169), .ZN(n20170) );
  OAI21_X1 U20250 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20170), .A(
        n18252), .ZN(n20183) );
  INV_X1 U20251 ( .A(n20183), .ZN(n18254) );
  AOI22_X1 U20252 ( .A1(n18256), .A2(n18255), .B1(n18254), .B2(n18253), .ZN(
        n18257) );
  OAI211_X1 U20253 ( .C1(n18285), .C2(n20882), .A(n18258), .B(n18257), .ZN(
        P3_U2827) );
  AOI21_X1 U20254 ( .B1(n20180), .B2(n20169), .A(n20170), .ZN(n18259) );
  INV_X1 U20255 ( .A(n18259), .ZN(n20173) );
  XOR2_X1 U20256 ( .A(n18261), .B(n18260), .Z(n18266) );
  AOI211_X1 U20257 ( .C1(n18264), .C2(n18263), .A(n18262), .B(n21210), .ZN(
        n18265) );
  AOI21_X1 U20258 ( .B1(n18266), .B2(n21203), .A(n18265), .ZN(n20866) );
  OAI22_X1 U20259 ( .A1(n18276), .A2(n20173), .B1(n20866), .B2(n21259), .ZN(
        n18267) );
  AOI21_X1 U20260 ( .B1(n10979), .B2(P3_REIP_REG_2__SCAN_IN), .A(n18267), .ZN(
        n18268) );
  OAI221_X1 U20261 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19083), .C1(
        n20180), .C2(n18280), .A(n18268), .ZN(P3_U2828) );
  AOI21_X1 U20262 ( .B1(n18270), .B2(n18278), .A(n18269), .ZN(n20855) );
  AOI21_X1 U20263 ( .B1(n18272), .B2(n18277), .A(n18271), .ZN(n20862) );
  OAI22_X1 U20264 ( .A1(n20862), .A2(n18285), .B1(n11764), .B2(n18357), .ZN(
        n18273) );
  AOI21_X1 U20265 ( .B1(n18279), .B2(n20855), .A(n18273), .ZN(n18274) );
  OAI221_X1 U20266 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18276), .C1(
        n20169), .C2(n18275), .A(n18274), .ZN(P3_U2829) );
  NAND2_X1 U20267 ( .A1(n18278), .A2(n18277), .ZN(n20849) );
  INV_X1 U20268 ( .A(n20849), .ZN(n20850) );
  INV_X1 U20269 ( .A(n18279), .ZN(n18284) );
  NAND3_X1 U20270 ( .A1(n20789), .A2(n18281), .A3(n18280), .ZN(n18282) );
  AOI22_X1 U20271 ( .A1(n10979), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18282), .ZN(n18283) );
  OAI221_X1 U20272 ( .B1(n20850), .B2(n18285), .C1(n20849), .C2(n18284), .A(
        n18283), .ZN(P3_U2830) );
  INV_X1 U20273 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21222) );
  NAND2_X1 U20274 ( .A1(n18795), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18778) );
  INV_X1 U20275 ( .A(n18778), .ZN(n18780) );
  NAND2_X1 U20276 ( .A1(n21222), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18803) );
  INV_X1 U20277 ( .A(n18803), .ZN(n18804) );
  NOR2_X1 U20278 ( .A1(n18780), .A2(n18804), .ZN(n18287) );
  OAI22_X1 U20279 ( .A1(n18288), .A2(n21222), .B1(n18287), .B2(n18286), .ZN(
        P3_U2866) );
  NAND2_X1 U20280 ( .A1(n18290), .A2(n18289), .ZN(n18293) );
  OAI21_X1 U20281 ( .B1(n18291), .B2(n18774), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18292) );
  OAI21_X1 U20282 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18293), .A(
        n18292), .ZN(P3_U2864) );
  NOR4_X1 U20283 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18297) );
  NOR4_X1 U20284 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18296) );
  NOR4_X1 U20285 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18295) );
  NOR4_X1 U20286 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18294) );
  NAND4_X1 U20287 ( .A1(n18297), .A2(n18296), .A3(n18295), .A4(n18294), .ZN(
        n18303) );
  NOR4_X1 U20288 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18301) );
  AOI211_X1 U20289 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18300) );
  NOR4_X1 U20290 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18299) );
  NOR4_X1 U20291 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18298) );
  NAND4_X1 U20292 ( .A1(n18301), .A2(n18300), .A3(n18299), .A4(n18298), .ZN(
        n18302) );
  NOR2_X1 U20293 ( .A1(n18303), .A2(n18302), .ZN(n18316) );
  INV_X1 U20294 ( .A(n18316), .ZN(n18313) );
  NOR2_X1 U20295 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18305) );
  NAND2_X1 U20296 ( .A1(n18313), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18304) );
  OAI21_X1 U20297 ( .B1(n18313), .B2(n18305), .A(n18304), .ZN(P3_U3293) );
  AOI211_X1 U20298 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18306) );
  AOI21_X1 U20299 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18306), .ZN(n18308) );
  INV_X1 U20300 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18307) );
  AOI22_X1 U20301 ( .A1(n18316), .A2(n18308), .B1(n18307), .B2(n18313), .ZN(
        P3_U3292) );
  INV_X1 U20302 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18310) );
  NOR3_X1 U20303 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18312) );
  NOR2_X1 U20304 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18312), .ZN(n18309) );
  MUX2_X1 U20305 ( .A(n18310), .B(n18309), .S(n18316), .Z(n18311) );
  INV_X1 U20306 ( .A(n18311), .ZN(P3_U2638) );
  INV_X1 U20307 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21604) );
  AOI21_X1 U20308 ( .B1(n18357), .B2(n21604), .A(n18312), .ZN(n18315) );
  INV_X1 U20309 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18314) );
  AOI22_X1 U20310 ( .A1(n18316), .A2(n18315), .B1(n18314), .B2(n18313), .ZN(
        P3_U2639) );
  OAI22_X1 U20311 ( .A1(n21651), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18364), .ZN(n18317) );
  INV_X1 U20312 ( .A(n18317), .ZN(P3_U3297) );
  INV_X1 U20313 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18318) );
  AOI22_X1 U20314 ( .A1(n18364), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18318), 
        .B2(n21651), .ZN(P3_U3294) );
  AOI21_X1 U20315 ( .B1(n21654), .B2(n21645), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18319) );
  AOI22_X1 U20316 ( .A1(n18364), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18319), 
        .B2(n21651), .ZN(P3_U2635) );
  INV_X1 U20317 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20785) );
  AOI22_X1 U20318 ( .A1(n18353), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18320) );
  OAI21_X1 U20319 ( .B1(n20785), .B2(n18336), .A(n18320), .ZN(P3_U2767) );
  INV_X1 U20320 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20141) );
  AOI22_X1 U20321 ( .A1(n18353), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18321) );
  OAI21_X1 U20322 ( .B1(n20141), .B2(n18336), .A(n18321), .ZN(P3_U2766) );
  INV_X1 U20323 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20648) );
  AOI22_X1 U20324 ( .A1(n18353), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18322) );
  OAI21_X1 U20325 ( .B1(n20648), .B2(n18336), .A(n18322), .ZN(P3_U2765) );
  INV_X1 U20326 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20144) );
  AOI22_X1 U20327 ( .A1(n18353), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18323) );
  OAI21_X1 U20328 ( .B1(n20144), .B2(n18336), .A(n18323), .ZN(P3_U2764) );
  INV_X1 U20329 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n20623) );
  AOI22_X1 U20330 ( .A1(n18353), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18324) );
  OAI21_X1 U20331 ( .B1(n20623), .B2(n18336), .A(n18324), .ZN(P3_U2763) );
  INV_X1 U20332 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20147) );
  AOI22_X1 U20333 ( .A1(n18353), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18325) );
  OAI21_X1 U20334 ( .B1(n20147), .B2(n18336), .A(n18325), .ZN(P3_U2762) );
  INV_X1 U20335 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20624) );
  AOI22_X1 U20336 ( .A1(n18353), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18326) );
  OAI21_X1 U20337 ( .B1(n20624), .B2(n18336), .A(n18326), .ZN(P3_U2761) );
  INV_X1 U20338 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20151) );
  AOI22_X1 U20339 ( .A1(n18353), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18327) );
  OAI21_X1 U20340 ( .B1(n20151), .B2(n18336), .A(n18327), .ZN(P3_U2760) );
  INV_X1 U20341 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20772) );
  AOI22_X1 U20342 ( .A1(n18353), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18328) );
  OAI21_X1 U20343 ( .B1(n20772), .B2(n18336), .A(n18328), .ZN(P3_U2759) );
  INV_X1 U20344 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20154) );
  AOI22_X1 U20345 ( .A1(n18353), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18329) );
  OAI21_X1 U20346 ( .B1(n20154), .B2(n18336), .A(n18329), .ZN(P3_U2758) );
  INV_X1 U20347 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20156) );
  AOI22_X1 U20348 ( .A1(n18353), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18330) );
  OAI21_X1 U20349 ( .B1(n20156), .B2(n18336), .A(n18330), .ZN(P3_U2757) );
  INV_X1 U20350 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20611) );
  AOI22_X1 U20351 ( .A1(n18353), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18331) );
  OAI21_X1 U20352 ( .B1(n20611), .B2(n18336), .A(n18331), .ZN(P3_U2756) );
  INV_X1 U20353 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20159) );
  AOI22_X1 U20354 ( .A1(n18353), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18332) );
  OAI21_X1 U20355 ( .B1(n20159), .B2(n18336), .A(n18332), .ZN(P3_U2755) );
  INV_X1 U20356 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20161) );
  AOI22_X1 U20357 ( .A1(n18353), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18333) );
  OAI21_X1 U20358 ( .B1(n20161), .B2(n18336), .A(n18333), .ZN(P3_U2754) );
  INV_X1 U20359 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20758) );
  AOI22_X1 U20360 ( .A1(n18353), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18334) );
  OAI21_X1 U20361 ( .B1(n20758), .B2(n18336), .A(n18334), .ZN(P3_U2753) );
  INV_X1 U20362 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20167) );
  AOI22_X1 U20363 ( .A1(n18353), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18335) );
  OAI21_X1 U20364 ( .B1(n20167), .B2(n18336), .A(n18335), .ZN(P3_U2752) );
  INV_X1 U20365 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20749) );
  AOI22_X1 U20366 ( .A1(n18353), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18338) );
  OAI21_X1 U20367 ( .B1(n20749), .B2(n18355), .A(n18338), .ZN(P3_U2751) );
  INV_X1 U20368 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20118) );
  AOI22_X1 U20369 ( .A1(n18353), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18339) );
  OAI21_X1 U20370 ( .B1(n20118), .B2(n18355), .A(n18339), .ZN(P3_U2750) );
  INV_X1 U20371 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20120) );
  AOI22_X1 U20372 ( .A1(n18353), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18340) );
  OAI21_X1 U20373 ( .B1(n20120), .B2(n18355), .A(n18340), .ZN(P3_U2749) );
  INV_X1 U20374 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20676) );
  AOI22_X1 U20375 ( .A1(n18353), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18341) );
  OAI21_X1 U20376 ( .B1(n20676), .B2(n18355), .A(n18341), .ZN(P3_U2748) );
  INV_X1 U20377 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20123) );
  AOI22_X1 U20378 ( .A1(n18353), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18342) );
  OAI21_X1 U20379 ( .B1(n20123), .B2(n18355), .A(n18342), .ZN(P3_U2747) );
  INV_X1 U20380 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20125) );
  AOI22_X1 U20381 ( .A1(n18353), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18343) );
  OAI21_X1 U20382 ( .B1(n20125), .B2(n18355), .A(n18343), .ZN(P3_U2746) );
  INV_X1 U20383 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20671) );
  AOI22_X1 U20384 ( .A1(n18353), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18344) );
  OAI21_X1 U20385 ( .B1(n20671), .B2(n18355), .A(n18344), .ZN(P3_U2745) );
  INV_X1 U20386 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20736) );
  AOI22_X1 U20387 ( .A1(n18353), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18345) );
  OAI21_X1 U20388 ( .B1(n20736), .B2(n18355), .A(n18345), .ZN(P3_U2744) );
  INV_X1 U20389 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20729) );
  AOI22_X1 U20390 ( .A1(n18353), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18346) );
  OAI21_X1 U20391 ( .B1(n20729), .B2(n18355), .A(n18346), .ZN(P3_U2743) );
  INV_X1 U20392 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20691) );
  AOI22_X1 U20393 ( .A1(n18353), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18347) );
  OAI21_X1 U20394 ( .B1(n20691), .B2(n18355), .A(n18347), .ZN(P3_U2742) );
  INV_X1 U20395 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20132) );
  AOI22_X1 U20396 ( .A1(n18353), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18349) );
  OAI21_X1 U20397 ( .B1(n20132), .B2(n18355), .A(n18349), .ZN(P3_U2741) );
  INV_X1 U20398 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20134) );
  AOI22_X1 U20399 ( .A1(n18353), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18350) );
  OAI21_X1 U20400 ( .B1(n20134), .B2(n18355), .A(n18350), .ZN(P3_U2740) );
  INV_X1 U20401 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20717) );
  AOI22_X1 U20402 ( .A1(n18353), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18351) );
  OAI21_X1 U20403 ( .B1(n20717), .B2(n18355), .A(n18351), .ZN(P3_U2739) );
  INV_X1 U20404 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20137) );
  AOI22_X1 U20405 ( .A1(n18353), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18352) );
  OAI21_X1 U20406 ( .B1(n20137), .B2(n18355), .A(n18352), .ZN(P3_U2738) );
  INV_X1 U20407 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20711) );
  AOI22_X1 U20408 ( .A1(n18353), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18348), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18354) );
  OAI21_X1 U20409 ( .B1(n20711), .B2(n18355), .A(n18354), .ZN(P3_U2737) );
  AOI21_X1 U20410 ( .B1(n21651), .B2(P3_ADS_N_REG_SCAN_IN), .A(n21605), .ZN(
        n18356) );
  INV_X1 U20411 ( .A(n18356), .ZN(P3_U2633) );
  NOR2_X1 U20412 ( .A1(n21651), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18358) );
  INV_X1 U20413 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20168) );
  INV_X1 U20414 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19822) );
  OAI222_X1 U20415 ( .A1(n18365), .A2(n20168), .B1(n19822), .B2(n18364), .C1(
        n18357), .C2(n18363), .ZN(P3_U3032) );
  AOI22_X1 U20416 ( .A1(n18358), .A2(P3_REIP_REG_3__SCAN_IN), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n21651), .ZN(n18359) );
  OAI21_X1 U20417 ( .B1(n18363), .B2(n20168), .A(n18359), .ZN(P3_U3033) );
  INV_X1 U20418 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U20419 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n18360), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n21651), .ZN(n18361) );
  OAI21_X1 U20420 ( .B1(n20890), .B2(n18365), .A(n18361), .ZN(P3_U3034) );
  INV_X1 U20421 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20219) );
  INV_X1 U20422 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19826) );
  OAI222_X1 U20423 ( .A1(n18365), .A2(n20219), .B1(n19826), .B2(n18364), .C1(
        n20890), .C2(n18363), .ZN(P3_U3035) );
  INV_X1 U20424 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20237) );
  INV_X1 U20425 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19828) );
  OAI222_X1 U20426 ( .A1(n18365), .A2(n20237), .B1(n19828), .B2(n18364), .C1(
        n20219), .C2(n18363), .ZN(P3_U3036) );
  INV_X1 U20427 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20245) );
  INV_X1 U20428 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19830) );
  OAI222_X1 U20429 ( .A1(n18365), .A2(n20245), .B1(n19830), .B2(n18364), .C1(
        n20237), .C2(n18363), .ZN(P3_U3037) );
  INV_X1 U20430 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19832) );
  OAI222_X1 U20431 ( .A1(n18365), .A2(n20266), .B1(n19832), .B2(n18364), .C1(
        n20245), .C2(n18363), .ZN(P3_U3038) );
  INV_X1 U20432 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19835) );
  OAI222_X1 U20433 ( .A1(n18365), .A2(n20289), .B1(n19835), .B2(n18364), .C1(
        n20266), .C2(n18363), .ZN(P3_U3039) );
  INV_X1 U20434 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20290) );
  INV_X1 U20435 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19837) );
  OAI222_X1 U20436 ( .A1(n18365), .A2(n20290), .B1(n19837), .B2(n18364), .C1(
        n20289), .C2(n18363), .ZN(P3_U3040) );
  INV_X1 U20437 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20295) );
  INV_X1 U20438 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19839) );
  OAI222_X1 U20439 ( .A1(n18365), .A2(n20295), .B1(n19839), .B2(n18364), .C1(
        n20290), .C2(n18363), .ZN(P3_U3041) );
  INV_X1 U20440 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19841) );
  OAI222_X1 U20441 ( .A1(n20295), .A2(n18363), .B1(n19841), .B2(n18364), .C1(
        n20321), .C2(n18365), .ZN(P3_U3042) );
  INV_X1 U20442 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19843) );
  OAI222_X1 U20443 ( .A1(n18365), .A2(n20331), .B1(n19843), .B2(n18364), .C1(
        n20321), .C2(n18363), .ZN(P3_U3043) );
  INV_X1 U20444 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19845) );
  OAI222_X1 U20445 ( .A1(n20331), .A2(n18363), .B1(n19845), .B2(n18364), .C1(
        n18362), .C2(n18365), .ZN(P3_U3044) );
  INV_X1 U20446 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19847) );
  OAI222_X1 U20447 ( .A1(n18365), .A2(n20371), .B1(n19847), .B2(n18364), .C1(
        n18362), .C2(n18363), .ZN(P3_U3045) );
  INV_X1 U20448 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20373) );
  INV_X1 U20449 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19849) );
  OAI222_X1 U20450 ( .A1(n18365), .A2(n20373), .B1(n19849), .B2(n18364), .C1(
        n20371), .C2(n18363), .ZN(P3_U3046) );
  INV_X1 U20451 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19851) );
  OAI222_X1 U20452 ( .A1(n18365), .A2(n21158), .B1(n19851), .B2(n18364), .C1(
        n20373), .C2(n18363), .ZN(P3_U3047) );
  INV_X1 U20453 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19853) );
  OAI222_X1 U20454 ( .A1(n18365), .A2(n21152), .B1(n19853), .B2(n18364), .C1(
        n21158), .C2(n18363), .ZN(P3_U3048) );
  INV_X1 U20455 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19855) );
  OAI222_X1 U20456 ( .A1(n18365), .A2(n20408), .B1(n19855), .B2(n18364), .C1(
        n21152), .C2(n18363), .ZN(P3_U3049) );
  INV_X1 U20457 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19857) );
  INV_X1 U20458 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n20425) );
  OAI222_X1 U20459 ( .A1(n20408), .A2(n18363), .B1(n19857), .B2(n18364), .C1(
        n20425), .C2(n18365), .ZN(P3_U3050) );
  INV_X1 U20460 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19859) );
  OAI222_X1 U20461 ( .A1(n18365), .A2(n20846), .B1(n19859), .B2(n18364), .C1(
        n20425), .C2(n18363), .ZN(P3_U3051) );
  INV_X1 U20462 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20463) );
  INV_X1 U20463 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19861) );
  OAI222_X1 U20464 ( .A1(n18365), .A2(n20463), .B1(n19861), .B2(n18364), .C1(
        n20846), .C2(n18363), .ZN(P3_U3052) );
  INV_X1 U20465 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19863) );
  OAI222_X1 U20466 ( .A1(n18365), .A2(n20474), .B1(n19863), .B2(n18364), .C1(
        n20463), .C2(n18363), .ZN(P3_U3053) );
  INV_X1 U20467 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19865) );
  INV_X1 U20468 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20488) );
  OAI222_X1 U20469 ( .A1(n20474), .A2(n18363), .B1(n19865), .B2(n18364), .C1(
        n20488), .C2(n18365), .ZN(P3_U3054) );
  INV_X1 U20470 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20500) );
  INV_X1 U20471 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19867) );
  OAI222_X1 U20472 ( .A1(n18365), .A2(n20500), .B1(n19867), .B2(n18364), .C1(
        n20488), .C2(n18363), .ZN(P3_U3055) );
  INV_X1 U20473 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19869) );
  INV_X1 U20474 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20499) );
  OAI222_X1 U20475 ( .A1(n20500), .A2(n18363), .B1(n19869), .B2(n18364), .C1(
        n20499), .C2(n18365), .ZN(P3_U3056) );
  INV_X1 U20476 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20529) );
  INV_X1 U20477 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19871) );
  OAI222_X1 U20478 ( .A1(n18365), .A2(n20529), .B1(n19871), .B2(n18364), .C1(
        n20499), .C2(n18363), .ZN(P3_U3057) );
  INV_X1 U20479 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19873) );
  OAI222_X1 U20480 ( .A1(n18365), .A2(n20539), .B1(n19873), .B2(n18364), .C1(
        n20529), .C2(n18363), .ZN(P3_U3058) );
  INV_X1 U20481 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19875) );
  OAI222_X1 U20482 ( .A1(n20539), .A2(n18363), .B1(n19875), .B2(n18364), .C1(
        n20552), .C2(n18365), .ZN(P3_U3059) );
  INV_X1 U20483 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n20569) );
  INV_X1 U20484 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19877) );
  OAI222_X1 U20485 ( .A1(n18365), .A2(n20569), .B1(n19877), .B2(n18364), .C1(
        n20552), .C2(n18363), .ZN(P3_U3060) );
  INV_X1 U20486 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19880) );
  OAI222_X1 U20487 ( .A1(n18365), .A2(n20575), .B1(n19880), .B2(n18364), .C1(
        n20569), .C2(n18363), .ZN(P3_U3061) );
  MUX2_X1 U20488 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .B(P3_BE_N_REG_0__SCAN_IN), .S(n21651), .Z(P3_U3277) );
  MUX2_X1 U20489 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .B(P3_BE_N_REG_1__SCAN_IN), .S(n21651), .Z(P3_U3276) );
  OAI22_X1 U20490 ( .A1(n21651), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18364), .ZN(n18366) );
  INV_X1 U20491 ( .A(n18366), .ZN(P3_U3275) );
  OAI22_X1 U20492 ( .A1(n21651), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18364), .ZN(n18367) );
  INV_X1 U20493 ( .A(n18367), .ZN(P3_U3274) );
  NOR4_X1 U20494 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18370)
         );
  INV_X1 U20495 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18368) );
  NOR4_X1 U20496 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18368), .ZN(n18369) );
  NAND3_X1 U20497 ( .A1(n18370), .A2(n18369), .A3(U215), .ZN(U213) );
  NAND2_X1 U20498 ( .A1(n18716), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n18375) );
  AOI21_X1 U20499 ( .B1(n18372), .B2(n18718), .A(n18371), .ZN(n18373) );
  OAI21_X1 U20500 ( .B1(n18374), .B2(n18375), .A(n18373), .ZN(n18383) );
  INV_X1 U20501 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21625) );
  INV_X1 U20502 ( .A(n18375), .ZN(n18376) );
  NOR2_X1 U20503 ( .A1(n18705), .A2(n18376), .ZN(n18381) );
  AOI21_X1 U20504 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n21630), .A(n18377), 
        .ZN(n18379) );
  NOR3_X1 U20505 ( .A1(n19703), .A2(n18711), .A3(n21630), .ZN(n18378) );
  MUX2_X1 U20506 ( .A(n18379), .B(n18378), .S(n12651), .Z(n18380) );
  OAI21_X1 U20507 ( .B1(n18381), .B2(n18380), .A(n18383), .ZN(n18382) );
  OAI21_X1 U20508 ( .B1(n18383), .B2(n21625), .A(n18382), .ZN(P2_U3610) );
  OR2_X1 U20509 ( .A1(n18386), .A2(n18385), .ZN(n18387) );
  NAND2_X1 U20510 ( .A1(n12658), .A2(n18387), .ZN(n19687) );
  INV_X1 U20511 ( .A(n19687), .ZN(n19693) );
  AOI22_X1 U20512 ( .A1(n18644), .A2(n19693), .B1(P2_EBX_REG_0__SCAN_IN), .B2(
        n18640), .ZN(n18389) );
  NAND2_X1 U20513 ( .A1(n18639), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n18388) );
  OAI211_X1 U20514 ( .C1(n18390), .C2(n18529), .A(n18389), .B(n18388), .ZN(
        n18392) );
  NOR2_X1 U20515 ( .A1(n19425), .A2(n18400), .ZN(n18391) );
  AOI211_X1 U20516 ( .C1(n18645), .C2(n18393), .A(n18392), .B(n18391), .ZN(
        n18395) );
  NAND2_X1 U20517 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18641), .ZN(
        n18394) );
  OAI211_X1 U20518 ( .C1(n15283), .C2(n18701), .A(n18395), .B(n18394), .ZN(
        P2_U2855) );
  INV_X1 U20519 ( .A(n19481), .ZN(n19432) );
  OAI22_X1 U20520 ( .A1(n18396), .A2(n18598), .B1(n12266), .B2(n18627), .ZN(
        n18397) );
  AOI211_X1 U20521 ( .C1(n18644), .C2(n19432), .A(n18532), .B(n18397), .ZN(
        n18410) );
  AOI22_X1 U20522 ( .A1(n18398), .A2(n18642), .B1(n18641), .B2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18409) );
  OAI22_X1 U20523 ( .A1(n19484), .A2(n18400), .B1(n18601), .B2(n18399), .ZN(
        n18401) );
  INV_X1 U20524 ( .A(n18401), .ZN(n18408) );
  INV_X1 U20525 ( .A(n18402), .ZN(n18406) );
  NOR2_X1 U20526 ( .A1(n18517), .A2(n18403), .ZN(n18405) );
  AOI21_X1 U20527 ( .B1(n18406), .B2(n18405), .A(n18701), .ZN(n18404) );
  OAI21_X1 U20528 ( .B1(n18406), .B2(n18405), .A(n18404), .ZN(n18407) );
  NAND4_X1 U20529 ( .A1(n18410), .A2(n18409), .A3(n18408), .A4(n18407), .ZN(
        P2_U2851) );
  NAND2_X1 U20530 ( .A1(n15429), .A2(n18411), .ZN(n18413) );
  XOR2_X1 U20531 ( .A(n18413), .B(n18412), .Z(n18420) );
  AOI22_X1 U20532 ( .A1(n18414), .A2(n18642), .B1(P2_REIP_REG_7__SCAN_IN), 
        .B2(n18639), .ZN(n18415) );
  OAI211_X1 U20533 ( .C1(n12401), .C2(n18598), .A(n18415), .B(n18680), .ZN(
        n18418) );
  OAI22_X1 U20534 ( .A1(n19221), .A2(n18638), .B1(n18416), .B2(n18601), .ZN(
        n18417) );
  AOI211_X1 U20535 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18641), .A(
        n18418), .B(n18417), .ZN(n18419) );
  OAI21_X1 U20536 ( .B1(n18420), .B2(n18701), .A(n18419), .ZN(P2_U2848) );
  AOI22_X1 U20537 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18641), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18639), .ZN(n18421) );
  OAI21_X1 U20538 ( .B1(n18422), .B2(n18529), .A(n18421), .ZN(n18423) );
  AOI211_X1 U20539 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n18640), .A(n18532), .B(
        n18423), .ZN(n18431) );
  NOR2_X1 U20540 ( .A1(n18517), .A2(n18424), .ZN(n18426) );
  XNOR2_X1 U20541 ( .A(n18426), .B(n18425), .ZN(n18429) );
  INV_X1 U20542 ( .A(n18427), .ZN(n18428) );
  AOI22_X1 U20543 ( .A1(n18429), .A2(n18617), .B1(n18428), .B2(n18645), .ZN(
        n18430) );
  OAI211_X1 U20544 ( .C1(n18638), .C2(n19217), .A(n18431), .B(n18430), .ZN(
        P2_U2847) );
  AOI211_X1 U20545 ( .C1(n18440), .C2(n18432), .A(n18449), .B(n18647), .ZN(
        n18439) );
  OAI22_X1 U20546 ( .A1(n18434), .A2(n18598), .B1(n18433), .B2(n18627), .ZN(
        n18435) );
  AOI211_X1 U20547 ( .C1(n19204), .C2(n18644), .A(n18500), .B(n18435), .ZN(
        n18436) );
  OAI21_X1 U20548 ( .B1(n18437), .B2(n18529), .A(n18436), .ZN(n18438) );
  AOI211_X1 U20549 ( .C1(n18641), .C2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n18439), .B(n18438), .ZN(n18445) );
  INV_X1 U20550 ( .A(n18440), .ZN(n18441) );
  OAI22_X1 U20551 ( .A1(n18442), .A2(n18601), .B1(n18441), .B2(n18509), .ZN(
        n18443) );
  INV_X1 U20552 ( .A(n18443), .ZN(n18444) );
  NAND2_X1 U20553 ( .A1(n18445), .A2(n18444), .ZN(P2_U2844) );
  AOI22_X1 U20554 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18641), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18639), .ZN(n18446) );
  OAI21_X1 U20555 ( .B1(n18447), .B2(n18529), .A(n18446), .ZN(n18448) );
  AOI211_X1 U20556 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n18640), .A(n18500), .B(
        n18448), .ZN(n18456) );
  NOR2_X1 U20557 ( .A1(n18517), .A2(n18449), .ZN(n18451) );
  XNOR2_X1 U20558 ( .A(n18451), .B(n18450), .ZN(n18454) );
  INV_X1 U20559 ( .A(n18452), .ZN(n18453) );
  AOI22_X1 U20560 ( .A1(n18454), .A2(n18617), .B1(n18453), .B2(n18645), .ZN(
        n18455) );
  OAI211_X1 U20561 ( .C1(n19202), .C2(n18638), .A(n18456), .B(n18455), .ZN(
        P2_U2843) );
  NAND2_X1 U20562 ( .A1(n18606), .A2(n18457), .ZN(n18458) );
  XOR2_X1 U20563 ( .A(n18459), .B(n18458), .Z(n18469) );
  OAI21_X1 U20564 ( .B1(n18460), .B2(n18598), .A(n18680), .ZN(n18464) );
  INV_X1 U20565 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18461) );
  OAI22_X1 U20566 ( .A1(n18462), .A2(n18529), .B1(n18461), .B2(n18596), .ZN(
        n18463) );
  AOI211_X1 U20567 ( .C1(P2_REIP_REG_13__SCAN_IN), .C2(n18639), .A(n18464), 
        .B(n18463), .ZN(n18468) );
  INV_X1 U20568 ( .A(n18465), .ZN(n19197) );
  AOI22_X1 U20569 ( .A1(n18466), .A2(n18645), .B1(n19197), .B2(n18644), .ZN(
        n18467) );
  OAI211_X1 U20570 ( .C1(n18701), .C2(n18469), .A(n18468), .B(n18467), .ZN(
        P2_U2842) );
  AOI22_X1 U20571 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18641), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18639), .ZN(n18470) );
  OAI21_X1 U20572 ( .B1(n18471), .B2(n18529), .A(n18470), .ZN(n18472) );
  AOI211_X1 U20573 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n18640), .A(n18532), .B(
        n18472), .ZN(n18480) );
  NOR2_X1 U20574 ( .A1(n18517), .A2(n18473), .ZN(n18475) );
  XNOR2_X1 U20575 ( .A(n18475), .B(n18474), .ZN(n18478) );
  INV_X1 U20576 ( .A(n18476), .ZN(n18477) );
  AOI22_X1 U20577 ( .A1(n18478), .A2(n18617), .B1(n18477), .B2(n18645), .ZN(
        n18479) );
  OAI211_X1 U20578 ( .C1(n19196), .C2(n18638), .A(n18480), .B(n18479), .ZN(
        P2_U2841) );
  OAI21_X1 U20579 ( .B1(n18481), .B2(n18598), .A(n18680), .ZN(n18486) );
  INV_X1 U20580 ( .A(n18482), .ZN(n18484) );
  INV_X1 U20581 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18483) );
  OAI22_X1 U20582 ( .A1(n18484), .A2(n18529), .B1(n18483), .B2(n18596), .ZN(
        n18485) );
  AOI211_X1 U20583 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n18639), .A(n18486), 
        .B(n18485), .ZN(n18494) );
  NOR2_X1 U20584 ( .A1(n18517), .A2(n18487), .ZN(n18489) );
  XNOR2_X1 U20585 ( .A(n18489), .B(n18488), .ZN(n18492) );
  INV_X1 U20586 ( .A(n18490), .ZN(n18491) );
  AOI22_X1 U20587 ( .A1(n18492), .A2(n18617), .B1(n18491), .B2(n18645), .ZN(
        n18493) );
  OAI211_X1 U20588 ( .C1(n18495), .C2(n18638), .A(n18494), .B(n18493), .ZN(
        P2_U2839) );
  INV_X1 U20589 ( .A(n18497), .ZN(n18510) );
  AOI211_X1 U20590 ( .C1(n18497), .C2(n18496), .A(n18516), .B(n18647), .ZN(
        n18504) );
  NOR2_X1 U20591 ( .A1(n18627), .A2(n18498), .ZN(n18499) );
  AOI211_X1 U20592 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n18640), .A(n18500), .B(
        n18499), .ZN(n18501) );
  OAI21_X1 U20593 ( .B1(n18502), .B2(n18529), .A(n18501), .ZN(n18503) );
  AOI211_X1 U20594 ( .C1(n18641), .C2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n18504), .B(n18503), .ZN(n18508) );
  AOI22_X1 U20595 ( .A1(n18506), .A2(n18645), .B1(n18644), .B2(n18505), .ZN(
        n18507) );
  OAI211_X1 U20596 ( .C1(n18510), .C2(n18509), .A(n18508), .B(n18507), .ZN(
        P2_U2838) );
  OAI21_X1 U20597 ( .B1(n12443), .B2(n18598), .A(n18680), .ZN(n18515) );
  INV_X1 U20598 ( .A(n18511), .ZN(n18513) );
  OAI22_X1 U20599 ( .A1(n18513), .A2(n18529), .B1(n18512), .B2(n18627), .ZN(
        n18514) );
  AOI211_X1 U20600 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18641), .A(
        n18515), .B(n18514), .ZN(n18523) );
  NOR2_X1 U20601 ( .A1(n18517), .A2(n18516), .ZN(n18519) );
  XNOR2_X1 U20602 ( .A(n18519), .B(n18518), .ZN(n18521) );
  AOI22_X1 U20603 ( .A1(n18521), .A2(n18617), .B1(n18520), .B2(n18645), .ZN(
        n18522) );
  OAI211_X1 U20604 ( .C1(n18524), .C2(n18638), .A(n18523), .B(n18522), .ZN(
        P2_U2837) );
  NAND2_X1 U20605 ( .A1(n18525), .A2(n18606), .ZN(n18526) );
  XOR2_X1 U20606 ( .A(n18527), .B(n18526), .Z(n18538) );
  AOI22_X1 U20607 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18641), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n18639), .ZN(n18528) );
  OAI21_X1 U20608 ( .B1(n18530), .B2(n18529), .A(n18528), .ZN(n18531) );
  AOI211_X1 U20609 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18640), .A(n18532), .B(
        n18531), .ZN(n18537) );
  OAI22_X1 U20610 ( .A1(n18534), .A2(n18601), .B1(n18533), .B2(n18638), .ZN(
        n18535) );
  INV_X1 U20611 ( .A(n18535), .ZN(n18536) );
  OAI211_X1 U20612 ( .C1(n18701), .C2(n18538), .A(n18537), .B(n18536), .ZN(
        P2_U2836) );
  OAI22_X1 U20613 ( .A1(n18598), .A2(n18539), .B1(n11299), .B2(n18596), .ZN(
        n18540) );
  AOI21_X1 U20614 ( .B1(P2_REIP_REG_20__SCAN_IN), .B2(n18639), .A(n18540), 
        .ZN(n18541) );
  OAI21_X1 U20615 ( .B1(n18542), .B2(n18601), .A(n18541), .ZN(n18543) );
  AOI21_X1 U20616 ( .B1(n18544), .B2(n18642), .A(n18543), .ZN(n18549) );
  OAI211_X1 U20617 ( .C1(n18547), .C2(n18546), .A(n18617), .B(n18545), .ZN(
        n18548) );
  OAI211_X1 U20618 ( .C1(n18638), .C2(n18550), .A(n18549), .B(n18548), .ZN(
        P2_U2835) );
  INV_X1 U20619 ( .A(n18551), .ZN(n18556) );
  OAI22_X1 U20620 ( .A1(n18598), .A2(n12495), .B1(n11301), .B2(n18596), .ZN(
        n18552) );
  AOI21_X1 U20621 ( .B1(P2_REIP_REG_22__SCAN_IN), .B2(n18639), .A(n18552), 
        .ZN(n18553) );
  OAI21_X1 U20622 ( .B1(n18554), .B2(n18601), .A(n18553), .ZN(n18555) );
  AOI21_X1 U20623 ( .B1(n18556), .B2(n18642), .A(n18555), .ZN(n18561) );
  OAI211_X1 U20624 ( .C1(n18559), .C2(n18558), .A(n18617), .B(n18557), .ZN(
        n18560) );
  OAI211_X1 U20625 ( .C1(n18638), .C2(n18562), .A(n18561), .B(n18560), .ZN(
        P2_U2833) );
  AOI22_X1 U20626 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n18640), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18639), .ZN(n18572) );
  AOI22_X1 U20627 ( .A1(n18563), .A2(n18642), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18641), .ZN(n18571) );
  AOI22_X1 U20628 ( .A1(n18565), .A2(n18645), .B1(n18564), .B2(n18644), .ZN(
        n18570) );
  OAI211_X1 U20629 ( .C1(n18568), .C2(n18567), .A(n18617), .B(n18566), .ZN(
        n18569) );
  NAND4_X1 U20630 ( .A1(n18572), .A2(n18571), .A3(n18570), .A4(n18569), .ZN(
        P2_U2832) );
  AOI22_X1 U20631 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n18640), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n18639), .ZN(n18583) );
  AOI22_X1 U20632 ( .A1(n18573), .A2(n18642), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18641), .ZN(n18582) );
  OAI22_X1 U20633 ( .A1(n18575), .A2(n18601), .B1(n18574), .B2(n18638), .ZN(
        n18576) );
  INV_X1 U20634 ( .A(n18576), .ZN(n18581) );
  OAI211_X1 U20635 ( .C1(n18579), .C2(n18578), .A(n18617), .B(n18577), .ZN(
        n18580) );
  NAND4_X1 U20636 ( .A1(n18583), .A2(n18582), .A3(n18581), .A4(n18580), .ZN(
        P2_U2830) );
  AOI22_X1 U20637 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n18640), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n18639), .ZN(n18594) );
  AOI22_X1 U20638 ( .A1(n18584), .A2(n18642), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18641), .ZN(n18593) );
  OAI22_X1 U20639 ( .A1(n18586), .A2(n18601), .B1(n18585), .B2(n18638), .ZN(
        n18587) );
  INV_X1 U20640 ( .A(n18587), .ZN(n18592) );
  OAI211_X1 U20641 ( .C1(n18590), .C2(n18589), .A(n18617), .B(n18588), .ZN(
        n18591) );
  NAND4_X1 U20642 ( .A1(n18594), .A2(n18593), .A3(n18592), .A4(n18591), .ZN(
        P2_U2829) );
  INV_X1 U20643 ( .A(n18595), .ZN(n18604) );
  OAI22_X1 U20644 ( .A1(n18598), .A2(n18597), .B1(n15750), .B2(n18596), .ZN(
        n18599) );
  AOI21_X1 U20645 ( .B1(P2_REIP_REG_28__SCAN_IN), .B2(n18639), .A(n18599), 
        .ZN(n18600) );
  OAI21_X1 U20646 ( .B1(n18602), .B2(n18601), .A(n18600), .ZN(n18603) );
  AOI21_X1 U20647 ( .B1(n18604), .B2(n18642), .A(n18603), .ZN(n18610) );
  NAND2_X1 U20648 ( .A1(n18606), .A2(n18605), .ZN(n18607) );
  OAI211_X1 U20649 ( .C1(n18608), .C2(n18607), .A(n18617), .B(n18616), .ZN(
        n18609) );
  OAI211_X1 U20650 ( .C1(n18638), .C2(n18611), .A(n18610), .B(n18609), .ZN(
        P2_U2827) );
  AOI22_X1 U20651 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n18640), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18639), .ZN(n18623) );
  AOI22_X1 U20652 ( .A1(n18612), .A2(n18642), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18641), .ZN(n18622) );
  INV_X1 U20653 ( .A(n18613), .ZN(n18615) );
  AOI22_X1 U20654 ( .A1(n18615), .A2(n18645), .B1(n18614), .B2(n18644), .ZN(
        n18621) );
  OAI211_X1 U20655 ( .C1(n18619), .C2(n18618), .A(n18617), .B(n18634), .ZN(
        n18620) );
  NAND4_X1 U20656 ( .A1(n18623), .A2(n18622), .A3(n18621), .A4(n18620), .ZN(
        P2_U2826) );
  NAND2_X1 U20657 ( .A1(n18624), .A2(n18645), .ZN(n18631) );
  AOI22_X1 U20658 ( .A1(n18640), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18641), .ZN(n18625) );
  INV_X1 U20659 ( .A(n18625), .ZN(n18629) );
  NOR2_X1 U20660 ( .A1(n18627), .A2(n18626), .ZN(n18628) );
  NOR2_X1 U20661 ( .A1(n18629), .A2(n18628), .ZN(n18630) );
  NAND2_X1 U20662 ( .A1(n18631), .A2(n18630), .ZN(n18632) );
  AOI21_X1 U20663 ( .B1(n18642), .B2(n18633), .A(n18632), .ZN(n18637) );
  OAI21_X1 U20664 ( .B1(n18649), .B2(n18648), .A(n18635), .ZN(n18636) );
  OAI211_X1 U20665 ( .C1(n18638), .C2(n15803), .A(n18637), .B(n18636), .ZN(
        P2_U2825) );
  AOI22_X1 U20666 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n18640), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n18639), .ZN(n18654) );
  AOI22_X1 U20667 ( .A1(n18643), .A2(n18642), .B1(n18641), .B2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n18653) );
  AOI22_X1 U20668 ( .A1(n18646), .A2(n18645), .B1(n18644), .B2(n11040), .ZN(
        n18652) );
  INV_X1 U20669 ( .A(n18647), .ZN(n18650) );
  NAND3_X1 U20670 ( .A1(n18650), .A2(n18649), .A3(n18648), .ZN(n18651) );
  NAND4_X1 U20671 ( .A1(n18654), .A2(n18653), .A3(n18652), .A4(n18651), .ZN(
        P2_U2824) );
  NOR4_X1 U20672 ( .A1(n18657), .A2(n18656), .A3(n18655), .A4(n18696), .ZN(
        n18658) );
  NAND2_X1 U20673 ( .A1(n18661), .A2(n18658), .ZN(n18659) );
  OAI21_X1 U20674 ( .B1(n18661), .B2(n18660), .A(n18659), .ZN(P2_U3595) );
  OAI22_X1 U20675 ( .A1(n18664), .A2(n18663), .B1(n18662), .B2(n19687), .ZN(
        n18670) );
  INV_X1 U20676 ( .A(n18665), .ZN(n18668) );
  OAI22_X1 U20677 ( .A1(n18668), .A2(n18667), .B1(n12950), .B2(n18666), .ZN(
        n18669) );
  AOI211_X1 U20678 ( .C1(n18667), .C2(n18671), .A(n18670), .B(n18669), .ZN(
        n18673) );
  OAI211_X1 U20679 ( .C1(n18674), .C2(n18688), .A(n18673), .B(n18672), .ZN(
        P2_U3046) );
  INV_X1 U20680 ( .A(n18675), .ZN(n18677) );
  AOI211_X1 U20681 ( .C1(n18678), .C2(n18693), .A(n18677), .B(n18676), .ZN(
        n18682) );
  NAND2_X1 U20682 ( .A1(n19420), .A2(n12928), .ZN(n18679) );
  OAI21_X1 U20683 ( .B1(n12270), .B2(n18680), .A(n18679), .ZN(n18681) );
  NOR2_X1 U20684 ( .A1(n18682), .A2(n18681), .ZN(n18692) );
  NAND2_X1 U20685 ( .A1(n18683), .A2(n13329), .ZN(n18687) );
  NAND2_X1 U20686 ( .A1(n18685), .A2(n18684), .ZN(n18686) );
  OAI211_X1 U20687 ( .C1(n18689), .C2(n18688), .A(n18687), .B(n18686), .ZN(
        n18690) );
  INV_X1 U20688 ( .A(n18690), .ZN(n18691) );
  OAI211_X1 U20689 ( .C1(n18694), .C2(n18693), .A(n18692), .B(n18691), .ZN(
        P2_U3041) );
  NAND2_X1 U20690 ( .A1(n18704), .A2(n18695), .ZN(n18707) );
  NAND2_X1 U20691 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18716), .ZN(n18697) );
  OAI21_X1 U20692 ( .B1(n18697), .B2(n18696), .A(n18718), .ZN(n18700) );
  NAND2_X1 U20693 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n21624), .ZN(n18698) );
  AOI21_X1 U20694 ( .B1(n18717), .B2(n18707), .A(n18698), .ZN(n18699) );
  AOI21_X1 U20695 ( .B1(n18707), .B2(n18700), .A(n18699), .ZN(n18702) );
  NAND2_X1 U20696 ( .A1(n18702), .A2(n18701), .ZN(P2_U3177) );
  NOR2_X1 U20697 ( .A1(n18704), .A2(n18703), .ZN(n18710) );
  AOI21_X1 U20698 ( .B1(n18711), .B2(n18706), .A(n18705), .ZN(n18709) );
  NOR2_X1 U20699 ( .A1(n18716), .A2(n18707), .ZN(n18708) );
  OAI222_X1 U20700 ( .A1(n18718), .A2(n18712), .B1(n18711), .B2(n18710), .C1(
        n18709), .C2(n18708), .ZN(n18713) );
  INV_X1 U20701 ( .A(n18713), .ZN(n18715) );
  OAI211_X1 U20702 ( .C1(n18717), .C2(n18716), .A(n18715), .B(n18714), .ZN(
        P2_U3176) );
  NOR2_X1 U20703 ( .A1(n18719), .A2(n18718), .ZN(n18722) );
  MUX2_X1 U20704 ( .A(P2_MORE_REG_SCAN_IN), .B(n18720), .S(n18722), .Z(
        P2_U3609) );
  OAI21_X1 U20705 ( .B1(n18722), .B2(n12247), .A(n18721), .ZN(P2_U2819) );
  INV_X1 U20706 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20099) );
  AOI22_X1 U20707 ( .A1(n19080), .A2(n20099), .B1(n20705), .B2(U215), .ZN(U282) );
  OAI22_X1 U20708 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19080), .ZN(n18723) );
  INV_X1 U20709 ( .A(n18723), .ZN(U281) );
  OAI22_X1 U20710 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19080), .ZN(n18724) );
  INV_X1 U20711 ( .A(n18724), .ZN(U280) );
  OAI22_X1 U20712 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19080), .ZN(n18725) );
  INV_X1 U20713 ( .A(n18725), .ZN(U279) );
  OAI22_X1 U20714 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19080), .ZN(n18726) );
  INV_X1 U20715 ( .A(n18726), .ZN(U278) );
  OAI22_X1 U20716 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19080), .ZN(n18727) );
  INV_X1 U20717 ( .A(n18727), .ZN(U277) );
  OAI22_X1 U20718 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19080), .ZN(n18728) );
  INV_X1 U20719 ( .A(n18728), .ZN(U276) );
  OAI22_X1 U20720 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19080), .ZN(n18729) );
  INV_X1 U20721 ( .A(n18729), .ZN(U275) );
  OAI22_X1 U20722 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19080), .ZN(n18730) );
  INV_X1 U20723 ( .A(n18730), .ZN(U274) );
  OAI22_X1 U20724 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n18745), .ZN(n18731) );
  INV_X1 U20725 ( .A(n18731), .ZN(U273) );
  OAI22_X1 U20726 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n18745), .ZN(n18732) );
  INV_X1 U20727 ( .A(n18732), .ZN(U272) );
  OAI22_X1 U20728 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18745), .ZN(n18733) );
  INV_X1 U20729 ( .A(n18733), .ZN(U271) );
  OAI22_X1 U20730 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18745), .ZN(n18734) );
  INV_X1 U20731 ( .A(n18734), .ZN(U270) );
  OAI22_X1 U20732 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18745), .ZN(n18735) );
  INV_X1 U20733 ( .A(n18735), .ZN(U269) );
  OAI22_X1 U20734 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18745), .ZN(n18736) );
  INV_X1 U20735 ( .A(n18736), .ZN(U268) );
  INV_X1 U20736 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n18737) );
  INV_X1 U20737 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n20753) );
  AOI22_X1 U20738 ( .A1(n19080), .A2(n18737), .B1(n20753), .B2(U215), .ZN(U267) );
  OAI22_X1 U20739 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18745), .ZN(n18738) );
  INV_X1 U20740 ( .A(n18738), .ZN(U266) );
  OAI22_X1 U20741 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n18745), .ZN(n18739) );
  INV_X1 U20742 ( .A(n18739), .ZN(U265) );
  OAI22_X1 U20743 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19080), .ZN(n18740) );
  INV_X1 U20744 ( .A(n18740), .ZN(U264) );
  OAI22_X1 U20745 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n18745), .ZN(n18741) );
  INV_X1 U20746 ( .A(n18741), .ZN(U263) );
  INV_X1 U20747 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n18743) );
  INV_X1 U20748 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n18742) );
  AOI22_X1 U20749 ( .A1(n19080), .A2(n18743), .B1(n18742), .B2(U215), .ZN(U262) );
  OAI22_X1 U20750 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n19080), .ZN(n18744) );
  INV_X1 U20751 ( .A(n18744), .ZN(U261) );
  OAI22_X1 U20752 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n18745), .ZN(n18746) );
  INV_X1 U20753 ( .A(n18746), .ZN(U260) );
  OAI22_X1 U20754 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19080), .ZN(n18747) );
  INV_X1 U20755 ( .A(n18747), .ZN(U259) );
  OAI22_X1 U20756 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19080), .ZN(n18748) );
  INV_X1 U20757 ( .A(n18748), .ZN(U258) );
  NAND3_X1 U20758 ( .A1(n18796), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18759) );
  NOR2_X2 U20759 ( .A1(n18802), .A2(n18759), .ZN(n19176) );
  INV_X1 U20760 ( .A(n19176), .ZN(n19037) );
  NAND2_X1 U20761 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19082), .ZN(n18794) );
  INV_X1 U20762 ( .A(n18759), .ZN(n18760) );
  NAND2_X1 U20763 ( .A1(n18802), .A2(n18760), .ZN(n19096) );
  INV_X1 U20764 ( .A(n19096), .ZN(n19102) );
  NOR2_X2 U20765 ( .A1(n20705), .A2(n19083), .ZN(n18829) );
  NOR2_X1 U20766 ( .A1(n21222), .A2(n18773), .ZN(n18824) );
  INV_X1 U20767 ( .A(n18824), .ZN(n18749) );
  NOR2_X1 U20768 ( .A1(n21239), .A2(n18749), .ZN(n19085) );
  INV_X1 U20769 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20741) );
  NOR2_X2 U20770 ( .A1(n20741), .A2(n18956), .ZN(n18828) );
  AOI22_X1 U20771 ( .A1(n19102), .A2(n18829), .B1(n19085), .B2(n18828), .ZN(
        n18754) );
  NOR2_X1 U20772 ( .A1(n18750), .A2(n18956), .ZN(n18779) );
  AOI22_X1 U20773 ( .A1(n19082), .A2(n18760), .B1(n18824), .B2(n18779), .ZN(
        n19088) );
  NAND2_X1 U20774 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18824), .ZN(
        n19164) );
  INV_X1 U20775 ( .A(n19164), .ZN(n19167) );
  NAND2_X1 U20776 ( .A1(n18752), .A2(n18751), .ZN(n19086) );
  NOR2_X1 U20777 ( .A1(n20768), .A2(n19086), .ZN(n18791) );
  AOI22_X1 U20778 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19088), .B1(
        n19167), .B2(n18791), .ZN(n18753) );
  OAI211_X1 U20779 ( .C1(n19037), .C2(n18794), .A(n18754), .B(n18753), .ZN(
        P3_U2995) );
  NOR2_X1 U20780 ( .A1(n18796), .A2(n18778), .ZN(n18767) );
  NAND2_X1 U20781 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18767), .ZN(
        n19045) );
  INV_X1 U20782 ( .A(n19045), .ZN(n19109) );
  NAND2_X1 U20783 ( .A1(n18802), .A2(n18824), .ZN(n19183) );
  NAND2_X1 U20784 ( .A1(n19037), .A2(n19183), .ZN(n18832) );
  INV_X1 U20785 ( .A(n18832), .ZN(n18755) );
  NOR2_X1 U20786 ( .A1(n21239), .A2(n18755), .ZN(n19091) );
  AOI22_X1 U20787 ( .A1(n18829), .A2(n19109), .B1(n18828), .B2(n19091), .ZN(
        n18758) );
  INV_X1 U20788 ( .A(n18956), .ZN(n19084) );
  NAND2_X1 U20789 ( .A1(n19096), .A2(n19045), .ZN(n18764) );
  INV_X1 U20790 ( .A(n18764), .ZN(n18763) );
  OAI21_X1 U20791 ( .B1(n18763), .B2(n18798), .A(n18755), .ZN(n18756) );
  OAI211_X1 U20792 ( .C1(n19092), .C2(n21246), .A(n19084), .B(n18756), .ZN(
        n19093) );
  AOI22_X1 U20793 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19093), .B1(
        n18791), .B2(n19092), .ZN(n18757) );
  OAI211_X1 U20794 ( .C1(n18794), .C2(n19096), .A(n18758), .B(n18757), .ZN(
        P3_U2987) );
  INV_X1 U20795 ( .A(n18794), .ZN(n18833) );
  NOR2_X1 U20796 ( .A1(n21239), .A2(n18759), .ZN(n19097) );
  AOI22_X1 U20797 ( .A1(n18833), .A2(n19109), .B1(n18828), .B2(n19097), .ZN(
        n18762) );
  AOI22_X1 U20798 ( .A1(n19082), .A2(n18767), .B1(n18760), .B2(n18779), .ZN(
        n19098) );
  NAND2_X1 U20799 ( .A1(n18802), .A2(n18767), .ZN(n19106) );
  AOI22_X1 U20800 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19098), .B1(
        n18829), .B2(n19114), .ZN(n18761) );
  OAI211_X1 U20801 ( .C1(n19037), .C2(n18836), .A(n18762), .B(n18761), .ZN(
        P3_U2979) );
  NOR2_X1 U20802 ( .A1(n18802), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18785) );
  NAND2_X1 U20803 ( .A1(n18780), .A2(n18785), .ZN(n19008) );
  NOR2_X1 U20804 ( .A1(n21239), .A2(n18763), .ZN(n19101) );
  AOI22_X1 U20805 ( .A1(n18829), .A2(n19120), .B1(n18828), .B2(n19101), .ZN(
        n18766) );
  NOR2_X1 U20806 ( .A1(n19114), .A2(n19120), .ZN(n18772) );
  INV_X1 U20807 ( .A(n18772), .ZN(n18775) );
  AOI21_X1 U20808 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18956), .ZN(n18831) );
  AOI22_X1 U20809 ( .A1(n19082), .A2(n18775), .B1(n18831), .B2(n18764), .ZN(
        n19103) );
  AOI22_X1 U20810 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19103), .B1(
        n18833), .B2(n19114), .ZN(n18765) );
  OAI211_X1 U20811 ( .C1(n18836), .C2(n19096), .A(n18766), .B(n18765), .ZN(
        P3_U2971) );
  INV_X1 U20812 ( .A(n18767), .ZN(n18768) );
  NOR2_X1 U20813 ( .A1(n21239), .A2(n18768), .ZN(n19107) );
  AOI22_X1 U20814 ( .A1(n18833), .A2(n19120), .B1(n18828), .B2(n19107), .ZN(
        n18771) );
  AOI21_X1 U20815 ( .B1(n18796), .B2(n18798), .A(n18956), .ZN(n18814) );
  NAND3_X1 U20816 ( .A1(n18780), .A2(n18814), .A3(n18769), .ZN(n19108) );
  NOR2_X1 U20817 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21215) );
  NAND2_X1 U20818 ( .A1(n21215), .A2(n18780), .ZN(n19112) );
  AOI22_X1 U20819 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19108), .B1(
        n18829), .B2(n19126), .ZN(n18770) );
  OAI211_X1 U20820 ( .C1(n18836), .C2(n19045), .A(n18771), .B(n18770), .ZN(
        P3_U2963) );
  NOR2_X1 U20821 ( .A1(n21239), .A2(n18772), .ZN(n19113) );
  AOI22_X1 U20822 ( .A1(n18833), .A2(n19126), .B1(n18828), .B2(n19113), .ZN(
        n18777) );
  NOR2_X1 U20823 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18773), .ZN(
        n18781) );
  INV_X1 U20824 ( .A(n18781), .ZN(n18790) );
  NOR2_X2 U20825 ( .A1(n18802), .A2(n18790), .ZN(n19132) );
  NOR2_X1 U20826 ( .A1(n19126), .A2(n19132), .ZN(n18784) );
  INV_X1 U20827 ( .A(n18784), .ZN(n18786) );
  OAI221_X1 U20828 ( .B1(n18775), .B2(n18774), .C1(n18775), .C2(n18786), .A(
        n18831), .ZN(n19115) );
  AOI22_X1 U20829 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19115), .B1(
        n18829), .B2(n19132), .ZN(n18776) );
  OAI211_X1 U20830 ( .C1(n18836), .C2(n19106), .A(n18777), .B(n18776), .ZN(
        P3_U2955) );
  AOI22_X1 U20831 ( .A1(n18833), .A2(n19132), .B1(n18828), .B2(n19119), .ZN(
        n18783) );
  AND2_X1 U20832 ( .A1(n18796), .A2(n18779), .ZN(n18823) );
  AOI22_X1 U20833 ( .A1(n19082), .A2(n18781), .B1(n18780), .B2(n18823), .ZN(
        n19121) );
  NAND2_X1 U20834 ( .A1(n18802), .A2(n18781), .ZN(n19124) );
  INV_X1 U20835 ( .A(n19124), .ZN(n19137) );
  AOI22_X1 U20836 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19121), .B1(
        n18829), .B2(n19137), .ZN(n18782) );
  OAI211_X1 U20837 ( .C1(n18836), .C2(n19008), .A(n18783), .B(n18782), .ZN(
        P3_U2947) );
  NOR2_X1 U20838 ( .A1(n21239), .A2(n18784), .ZN(n19125) );
  AOI22_X1 U20839 ( .A1(n18833), .A2(n19137), .B1(n18828), .B2(n19125), .ZN(
        n18789) );
  INV_X1 U20840 ( .A(n18785), .ZN(n18808) );
  NOR2_X2 U20841 ( .A1(n18808), .A2(n18803), .ZN(n19143) );
  NOR2_X1 U20842 ( .A1(n19137), .A2(n19143), .ZN(n18797) );
  INV_X1 U20843 ( .A(n18797), .ZN(n18787) );
  AOI22_X1 U20844 ( .A1(n19082), .A2(n18787), .B1(n18831), .B2(n18786), .ZN(
        n19127) );
  AOI22_X1 U20845 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19127), .B1(
        n18829), .B2(n19143), .ZN(n18788) );
  OAI211_X1 U20846 ( .C1(n18836), .C2(n19112), .A(n18789), .B(n18788), .ZN(
        P3_U2939) );
  OAI211_X1 U20847 ( .C1(n19132), .C2(n21246), .A(n18814), .B(n18804), .ZN(
        n19133) );
  NOR2_X1 U20848 ( .A1(n21239), .A2(n18790), .ZN(n19131) );
  AOI22_X1 U20849 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19133), .B1(
        n18828), .B2(n19131), .ZN(n18793) );
  NAND2_X1 U20850 ( .A1(n21215), .A2(n18804), .ZN(n19141) );
  AOI22_X1 U20851 ( .A1(n18791), .A2(n19132), .B1(n18829), .B2(n19148), .ZN(
        n18792) );
  OAI211_X1 U20852 ( .C1(n18794), .C2(n19130), .A(n18793), .B(n18792), .ZN(
        P3_U2931) );
  NAND2_X1 U20853 ( .A1(n18795), .A2(n21222), .ZN(n18821) );
  NOR2_X1 U20854 ( .A1(n18796), .A2(n18821), .ZN(n18812) );
  NAND2_X1 U20855 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18812), .ZN(
        n19062) );
  INV_X1 U20856 ( .A(n19062), .ZN(n19155) );
  NOR2_X1 U20857 ( .A1(n21239), .A2(n18797), .ZN(n19136) );
  AOI22_X1 U20858 ( .A1(n18829), .A2(n19155), .B1(n18828), .B2(n19136), .ZN(
        n18801) );
  NAND2_X1 U20859 ( .A1(n19141), .A2(n19062), .ZN(n18809) );
  INV_X1 U20860 ( .A(n18809), .ZN(n18807) );
  OAI21_X1 U20861 ( .B1(n18807), .B2(n18798), .A(n18797), .ZN(n18799) );
  OAI211_X1 U20862 ( .C1(n19137), .C2(n21246), .A(n19084), .B(n18799), .ZN(
        n19138) );
  AOI22_X1 U20863 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19138), .B1(
        n18833), .B2(n19148), .ZN(n18800) );
  OAI211_X1 U20864 ( .C1(n18836), .C2(n19124), .A(n18801), .B(n18800), .ZN(
        P3_U2923) );
  NAND2_X1 U20865 ( .A1(n18802), .A2(n18812), .ZN(n19152) );
  AOI22_X1 U20866 ( .A1(n18829), .A2(n19160), .B1(n18828), .B2(n19142), .ZN(
        n18806) );
  AOI22_X1 U20867 ( .A1(n19082), .A2(n18812), .B1(n18823), .B2(n18804), .ZN(
        n19144) );
  AOI22_X1 U20868 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19144), .B1(
        n18833), .B2(n19155), .ZN(n18805) );
  OAI211_X1 U20869 ( .C1(n18836), .C2(n19130), .A(n18806), .B(n18805), .ZN(
        P3_U2915) );
  NOR2_X1 U20870 ( .A1(n21239), .A2(n18807), .ZN(n19147) );
  AOI22_X1 U20871 ( .A1(n18833), .A2(n19160), .B1(n18828), .B2(n19147), .ZN(
        n18811) );
  NOR2_X1 U20872 ( .A1(n19160), .A2(n19168), .ZN(n18817) );
  INV_X1 U20873 ( .A(n18817), .ZN(n18818) );
  AOI22_X1 U20874 ( .A1(n19082), .A2(n18818), .B1(n18831), .B2(n18809), .ZN(
        n19149) );
  AOI22_X1 U20875 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19149), .B1(
        n18829), .B2(n19168), .ZN(n18810) );
  OAI211_X1 U20876 ( .C1(n18836), .C2(n19141), .A(n18811), .B(n18810), .ZN(
        P3_U2907) );
  INV_X1 U20877 ( .A(n18812), .ZN(n18813) );
  NOR2_X1 U20878 ( .A1(n21239), .A2(n18813), .ZN(n19153) );
  AOI22_X1 U20879 ( .A1(n18833), .A2(n19168), .B1(n18828), .B2(n19153), .ZN(
        n18816) );
  INV_X1 U20880 ( .A(n18821), .ZN(n18822) );
  OAI211_X1 U20881 ( .C1(n19155), .C2(n21246), .A(n18822), .B(n18814), .ZN(
        n19154) );
  NAND2_X1 U20882 ( .A1(n21215), .A2(n18822), .ZN(n19067) );
  AOI22_X1 U20883 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19154), .B1(
        n18829), .B2(n19178), .ZN(n18815) );
  OAI211_X1 U20884 ( .C1(n18836), .C2(n19062), .A(n18816), .B(n18815), .ZN(
        P3_U2899) );
  NOR2_X1 U20885 ( .A1(n21239), .A2(n18817), .ZN(n19159) );
  AOI22_X1 U20886 ( .A1(n18833), .A2(n19178), .B1(n18828), .B2(n19159), .ZN(
        n18820) );
  NOR2_X1 U20887 ( .A1(n19167), .A2(n19178), .ZN(n18827) );
  INV_X1 U20888 ( .A(n18827), .ZN(n18830) );
  AOI22_X1 U20889 ( .A1(n19082), .A2(n18830), .B1(n18831), .B2(n18818), .ZN(
        n19161) );
  AOI22_X1 U20890 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19161), .B1(
        n19167), .B2(n18829), .ZN(n18819) );
  OAI211_X1 U20891 ( .C1(n18836), .C2(n19152), .A(n18820), .B(n18819), .ZN(
        P3_U2891) );
  INV_X1 U20892 ( .A(n19168), .ZN(n19158) );
  AOI22_X1 U20893 ( .A1(n18833), .A2(n19167), .B1(n18828), .B2(n19165), .ZN(
        n18826) );
  AOI22_X1 U20894 ( .A1(n19082), .A2(n18824), .B1(n18823), .B2(n18822), .ZN(
        n19169) );
  AOI22_X1 U20895 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19169), .B1(
        n18829), .B2(n19092), .ZN(n18825) );
  OAI211_X1 U20896 ( .C1(n18836), .C2(n19158), .A(n18826), .B(n18825), .ZN(
        P3_U2883) );
  NOR2_X1 U20897 ( .A1(n21239), .A2(n18827), .ZN(n19174) );
  AOI22_X1 U20898 ( .A1(n19176), .A2(n18829), .B1(n18828), .B2(n19174), .ZN(
        n18835) );
  AOI22_X1 U20899 ( .A1(n19082), .A2(n18832), .B1(n18831), .B2(n18830), .ZN(
        n19179) );
  AOI22_X1 U20900 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19179), .B1(
        n18833), .B2(n19092), .ZN(n18834) );
  OAI211_X1 U20901 ( .C1(n18836), .C2(n19067), .A(n18835), .B(n18834), .ZN(
        P3_U2875) );
  OAI22_X1 U20902 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19080), .ZN(n18837) );
  INV_X1 U20903 ( .A(n18837), .ZN(U257) );
  INV_X1 U20904 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n20665) );
  NOR2_X1 U20905 ( .A1(n20665), .A2(n19083), .ZN(n18866) );
  INV_X1 U20906 ( .A(n18866), .ZN(n18875) );
  NAND2_X1 U20907 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19082), .ZN(n18869) );
  INV_X1 U20908 ( .A(n18869), .ZN(n18871) );
  INV_X1 U20909 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20674) );
  NOR2_X2 U20910 ( .A1(n20674), .A2(n18956), .ZN(n18870) );
  AOI22_X1 U20911 ( .A1(n19102), .A2(n18871), .B1(n19085), .B2(n18870), .ZN(
        n18839) );
  NOR2_X2 U20912 ( .A1(n20652), .A2(n19086), .ZN(n18872) );
  AOI22_X1 U20913 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19088), .B1(
        n19167), .B2(n18872), .ZN(n18838) );
  OAI211_X1 U20914 ( .C1(n19037), .C2(n18875), .A(n18839), .B(n18838), .ZN(
        P3_U2994) );
  AOI22_X1 U20915 ( .A1(n19109), .A2(n18871), .B1(n19091), .B2(n18870), .ZN(
        n18841) );
  AOI22_X1 U20916 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19093), .B1(
        n19092), .B2(n18872), .ZN(n18840) );
  OAI211_X1 U20917 ( .C1(n19096), .C2(n18875), .A(n18841), .B(n18840), .ZN(
        P3_U2986) );
  AOI22_X1 U20918 ( .A1(n19114), .A2(n18871), .B1(n19097), .B2(n18870), .ZN(
        n18843) );
  AOI22_X1 U20919 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19098), .B1(
        n19176), .B2(n18872), .ZN(n18842) );
  OAI211_X1 U20920 ( .C1(n19045), .C2(n18875), .A(n18843), .B(n18842), .ZN(
        P3_U2978) );
  AOI22_X1 U20921 ( .A1(n19114), .A2(n18866), .B1(n19101), .B2(n18870), .ZN(
        n18845) );
  AOI22_X1 U20922 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19103), .B1(
        n19102), .B2(n18872), .ZN(n18844) );
  OAI211_X1 U20923 ( .C1(n19008), .C2(n18869), .A(n18845), .B(n18844), .ZN(
        P3_U2970) );
  AOI22_X1 U20924 ( .A1(n19120), .A2(n18866), .B1(n19107), .B2(n18870), .ZN(
        n18847) );
  AOI22_X1 U20925 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19108), .B1(
        n19109), .B2(n18872), .ZN(n18846) );
  OAI211_X1 U20926 ( .C1(n19112), .C2(n18869), .A(n18847), .B(n18846), .ZN(
        P3_U2962) );
  AOI22_X1 U20927 ( .A1(n19132), .A2(n18871), .B1(n19113), .B2(n18870), .ZN(
        n18849) );
  AOI22_X1 U20928 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19115), .B1(
        n19114), .B2(n18872), .ZN(n18848) );
  OAI211_X1 U20929 ( .C1(n19112), .C2(n18875), .A(n18849), .B(n18848), .ZN(
        P3_U2954) );
  INV_X1 U20930 ( .A(n19132), .ZN(n19118) );
  AOI22_X1 U20931 ( .A1(n19137), .A2(n18871), .B1(n19119), .B2(n18870), .ZN(
        n18851) );
  AOI22_X1 U20932 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19121), .B1(
        n19120), .B2(n18872), .ZN(n18850) );
  OAI211_X1 U20933 ( .C1(n19118), .C2(n18875), .A(n18851), .B(n18850), .ZN(
        P3_U2946) );
  AOI22_X1 U20934 ( .A1(n19143), .A2(n18871), .B1(n19125), .B2(n18870), .ZN(
        n18853) );
  AOI22_X1 U20935 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19127), .B1(
        n19126), .B2(n18872), .ZN(n18852) );
  OAI211_X1 U20936 ( .C1(n19124), .C2(n18875), .A(n18853), .B(n18852), .ZN(
        P3_U2938) );
  AOI22_X1 U20937 ( .A1(n19143), .A2(n18866), .B1(n19131), .B2(n18870), .ZN(
        n18855) );
  AOI22_X1 U20938 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19133), .B1(
        n19132), .B2(n18872), .ZN(n18854) );
  OAI211_X1 U20939 ( .C1(n19141), .C2(n18869), .A(n18855), .B(n18854), .ZN(
        P3_U2930) );
  AOI22_X1 U20940 ( .A1(n19148), .A2(n18866), .B1(n19136), .B2(n18870), .ZN(
        n18857) );
  AOI22_X1 U20941 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19138), .B1(
        n19137), .B2(n18872), .ZN(n18856) );
  OAI211_X1 U20942 ( .C1(n19062), .C2(n18869), .A(n18857), .B(n18856), .ZN(
        P3_U2922) );
  AOI22_X1 U20943 ( .A1(n19142), .A2(n18870), .B1(n19160), .B2(n18871), .ZN(
        n18859) );
  AOI22_X1 U20944 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19144), .B1(
        n19143), .B2(n18872), .ZN(n18858) );
  OAI211_X1 U20945 ( .C1(n19062), .C2(n18875), .A(n18859), .B(n18858), .ZN(
        P3_U2914) );
  AOI22_X1 U20946 ( .A1(n19168), .A2(n18871), .B1(n19147), .B2(n18870), .ZN(
        n18861) );
  AOI22_X1 U20947 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19149), .B1(
        n19148), .B2(n18872), .ZN(n18860) );
  OAI211_X1 U20948 ( .C1(n19152), .C2(n18875), .A(n18861), .B(n18860), .ZN(
        P3_U2906) );
  AOI22_X1 U20949 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n18870), .ZN(n18863) );
  AOI22_X1 U20950 ( .A1(n19155), .A2(n18872), .B1(n19168), .B2(n18866), .ZN(
        n18862) );
  OAI211_X1 U20951 ( .C1(n19067), .C2(n18869), .A(n18863), .B(n18862), .ZN(
        P3_U2898) );
  AOI22_X1 U20952 ( .A1(n19178), .A2(n18866), .B1(n19159), .B2(n18870), .ZN(
        n18865) );
  AOI22_X1 U20953 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19161), .B1(
        n19160), .B2(n18872), .ZN(n18864) );
  OAI211_X1 U20954 ( .C1(n19164), .C2(n18869), .A(n18865), .B(n18864), .ZN(
        P3_U2890) );
  AOI22_X1 U20955 ( .A1(n19167), .A2(n18866), .B1(n19165), .B2(n18870), .ZN(
        n18868) );
  AOI22_X1 U20956 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19169), .B1(
        n19168), .B2(n18872), .ZN(n18867) );
  OAI211_X1 U20957 ( .C1(n19183), .C2(n18869), .A(n18868), .B(n18867), .ZN(
        P3_U2882) );
  AOI22_X1 U20958 ( .A1(n19176), .A2(n18871), .B1(n19174), .B2(n18870), .ZN(
        n18874) );
  AOI22_X1 U20959 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19179), .B1(
        n19178), .B2(n18872), .ZN(n18873) );
  OAI211_X1 U20960 ( .C1(n19183), .C2(n18875), .A(n18874), .B(n18873), .ZN(
        P3_U2874) );
  OAI22_X1 U20961 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19080), .ZN(n18876) );
  INV_X1 U20962 ( .A(n18876), .ZN(U256) );
  INV_X1 U20963 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n20660) );
  NOR2_X1 U20964 ( .A1(n20660), .A2(n19083), .ZN(n18910) );
  NAND2_X1 U20965 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19082), .ZN(n18914) );
  INV_X1 U20966 ( .A(n18914), .ZN(n18905) );
  INV_X1 U20967 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n20636) );
  NOR2_X2 U20968 ( .A1(n20636), .A2(n18956), .ZN(n18909) );
  AOI22_X1 U20969 ( .A1(n19102), .A2(n18905), .B1(n19085), .B2(n18909), .ZN(
        n18878) );
  NOR2_X2 U20970 ( .A1(n20653), .A2(n19086), .ZN(n18911) );
  AOI22_X1 U20971 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19088), .B1(
        n19167), .B2(n18911), .ZN(n18877) );
  OAI211_X1 U20972 ( .C1(n19037), .C2(n18908), .A(n18878), .B(n18877), .ZN(
        P3_U2993) );
  AOI22_X1 U20973 ( .A1(n19109), .A2(n18905), .B1(n19091), .B2(n18909), .ZN(
        n18880) );
  AOI22_X1 U20974 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19093), .B1(
        n19092), .B2(n18911), .ZN(n18879) );
  OAI211_X1 U20975 ( .C1(n19096), .C2(n18908), .A(n18880), .B(n18879), .ZN(
        P3_U2985) );
  AOI22_X1 U20976 ( .A1(n19109), .A2(n18910), .B1(n19097), .B2(n18909), .ZN(
        n18882) );
  AOI22_X1 U20977 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19098), .B1(
        n19176), .B2(n18911), .ZN(n18881) );
  OAI211_X1 U20978 ( .C1(n19106), .C2(n18914), .A(n18882), .B(n18881), .ZN(
        P3_U2977) );
  AOI22_X1 U20979 ( .A1(n19120), .A2(n18905), .B1(n19101), .B2(n18909), .ZN(
        n18884) );
  AOI22_X1 U20980 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19103), .B1(
        n19102), .B2(n18911), .ZN(n18883) );
  OAI211_X1 U20981 ( .C1(n19106), .C2(n18908), .A(n18884), .B(n18883), .ZN(
        P3_U2969) );
  AOI22_X1 U20982 ( .A1(n19126), .A2(n18905), .B1(n19107), .B2(n18909), .ZN(
        n18886) );
  AOI22_X1 U20983 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19108), .B1(
        n19109), .B2(n18911), .ZN(n18885) );
  OAI211_X1 U20984 ( .C1(n19008), .C2(n18908), .A(n18886), .B(n18885), .ZN(
        P3_U2961) );
  AOI22_X1 U20985 ( .A1(n19126), .A2(n18910), .B1(n19113), .B2(n18909), .ZN(
        n18888) );
  AOI22_X1 U20986 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19115), .B1(
        n19114), .B2(n18911), .ZN(n18887) );
  OAI211_X1 U20987 ( .C1(n19118), .C2(n18914), .A(n18888), .B(n18887), .ZN(
        P3_U2953) );
  AOI22_X1 U20988 ( .A1(n19137), .A2(n18905), .B1(n19119), .B2(n18909), .ZN(
        n18890) );
  AOI22_X1 U20989 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19121), .B1(
        n19120), .B2(n18911), .ZN(n18889) );
  OAI211_X1 U20990 ( .C1(n19118), .C2(n18908), .A(n18890), .B(n18889), .ZN(
        P3_U2945) );
  AOI22_X1 U20991 ( .A1(n19137), .A2(n18910), .B1(n19125), .B2(n18909), .ZN(
        n18892) );
  AOI22_X1 U20992 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19127), .B1(
        n19126), .B2(n18911), .ZN(n18891) );
  OAI211_X1 U20993 ( .C1(n19130), .C2(n18914), .A(n18892), .B(n18891), .ZN(
        P3_U2937) );
  AOI22_X1 U20994 ( .A1(n19148), .A2(n18905), .B1(n19131), .B2(n18909), .ZN(
        n18894) );
  AOI22_X1 U20995 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19133), .B1(
        n19132), .B2(n18911), .ZN(n18893) );
  OAI211_X1 U20996 ( .C1(n19130), .C2(n18908), .A(n18894), .B(n18893), .ZN(
        P3_U2929) );
  AOI22_X1 U20997 ( .A1(n19155), .A2(n18905), .B1(n19136), .B2(n18909), .ZN(
        n18896) );
  AOI22_X1 U20998 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19138), .B1(
        n19137), .B2(n18911), .ZN(n18895) );
  OAI211_X1 U20999 ( .C1(n19141), .C2(n18908), .A(n18896), .B(n18895), .ZN(
        P3_U2921) );
  AOI22_X1 U21000 ( .A1(n19155), .A2(n18910), .B1(n19142), .B2(n18909), .ZN(
        n18898) );
  AOI22_X1 U21001 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19144), .B1(
        n19143), .B2(n18911), .ZN(n18897) );
  OAI211_X1 U21002 ( .C1(n19152), .C2(n18914), .A(n18898), .B(n18897), .ZN(
        P3_U2913) );
  AOI22_X1 U21003 ( .A1(n19160), .A2(n18910), .B1(n19147), .B2(n18909), .ZN(
        n18900) );
  AOI22_X1 U21004 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19149), .B1(
        n19148), .B2(n18911), .ZN(n18899) );
  OAI211_X1 U21005 ( .C1(n19158), .C2(n18914), .A(n18900), .B(n18899), .ZN(
        P3_U2905) );
  AOI22_X1 U21006 ( .A1(n19178), .A2(n18905), .B1(n19153), .B2(n18909), .ZN(
        n18902) );
  AOI22_X1 U21007 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19154), .B1(
        n19155), .B2(n18911), .ZN(n18901) );
  OAI211_X1 U21008 ( .C1(n19158), .C2(n18908), .A(n18902), .B(n18901), .ZN(
        P3_U2897) );
  AOI22_X1 U21009 ( .A1(n19178), .A2(n18910), .B1(n19159), .B2(n18909), .ZN(
        n18904) );
  AOI22_X1 U21010 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19161), .B1(
        n19160), .B2(n18911), .ZN(n18903) );
  OAI211_X1 U21011 ( .C1(n19164), .C2(n18914), .A(n18904), .B(n18903), .ZN(
        P3_U2889) );
  AOI22_X1 U21012 ( .A1(n19092), .A2(n18905), .B1(n19165), .B2(n18909), .ZN(
        n18907) );
  AOI22_X1 U21013 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19169), .B1(
        n19168), .B2(n18911), .ZN(n18906) );
  OAI211_X1 U21014 ( .C1(n19164), .C2(n18908), .A(n18907), .B(n18906), .ZN(
        P3_U2881) );
  AOI22_X1 U21015 ( .A1(n19092), .A2(n18910), .B1(n19174), .B2(n18909), .ZN(
        n18913) );
  AOI22_X1 U21016 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19179), .B1(
        n19178), .B2(n18911), .ZN(n18912) );
  OAI211_X1 U21017 ( .C1(n19037), .C2(n18914), .A(n18913), .B(n18912), .ZN(
        P3_U2873) );
  OAI22_X1 U21018 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19080), .ZN(n18915) );
  INV_X1 U21019 ( .A(n18915), .ZN(U255) );
  NAND2_X1 U21020 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19082), .ZN(n18954) );
  NAND2_X1 U21021 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n19082), .ZN(n18942) );
  INV_X1 U21022 ( .A(n18942), .ZN(n18950) );
  INV_X1 U21023 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n20641) );
  NOR2_X2 U21024 ( .A1(n20641), .A2(n18956), .ZN(n18949) );
  AOI22_X1 U21025 ( .A1(n19176), .A2(n18950), .B1(n19085), .B2(n18949), .ZN(
        n18918) );
  NOR2_X2 U21026 ( .A1(n18916), .A2(n19086), .ZN(n18951) );
  AOI22_X1 U21027 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19088), .B1(
        n19167), .B2(n18951), .ZN(n18917) );
  OAI211_X1 U21028 ( .C1(n19096), .C2(n18954), .A(n18918), .B(n18917), .ZN(
        P3_U2992) );
  INV_X1 U21029 ( .A(n18954), .ZN(n18939) );
  AOI22_X1 U21030 ( .A1(n19109), .A2(n18939), .B1(n19091), .B2(n18949), .ZN(
        n18920) );
  AOI22_X1 U21031 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19093), .B1(
        n19092), .B2(n18951), .ZN(n18919) );
  OAI211_X1 U21032 ( .C1(n19096), .C2(n18942), .A(n18920), .B(n18919), .ZN(
        P3_U2984) );
  AOI22_X1 U21033 ( .A1(n19114), .A2(n18939), .B1(n19097), .B2(n18949), .ZN(
        n18922) );
  AOI22_X1 U21034 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19098), .B1(
        n19176), .B2(n18951), .ZN(n18921) );
  OAI211_X1 U21035 ( .C1(n19045), .C2(n18942), .A(n18922), .B(n18921), .ZN(
        P3_U2976) );
  AOI22_X1 U21036 ( .A1(n19114), .A2(n18950), .B1(n19101), .B2(n18949), .ZN(
        n18924) );
  AOI22_X1 U21037 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19103), .B1(
        n19102), .B2(n18951), .ZN(n18923) );
  OAI211_X1 U21038 ( .C1(n19008), .C2(n18954), .A(n18924), .B(n18923), .ZN(
        P3_U2968) );
  AOI22_X1 U21039 ( .A1(n19126), .A2(n18939), .B1(n19107), .B2(n18949), .ZN(
        n18926) );
  AOI22_X1 U21040 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19108), .B1(
        n19109), .B2(n18951), .ZN(n18925) );
  OAI211_X1 U21041 ( .C1(n19008), .C2(n18942), .A(n18926), .B(n18925), .ZN(
        P3_U2960) );
  AOI22_X1 U21042 ( .A1(n19132), .A2(n18939), .B1(n19113), .B2(n18949), .ZN(
        n18928) );
  AOI22_X1 U21043 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19115), .B1(
        n19114), .B2(n18951), .ZN(n18927) );
  OAI211_X1 U21044 ( .C1(n19112), .C2(n18942), .A(n18928), .B(n18927), .ZN(
        P3_U2952) );
  AOI22_X1 U21045 ( .A1(n19137), .A2(n18939), .B1(n19119), .B2(n18949), .ZN(
        n18930) );
  AOI22_X1 U21046 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19121), .B1(
        n19120), .B2(n18951), .ZN(n18929) );
  OAI211_X1 U21047 ( .C1(n19118), .C2(n18942), .A(n18930), .B(n18929), .ZN(
        P3_U2944) );
  AOI22_X1 U21048 ( .A1(n19137), .A2(n18950), .B1(n19125), .B2(n18949), .ZN(
        n18932) );
  AOI22_X1 U21049 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19127), .B1(
        n19126), .B2(n18951), .ZN(n18931) );
  OAI211_X1 U21050 ( .C1(n19130), .C2(n18954), .A(n18932), .B(n18931), .ZN(
        P3_U2936) );
  AOI22_X1 U21051 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19133), .B1(
        n19131), .B2(n18949), .ZN(n18934) );
  AOI22_X1 U21052 ( .A1(n19132), .A2(n18951), .B1(n19143), .B2(n18950), .ZN(
        n18933) );
  OAI211_X1 U21053 ( .C1(n19141), .C2(n18954), .A(n18934), .B(n18933), .ZN(
        P3_U2928) );
  AOI22_X1 U21054 ( .A1(n19155), .A2(n18939), .B1(n19136), .B2(n18949), .ZN(
        n18936) );
  AOI22_X1 U21055 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19138), .B1(
        n19137), .B2(n18951), .ZN(n18935) );
  OAI211_X1 U21056 ( .C1(n19141), .C2(n18942), .A(n18936), .B(n18935), .ZN(
        P3_U2920) );
  AOI22_X1 U21057 ( .A1(n19155), .A2(n18950), .B1(n19142), .B2(n18949), .ZN(
        n18938) );
  AOI22_X1 U21058 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19144), .B1(
        n19143), .B2(n18951), .ZN(n18937) );
  OAI211_X1 U21059 ( .C1(n19152), .C2(n18954), .A(n18938), .B(n18937), .ZN(
        P3_U2912) );
  AOI22_X1 U21060 ( .A1(n19168), .A2(n18939), .B1(n19147), .B2(n18949), .ZN(
        n18941) );
  AOI22_X1 U21061 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19149), .B1(
        n19148), .B2(n18951), .ZN(n18940) );
  OAI211_X1 U21062 ( .C1(n19152), .C2(n18942), .A(n18941), .B(n18940), .ZN(
        P3_U2904) );
  AOI22_X1 U21063 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n18949), .ZN(n18944) );
  AOI22_X1 U21064 ( .A1(n19155), .A2(n18951), .B1(n19168), .B2(n18950), .ZN(
        n18943) );
  OAI211_X1 U21065 ( .C1(n19067), .C2(n18954), .A(n18944), .B(n18943), .ZN(
        P3_U2896) );
  AOI22_X1 U21066 ( .A1(n19178), .A2(n18950), .B1(n19159), .B2(n18949), .ZN(
        n18946) );
  AOI22_X1 U21067 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19161), .B1(
        n19160), .B2(n18951), .ZN(n18945) );
  OAI211_X1 U21068 ( .C1(n19164), .C2(n18954), .A(n18946), .B(n18945), .ZN(
        P3_U2888) );
  AOI22_X1 U21069 ( .A1(n19167), .A2(n18950), .B1(n19165), .B2(n18949), .ZN(
        n18948) );
  AOI22_X1 U21070 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19169), .B1(
        n19168), .B2(n18951), .ZN(n18947) );
  OAI211_X1 U21071 ( .C1(n19183), .C2(n18954), .A(n18948), .B(n18947), .ZN(
        P3_U2880) );
  AOI22_X1 U21072 ( .A1(n19092), .A2(n18950), .B1(n19174), .B2(n18949), .ZN(
        n18953) );
  AOI22_X1 U21073 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19179), .B1(
        n19178), .B2(n18951), .ZN(n18952) );
  OAI211_X1 U21074 ( .C1(n19037), .C2(n18954), .A(n18953), .B(n18952), .ZN(
        P3_U2872) );
  OAI22_X1 U21075 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19080), .ZN(n18955) );
  INV_X1 U21076 ( .A(n18955), .ZN(U254) );
  NAND2_X1 U21077 ( .A1(n19082), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18985) );
  NAND2_X1 U21078 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19082), .ZN(n18995) );
  INV_X1 U21079 ( .A(n18995), .ZN(n18982) );
  INV_X1 U21080 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n20646) );
  NOR2_X2 U21081 ( .A1(n18956), .A2(n20646), .ZN(n18990) );
  AOI22_X1 U21082 ( .A1(n19102), .A2(n18982), .B1(n19085), .B2(n18990), .ZN(
        n18959) );
  NOR2_X2 U21083 ( .A1(n18957), .A2(n19086), .ZN(n18992) );
  AOI22_X1 U21084 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19088), .B1(
        n19167), .B2(n18992), .ZN(n18958) );
  OAI211_X1 U21085 ( .C1(n19037), .C2(n18985), .A(n18959), .B(n18958), .ZN(
        P3_U2991) );
  AOI22_X1 U21086 ( .A1(n19109), .A2(n18982), .B1(n19091), .B2(n18990), .ZN(
        n18961) );
  AOI22_X1 U21087 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19093), .B1(
        n19092), .B2(n18992), .ZN(n18960) );
  OAI211_X1 U21088 ( .C1(n19096), .C2(n18985), .A(n18961), .B(n18960), .ZN(
        P3_U2983) );
  AOI22_X1 U21089 ( .A1(n19114), .A2(n18982), .B1(n19097), .B2(n18990), .ZN(
        n18963) );
  AOI22_X1 U21090 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19098), .B1(
        n19176), .B2(n18992), .ZN(n18962) );
  OAI211_X1 U21091 ( .C1(n19045), .C2(n18985), .A(n18963), .B(n18962), .ZN(
        P3_U2975) );
  AOI22_X1 U21092 ( .A1(n19120), .A2(n18982), .B1(n19101), .B2(n18990), .ZN(
        n18965) );
  AOI22_X1 U21093 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19103), .B1(
        n19102), .B2(n18992), .ZN(n18964) );
  OAI211_X1 U21094 ( .C1(n19106), .C2(n18985), .A(n18965), .B(n18964), .ZN(
        P3_U2967) );
  AOI22_X1 U21095 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19108), .B1(
        n19107), .B2(n18990), .ZN(n18967) );
  AOI22_X1 U21096 ( .A1(n19109), .A2(n18992), .B1(n19126), .B2(n18982), .ZN(
        n18966) );
  OAI211_X1 U21097 ( .C1(n19008), .C2(n18985), .A(n18967), .B(n18966), .ZN(
        P3_U2959) );
  INV_X1 U21098 ( .A(n18985), .ZN(n18991) );
  AOI22_X1 U21099 ( .A1(n19126), .A2(n18991), .B1(n19113), .B2(n18990), .ZN(
        n18969) );
  AOI22_X1 U21100 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19115), .B1(
        n19114), .B2(n18992), .ZN(n18968) );
  OAI211_X1 U21101 ( .C1(n19118), .C2(n18995), .A(n18969), .B(n18968), .ZN(
        P3_U2951) );
  AOI22_X1 U21102 ( .A1(n19137), .A2(n18982), .B1(n19119), .B2(n18990), .ZN(
        n18971) );
  AOI22_X1 U21103 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19121), .B1(
        n19120), .B2(n18992), .ZN(n18970) );
  OAI211_X1 U21104 ( .C1(n19118), .C2(n18985), .A(n18971), .B(n18970), .ZN(
        P3_U2943) );
  AOI22_X1 U21105 ( .A1(n19143), .A2(n18982), .B1(n19125), .B2(n18990), .ZN(
        n18973) );
  AOI22_X1 U21106 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19127), .B1(
        n19126), .B2(n18992), .ZN(n18972) );
  OAI211_X1 U21107 ( .C1(n19124), .C2(n18985), .A(n18973), .B(n18972), .ZN(
        P3_U2935) );
  AOI22_X1 U21108 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19133), .B1(
        n19131), .B2(n18990), .ZN(n18975) );
  AOI22_X1 U21109 ( .A1(n19132), .A2(n18992), .B1(n19148), .B2(n18982), .ZN(
        n18974) );
  OAI211_X1 U21110 ( .C1(n19130), .C2(n18985), .A(n18975), .B(n18974), .ZN(
        P3_U2927) );
  AOI22_X1 U21111 ( .A1(n19148), .A2(n18991), .B1(n19136), .B2(n18990), .ZN(
        n18977) );
  AOI22_X1 U21112 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19138), .B1(
        n19137), .B2(n18992), .ZN(n18976) );
  OAI211_X1 U21113 ( .C1(n19062), .C2(n18995), .A(n18977), .B(n18976), .ZN(
        P3_U2919) );
  AOI22_X1 U21114 ( .A1(n19155), .A2(n18991), .B1(n19142), .B2(n18990), .ZN(
        n18979) );
  AOI22_X1 U21115 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19144), .B1(
        n19143), .B2(n18992), .ZN(n18978) );
  OAI211_X1 U21116 ( .C1(n19152), .C2(n18995), .A(n18979), .B(n18978), .ZN(
        P3_U2911) );
  AOI22_X1 U21117 ( .A1(n19168), .A2(n18982), .B1(n19147), .B2(n18990), .ZN(
        n18981) );
  AOI22_X1 U21118 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19149), .B1(
        n19148), .B2(n18992), .ZN(n18980) );
  OAI211_X1 U21119 ( .C1(n19152), .C2(n18985), .A(n18981), .B(n18980), .ZN(
        P3_U2903) );
  AOI22_X1 U21120 ( .A1(n19178), .A2(n18982), .B1(n19153), .B2(n18990), .ZN(
        n18984) );
  AOI22_X1 U21121 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19154), .B1(
        n19155), .B2(n18992), .ZN(n18983) );
  OAI211_X1 U21122 ( .C1(n19158), .C2(n18985), .A(n18984), .B(n18983), .ZN(
        P3_U2895) );
  AOI22_X1 U21123 ( .A1(n19178), .A2(n18991), .B1(n19159), .B2(n18990), .ZN(
        n18987) );
  AOI22_X1 U21124 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19161), .B1(
        n19160), .B2(n18992), .ZN(n18986) );
  OAI211_X1 U21125 ( .C1(n19164), .C2(n18995), .A(n18987), .B(n18986), .ZN(
        P3_U2887) );
  AOI22_X1 U21126 ( .A1(n19167), .A2(n18991), .B1(n19165), .B2(n18990), .ZN(
        n18989) );
  AOI22_X1 U21127 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19169), .B1(
        n19168), .B2(n18992), .ZN(n18988) );
  OAI211_X1 U21128 ( .C1(n19183), .C2(n18995), .A(n18989), .B(n18988), .ZN(
        P3_U2879) );
  AOI22_X1 U21129 ( .A1(n19092), .A2(n18991), .B1(n19174), .B2(n18990), .ZN(
        n18994) );
  AOI22_X1 U21130 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19179), .B1(
        n19178), .B2(n18992), .ZN(n18993) );
  OAI211_X1 U21131 ( .C1(n19037), .C2(n18995), .A(n18994), .B(n18993), .ZN(
        P3_U2871) );
  OAI22_X1 U21132 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19080), .ZN(n18996) );
  INV_X1 U21133 ( .A(n18996), .ZN(U253) );
  NAND2_X1 U21134 ( .A1(n19082), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19030) );
  NAND2_X1 U21135 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19082), .ZN(n19036) );
  INV_X1 U21136 ( .A(n19036), .ZN(n19027) );
  AND2_X1 U21137 ( .A1(n19084), .A2(BUF2_REG_2__SCAN_IN), .ZN(n19031) );
  AOI22_X1 U21138 ( .A1(n19102), .A2(n19027), .B1(n19085), .B2(n19031), .ZN(
        n18999) );
  NOR2_X2 U21139 ( .A1(n18997), .A2(n19086), .ZN(n19033) );
  AOI22_X1 U21140 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19088), .B1(
        n19167), .B2(n19033), .ZN(n18998) );
  OAI211_X1 U21141 ( .C1(n19037), .C2(n19030), .A(n18999), .B(n18998), .ZN(
        P3_U2990) );
  INV_X1 U21142 ( .A(n19030), .ZN(n19032) );
  AOI22_X1 U21143 ( .A1(n19102), .A2(n19032), .B1(n19091), .B2(n19031), .ZN(
        n19001) );
  AOI22_X1 U21144 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19093), .B1(
        n19092), .B2(n19033), .ZN(n19000) );
  OAI211_X1 U21145 ( .C1(n19045), .C2(n19036), .A(n19001), .B(n19000), .ZN(
        P3_U2982) );
  AOI22_X1 U21146 ( .A1(n19109), .A2(n19032), .B1(n19097), .B2(n19031), .ZN(
        n19003) );
  AOI22_X1 U21147 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19098), .B1(
        n19176), .B2(n19033), .ZN(n19002) );
  OAI211_X1 U21148 ( .C1(n19106), .C2(n19036), .A(n19003), .B(n19002), .ZN(
        P3_U2974) );
  AOI22_X1 U21149 ( .A1(n19120), .A2(n19027), .B1(n19101), .B2(n19031), .ZN(
        n19005) );
  AOI22_X1 U21150 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19103), .B1(
        n19102), .B2(n19033), .ZN(n19004) );
  OAI211_X1 U21151 ( .C1(n19106), .C2(n19030), .A(n19005), .B(n19004), .ZN(
        P3_U2966) );
  AOI22_X1 U21152 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19108), .B1(
        n19107), .B2(n19031), .ZN(n19007) );
  AOI22_X1 U21153 ( .A1(n19109), .A2(n19033), .B1(n19126), .B2(n19027), .ZN(
        n19006) );
  OAI211_X1 U21154 ( .C1(n19008), .C2(n19030), .A(n19007), .B(n19006), .ZN(
        P3_U2958) );
  AOI22_X1 U21155 ( .A1(n19126), .A2(n19032), .B1(n19113), .B2(n19031), .ZN(
        n19010) );
  AOI22_X1 U21156 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19115), .B1(
        n19114), .B2(n19033), .ZN(n19009) );
  OAI211_X1 U21157 ( .C1(n19118), .C2(n19036), .A(n19010), .B(n19009), .ZN(
        P3_U2950) );
  AOI22_X1 U21158 ( .A1(n19137), .A2(n19027), .B1(n19119), .B2(n19031), .ZN(
        n19012) );
  AOI22_X1 U21159 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19121), .B1(
        n19120), .B2(n19033), .ZN(n19011) );
  OAI211_X1 U21160 ( .C1(n19118), .C2(n19030), .A(n19012), .B(n19011), .ZN(
        P3_U2942) );
  AOI22_X1 U21161 ( .A1(n19137), .A2(n19032), .B1(n19125), .B2(n19031), .ZN(
        n19014) );
  AOI22_X1 U21162 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19127), .B1(
        n19126), .B2(n19033), .ZN(n19013) );
  OAI211_X1 U21163 ( .C1(n19130), .C2(n19036), .A(n19014), .B(n19013), .ZN(
        P3_U2934) );
  AOI22_X1 U21164 ( .A1(n19148), .A2(n19027), .B1(n19131), .B2(n19031), .ZN(
        n19016) );
  AOI22_X1 U21165 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19133), .B1(
        n19132), .B2(n19033), .ZN(n19015) );
  OAI211_X1 U21166 ( .C1(n19130), .C2(n19030), .A(n19016), .B(n19015), .ZN(
        P3_U2926) );
  AOI22_X1 U21167 ( .A1(n19148), .A2(n19032), .B1(n19136), .B2(n19031), .ZN(
        n19018) );
  AOI22_X1 U21168 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19138), .B1(
        n19137), .B2(n19033), .ZN(n19017) );
  OAI211_X1 U21169 ( .C1(n19062), .C2(n19036), .A(n19018), .B(n19017), .ZN(
        P3_U2918) );
  AOI22_X1 U21170 ( .A1(n19142), .A2(n19031), .B1(n19160), .B2(n19027), .ZN(
        n19020) );
  AOI22_X1 U21171 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19144), .B1(
        n19143), .B2(n19033), .ZN(n19019) );
  OAI211_X1 U21172 ( .C1(n19062), .C2(n19030), .A(n19020), .B(n19019), .ZN(
        P3_U2910) );
  AOI22_X1 U21173 ( .A1(n19168), .A2(n19027), .B1(n19147), .B2(n19031), .ZN(
        n19022) );
  AOI22_X1 U21174 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19149), .B1(
        n19148), .B2(n19033), .ZN(n19021) );
  OAI211_X1 U21175 ( .C1(n19152), .C2(n19030), .A(n19022), .B(n19021), .ZN(
        P3_U2902) );
  AOI22_X1 U21176 ( .A1(n19168), .A2(n19032), .B1(n19153), .B2(n19031), .ZN(
        n19024) );
  AOI22_X1 U21177 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19154), .B1(
        n19155), .B2(n19033), .ZN(n19023) );
  OAI211_X1 U21178 ( .C1(n19067), .C2(n19036), .A(n19024), .B(n19023), .ZN(
        P3_U2894) );
  AOI22_X1 U21179 ( .A1(n19178), .A2(n19032), .B1(n19159), .B2(n19031), .ZN(
        n19026) );
  AOI22_X1 U21180 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19161), .B1(
        n19160), .B2(n19033), .ZN(n19025) );
  OAI211_X1 U21181 ( .C1(n19164), .C2(n19036), .A(n19026), .B(n19025), .ZN(
        P3_U2886) );
  AOI22_X1 U21182 ( .A1(n19092), .A2(n19027), .B1(n19165), .B2(n19031), .ZN(
        n19029) );
  AOI22_X1 U21183 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19169), .B1(
        n19168), .B2(n19033), .ZN(n19028) );
  OAI211_X1 U21184 ( .C1(n19164), .C2(n19030), .A(n19029), .B(n19028), .ZN(
        P3_U2878) );
  AOI22_X1 U21185 ( .A1(n19092), .A2(n19032), .B1(n19174), .B2(n19031), .ZN(
        n19035) );
  AOI22_X1 U21186 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19179), .B1(
        n19178), .B2(n19033), .ZN(n19034) );
  OAI211_X1 U21187 ( .C1(n19037), .C2(n19036), .A(n19035), .B(n19034), .ZN(
        P3_U2870) );
  OAI22_X1 U21188 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19080), .ZN(n19038) );
  INV_X1 U21189 ( .A(n19038), .ZN(U252) );
  NOR2_X1 U21190 ( .A1(n16551), .A2(n19083), .ZN(n19075) );
  INV_X1 U21191 ( .A(n19075), .ZN(n19073) );
  NAND2_X1 U21192 ( .A1(n19082), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19079) );
  INV_X1 U21193 ( .A(n19079), .ZN(n19070) );
  AOI22_X1 U21194 ( .A1(n19176), .A2(n19070), .B1(n19085), .B2(n19074), .ZN(
        n19040) );
  NOR2_X2 U21195 ( .A1(n20106), .A2(n19086), .ZN(n19076) );
  AOI22_X1 U21196 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19088), .B1(
        n19167), .B2(n19076), .ZN(n19039) );
  OAI211_X1 U21197 ( .C1(n19096), .C2(n19073), .A(n19040), .B(n19039), .ZN(
        P3_U2989) );
  AOI22_X1 U21198 ( .A1(n19102), .A2(n19070), .B1(n19091), .B2(n19074), .ZN(
        n19042) );
  AOI22_X1 U21199 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19093), .B1(
        n19092), .B2(n19076), .ZN(n19041) );
  OAI211_X1 U21200 ( .C1(n19045), .C2(n19073), .A(n19042), .B(n19041), .ZN(
        P3_U2981) );
  AOI22_X1 U21201 ( .A1(n19114), .A2(n19075), .B1(n19097), .B2(n19074), .ZN(
        n19044) );
  AOI22_X1 U21202 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19098), .B1(
        n19176), .B2(n19076), .ZN(n19043) );
  OAI211_X1 U21203 ( .C1(n19045), .C2(n19079), .A(n19044), .B(n19043), .ZN(
        P3_U2973) );
  AOI22_X1 U21204 ( .A1(n19120), .A2(n19075), .B1(n19101), .B2(n19074), .ZN(
        n19047) );
  AOI22_X1 U21205 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19103), .B1(
        n19102), .B2(n19076), .ZN(n19046) );
  OAI211_X1 U21206 ( .C1(n19106), .C2(n19079), .A(n19047), .B(n19046), .ZN(
        P3_U2965) );
  AOI22_X1 U21207 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19108), .B1(
        n19107), .B2(n19074), .ZN(n19049) );
  AOI22_X1 U21208 ( .A1(n19109), .A2(n19076), .B1(n19120), .B2(n19070), .ZN(
        n19048) );
  OAI211_X1 U21209 ( .C1(n19112), .C2(n19073), .A(n19049), .B(n19048), .ZN(
        P3_U2957) );
  AOI22_X1 U21210 ( .A1(n19132), .A2(n19075), .B1(n19113), .B2(n19074), .ZN(
        n19051) );
  AOI22_X1 U21211 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19115), .B1(
        n19114), .B2(n19076), .ZN(n19050) );
  OAI211_X1 U21212 ( .C1(n19112), .C2(n19079), .A(n19051), .B(n19050), .ZN(
        P3_U2949) );
  AOI22_X1 U21213 ( .A1(n19132), .A2(n19070), .B1(n19119), .B2(n19074), .ZN(
        n19053) );
  AOI22_X1 U21214 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19121), .B1(
        n19120), .B2(n19076), .ZN(n19052) );
  OAI211_X1 U21215 ( .C1(n19124), .C2(n19073), .A(n19053), .B(n19052), .ZN(
        P3_U2941) );
  AOI22_X1 U21216 ( .A1(n19143), .A2(n19075), .B1(n19125), .B2(n19074), .ZN(
        n19055) );
  AOI22_X1 U21217 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19127), .B1(
        n19126), .B2(n19076), .ZN(n19054) );
  OAI211_X1 U21218 ( .C1(n19124), .C2(n19079), .A(n19055), .B(n19054), .ZN(
        P3_U2933) );
  AOI22_X1 U21219 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19133), .B1(
        n19131), .B2(n19074), .ZN(n19057) );
  AOI22_X1 U21220 ( .A1(n19132), .A2(n19076), .B1(n19148), .B2(n19075), .ZN(
        n19056) );
  OAI211_X1 U21221 ( .C1(n19130), .C2(n19079), .A(n19057), .B(n19056), .ZN(
        P3_U2925) );
  AOI22_X1 U21222 ( .A1(n19155), .A2(n19075), .B1(n19136), .B2(n19074), .ZN(
        n19059) );
  AOI22_X1 U21223 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19138), .B1(
        n19137), .B2(n19076), .ZN(n19058) );
  OAI211_X1 U21224 ( .C1(n19141), .C2(n19079), .A(n19059), .B(n19058), .ZN(
        P3_U2917) );
  AOI22_X1 U21225 ( .A1(n19142), .A2(n19074), .B1(n19160), .B2(n19075), .ZN(
        n19061) );
  AOI22_X1 U21226 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19144), .B1(
        n19143), .B2(n19076), .ZN(n19060) );
  OAI211_X1 U21227 ( .C1(n19062), .C2(n19079), .A(n19061), .B(n19060), .ZN(
        P3_U2909) );
  AOI22_X1 U21228 ( .A1(n19168), .A2(n19075), .B1(n19147), .B2(n19074), .ZN(
        n19064) );
  AOI22_X1 U21229 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19149), .B1(
        n19148), .B2(n19076), .ZN(n19063) );
  OAI211_X1 U21230 ( .C1(n19152), .C2(n19079), .A(n19064), .B(n19063), .ZN(
        P3_U2901) );
  AOI22_X1 U21231 ( .A1(n19168), .A2(n19070), .B1(n19153), .B2(n19074), .ZN(
        n19066) );
  AOI22_X1 U21232 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19154), .B1(
        n19155), .B2(n19076), .ZN(n19065) );
  OAI211_X1 U21233 ( .C1(n19067), .C2(n19073), .A(n19066), .B(n19065), .ZN(
        P3_U2893) );
  AOI22_X1 U21234 ( .A1(n19178), .A2(n19070), .B1(n19159), .B2(n19074), .ZN(
        n19069) );
  AOI22_X1 U21235 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19161), .B1(
        n19160), .B2(n19076), .ZN(n19068) );
  OAI211_X1 U21236 ( .C1(n19164), .C2(n19073), .A(n19069), .B(n19068), .ZN(
        P3_U2885) );
  AOI22_X1 U21237 ( .A1(n19167), .A2(n19070), .B1(n19165), .B2(n19074), .ZN(
        n19072) );
  AOI22_X1 U21238 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19169), .B1(
        n19168), .B2(n19076), .ZN(n19071) );
  OAI211_X1 U21239 ( .C1(n19183), .C2(n19073), .A(n19072), .B(n19071), .ZN(
        P3_U2877) );
  AOI22_X1 U21240 ( .A1(n19176), .A2(n19075), .B1(n19174), .B2(n19074), .ZN(
        n19078) );
  AOI22_X1 U21241 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19179), .B1(
        n19178), .B2(n19076), .ZN(n19077) );
  OAI211_X1 U21242 ( .C1(n19183), .C2(n19079), .A(n19078), .B(n19077), .ZN(
        P3_U2869) );
  OAI22_X1 U21243 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19080), .ZN(n19081) );
  INV_X1 U21244 ( .A(n19081), .ZN(U251) );
  NAND2_X1 U21245 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19082), .ZN(n19172) );
  NOR2_X1 U21246 ( .A1(n19083), .A2(n20753), .ZN(n19166) );
  AND2_X1 U21247 ( .A1(n19084), .A2(BUF2_REG_0__SCAN_IN), .ZN(n19173) );
  AOI22_X1 U21248 ( .A1(n19176), .A2(n19166), .B1(n19085), .B2(n19173), .ZN(
        n19090) );
  NOR2_X2 U21249 ( .A1(n19087), .A2(n19086), .ZN(n19177) );
  AOI22_X1 U21250 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19088), .B1(
        n19167), .B2(n19177), .ZN(n19089) );
  OAI211_X1 U21251 ( .C1(n19096), .C2(n19172), .A(n19090), .B(n19089), .ZN(
        P3_U2988) );
  INV_X1 U21252 ( .A(n19166), .ZN(n19182) );
  INV_X1 U21253 ( .A(n19172), .ZN(n19175) );
  AOI22_X1 U21254 ( .A1(n19109), .A2(n19175), .B1(n19091), .B2(n19173), .ZN(
        n19095) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19093), .B1(
        n19092), .B2(n19177), .ZN(n19094) );
  OAI211_X1 U21256 ( .C1(n19096), .C2(n19182), .A(n19095), .B(n19094), .ZN(
        P3_U2980) );
  AOI22_X1 U21257 ( .A1(n19109), .A2(n19166), .B1(n19097), .B2(n19173), .ZN(
        n19100) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19098), .B1(
        n19176), .B2(n19177), .ZN(n19099) );
  OAI211_X1 U21259 ( .C1(n19106), .C2(n19172), .A(n19100), .B(n19099), .ZN(
        P3_U2972) );
  AOI22_X1 U21260 ( .A1(n19120), .A2(n19175), .B1(n19101), .B2(n19173), .ZN(
        n19105) );
  AOI22_X1 U21261 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19103), .B1(
        n19102), .B2(n19177), .ZN(n19104) );
  OAI211_X1 U21262 ( .C1(n19106), .C2(n19182), .A(n19105), .B(n19104), .ZN(
        P3_U2964) );
  AOI22_X1 U21263 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19108), .B1(
        n19107), .B2(n19173), .ZN(n19111) );
  AOI22_X1 U21264 ( .A1(n19109), .A2(n19177), .B1(n19120), .B2(n19166), .ZN(
        n19110) );
  OAI211_X1 U21265 ( .C1(n19112), .C2(n19172), .A(n19111), .B(n19110), .ZN(
        P3_U2956) );
  AOI22_X1 U21266 ( .A1(n19126), .A2(n19166), .B1(n19113), .B2(n19173), .ZN(
        n19117) );
  AOI22_X1 U21267 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19115), .B1(
        n19114), .B2(n19177), .ZN(n19116) );
  OAI211_X1 U21268 ( .C1(n19118), .C2(n19172), .A(n19117), .B(n19116), .ZN(
        P3_U2948) );
  AOI22_X1 U21269 ( .A1(n19132), .A2(n19166), .B1(n19119), .B2(n19173), .ZN(
        n19123) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19121), .B1(
        n19120), .B2(n19177), .ZN(n19122) );
  OAI211_X1 U21271 ( .C1(n19124), .C2(n19172), .A(n19123), .B(n19122), .ZN(
        P3_U2940) );
  AOI22_X1 U21272 ( .A1(n19137), .A2(n19166), .B1(n19125), .B2(n19173), .ZN(
        n19129) );
  AOI22_X1 U21273 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19127), .B1(
        n19126), .B2(n19177), .ZN(n19128) );
  OAI211_X1 U21274 ( .C1(n19130), .C2(n19172), .A(n19129), .B(n19128), .ZN(
        P3_U2932) );
  AOI22_X1 U21275 ( .A1(n19143), .A2(n19166), .B1(n19131), .B2(n19173), .ZN(
        n19135) );
  AOI22_X1 U21276 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19133), .B1(
        n19132), .B2(n19177), .ZN(n19134) );
  OAI211_X1 U21277 ( .C1(n19141), .C2(n19172), .A(n19135), .B(n19134), .ZN(
        P3_U2924) );
  AOI22_X1 U21278 ( .A1(n19155), .A2(n19175), .B1(n19136), .B2(n19173), .ZN(
        n19140) );
  AOI22_X1 U21279 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19138), .B1(
        n19137), .B2(n19177), .ZN(n19139) );
  OAI211_X1 U21280 ( .C1(n19141), .C2(n19182), .A(n19140), .B(n19139), .ZN(
        P3_U2916) );
  AOI22_X1 U21281 ( .A1(n19155), .A2(n19166), .B1(n19142), .B2(n19173), .ZN(
        n19146) );
  AOI22_X1 U21282 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19144), .B1(
        n19143), .B2(n19177), .ZN(n19145) );
  OAI211_X1 U21283 ( .C1(n19152), .C2(n19172), .A(n19146), .B(n19145), .ZN(
        P3_U2908) );
  AOI22_X1 U21284 ( .A1(n19168), .A2(n19175), .B1(n19147), .B2(n19173), .ZN(
        n19151) );
  AOI22_X1 U21285 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19149), .B1(
        n19148), .B2(n19177), .ZN(n19150) );
  OAI211_X1 U21286 ( .C1(n19152), .C2(n19182), .A(n19151), .B(n19150), .ZN(
        P3_U2900) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19173), .ZN(n19157) );
  AOI22_X1 U21288 ( .A1(n19155), .A2(n19177), .B1(n19178), .B2(n19175), .ZN(
        n19156) );
  OAI211_X1 U21289 ( .C1(n19158), .C2(n19182), .A(n19157), .B(n19156), .ZN(
        P3_U2892) );
  AOI22_X1 U21290 ( .A1(n19178), .A2(n19166), .B1(n19159), .B2(n19173), .ZN(
        n19163) );
  AOI22_X1 U21291 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19161), .B1(
        n19160), .B2(n19177), .ZN(n19162) );
  OAI211_X1 U21292 ( .C1(n19164), .C2(n19172), .A(n19163), .B(n19162), .ZN(
        P3_U2884) );
  AOI22_X1 U21293 ( .A1(n19167), .A2(n19166), .B1(n19165), .B2(n19173), .ZN(
        n19171) );
  AOI22_X1 U21294 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19169), .B1(
        n19168), .B2(n19177), .ZN(n19170) );
  OAI211_X1 U21295 ( .C1(n19183), .C2(n19172), .A(n19171), .B(n19170), .ZN(
        P3_U2876) );
  AOI22_X1 U21296 ( .A1(n19176), .A2(n19175), .B1(n19174), .B2(n19173), .ZN(
        n19181) );
  AOI22_X1 U21297 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19179), .B1(
        n19178), .B2(n19177), .ZN(n19180) );
  OAI211_X1 U21298 ( .C1(n19183), .C2(n19182), .A(n19181), .B(n19180), .ZN(
        P3_U2868) );
  AOI22_X1 U21299 ( .A1(n11040), .A2(n19633), .B1(n19184), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19187) );
  AOI22_X1 U21300 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19631), .B1(n19185), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19186) );
  NAND2_X1 U21301 ( .A1(n19187), .A2(n19186), .ZN(P2_U2888) );
  INV_X1 U21302 ( .A(n19188), .ZN(n19190) );
  AOI22_X1 U21303 ( .A1(P2_EAX_REG_15__SCAN_IN), .A2(n19631), .B1(n19191), 
        .B2(n19419), .ZN(n19192) );
  OAI21_X1 U21304 ( .B1(n19697), .B2(n19193), .A(n19192), .ZN(P2_U2904) );
  OAI222_X1 U21305 ( .A1(n19196), .A2(n19220), .B1(n19195), .B2(n19686), .C1(
        n19697), .C2(n19194), .ZN(P2_U2905) );
  AOI22_X1 U21306 ( .A1(P2_EAX_REG_13__SCAN_IN), .A2(n19631), .B1(n19197), 
        .B2(n19419), .ZN(n19198) );
  OAI21_X1 U21307 ( .B1(n19199), .B2(n19697), .A(n19198), .ZN(P2_U2906) );
  OAI222_X1 U21308 ( .A1(n19202), .A2(n19220), .B1(n19201), .B2(n19686), .C1(
        n19697), .C2(n19200), .ZN(P2_U2907) );
  INV_X1 U21309 ( .A(n19697), .ZN(n19210) );
  AOI22_X1 U21310 ( .A1(n19204), .A2(n19419), .B1(n19203), .B2(n19210), .ZN(
        n19205) );
  OAI21_X1 U21311 ( .B1(n19686), .B2(n19206), .A(n19205), .ZN(P2_U2908) );
  AOI22_X1 U21312 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19631), .B1(n19207), 
        .B2(n19419), .ZN(n19208) );
  OAI21_X1 U21313 ( .B1(n19209), .B2(n19697), .A(n19208), .ZN(P2_U2909) );
  AOI22_X1 U21314 ( .A1(n19212), .A2(n19419), .B1(n19211), .B2(n19210), .ZN(
        n19213) );
  OAI21_X1 U21315 ( .B1(n19686), .B2(n19214), .A(n19213), .ZN(P2_U2910) );
  OAI222_X1 U21316 ( .A1(n19217), .A2(n19220), .B1(n19216), .B2(n19686), .C1(
        n19697), .C2(n19215), .ZN(P2_U2911) );
  OAI222_X1 U21317 ( .A1(n19221), .A2(n19220), .B1(n19219), .B2(n19686), .C1(
        n19697), .C2(n19218), .ZN(P2_U2912) );
  NAND3_X1 U21318 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19233) );
  OAI21_X1 U21319 ( .B1(n19226), .B2(n19704), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19222) );
  OAI21_X1 U21320 ( .B1(n19233), .B2(n19355), .A(n19222), .ZN(n19705) );
  AOI22_X1 U21321 ( .A1(n19705), .A2(n15143), .B1(n19704), .B2(n19357), .ZN(
        n19232) );
  OAI21_X1 U21322 ( .B1(n19225), .B2(n19224), .A(n19233), .ZN(n19230) );
  INV_X1 U21323 ( .A(n19226), .ZN(n19228) );
  OAI21_X1 U21324 ( .B1(n19346), .B2(n19704), .A(n19362), .ZN(n19227) );
  OAI21_X1 U21325 ( .B1(n19228), .B2(n19364), .A(n19227), .ZN(n19229) );
  NAND2_X1 U21326 ( .A1(n19230), .A2(n19229), .ZN(n19708) );
  AOI22_X1 U21327 ( .A1(n19714), .A2(n19369), .B1(n19708), .B2(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19231) );
  OAI211_X1 U21328 ( .C1(n19372), .C2(n19817), .A(n19232), .B(n19231), .ZN(
        P2_U3175) );
  NOR2_X1 U21329 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19233), .ZN(
        n19713) );
  AOI22_X1 U21330 ( .A1(n19590), .A2(n19369), .B1(n19357), .B2(n19713), .ZN(
        n19243) );
  NAND2_X1 U21331 ( .A1(n19712), .A2(n19724), .ZN(n19234) );
  AOI21_X1 U21332 ( .B1(n19234), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19355), 
        .ZN(n19239) );
  AOI21_X1 U21333 ( .B1(n12099), .B2(n19235), .A(n19361), .ZN(n19236) );
  AOI21_X1 U21334 ( .B1(n19239), .B2(n19237), .A(n19236), .ZN(n19238) );
  AOI21_X1 U21335 ( .B1(n19713), .B2(n19362), .A(n19238), .ZN(n19716) );
  OAI21_X1 U21336 ( .B1(n19713), .B2(n19719), .A(n19239), .ZN(n19241) );
  OAI21_X1 U21337 ( .B1(n12099), .B2(n19713), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19240) );
  AOI22_X1 U21338 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19716), .B1(
        n15143), .B2(n19715), .ZN(n19242) );
  OAI211_X1 U21339 ( .C1(n19372), .C2(n19712), .A(n19243), .B(n19242), .ZN(
        P2_U3167) );
  NAND2_X1 U21340 ( .A1(n19244), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19251) );
  NOR2_X1 U21341 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19245), .ZN(
        n19725) );
  OAI21_X1 U21342 ( .B1(n12106), .B2(n19725), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19246) );
  OAI21_X1 U21343 ( .B1(n19355), .B2(n19251), .A(n19246), .ZN(n19726) );
  AOI22_X1 U21344 ( .A1(n19726), .A2(n15143), .B1(n19357), .B2(n19725), .ZN(
        n19256) );
  INV_X1 U21345 ( .A(n12106), .ZN(n19249) );
  NOR2_X1 U21346 ( .A1(n19249), .A2(n19364), .ZN(n19254) );
  INV_X1 U21347 ( .A(n19725), .ZN(n19250) );
  AOI21_X1 U21348 ( .B1(n19250), .B2(n19355), .A(n19700), .ZN(n19253) );
  OAI221_X1 U21349 ( .B1(n21597), .B2(n19737), .C1(n21597), .C2(n19495), .A(
        n19251), .ZN(n19252) );
  AOI22_X1 U21350 ( .A1(n19651), .A2(n19369), .B1(
        P2_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n19727), .ZN(n19255) );
  OAI211_X1 U21351 ( .C1(n19372), .C2(n19495), .A(n19256), .B(n19255), .ZN(
        P2_U3151) );
  NAND3_X1 U21352 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19257), .ZN(n19267) );
  NOR2_X1 U21353 ( .A1(n19353), .A2(n19267), .ZN(n19731) );
  OAI21_X1 U21354 ( .B1(n19259), .B2(n19731), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19258) );
  OAI21_X1 U21355 ( .B1(n19267), .B2(n19355), .A(n19258), .ZN(n19732) );
  AOI22_X1 U21356 ( .A1(n19732), .A2(n15143), .B1(n19357), .B2(n19731), .ZN(
        n19266) );
  OAI21_X1 U21357 ( .B1(n19431), .B2(n19328), .A(n19267), .ZN(n19263) );
  INV_X1 U21358 ( .A(n19259), .ZN(n19261) );
  AOI21_X1 U21359 ( .B1(n19731), .B2(n19362), .A(n19361), .ZN(n19260) );
  OAI21_X1 U21360 ( .B1(n19261), .B2(n19364), .A(n19260), .ZN(n19262) );
  NAND2_X1 U21361 ( .A1(n19263), .A2(n19262), .ZN(n19734) );
  AOI22_X1 U21362 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n19369), .ZN(n19265) );
  OAI211_X1 U21363 ( .C1(n19372), .C2(n19737), .A(n19266), .B(n19265), .ZN(
        P2_U3143) );
  NOR2_X1 U21364 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19267), .ZN(
        n19738) );
  INV_X1 U21365 ( .A(n19738), .ZN(n19388) );
  OAI22_X1 U21366 ( .A1(n19746), .A2(n19282), .B1(n19281), .B2(n19388), .ZN(
        n19268) );
  INV_X1 U21367 ( .A(n19268), .ZN(n19278) );
  OAI21_X1 U21368 ( .B1(n19739), .B2(n19733), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19269) );
  NAND2_X1 U21369 ( .A1(n19269), .A2(n19346), .ZN(n19276) );
  NOR2_X1 U21370 ( .A1(n19656), .A2(n19738), .ZN(n19275) );
  INV_X1 U21371 ( .A(n19275), .ZN(n19272) );
  INV_X1 U21372 ( .A(n19273), .ZN(n19270) );
  OAI211_X1 U21373 ( .C1(n19270), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19388), 
        .B(n19355), .ZN(n19271) );
  OAI211_X1 U21374 ( .C1(n19276), .C2(n19272), .A(n19362), .B(n19271), .ZN(
        n19741) );
  OAI21_X1 U21375 ( .B1(n19273), .B2(n19738), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19274) );
  AOI22_X1 U21376 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19741), .B1(
        n15143), .B2(n19740), .ZN(n19277) );
  OAI211_X1 U21377 ( .C1(n19372), .C2(n19744), .A(n19278), .B(n19277), .ZN(
        P2_U3135) );
  INV_X1 U21378 ( .A(n19298), .ZN(n19279) );
  NOR2_X1 U21379 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19280), .ZN(
        n19659) );
  INV_X1 U21380 ( .A(n19659), .ZN(n19753) );
  OAI22_X1 U21381 ( .A1(n19760), .A2(n19282), .B1(n19281), .B2(n19753), .ZN(
        n19283) );
  INV_X1 U21382 ( .A(n19283), .ZN(n19292) );
  NAND2_X1 U21383 ( .A1(n19760), .A2(n19754), .ZN(n19284) );
  AOI21_X1 U21384 ( .B1(n19284), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19355), 
        .ZN(n19287) );
  NAND2_X1 U21385 ( .A1(n19327), .A2(n19312), .ZN(n19294) );
  OAI21_X1 U21386 ( .B1(n19288), .B2(n19293), .A(n12654), .ZN(n19285) );
  AOI21_X1 U21387 ( .B1(n19287), .B2(n19294), .A(n19285), .ZN(n19286) );
  OAI21_X1 U21388 ( .B1(n19659), .B2(n19286), .A(n19362), .ZN(n19757) );
  INV_X1 U21389 ( .A(n19294), .ZN(n19761) );
  OAI21_X1 U21390 ( .B1(n19761), .B2(n19659), .A(n19287), .ZN(n19290) );
  OAI21_X1 U21391 ( .B1(n19288), .B2(n19659), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19289) );
  NAND2_X1 U21392 ( .A1(n19290), .A2(n19289), .ZN(n19756) );
  AOI22_X1 U21393 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n15143), .ZN(n19291) );
  OAI211_X1 U21394 ( .C1(n19372), .C2(n19754), .A(n19292), .B(n19291), .ZN(
        P2_U3119) );
  NOR2_X1 U21395 ( .A1(n12096), .A2(n19761), .ZN(n19295) );
  NAND2_X1 U21396 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19312), .ZN(
        n19303) );
  OAI22_X1 U21397 ( .A1(n19295), .A2(n19293), .B1(n19303), .B2(n19355), .ZN(
        n19762) );
  AOI22_X1 U21398 ( .A1(n19762), .A2(n15143), .B1(n19357), .B2(n19761), .ZN(
        n19300) );
  OAI22_X1 U21399 ( .A1(n19295), .A2(n19364), .B1(n19700), .B2(n19294), .ZN(
        n19297) );
  OAI21_X1 U21400 ( .B1(n21597), .B2(n19298), .A(n19303), .ZN(n19296) );
  OAI21_X1 U21401 ( .B1(n19361), .B2(n19297), .A(n19296), .ZN(n19764) );
  AOI22_X1 U21402 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19764), .B1(
        n19608), .B2(n19369), .ZN(n19299) );
  OAI211_X1 U21403 ( .C1(n19372), .C2(n19760), .A(n19300), .B(n19299), .ZN(
        P2_U3111) );
  NAND3_X1 U21404 ( .A1(n19302), .A2(n19312), .A3(n19301), .ZN(n19307) );
  NOR2_X1 U21405 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19303), .ZN(
        n19767) );
  OAI21_X1 U21406 ( .B1(n12104), .B2(n19767), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19304) );
  OAI21_X1 U21407 ( .B1(n19355), .B2(n19307), .A(n19304), .ZN(n19768) );
  AOI22_X1 U21408 ( .A1(n19768), .A2(n15143), .B1(n19357), .B2(n19767), .ZN(
        n19311) );
  INV_X1 U21409 ( .A(n12104), .ZN(n19306) );
  OAI21_X1 U21410 ( .B1(n19346), .B2(n19767), .A(n19362), .ZN(n19305) );
  OAI21_X1 U21411 ( .B1(n19306), .B2(n19364), .A(n19305), .ZN(n19309) );
  OAI221_X1 U21412 ( .B1(n21597), .B2(n19613), .C1(n21597), .C2(n19772), .A(
        n19307), .ZN(n19308) );
  AOI22_X1 U21413 ( .A1(n19774), .A2(n19369), .B1(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n19769), .ZN(n19310) );
  OAI211_X1 U21414 ( .C1(n19372), .C2(n19772), .A(n19311), .B(n19310), .ZN(
        P2_U3103) );
  NAND2_X1 U21415 ( .A1(n19312), .A2(n14986), .ZN(n19320) );
  NOR2_X1 U21416 ( .A1(n19353), .A2(n19320), .ZN(n19773) );
  AOI22_X1 U21417 ( .A1(n19781), .A2(n19369), .B1(n19357), .B2(n19773), .ZN(
        n19323) );
  OAI21_X1 U21418 ( .B1(n19314), .B2(n19313), .A(n19346), .ZN(n19321) );
  INV_X1 U21419 ( .A(n19320), .ZN(n19318) );
  INV_X1 U21420 ( .A(n12098), .ZN(n19316) );
  OAI21_X1 U21421 ( .B1(n19346), .B2(n19773), .A(n19362), .ZN(n19315) );
  OAI21_X1 U21422 ( .B1(n19316), .B2(n19364), .A(n19315), .ZN(n19317) );
  OAI21_X1 U21423 ( .B1(n19321), .B2(n19318), .A(n19317), .ZN(n19776) );
  OAI21_X1 U21424 ( .B1(n12098), .B2(n19773), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19319) );
  OAI21_X1 U21425 ( .B1(n19321), .B2(n19320), .A(n19319), .ZN(n19775) );
  AOI22_X1 U21426 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19776), .B1(
        n15143), .B2(n19775), .ZN(n19322) );
  OAI211_X1 U21427 ( .C1(n19372), .C2(n19613), .A(n19323), .B(n19322), .ZN(
        P2_U3095) );
  INV_X1 U21428 ( .A(n19324), .ZN(n19325) );
  AND2_X1 U21429 ( .A1(n19327), .A2(n19326), .ZN(n19787) );
  AOI22_X1 U21430 ( .A1(n19617), .A2(n19369), .B1(n19357), .B2(n19787), .ZN(
        n19337) );
  OAI21_X1 U21431 ( .B1(n19359), .B2(n19328), .A(n19346), .ZN(n19335) );
  NOR2_X1 U21432 ( .A1(n14986), .A2(n19352), .ZN(n19332) );
  INV_X1 U21433 ( .A(n19333), .ZN(n19330) );
  AOI21_X1 U21434 ( .B1(n19787), .B2(n19362), .A(n19361), .ZN(n19329) );
  OAI21_X1 U21435 ( .B1(n19330), .B2(n19364), .A(n19329), .ZN(n19331) );
  OAI21_X1 U21436 ( .B1(n19335), .B2(n19332), .A(n19331), .ZN(n19790) );
  INV_X1 U21437 ( .A(n19332), .ZN(n19338) );
  OAI21_X1 U21438 ( .B1(n19333), .B2(n19787), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19334) );
  OAI21_X1 U21439 ( .B1(n19335), .B2(n19338), .A(n19334), .ZN(n19789) );
  AOI22_X1 U21440 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19790), .B1(
        n15143), .B2(n19789), .ZN(n19336) );
  OAI211_X1 U21441 ( .C1(n19372), .C2(n19620), .A(n19337), .B(n19336), .ZN(
        P2_U3079) );
  NOR2_X1 U21442 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19338), .ZN(
        n19793) );
  OAI21_X1 U21443 ( .B1(n19344), .B2(n19793), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19340) );
  OR2_X1 U21444 ( .A1(n19339), .A2(n19352), .ZN(n19345) );
  NAND2_X1 U21445 ( .A1(n19340), .A2(n19345), .ZN(n19794) );
  AOI22_X1 U21446 ( .A1(n19794), .A2(n15143), .B1(n19357), .B2(n19793), .ZN(
        n19351) );
  NOR2_X2 U21447 ( .A1(n19342), .A2(n19341), .ZN(n19803) );
  INV_X1 U21448 ( .A(n19803), .ZN(n19522) );
  AOI21_X1 U21449 ( .B1(n19522), .B2(n19799), .A(n19343), .ZN(n19349) );
  AOI21_X1 U21450 ( .B1(n19344), .B2(n12654), .A(n19793), .ZN(n19347) );
  OAI21_X1 U21451 ( .B1(n19347), .B2(n19346), .A(n19345), .ZN(n19348) );
  OAI21_X1 U21452 ( .B1(n19349), .B2(n19348), .A(n19362), .ZN(n19796) );
  AOI22_X1 U21453 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19796), .B1(
        n19803), .B2(n19369), .ZN(n19350) );
  OAI211_X1 U21454 ( .C1(n19372), .C2(n19799), .A(n19351), .B(n19350), .ZN(
        P2_U3071) );
  NOR2_X1 U21455 ( .A1(n19352), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19367) );
  INV_X1 U21456 ( .A(n19367), .ZN(n19356) );
  NOR2_X1 U21457 ( .A1(n19353), .A2(n19356), .ZN(n19801) );
  OAI21_X1 U21458 ( .B1(n19360), .B2(n19801), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19354) );
  OAI21_X1 U21459 ( .B1(n19356), .B2(n19355), .A(n19354), .ZN(n19802) );
  AOI22_X1 U21460 ( .A1(n19802), .A2(n15143), .B1(n19357), .B2(n19801), .ZN(
        n19371) );
  NOR2_X1 U21461 ( .A1(n19359), .A2(n19358), .ZN(n19368) );
  INV_X1 U21462 ( .A(n19360), .ZN(n19365) );
  AOI21_X1 U21463 ( .B1(n19801), .B2(n19362), .A(n19361), .ZN(n19363) );
  OAI21_X1 U21464 ( .B1(n19365), .B2(n19364), .A(n19363), .ZN(n19366) );
  OAI21_X1 U21465 ( .B1(n19368), .B2(n19367), .A(n19366), .ZN(n19804) );
  AOI22_X1 U21466 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19804), .B1(
        n19811), .B2(n19369), .ZN(n19370) );
  OAI211_X1 U21467 ( .C1(n19372), .C2(n19522), .A(n19371), .B(n19370), .ZN(
        P2_U3063) );
  AOI22_X1 U21468 ( .A1(P2_EAX_REG_6__SCAN_IN), .A2(n19631), .B1(n11076), .B2(
        n19419), .ZN(n19373) );
  OAI21_X1 U21469 ( .B1(n19374), .B2(n19697), .A(n19373), .ZN(P2_U2913) );
  INV_X1 U21470 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n22166) );
  INV_X1 U21471 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n20706) );
  AOI22_X1 U21472 ( .A1(n19705), .A2(n19375), .B1(n19704), .B2(n19413), .ZN(
        n19378) );
  AOI22_X1 U21473 ( .A1(n19709), .A2(n19414), .B1(n19708), .B2(
        P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n19377) );
  OAI211_X1 U21474 ( .C1(n19412), .C2(n19712), .A(n19378), .B(n19377), .ZN(
        P2_U3174) );
  AOI22_X1 U21475 ( .A1(n19590), .A2(n19415), .B1(n19413), .B2(n19713), .ZN(
        n19380) );
  AOI22_X1 U21476 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19716), .B1(
        n19375), .B2(n19715), .ZN(n19379) );
  OAI211_X1 U21477 ( .C1(n19409), .C2(n19712), .A(n19380), .B(n19379), .ZN(
        P2_U3166) );
  AOI22_X1 U21478 ( .A1(n19720), .A2(n19375), .B1(n19413), .B2(n19719), .ZN(
        n19382) );
  AOI22_X1 U21479 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19721), .B1(
        n19590), .B2(n19414), .ZN(n19381) );
  OAI211_X1 U21480 ( .C1(n19412), .C2(n19495), .A(n19382), .B(n19381), .ZN(
        P2_U3158) );
  AOI22_X1 U21481 ( .A1(n19726), .A2(n19375), .B1(n19413), .B2(n19725), .ZN(
        n19384) );
  AOI22_X1 U21482 ( .A1(n19651), .A2(n19415), .B1(
        P2_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n19727), .ZN(n19383) );
  OAI211_X1 U21483 ( .C1(n19409), .C2(n19495), .A(n19384), .B(n19383), .ZN(
        P2_U3150) );
  AOI22_X1 U21484 ( .A1(n19732), .A2(n19375), .B1(n19413), .B2(n19731), .ZN(
        n19386) );
  AOI22_X1 U21485 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19734), .B1(
        n19651), .B2(n19414), .ZN(n19385) );
  OAI211_X1 U21486 ( .C1(n19412), .C2(n19744), .A(n19386), .B(n19385), .ZN(
        P2_U3142) );
  INV_X1 U21487 ( .A(n19413), .ZN(n19387) );
  OAI22_X1 U21488 ( .A1(n19746), .A2(n19412), .B1(n19388), .B2(n19387), .ZN(
        n19389) );
  INV_X1 U21489 ( .A(n19389), .ZN(n19391) );
  AOI22_X1 U21490 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19741), .B1(
        n19375), .B2(n19740), .ZN(n19390) );
  OAI211_X1 U21491 ( .C1(n19409), .C2(n19744), .A(n19391), .B(n19390), .ZN(
        P2_U3134) );
  AOI22_X1 U21492 ( .A1(n19739), .A2(n19414), .B1(n19656), .B2(n19413), .ZN(
        n19393) );
  AOI22_X1 U21493 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19749), .B1(
        n19375), .B2(n19748), .ZN(n19392) );
  OAI211_X1 U21494 ( .C1(n19412), .C2(n19754), .A(n19393), .B(n19392), .ZN(
        P2_U3126) );
  INV_X1 U21495 ( .A(n19754), .ZN(n19601) );
  AOI22_X1 U21496 ( .A1(n19601), .A2(n19414), .B1(n19659), .B2(n19413), .ZN(
        n19395) );
  AOI22_X1 U21497 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n19375), .ZN(n19394) );
  OAI211_X1 U21498 ( .C1(n19412), .C2(n19760), .A(n19395), .B(n19394), .ZN(
        P2_U3118) );
  AOI22_X1 U21499 ( .A1(n19762), .A2(n19375), .B1(n19761), .B2(n19413), .ZN(
        n19397) );
  AOI22_X1 U21500 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n19414), .ZN(n19396) );
  OAI211_X1 U21501 ( .C1(n19412), .C2(n19772), .A(n19397), .B(n19396), .ZN(
        P2_U3110) );
  AOI22_X1 U21502 ( .A1(n19768), .A2(n19375), .B1(n19413), .B2(n19767), .ZN(
        n19399) );
  AOI22_X1 U21503 ( .A1(n19774), .A2(n19415), .B1(
        P2_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n19769), .ZN(n19398) );
  OAI211_X1 U21504 ( .C1(n19409), .C2(n19772), .A(n19399), .B(n19398), .ZN(
        P2_U3102) );
  AOI22_X1 U21505 ( .A1(n19781), .A2(n19415), .B1(n19413), .B2(n19773), .ZN(
        n19401) );
  AOI22_X1 U21506 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19776), .B1(
        n19375), .B2(n19775), .ZN(n19400) );
  OAI211_X1 U21507 ( .C1(n19409), .C2(n19613), .A(n19401), .B(n19400), .ZN(
        P2_U3094) );
  INV_X1 U21508 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n19404) );
  AOI22_X1 U21509 ( .A1(n19414), .A2(n19781), .B1(n19780), .B2(n19413), .ZN(
        n19403) );
  AOI22_X1 U21510 ( .A1(n19375), .A2(n19782), .B1(n19788), .B2(n19415), .ZN(
        n19402) );
  OAI211_X1 U21511 ( .C1(n19786), .C2(n19404), .A(n19403), .B(n19402), .ZN(
        P2_U3086) );
  AOI22_X1 U21512 ( .A1(n19617), .A2(n19415), .B1(n19413), .B2(n19787), .ZN(
        n19406) );
  AOI22_X1 U21513 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19790), .B1(
        n19375), .B2(n19789), .ZN(n19405) );
  OAI211_X1 U21514 ( .C1(n19409), .C2(n19620), .A(n19406), .B(n19405), .ZN(
        P2_U3078) );
  AOI22_X1 U21515 ( .A1(n19794), .A2(n19375), .B1(n19413), .B2(n19793), .ZN(
        n19408) );
  AOI22_X1 U21516 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19796), .B1(
        n19803), .B2(n19415), .ZN(n19407) );
  OAI211_X1 U21517 ( .C1(n19409), .C2(n19799), .A(n19408), .B(n19407), .ZN(
        P2_U3070) );
  AOI22_X1 U21518 ( .A1(n19802), .A2(n19375), .B1(n19413), .B2(n19801), .ZN(
        n19411) );
  AOI22_X1 U21519 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19804), .B1(
        n19803), .B2(n19414), .ZN(n19410) );
  OAI211_X1 U21520 ( .C1(n19412), .C2(n19807), .A(n19411), .B(n19410), .ZN(
        P2_U3062) );
  AOI22_X1 U21521 ( .A1(n19414), .A2(n19811), .B1(n19809), .B2(n19413), .ZN(
        n19417) );
  AOI22_X1 U21522 ( .A1(n19709), .A2(n19415), .B1(n19813), .B2(n19375), .ZN(
        n19416) );
  OAI211_X1 U21523 ( .C1(n19680), .C2(n19418), .A(n19417), .B(n19416), .ZN(
        P2_U3054) );
  AOI22_X1 U21524 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19631), .B1(n19420), .B2(
        n19419), .ZN(n19435) );
  NOR2_X1 U21525 ( .A1(n19421), .A2(n19632), .ZN(n19426) );
  INV_X1 U21526 ( .A(n19426), .ZN(n19422) );
  OAI21_X1 U21527 ( .B1(n19424), .B2(n19423), .A(n19422), .ZN(n19635) );
  NOR2_X1 U21528 ( .A1(n19425), .A2(n19687), .ZN(n19690) );
  NOR2_X1 U21529 ( .A1(n19635), .A2(n19690), .ZN(n19634) );
  NOR2_X1 U21530 ( .A1(n19426), .A2(n19634), .ZN(n19427) );
  XOR2_X1 U21531 ( .A(n19578), .B(n19427), .Z(n19580) );
  INV_X1 U21532 ( .A(n19580), .ZN(n19429) );
  NAND2_X1 U21533 ( .A1(n19427), .A2(n19578), .ZN(n19428) );
  OAI21_X1 U21534 ( .B1(n19429), .B2(n19579), .A(n19428), .ZN(n19533) );
  XNOR2_X1 U21535 ( .A(n19431), .B(n19430), .ZN(n19534) );
  NOR2_X1 U21536 ( .A1(n19533), .A2(n19534), .ZN(n19532) );
  AOI21_X1 U21537 ( .B1(n19431), .B2(n19430), .A(n19532), .ZN(n19433) );
  NOR2_X1 U21538 ( .A1(n19433), .A2(n19432), .ZN(n19483) );
  OR3_X1 U21539 ( .A1(n19483), .A2(n19484), .A3(n19636), .ZN(n19434) );
  OAI211_X1 U21540 ( .C1(n19436), .C2(n19697), .A(n19435), .B(n19434), .ZN(
        P2_U2914) );
  INV_X1 U21541 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n22119) );
  NOR2_X2 U21542 ( .A1(n19436), .A2(n19700), .ZN(n19475) );
  NAND2_X1 U21543 ( .A1(n12357), .A2(n19702), .ZN(n19452) );
  AOI22_X1 U21544 ( .A1(n19705), .A2(n19475), .B1(n19704), .B2(n19473), .ZN(
        n19438) );
  AOI22_X1 U21545 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19698), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19699), .ZN(n19462) );
  AOI22_X1 U21546 ( .A1(n19714), .A2(n19474), .B1(n19708), .B2(
        P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n19437) );
  OAI211_X1 U21547 ( .C1(n19472), .C2(n19817), .A(n19438), .B(n19437), .ZN(
        P2_U3173) );
  AOI22_X1 U21548 ( .A1(n19714), .A2(n19476), .B1(n19473), .B2(n19713), .ZN(
        n19440) );
  AOI22_X1 U21549 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19716), .B1(
        n19475), .B2(n19715), .ZN(n19439) );
  OAI211_X1 U21550 ( .C1(n19462), .C2(n19724), .A(n19440), .B(n19439), .ZN(
        P2_U3165) );
  AOI22_X1 U21551 ( .A1(n19720), .A2(n19475), .B1(n19473), .B2(n19719), .ZN(
        n19442) );
  AOI22_X1 U21552 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19721), .B1(
        n19728), .B2(n19474), .ZN(n19441) );
  OAI211_X1 U21553 ( .C1(n19472), .C2(n19724), .A(n19442), .B(n19441), .ZN(
        P2_U3157) );
  AOI22_X1 U21554 ( .A1(n19726), .A2(n19475), .B1(n19473), .B2(n19725), .ZN(
        n19444) );
  AOI22_X1 U21555 ( .A1(n19651), .A2(n19474), .B1(
        P2_INSTQUEUE_REG_12__5__SCAN_IN), .B2(n19727), .ZN(n19443) );
  OAI211_X1 U21556 ( .C1(n19472), .C2(n19495), .A(n19444), .B(n19443), .ZN(
        P2_U3149) );
  AOI22_X1 U21557 ( .A1(n19732), .A2(n19475), .B1(n19473), .B2(n19731), .ZN(
        n19446) );
  AOI22_X1 U21558 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n19474), .ZN(n19445) );
  OAI211_X1 U21559 ( .C1(n19472), .C2(n19737), .A(n19446), .B(n19445), .ZN(
        P2_U3141) );
  AOI22_X1 U21560 ( .A1(n19739), .A2(n19474), .B1(n19473), .B2(n19738), .ZN(
        n19448) );
  AOI22_X1 U21561 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19741), .B1(
        n19475), .B2(n19740), .ZN(n19447) );
  OAI211_X1 U21562 ( .C1(n19472), .C2(n19744), .A(n19448), .B(n19447), .ZN(
        P2_U3133) );
  OAI22_X1 U21563 ( .A1(n19746), .A2(n19472), .B1(n19745), .B2(n19452), .ZN(
        n19449) );
  INV_X1 U21564 ( .A(n19449), .ZN(n19451) );
  AOI22_X1 U21565 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19749), .B1(
        n19475), .B2(n19748), .ZN(n19450) );
  OAI211_X1 U21566 ( .C1(n19462), .C2(n19754), .A(n19451), .B(n19450), .ZN(
        P2_U3125) );
  OAI22_X1 U21567 ( .A1(n19760), .A2(n19462), .B1(n19753), .B2(n19452), .ZN(
        n19453) );
  INV_X1 U21568 ( .A(n19453), .ZN(n19455) );
  AOI22_X1 U21569 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n19475), .ZN(n19454) );
  OAI211_X1 U21570 ( .C1(n19472), .C2(n19754), .A(n19455), .B(n19454), .ZN(
        P2_U3117) );
  AOI22_X1 U21571 ( .A1(n19762), .A2(n19475), .B1(n19761), .B2(n19473), .ZN(
        n19457) );
  AOI22_X1 U21572 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n19476), .ZN(n19456) );
  OAI211_X1 U21573 ( .C1(n19462), .C2(n19772), .A(n19457), .B(n19456), .ZN(
        P2_U3109) );
  AOI22_X1 U21574 ( .A1(n19768), .A2(n19475), .B1(n19473), .B2(n19767), .ZN(
        n19459) );
  AOI22_X1 U21575 ( .A1(n19774), .A2(n19474), .B1(
        P2_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n19769), .ZN(n19458) );
  OAI211_X1 U21576 ( .C1(n19472), .C2(n19772), .A(n19459), .B(n19458), .ZN(
        P2_U3101) );
  AOI22_X1 U21577 ( .A1(n19774), .A2(n19476), .B1(n19473), .B2(n19773), .ZN(
        n19461) );
  AOI22_X1 U21578 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19776), .B1(
        n19475), .B2(n19775), .ZN(n19460) );
  OAI211_X1 U21579 ( .C1(n19462), .C2(n19779), .A(n19461), .B(n19460), .ZN(
        P2_U3093) );
  INV_X1 U21580 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n19465) );
  AOI22_X1 U21581 ( .A1(n19781), .A2(n19476), .B1(n19780), .B2(n19473), .ZN(
        n19464) );
  AOI22_X1 U21582 ( .A1(n19475), .A2(n19782), .B1(n19788), .B2(n19474), .ZN(
        n19463) );
  OAI211_X1 U21583 ( .C1(n19786), .C2(n19465), .A(n19464), .B(n19463), .ZN(
        P2_U3085) );
  AOI22_X1 U21584 ( .A1(n19617), .A2(n19474), .B1(n19473), .B2(n19787), .ZN(
        n19467) );
  AOI22_X1 U21585 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19790), .B1(
        n19475), .B2(n19789), .ZN(n19466) );
  OAI211_X1 U21586 ( .C1(n19472), .C2(n19620), .A(n19467), .B(n19466), .ZN(
        P2_U3077) );
  AOI22_X1 U21587 ( .A1(n19794), .A2(n19475), .B1(n19473), .B2(n19793), .ZN(
        n19469) );
  AOI22_X1 U21588 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19796), .B1(
        n19803), .B2(n19474), .ZN(n19468) );
  OAI211_X1 U21589 ( .C1(n19472), .C2(n19799), .A(n19469), .B(n19468), .ZN(
        P2_U3069) );
  AOI22_X1 U21590 ( .A1(n19802), .A2(n19475), .B1(n19473), .B2(n19801), .ZN(
        n19471) );
  AOI22_X1 U21591 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19804), .B1(
        n19811), .B2(n19474), .ZN(n19470) );
  OAI211_X1 U21592 ( .C1(n19472), .C2(n19522), .A(n19471), .B(n19470), .ZN(
        P2_U3061) );
  AOI22_X1 U21593 ( .A1(n19709), .A2(n19474), .B1(n19809), .B2(n19473), .ZN(
        n19478) );
  AOI22_X1 U21594 ( .A1(n19811), .A2(n19476), .B1(n19813), .B2(n19475), .ZN(
        n19477) );
  OAI211_X1 U21595 ( .C1(n19680), .C2(n19479), .A(n19478), .B(n19477), .ZN(
        P2_U3053) );
  OAI22_X1 U21596 ( .A1(n19481), .A2(n19688), .B1(n19686), .B2(n19480), .ZN(
        n19482) );
  INV_X1 U21597 ( .A(n19482), .ZN(n19487) );
  XOR2_X1 U21598 ( .A(n19484), .B(n19483), .Z(n19485) );
  INV_X1 U21599 ( .A(n19636), .ZN(n19691) );
  NAND2_X1 U21600 ( .A1(n19485), .A2(n19691), .ZN(n19486) );
  OAI211_X1 U21601 ( .C1(n19488), .C2(n19697), .A(n19487), .B(n19486), .ZN(
        P2_U2915) );
  NOR2_X2 U21602 ( .A1(n19488), .A2(n19700), .ZN(n19526) );
  NOR2_X2 U21603 ( .A1(n11867), .A2(n19641), .ZN(n19524) );
  AOI22_X1 U21604 ( .A1(n19705), .A2(n19526), .B1(n19704), .B2(n19524), .ZN(
        n19490) );
  AOI22_X1 U21605 ( .A1(n19714), .A2(n19527), .B1(n19708), .B2(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n19489) );
  OAI211_X1 U21606 ( .C1(n19523), .C2(n19817), .A(n19490), .B(n19489), .ZN(
        P2_U3172) );
  AOI22_X1 U21607 ( .A1(n19714), .A2(n19525), .B1(n19524), .B2(n19713), .ZN(
        n19492) );
  AOI22_X1 U21608 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19716), .B1(
        n19526), .B2(n19715), .ZN(n19491) );
  OAI211_X1 U21609 ( .C1(n19517), .C2(n19724), .A(n19492), .B(n19491), .ZN(
        P2_U3164) );
  AOI22_X1 U21610 ( .A1(n19720), .A2(n19526), .B1(n19524), .B2(n19719), .ZN(
        n19494) );
  AOI22_X1 U21611 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19721), .B1(
        n19590), .B2(n19525), .ZN(n19493) );
  OAI211_X1 U21612 ( .C1(n19517), .C2(n19495), .A(n19494), .B(n19493), .ZN(
        P2_U3156) );
  AOI22_X1 U21613 ( .A1(n19726), .A2(n19526), .B1(n19524), .B2(n19725), .ZN(
        n19497) );
  AOI22_X1 U21614 ( .A1(n19525), .A2(n19728), .B1(
        P2_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n19727), .ZN(n19496) );
  OAI211_X1 U21615 ( .C1(n19517), .C2(n19737), .A(n19497), .B(n19496), .ZN(
        P2_U3148) );
  AOI22_X1 U21616 ( .A1(n19732), .A2(n19526), .B1(n19524), .B2(n19731), .ZN(
        n19499) );
  AOI22_X1 U21617 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19734), .B1(
        n19651), .B2(n19525), .ZN(n19498) );
  OAI211_X1 U21618 ( .C1(n19517), .C2(n19744), .A(n19499), .B(n19498), .ZN(
        P2_U3140) );
  AOI22_X1 U21619 ( .A1(n19733), .A2(n19525), .B1(n19738), .B2(n19524), .ZN(
        n19501) );
  AOI22_X1 U21620 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19741), .B1(
        n19526), .B2(n19740), .ZN(n19500) );
  OAI211_X1 U21621 ( .C1(n19517), .C2(n19746), .A(n19501), .B(n19500), .ZN(
        P2_U3132) );
  AOI22_X1 U21622 ( .A1(n19601), .A2(n19527), .B1(n19656), .B2(n19524), .ZN(
        n19503) );
  AOI22_X1 U21623 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19749), .B1(
        n19526), .B2(n19748), .ZN(n19502) );
  OAI211_X1 U21624 ( .C1(n19523), .C2(n19746), .A(n19503), .B(n19502), .ZN(
        P2_U3124) );
  AOI22_X1 U21625 ( .A1(n19601), .A2(n19525), .B1(n19659), .B2(n19524), .ZN(
        n19505) );
  AOI22_X1 U21626 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n19526), .ZN(n19504) );
  OAI211_X1 U21627 ( .C1(n19517), .C2(n19760), .A(n19505), .B(n19504), .ZN(
        P2_U3116) );
  AOI22_X1 U21628 ( .A1(n19762), .A2(n19526), .B1(n19761), .B2(n19524), .ZN(
        n19507) );
  AOI22_X1 U21629 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19764), .B1(
        n19608), .B2(n19527), .ZN(n19506) );
  OAI211_X1 U21630 ( .C1(n19523), .C2(n19760), .A(n19507), .B(n19506), .ZN(
        P2_U3108) );
  AOI22_X1 U21631 ( .A1(n19768), .A2(n19526), .B1(n19524), .B2(n19767), .ZN(
        n19509) );
  AOI22_X1 U21632 ( .A1(n19608), .A2(n19525), .B1(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n19769), .ZN(n19508) );
  OAI211_X1 U21633 ( .C1(n19517), .C2(n19613), .A(n19509), .B(n19508), .ZN(
        P2_U3100) );
  AOI22_X1 U21634 ( .A1(n19527), .A2(n19781), .B1(n19524), .B2(n19773), .ZN(
        n19511) );
  AOI22_X1 U21635 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19776), .B1(
        n19526), .B2(n19775), .ZN(n19510) );
  OAI211_X1 U21636 ( .C1(n19523), .C2(n19613), .A(n19511), .B(n19510), .ZN(
        P2_U3092) );
  INV_X1 U21637 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n19514) );
  AOI22_X1 U21638 ( .A1(n19525), .A2(n19781), .B1(n19780), .B2(n19524), .ZN(
        n19513) );
  AOI22_X1 U21639 ( .A1(n19526), .A2(n19782), .B1(n19788), .B2(n19527), .ZN(
        n19512) );
  OAI211_X1 U21640 ( .C1(n19786), .C2(n19514), .A(n19513), .B(n19512), .ZN(
        P2_U3084) );
  AOI22_X1 U21641 ( .A1(n19525), .A2(n19788), .B1(n19524), .B2(n19787), .ZN(
        n19516) );
  AOI22_X1 U21642 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19790), .B1(
        n19526), .B2(n19789), .ZN(n19515) );
  OAI211_X1 U21643 ( .C1(n19517), .C2(n19799), .A(n19516), .B(n19515), .ZN(
        P2_U3076) );
  AOI22_X1 U21644 ( .A1(n19794), .A2(n19526), .B1(n19524), .B2(n19793), .ZN(
        n19519) );
  AOI22_X1 U21645 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19796), .B1(
        n19803), .B2(n19527), .ZN(n19518) );
  OAI211_X1 U21646 ( .C1(n19523), .C2(n19799), .A(n19519), .B(n19518), .ZN(
        P2_U3068) );
  AOI22_X1 U21647 ( .A1(n19802), .A2(n19526), .B1(n19524), .B2(n19801), .ZN(
        n19521) );
  AOI22_X1 U21648 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19804), .B1(
        n19811), .B2(n19527), .ZN(n19520) );
  OAI211_X1 U21649 ( .C1(n19523), .C2(n19522), .A(n19521), .B(n19520), .ZN(
        P2_U3060) );
  AOI22_X1 U21650 ( .A1(n19525), .A2(n19811), .B1(n19809), .B2(n19524), .ZN(
        n19529) );
  AOI22_X1 U21651 ( .A1(n19709), .A2(n19527), .B1(n19813), .B2(n19526), .ZN(
        n19528) );
  OAI211_X1 U21652 ( .C1(n19680), .C2(n19530), .A(n19529), .B(n19528), .ZN(
        P2_U3052) );
  AOI22_X1 U21653 ( .A1(n19633), .A2(n19531), .B1(n19631), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19537) );
  AOI21_X1 U21654 ( .B1(n19534), .B2(n19533), .A(n19532), .ZN(n19535) );
  OR2_X1 U21655 ( .A1(n19535), .A2(n19636), .ZN(n19536) );
  OAI211_X1 U21656 ( .C1(n19538), .C2(n19697), .A(n19537), .B(n19536), .ZN(
        P2_U2916) );
  NOR2_X2 U21657 ( .A1(n19538), .A2(n19700), .ZN(n19574) );
  NOR2_X2 U21658 ( .A1(n11880), .A2(n19641), .ZN(n19572) );
  AOI22_X1 U21659 ( .A1(n19705), .A2(n19574), .B1(n19704), .B2(n19572), .ZN(
        n19540) );
  AOI22_X1 U21660 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19699), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19698), .ZN(n19568) );
  AOI22_X1 U21661 ( .A1(n19709), .A2(n19573), .B1(n19708), .B2(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n19539) );
  OAI211_X1 U21662 ( .C1(n19571), .C2(n19712), .A(n19540), .B(n19539), .ZN(
        P2_U3171) );
  AOI22_X1 U21663 ( .A1(n19714), .A2(n19573), .B1(n19572), .B2(n19713), .ZN(
        n19542) );
  AOI22_X1 U21664 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19716), .B1(
        n19574), .B2(n19715), .ZN(n19541) );
  OAI211_X1 U21665 ( .C1(n19571), .C2(n19724), .A(n19542), .B(n19541), .ZN(
        P2_U3163) );
  AOI22_X1 U21666 ( .A1(n19720), .A2(n19574), .B1(n19572), .B2(n19719), .ZN(
        n19544) );
  AOI22_X1 U21667 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19721), .B1(
        n19728), .B2(n19575), .ZN(n19543) );
  OAI211_X1 U21668 ( .C1(n19568), .C2(n19724), .A(n19544), .B(n19543), .ZN(
        P2_U3155) );
  AOI22_X1 U21669 ( .A1(n19726), .A2(n19574), .B1(n19572), .B2(n19725), .ZN(
        n19546) );
  AOI22_X1 U21670 ( .A1(n19728), .A2(n19573), .B1(
        P2_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n19727), .ZN(n19545) );
  OAI211_X1 U21671 ( .C1(n19571), .C2(n19737), .A(n19546), .B(n19545), .ZN(
        P2_U3147) );
  AOI22_X1 U21672 ( .A1(n19732), .A2(n19574), .B1(n19572), .B2(n19731), .ZN(
        n19548) );
  AOI22_X1 U21673 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19734), .B1(
        n19651), .B2(n19573), .ZN(n19547) );
  OAI211_X1 U21674 ( .C1(n19571), .C2(n19744), .A(n19548), .B(n19547), .ZN(
        P2_U3139) );
  AOI22_X1 U21675 ( .A1(n19733), .A2(n19573), .B1(n19572), .B2(n19738), .ZN(
        n19550) );
  AOI22_X1 U21676 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19741), .B1(
        n19574), .B2(n19740), .ZN(n19549) );
  OAI211_X1 U21677 ( .C1(n19571), .C2(n19746), .A(n19550), .B(n19549), .ZN(
        P2_U3131) );
  AOI22_X1 U21678 ( .A1(n19739), .A2(n19573), .B1(n19656), .B2(n19572), .ZN(
        n19552) );
  AOI22_X1 U21679 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19749), .B1(
        n19574), .B2(n19748), .ZN(n19551) );
  OAI211_X1 U21680 ( .C1(n19571), .C2(n19754), .A(n19552), .B(n19551), .ZN(
        P2_U3123) );
  AOI22_X1 U21681 ( .A1(n19763), .A2(n19575), .B1(n19659), .B2(n19572), .ZN(
        n19554) );
  AOI22_X1 U21682 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n19574), .ZN(n19553) );
  OAI211_X1 U21683 ( .C1(n19568), .C2(n19754), .A(n19554), .B(n19553), .ZN(
        P2_U3115) );
  AOI22_X1 U21684 ( .A1(n19762), .A2(n19574), .B1(n19761), .B2(n19572), .ZN(
        n19556) );
  AOI22_X1 U21685 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19764), .B1(
        n19608), .B2(n19575), .ZN(n19555) );
  OAI211_X1 U21686 ( .C1(n19568), .C2(n19760), .A(n19556), .B(n19555), .ZN(
        P2_U3107) );
  AOI22_X1 U21687 ( .A1(n19768), .A2(n19574), .B1(n19572), .B2(n19767), .ZN(
        n19558) );
  AOI22_X1 U21688 ( .A1(n19575), .A2(n19774), .B1(
        P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n19769), .ZN(n19557) );
  OAI211_X1 U21689 ( .C1(n19568), .C2(n19772), .A(n19558), .B(n19557), .ZN(
        P2_U3099) );
  AOI22_X1 U21690 ( .A1(n19774), .A2(n19573), .B1(n19572), .B2(n19773), .ZN(
        n19560) );
  AOI22_X1 U21691 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19776), .B1(
        n19574), .B2(n19775), .ZN(n19559) );
  OAI211_X1 U21692 ( .C1(n19571), .C2(n19779), .A(n19560), .B(n19559), .ZN(
        P2_U3091) );
  INV_X1 U21693 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n19563) );
  AOI22_X1 U21694 ( .A1(n19781), .A2(n19573), .B1(n19780), .B2(n19572), .ZN(
        n19562) );
  AOI22_X1 U21695 ( .A1(n19574), .A2(n19782), .B1(n19788), .B2(n19575), .ZN(
        n19561) );
  OAI211_X1 U21696 ( .C1(n19786), .C2(n19563), .A(n19562), .B(n19561), .ZN(
        P2_U3083) );
  AOI22_X1 U21697 ( .A1(n19788), .A2(n19573), .B1(n19572), .B2(n19787), .ZN(
        n19565) );
  AOI22_X1 U21698 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19790), .B1(
        n19574), .B2(n19789), .ZN(n19564) );
  OAI211_X1 U21699 ( .C1(n19571), .C2(n19799), .A(n19565), .B(n19564), .ZN(
        P2_U3075) );
  AOI22_X1 U21700 ( .A1(n19794), .A2(n19574), .B1(n19572), .B2(n19793), .ZN(
        n19567) );
  AOI22_X1 U21701 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19796), .B1(
        n19803), .B2(n19575), .ZN(n19566) );
  OAI211_X1 U21702 ( .C1(n19568), .C2(n19799), .A(n19567), .B(n19566), .ZN(
        P2_U3067) );
  AOI22_X1 U21703 ( .A1(n19802), .A2(n19574), .B1(n19572), .B2(n19801), .ZN(
        n19570) );
  AOI22_X1 U21704 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19804), .B1(
        n19803), .B2(n19573), .ZN(n19569) );
  OAI211_X1 U21705 ( .C1(n19571), .C2(n19807), .A(n19570), .B(n19569), .ZN(
        P2_U3059) );
  AOI22_X1 U21706 ( .A1(n19811), .A2(n19573), .B1(n19809), .B2(n19572), .ZN(
        n19577) );
  AOI22_X1 U21707 ( .A1(n19709), .A2(n19575), .B1(n19813), .B2(n19574), .ZN(
        n19576) );
  OAI211_X1 U21708 ( .C1(n19680), .C2(n13172), .A(n19577), .B(n19576), .ZN(
        P2_U3051) );
  AOI22_X1 U21709 ( .A1(n19578), .A2(n19633), .B1(n19631), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n19583) );
  XNOR2_X1 U21710 ( .A(n19580), .B(n19579), .ZN(n19581) );
  NAND2_X1 U21711 ( .A1(n19581), .A2(n19691), .ZN(n19582) );
  OAI211_X1 U21712 ( .C1(n19584), .C2(n19697), .A(n19583), .B(n19582), .ZN(
        P2_U2917) );
  AOI22_X1 U21713 ( .A1(n19705), .A2(n19626), .B1(n19704), .B2(n19625), .ZN(
        n19587) );
  AOI22_X1 U21714 ( .A1(n19709), .A2(n19627), .B1(n19708), .B2(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n19586) );
  OAI211_X1 U21715 ( .C1(n19630), .C2(n19712), .A(n19587), .B(n19586), .ZN(
        P2_U3170) );
  AOI22_X1 U21716 ( .A1(n19714), .A2(n19627), .B1(n19625), .B2(n19713), .ZN(
        n19589) );
  AOI22_X1 U21717 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19716), .B1(
        n19626), .B2(n19715), .ZN(n19588) );
  OAI211_X1 U21718 ( .C1(n19630), .C2(n19724), .A(n19589), .B(n19588), .ZN(
        P2_U3162) );
  INV_X1 U21719 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n19593) );
  AOI22_X1 U21720 ( .A1(n19720), .A2(n19626), .B1(n19625), .B2(n19719), .ZN(
        n19592) );
  AOI22_X1 U21721 ( .A1(n19728), .A2(n19621), .B1(n19590), .B2(n19627), .ZN(
        n19591) );
  OAI211_X1 U21722 ( .C1(n19594), .C2(n19593), .A(n19592), .B(n19591), .ZN(
        P2_U3154) );
  AOI22_X1 U21723 ( .A1(n19726), .A2(n19626), .B1(n19625), .B2(n19725), .ZN(
        n19596) );
  AOI22_X1 U21724 ( .A1(n19627), .A2(n19728), .B1(
        P2_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n19727), .ZN(n19595) );
  OAI211_X1 U21725 ( .C1(n19630), .C2(n19737), .A(n19596), .B(n19595), .ZN(
        P2_U3146) );
  AOI22_X1 U21726 ( .A1(n19732), .A2(n19626), .B1(n19625), .B2(n19731), .ZN(
        n19598) );
  AOI22_X1 U21727 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n19621), .ZN(n19597) );
  OAI211_X1 U21728 ( .C1(n19624), .C2(n19737), .A(n19598), .B(n19597), .ZN(
        P2_U3138) );
  AOI22_X1 U21729 ( .A1(n19739), .A2(n19621), .B1(n19625), .B2(n19738), .ZN(
        n19600) );
  AOI22_X1 U21730 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19741), .B1(
        n19626), .B2(n19740), .ZN(n19599) );
  OAI211_X1 U21731 ( .C1(n19624), .C2(n19744), .A(n19600), .B(n19599), .ZN(
        P2_U3130) );
  AOI22_X1 U21732 ( .A1(n19601), .A2(n19621), .B1(n19625), .B2(n19656), .ZN(
        n19603) );
  AOI22_X1 U21733 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19749), .B1(
        n19626), .B2(n19748), .ZN(n19602) );
  OAI211_X1 U21734 ( .C1(n19624), .C2(n19746), .A(n19603), .B(n19602), .ZN(
        P2_U3122) );
  AOI22_X1 U21735 ( .A1(n19763), .A2(n19621), .B1(n19625), .B2(n19659), .ZN(
        n19605) );
  AOI22_X1 U21736 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n19626), .ZN(n19604) );
  OAI211_X1 U21737 ( .C1(n19624), .C2(n19754), .A(n19605), .B(n19604), .ZN(
        P2_U3114) );
  AOI22_X1 U21738 ( .A1(n19762), .A2(n19626), .B1(n19625), .B2(n19761), .ZN(
        n19607) );
  AOI22_X1 U21739 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n19627), .ZN(n19606) );
  OAI211_X1 U21740 ( .C1(n19630), .C2(n19772), .A(n19607), .B(n19606), .ZN(
        P2_U3106) );
  AOI22_X1 U21741 ( .A1(n19768), .A2(n19626), .B1(n19625), .B2(n19767), .ZN(
        n19610) );
  AOI22_X1 U21742 ( .A1(n19608), .A2(n19627), .B1(
        P2_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n19769), .ZN(n19609) );
  OAI211_X1 U21743 ( .C1(n19630), .C2(n19613), .A(n19610), .B(n19609), .ZN(
        P2_U3098) );
  AOI22_X1 U21744 ( .A1(n19621), .A2(n19781), .B1(n19625), .B2(n19773), .ZN(
        n19612) );
  AOI22_X1 U21745 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19776), .B1(
        n19626), .B2(n19775), .ZN(n19611) );
  OAI211_X1 U21746 ( .C1(n19624), .C2(n19613), .A(n19612), .B(n19611), .ZN(
        P2_U3090) );
  INV_X1 U21747 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n19616) );
  AOI22_X1 U21748 ( .A1(n19627), .A2(n19781), .B1(n19625), .B2(n19780), .ZN(
        n19615) );
  AOI22_X1 U21749 ( .A1(n19626), .A2(n19782), .B1(n19788), .B2(n19621), .ZN(
        n19614) );
  OAI211_X1 U21750 ( .C1(n19786), .C2(n19616), .A(n19615), .B(n19614), .ZN(
        P2_U3082) );
  AOI22_X1 U21751 ( .A1(n19621), .A2(n19617), .B1(n19625), .B2(n19787), .ZN(
        n19619) );
  AOI22_X1 U21752 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19790), .B1(
        n19626), .B2(n19789), .ZN(n19618) );
  OAI211_X1 U21753 ( .C1(n19624), .C2(n19620), .A(n19619), .B(n19618), .ZN(
        P2_U3074) );
  AOI22_X1 U21754 ( .A1(n19794), .A2(n19626), .B1(n19625), .B2(n19793), .ZN(
        n19623) );
  AOI22_X1 U21755 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19796), .B1(
        n19803), .B2(n19621), .ZN(n19622) );
  OAI211_X1 U21756 ( .C1(n19624), .C2(n19799), .A(n19623), .B(n19622), .ZN(
        P2_U3066) );
  AOI22_X1 U21757 ( .A1(n19802), .A2(n19626), .B1(n19625), .B2(n19801), .ZN(
        n19629) );
  AOI22_X1 U21758 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19804), .B1(
        n19803), .B2(n19627), .ZN(n19628) );
  OAI211_X1 U21759 ( .C1(n19630), .C2(n19807), .A(n19629), .B(n19628), .ZN(
        P2_U3058) );
  AOI22_X1 U21760 ( .A1(n19633), .A2(n19632), .B1(n19631), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19639) );
  AOI21_X1 U21761 ( .B1(n19690), .B2(n19635), .A(n19634), .ZN(n19637) );
  OR2_X1 U21762 ( .A1(n19637), .A2(n19636), .ZN(n19638) );
  OAI211_X1 U21763 ( .C1(n19640), .C2(n19697), .A(n19639), .B(n19638), .ZN(
        P2_U2918) );
  NOR2_X2 U21764 ( .A1(n19640), .A2(n19700), .ZN(n19681) );
  NOR2_X2 U21765 ( .A1(n19642), .A2(n19641), .ZN(n19678) );
  AOI22_X1 U21766 ( .A1(n19705), .A2(n19681), .B1(n19704), .B2(n19678), .ZN(
        n19644) );
  AOI22_X1 U21767 ( .A1(n19714), .A2(n19679), .B1(n19708), .B2(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n19643) );
  OAI211_X1 U21768 ( .C1(n19684), .C2(n19817), .A(n19644), .B(n19643), .ZN(
        P2_U3169) );
  AOI22_X1 U21769 ( .A1(n19714), .A2(n19674), .B1(n19678), .B2(n19713), .ZN(
        n19646) );
  AOI22_X1 U21770 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19716), .B1(
        n19681), .B2(n19715), .ZN(n19645) );
  OAI211_X1 U21771 ( .C1(n19677), .C2(n19724), .A(n19646), .B(n19645), .ZN(
        P2_U3161) );
  AOI22_X1 U21772 ( .A1(n19720), .A2(n19681), .B1(n19678), .B2(n19719), .ZN(
        n19648) );
  AOI22_X1 U21773 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19721), .B1(
        n19728), .B2(n19679), .ZN(n19647) );
  OAI211_X1 U21774 ( .C1(n19684), .C2(n19724), .A(n19648), .B(n19647), .ZN(
        P2_U3153) );
  AOI22_X1 U21775 ( .A1(n19726), .A2(n19681), .B1(n19678), .B2(n19725), .ZN(
        n19650) );
  AOI22_X1 U21776 ( .A1(n19674), .A2(n19728), .B1(
        P2_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n19727), .ZN(n19649) );
  OAI211_X1 U21777 ( .C1(n19677), .C2(n19737), .A(n19650), .B(n19649), .ZN(
        P2_U3145) );
  AOI22_X1 U21778 ( .A1(n19732), .A2(n19681), .B1(n19678), .B2(n19731), .ZN(
        n19653) );
  AOI22_X1 U21779 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19734), .B1(
        n19651), .B2(n19674), .ZN(n19652) );
  OAI211_X1 U21780 ( .C1(n19677), .C2(n19744), .A(n19653), .B(n19652), .ZN(
        P2_U3137) );
  AOI22_X1 U21781 ( .A1(n19739), .A2(n19679), .B1(n19678), .B2(n19738), .ZN(
        n19655) );
  AOI22_X1 U21782 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19741), .B1(
        n19681), .B2(n19740), .ZN(n19654) );
  OAI211_X1 U21783 ( .C1(n19684), .C2(n19744), .A(n19655), .B(n19654), .ZN(
        P2_U3129) );
  AOI22_X1 U21784 ( .A1(n19739), .A2(n19674), .B1(n19656), .B2(n19678), .ZN(
        n19658) );
  AOI22_X1 U21785 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19749), .B1(
        n19681), .B2(n19748), .ZN(n19657) );
  OAI211_X1 U21786 ( .C1(n19677), .C2(n19754), .A(n19658), .B(n19657), .ZN(
        P2_U3121) );
  AOI22_X1 U21787 ( .A1(n19763), .A2(n19679), .B1(n19659), .B2(n19678), .ZN(
        n19661) );
  AOI22_X1 U21788 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n19681), .ZN(n19660) );
  OAI211_X1 U21789 ( .C1(n19684), .C2(n19754), .A(n19661), .B(n19660), .ZN(
        P2_U3113) );
  AOI22_X1 U21790 ( .A1(n19762), .A2(n19681), .B1(n19761), .B2(n19678), .ZN(
        n19663) );
  AOI22_X1 U21791 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n19674), .ZN(n19662) );
  OAI211_X1 U21792 ( .C1(n19677), .C2(n19772), .A(n19663), .B(n19662), .ZN(
        P2_U3105) );
  AOI22_X1 U21793 ( .A1(n19768), .A2(n19681), .B1(n19678), .B2(n19767), .ZN(
        n19665) );
  AOI22_X1 U21794 ( .A1(n19679), .A2(n19774), .B1(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n19769), .ZN(n19664) );
  OAI211_X1 U21795 ( .C1(n19684), .C2(n19772), .A(n19665), .B(n19664), .ZN(
        P2_U3097) );
  AOI22_X1 U21796 ( .A1(n19674), .A2(n19774), .B1(n19678), .B2(n19773), .ZN(
        n19667) );
  AOI22_X1 U21797 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19776), .B1(
        n19681), .B2(n19775), .ZN(n19666) );
  OAI211_X1 U21798 ( .C1(n19677), .C2(n19779), .A(n19667), .B(n19666), .ZN(
        P2_U3089) );
  AOI22_X1 U21799 ( .A1(n19674), .A2(n19781), .B1(n19780), .B2(n19678), .ZN(
        n19669) );
  AOI22_X1 U21800 ( .A1(n19681), .A2(n19782), .B1(n19788), .B2(n19679), .ZN(
        n19668) );
  OAI211_X1 U21801 ( .C1(n19786), .C2(n13130), .A(n19669), .B(n19668), .ZN(
        P2_U3081) );
  AOI22_X1 U21802 ( .A1(n19674), .A2(n19788), .B1(n19678), .B2(n19787), .ZN(
        n19671) );
  AOI22_X1 U21803 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19790), .B1(
        n19681), .B2(n19789), .ZN(n19670) );
  OAI211_X1 U21804 ( .C1(n19677), .C2(n19799), .A(n19671), .B(n19670), .ZN(
        P2_U3073) );
  AOI22_X1 U21805 ( .A1(n19794), .A2(n19681), .B1(n19678), .B2(n19793), .ZN(
        n19673) );
  AOI22_X1 U21806 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19796), .B1(
        n19803), .B2(n19679), .ZN(n19672) );
  OAI211_X1 U21807 ( .C1(n19684), .C2(n19799), .A(n19673), .B(n19672), .ZN(
        P2_U3065) );
  AOI22_X1 U21808 ( .A1(n19802), .A2(n19681), .B1(n19678), .B2(n19801), .ZN(
        n19676) );
  AOI22_X1 U21809 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19804), .B1(
        n19803), .B2(n19674), .ZN(n19675) );
  OAI211_X1 U21810 ( .C1(n19677), .C2(n19807), .A(n19676), .B(n19675), .ZN(
        P2_U3057) );
  AOI22_X1 U21811 ( .A1(n19709), .A2(n19679), .B1(n19809), .B2(n19678), .ZN(
        n19683) );
  INV_X1 U21812 ( .A(n19680), .ZN(n19814) );
  AOI22_X1 U21813 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19814), .B1(
        n19813), .B2(n19681), .ZN(n19682) );
  OAI211_X1 U21814 ( .C1(n19684), .C2(n19807), .A(n19683), .B(n19682), .ZN(
        P2_U3049) );
  OAI22_X1 U21815 ( .A1(n19688), .A2(n19687), .B1(n19686), .B2(n19685), .ZN(
        n19689) );
  INV_X1 U21816 ( .A(n19689), .ZN(n19696) );
  INV_X1 U21817 ( .A(n19690), .ZN(n19692) );
  OAI211_X1 U21818 ( .C1(n19694), .C2(n19693), .A(n19692), .B(n19691), .ZN(
        n19695) );
  OAI211_X1 U21819 ( .C1(n19701), .C2(n19697), .A(n19696), .B(n19695), .ZN(
        P2_U2919) );
  NOR2_X2 U21820 ( .A1(n19701), .A2(n19700), .ZN(n19812) );
  AND2_X1 U21821 ( .A1(n19703), .A2(n19702), .ZN(n19808) );
  AOI22_X1 U21822 ( .A1(n19705), .A2(n19812), .B1(n19704), .B2(n19808), .ZN(
        n19711) );
  INV_X1 U21823 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n21747) );
  AOI22_X1 U21824 ( .A1(n19709), .A2(n19810), .B1(n19708), .B2(
        P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n19710) );
  OAI211_X1 U21825 ( .C1(n19818), .C2(n19712), .A(n19711), .B(n19710), .ZN(
        P2_U3168) );
  AOI22_X1 U21826 ( .A1(n19714), .A2(n19810), .B1(n19808), .B2(n19713), .ZN(
        n19718) );
  AOI22_X1 U21827 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19716), .B1(
        n19812), .B2(n19715), .ZN(n19717) );
  OAI211_X1 U21828 ( .C1(n19818), .C2(n19724), .A(n19718), .B(n19717), .ZN(
        P2_U3160) );
  AOI22_X1 U21829 ( .A1(n19720), .A2(n19812), .B1(n19808), .B2(n19719), .ZN(
        n19723) );
  INV_X1 U21830 ( .A(n19818), .ZN(n19795) );
  AOI22_X1 U21831 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19721), .B1(
        n19728), .B2(n19795), .ZN(n19722) );
  OAI211_X1 U21832 ( .C1(n19800), .C2(n19724), .A(n19723), .B(n19722), .ZN(
        P2_U3152) );
  AOI22_X1 U21833 ( .A1(n19726), .A2(n19812), .B1(n19808), .B2(n19725), .ZN(
        n19730) );
  AOI22_X1 U21834 ( .A1(n19728), .A2(n19810), .B1(
        P2_INSTQUEUE_REG_12__0__SCAN_IN), .B2(n19727), .ZN(n19729) );
  OAI211_X1 U21835 ( .C1(n19818), .C2(n19737), .A(n19730), .B(n19729), .ZN(
        P2_U3144) );
  AOI22_X1 U21836 ( .A1(n19732), .A2(n19812), .B1(n19808), .B2(n19731), .ZN(
        n19736) );
  AOI22_X1 U21837 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19734), .B1(
        n19733), .B2(n19795), .ZN(n19735) );
  OAI211_X1 U21838 ( .C1(n19800), .C2(n19737), .A(n19736), .B(n19735), .ZN(
        P2_U3136) );
  AOI22_X1 U21839 ( .A1(n19739), .A2(n19795), .B1(n19738), .B2(n19808), .ZN(
        n19743) );
  AOI22_X1 U21840 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19741), .B1(
        n19812), .B2(n19740), .ZN(n19742) );
  OAI211_X1 U21841 ( .C1(n19800), .C2(n19744), .A(n19743), .B(n19742), .ZN(
        P2_U3128) );
  INV_X1 U21842 ( .A(n19808), .ZN(n19752) );
  OAI22_X1 U21843 ( .A1(n19746), .A2(n19800), .B1(n19745), .B2(n19752), .ZN(
        n19747) );
  INV_X1 U21844 ( .A(n19747), .ZN(n19751) );
  AOI22_X1 U21845 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19749), .B1(
        n19812), .B2(n19748), .ZN(n19750) );
  OAI211_X1 U21846 ( .C1(n19818), .C2(n19754), .A(n19751), .B(n19750), .ZN(
        P2_U3120) );
  OAI22_X1 U21847 ( .A1(n19754), .A2(n19800), .B1(n19753), .B2(n19752), .ZN(
        n19755) );
  INV_X1 U21848 ( .A(n19755), .ZN(n19759) );
  AOI22_X1 U21849 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19757), .B1(
        n19756), .B2(n19812), .ZN(n19758) );
  OAI211_X1 U21850 ( .C1(n19818), .C2(n19760), .A(n19759), .B(n19758), .ZN(
        P2_U3112) );
  AOI22_X1 U21851 ( .A1(n19762), .A2(n19812), .B1(n19761), .B2(n19808), .ZN(
        n19766) );
  AOI22_X1 U21852 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19764), .B1(
        n19763), .B2(n19810), .ZN(n19765) );
  OAI211_X1 U21853 ( .C1(n19818), .C2(n19772), .A(n19766), .B(n19765), .ZN(
        P2_U3104) );
  AOI22_X1 U21854 ( .A1(n19768), .A2(n19812), .B1(n19808), .B2(n19767), .ZN(
        n19771) );
  AOI22_X1 U21855 ( .A1(n19795), .A2(n19774), .B1(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n19769), .ZN(n19770) );
  OAI211_X1 U21856 ( .C1(n19800), .C2(n19772), .A(n19771), .B(n19770), .ZN(
        P2_U3096) );
  AOI22_X1 U21857 ( .A1(n19774), .A2(n19810), .B1(n19808), .B2(n19773), .ZN(
        n19778) );
  AOI22_X1 U21858 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19776), .B1(
        n19812), .B2(n19775), .ZN(n19777) );
  OAI211_X1 U21859 ( .C1(n19818), .C2(n19779), .A(n19778), .B(n19777), .ZN(
        P2_U3088) );
  INV_X1 U21860 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U21861 ( .A1(n19781), .A2(n19810), .B1(n19780), .B2(n19808), .ZN(
        n19784) );
  AOI22_X1 U21862 ( .A1(n19812), .A2(n19782), .B1(n19788), .B2(n19795), .ZN(
        n19783) );
  OAI211_X1 U21863 ( .C1(n19786), .C2(n19785), .A(n19784), .B(n19783), .ZN(
        P2_U3080) );
  AOI22_X1 U21864 ( .A1(n19788), .A2(n19810), .B1(n19808), .B2(n19787), .ZN(
        n19792) );
  AOI22_X1 U21865 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19790), .B1(
        n19812), .B2(n19789), .ZN(n19791) );
  OAI211_X1 U21866 ( .C1(n19818), .C2(n19799), .A(n19792), .B(n19791), .ZN(
        P2_U3072) );
  AOI22_X1 U21867 ( .A1(n19794), .A2(n19812), .B1(n19808), .B2(n19793), .ZN(
        n19798) );
  AOI22_X1 U21868 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19796), .B1(
        n19803), .B2(n19795), .ZN(n19797) );
  OAI211_X1 U21869 ( .C1(n19800), .C2(n19799), .A(n19798), .B(n19797), .ZN(
        P2_U3064) );
  AOI22_X1 U21870 ( .A1(n19802), .A2(n19812), .B1(n19808), .B2(n19801), .ZN(
        n19806) );
  AOI22_X1 U21871 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19804), .B1(
        n19803), .B2(n19810), .ZN(n19805) );
  OAI211_X1 U21872 ( .C1(n19818), .C2(n19807), .A(n19806), .B(n19805), .ZN(
        P2_U3056) );
  AOI22_X1 U21873 ( .A1(n19811), .A2(n19810), .B1(n19809), .B2(n19808), .ZN(
        n19816) );
  AOI22_X1 U21874 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19814), .B1(
        n19813), .B2(n19812), .ZN(n19815) );
  OAI211_X1 U21875 ( .C1(n19818), .C2(n19817), .A(n19816), .B(n19815), .ZN(
        P2_U3048) );
  INV_X1 U21876 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20097) );
  INV_X1 U21877 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n19819) );
  AOI222_X1 U21878 ( .A1(n20097), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20099), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n19819), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n19820) );
  INV_X1 U21879 ( .A(n19878), .ZN(n19881) );
  AOI22_X1 U21880 ( .A1(n19881), .A2(n19822), .B1(n19821), .B2(n19878), .ZN(
        U376) );
  INV_X1 U21881 ( .A(n19878), .ZN(n19833) );
  OAI22_X1 U21882 ( .A1(n19878), .A2(P3_ADDRESS_REG_1__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n19833), .ZN(n19823) );
  INV_X1 U21883 ( .A(n19823), .ZN(U365) );
  OAI22_X1 U21884 ( .A1(n19878), .A2(P3_ADDRESS_REG_2__SCAN_IN), .B1(
        P2_ADDRESS_REG_2__SCAN_IN), .B2(n19833), .ZN(n19824) );
  INV_X1 U21885 ( .A(n19824), .ZN(U354) );
  AOI22_X1 U21886 ( .A1(n19833), .A2(n19826), .B1(n19825), .B2(n19878), .ZN(
        U353) );
  AOI22_X1 U21887 ( .A1(n19833), .A2(n19828), .B1(n19827), .B2(n19878), .ZN(
        U352) );
  AOI22_X1 U21888 ( .A1(n19833), .A2(n19830), .B1(n19829), .B2(n19878), .ZN(
        U351) );
  AOI22_X1 U21889 ( .A1(n19833), .A2(n19832), .B1(n19831), .B2(n19878), .ZN(
        U350) );
  AOI22_X1 U21890 ( .A1(n19881), .A2(n19835), .B1(n19834), .B2(n19878), .ZN(
        U349) );
  AOI22_X1 U21891 ( .A1(n19881), .A2(n19837), .B1(n19836), .B2(n19878), .ZN(
        U348) );
  AOI22_X1 U21892 ( .A1(n19881), .A2(n19839), .B1(n19838), .B2(n19878), .ZN(
        U347) );
  AOI22_X1 U21893 ( .A1(n19881), .A2(n19841), .B1(n19840), .B2(n19878), .ZN(
        U375) );
  AOI22_X1 U21894 ( .A1(n19881), .A2(n19843), .B1(n19842), .B2(n19878), .ZN(
        U374) );
  AOI22_X1 U21895 ( .A1(n19881), .A2(n19845), .B1(n19844), .B2(n19878), .ZN(
        U373) );
  AOI22_X1 U21896 ( .A1(n19881), .A2(n19847), .B1(n19846), .B2(n19878), .ZN(
        U372) );
  AOI22_X1 U21897 ( .A1(n19881), .A2(n19849), .B1(n19848), .B2(n19878), .ZN(
        U371) );
  AOI22_X1 U21898 ( .A1(n19881), .A2(n19851), .B1(n19850), .B2(n19878), .ZN(
        U370) );
  AOI22_X1 U21899 ( .A1(n19881), .A2(n19853), .B1(n19852), .B2(n19878), .ZN(
        U369) );
  AOI22_X1 U21900 ( .A1(n19881), .A2(n19855), .B1(n19854), .B2(n19878), .ZN(
        U368) );
  AOI22_X1 U21901 ( .A1(n19881), .A2(n19857), .B1(n19856), .B2(n19878), .ZN(
        U367) );
  AOI22_X1 U21902 ( .A1(n19881), .A2(n19859), .B1(n19858), .B2(n19878), .ZN(
        U366) );
  AOI22_X1 U21903 ( .A1(n19881), .A2(n19861), .B1(n19860), .B2(n19878), .ZN(
        U364) );
  AOI22_X1 U21904 ( .A1(n19881), .A2(n19863), .B1(n19862), .B2(n19878), .ZN(
        U363) );
  AOI22_X1 U21905 ( .A1(n19881), .A2(n19865), .B1(n19864), .B2(n19878), .ZN(
        U362) );
  AOI22_X1 U21906 ( .A1(n19881), .A2(n19867), .B1(n19866), .B2(n19878), .ZN(
        U361) );
  AOI22_X1 U21907 ( .A1(n19881), .A2(n19869), .B1(n19868), .B2(n19878), .ZN(
        U360) );
  AOI22_X1 U21908 ( .A1(n19881), .A2(n19871), .B1(n19870), .B2(n19878), .ZN(
        U359) );
  AOI22_X1 U21909 ( .A1(n19881), .A2(n19873), .B1(n19872), .B2(n19878), .ZN(
        U358) );
  AOI22_X1 U21910 ( .A1(n19881), .A2(n19875), .B1(n19874), .B2(n19878), .ZN(
        U357) );
  AOI22_X1 U21911 ( .A1(n19881), .A2(n19877), .B1(n19876), .B2(n19878), .ZN(
        U356) );
  AOI22_X1 U21912 ( .A1(n19881), .A2(n19880), .B1(n19879), .B2(n19878), .ZN(
        U355) );
  AOI22_X1 U21913 ( .A1(n21264), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19883) );
  OAI21_X1 U21914 ( .B1(n19884), .B2(n19907), .A(n19883), .ZN(P1_U2936) );
  AOI22_X1 U21915 ( .A1(n19897), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19885) );
  OAI21_X1 U21916 ( .B1(n19886), .B2(n19907), .A(n19885), .ZN(P1_U2935) );
  AOI22_X1 U21917 ( .A1(n19897), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19894), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19887) );
  OAI21_X1 U21918 ( .B1(n19888), .B2(n19907), .A(n19887), .ZN(P1_U2934) );
  AOI22_X1 U21919 ( .A1(n19897), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19894), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19889) );
  OAI21_X1 U21920 ( .B1(n19890), .B2(n19907), .A(n19889), .ZN(P1_U2933) );
  AOI22_X1 U21921 ( .A1(n19897), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19894), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19891) );
  OAI21_X1 U21922 ( .B1(n19892), .B2(n19907), .A(n19891), .ZN(P1_U2932) );
  AOI22_X1 U21923 ( .A1(n19897), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19894), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19893) );
  OAI21_X1 U21924 ( .B1(n14070), .B2(n19907), .A(n19893), .ZN(P1_U2931) );
  AOI22_X1 U21925 ( .A1(n19897), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19894), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19895) );
  OAI21_X1 U21926 ( .B1(n14080), .B2(n19907), .A(n19895), .ZN(P1_U2930) );
  AOI22_X1 U21927 ( .A1(n21264), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19896) );
  OAI21_X1 U21928 ( .B1(n14018), .B2(n19907), .A(n19896), .ZN(P1_U2929) );
  AOI22_X1 U21929 ( .A1(n19897), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19898) );
  OAI21_X1 U21930 ( .B1(n15351), .B2(n19907), .A(n19898), .ZN(P1_U2928) );
  AOI22_X1 U21931 ( .A1(n21264), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19899) );
  OAI21_X1 U21932 ( .B1(n15449), .B2(n19907), .A(n19899), .ZN(P1_U2927) );
  AOI22_X1 U21933 ( .A1(n21264), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19900) );
  OAI21_X1 U21934 ( .B1(n15462), .B2(n19907), .A(n19900), .ZN(P1_U2926) );
  AOI22_X1 U21935 ( .A1(n21264), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19901) );
  OAI21_X1 U21936 ( .B1(n15550), .B2(n19907), .A(n19901), .ZN(P1_U2925) );
  AOI22_X1 U21937 ( .A1(n21264), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19902) );
  OAI21_X1 U21938 ( .B1(n15597), .B2(n19907), .A(n19902), .ZN(P1_U2924) );
  AOI22_X1 U21939 ( .A1(n21264), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19903) );
  OAI21_X1 U21940 ( .B1(n15590), .B2(n19907), .A(n19903), .ZN(P1_U2923) );
  AOI22_X1 U21941 ( .A1(n21264), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19904) );
  OAI21_X1 U21942 ( .B1(n15621), .B2(n19907), .A(n19904), .ZN(P1_U2922) );
  AOI22_X1 U21943 ( .A1(n21264), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n19905), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19906) );
  OAI21_X1 U21944 ( .B1(n19908), .B2(n19907), .A(n19906), .ZN(P1_U2921) );
  OR2_X1 U21945 ( .A1(n21611), .A2(n22329), .ZN(n19942) );
  INV_X1 U21946 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21369) );
  OAI222_X1 U21947 ( .A1(n19942), .A2(n15268), .B1(n19909), .B2(n22328), .C1(
        n21369), .C2(n19946), .ZN(P1_U3197) );
  INV_X1 U21948 ( .A(n19942), .ZN(n19944) );
  AOI222_X1 U21949 ( .A1(n19940), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(n19944), .ZN(n19910) );
  INV_X1 U21950 ( .A(n19910), .ZN(P1_U3198) );
  AOI222_X1 U21951 ( .A1(n19940), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n19944), .ZN(n19911) );
  INV_X1 U21952 ( .A(n19911), .ZN(P1_U3199) );
  AOI22_X1 U21953 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19940), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n19938), .ZN(n19912) );
  OAI21_X1 U21954 ( .B1(n21376), .B2(n19942), .A(n19912), .ZN(P1_U3200) );
  AOI22_X1 U21955 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19944), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n19938), .ZN(n19913) );
  OAI21_X1 U21956 ( .B1(n21401), .B2(n19946), .A(n19913), .ZN(P1_U3201) );
  AOI222_X1 U21957 ( .A1(n19940), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n19944), .ZN(n19914) );
  INV_X1 U21958 ( .A(n19914), .ZN(P1_U3202) );
  INV_X1 U21959 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21410) );
  AOI22_X1 U21960 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19940), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n19938), .ZN(n19915) );
  OAI21_X1 U21961 ( .B1(n21410), .B2(n19942), .A(n19915), .ZN(P1_U3203) );
  AOI22_X1 U21962 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19944), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n19938), .ZN(n19916) );
  OAI21_X1 U21963 ( .B1(n21431), .B2(n19946), .A(n19916), .ZN(P1_U3204) );
  AOI222_X1 U21964 ( .A1(n19940), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n19944), .ZN(n19917) );
  INV_X1 U21965 ( .A(n19917), .ZN(P1_U3205) );
  AOI222_X1 U21966 ( .A1(n19940), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n19944), .ZN(n19918) );
  INV_X1 U21967 ( .A(n19918), .ZN(P1_U3206) );
  AOI222_X1 U21968 ( .A1(n19940), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n19944), .ZN(n19919) );
  INV_X1 U21969 ( .A(n19919), .ZN(P1_U3207) );
  AOI222_X1 U21970 ( .A1(n19940), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n19944), .ZN(n19920) );
  INV_X1 U21971 ( .A(n19920), .ZN(P1_U3208) );
  AOI22_X1 U21972 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n19940), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n19938), .ZN(n19921) );
  OAI21_X1 U21973 ( .B1(n19922), .B2(n19942), .A(n19921), .ZN(P1_U3209) );
  AOI22_X1 U21974 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n19944), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n19938), .ZN(n19923) );
  OAI21_X1 U21975 ( .B1(n21474), .B2(n19946), .A(n19923), .ZN(P1_U3210) );
  AOI22_X1 U21976 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n19940), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n19938), .ZN(n19924) );
  OAI21_X1 U21977 ( .B1(n21474), .B2(n19942), .A(n19924), .ZN(P1_U3211) );
  AOI22_X1 U21978 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n19944), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n22329), .ZN(n19925) );
  OAI21_X1 U21979 ( .B1(n19927), .B2(n19946), .A(n19925), .ZN(P1_U3212) );
  AOI22_X1 U21980 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n19940), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n22329), .ZN(n19926) );
  OAI21_X1 U21981 ( .B1(n19927), .B2(n19942), .A(n19926), .ZN(P1_U3213) );
  AOI22_X1 U21982 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n19944), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n22329), .ZN(n19928) );
  OAI21_X1 U21983 ( .B1(n21487), .B2(n19946), .A(n19928), .ZN(P1_U3214) );
  AOI222_X1 U21984 ( .A1(n19944), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n19940), .ZN(n19929) );
  INV_X1 U21985 ( .A(n19929), .ZN(P1_U3215) );
  AOI222_X1 U21986 ( .A1(n19940), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n19944), .ZN(n19930) );
  INV_X1 U21987 ( .A(n19930), .ZN(P1_U3216) );
  AOI222_X1 U21988 ( .A1(n19940), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n19944), .ZN(n19931) );
  INV_X1 U21989 ( .A(n19931), .ZN(P1_U3217) );
  AOI222_X1 U21990 ( .A1(n19944), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n19940), .ZN(n19932) );
  INV_X1 U21991 ( .A(n19932), .ZN(P1_U3218) );
  AOI222_X1 U21992 ( .A1(n19944), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n19940), .ZN(n19933) );
  INV_X1 U21993 ( .A(n19933), .ZN(P1_U3219) );
  AOI222_X1 U21994 ( .A1(n19944), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n19940), .ZN(n19934) );
  INV_X1 U21995 ( .A(n19934), .ZN(P1_U3220) );
  AOI222_X1 U21996 ( .A1(n19944), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n19940), .ZN(n19935) );
  INV_X1 U21997 ( .A(n19935), .ZN(P1_U3221) );
  AOI222_X1 U21998 ( .A1(n19944), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n19940), .ZN(n19936) );
  INV_X1 U21999 ( .A(n19936), .ZN(P1_U3222) );
  AOI222_X1 U22000 ( .A1(n19940), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n19944), .ZN(n19937) );
  INV_X1 U22001 ( .A(n19937), .ZN(P1_U3223) );
  AOI222_X1 U22002 ( .A1(n19944), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n19938), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n19940), .ZN(n19939) );
  INV_X1 U22003 ( .A(n19939), .ZN(P1_U3224) );
  AOI22_X1 U22004 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n19940), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n22329), .ZN(n19941) );
  OAI21_X1 U22005 ( .B1(n19943), .B2(n19942), .A(n19941), .ZN(P1_U3225) );
  AOI22_X1 U22006 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n19944), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n22329), .ZN(n19945) );
  OAI21_X1 U22007 ( .B1(n19947), .B2(n19946), .A(n19945), .ZN(P1_U3226) );
  OAI22_X1 U22008 ( .A1(n22329), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22328), .ZN(n19948) );
  INV_X1 U22009 ( .A(n19948), .ZN(P1_U3458) );
  AOI221_X1 U22010 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19959) );
  NOR4_X1 U22011 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19952) );
  NOR4_X1 U22012 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19951) );
  NOR4_X1 U22013 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19950) );
  NOR4_X1 U22014 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19949) );
  NAND4_X1 U22015 ( .A1(n19952), .A2(n19951), .A3(n19950), .A4(n19949), .ZN(
        n19958) );
  NOR4_X1 U22016 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19956) );
  AOI211_X1 U22017 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19955) );
  NOR4_X1 U22018 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19954) );
  NOR4_X1 U22019 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19953) );
  NAND4_X1 U22020 ( .A1(n19956), .A2(n19955), .A3(n19954), .A4(n19953), .ZN(
        n19957) );
  NOR2_X1 U22021 ( .A1(n19958), .A2(n19957), .ZN(n19971) );
  MUX2_X1 U22022 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(n19959), .S(n19971), 
        .Z(P1_U2808) );
  OAI22_X1 U22023 ( .A1(n22329), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22328), .ZN(n19960) );
  INV_X1 U22024 ( .A(n19960), .ZN(P1_U3459) );
  AOI21_X1 U22025 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19961) );
  OAI221_X1 U22026 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19961), .C1(n15268), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n19971), .ZN(n19962) );
  OAI21_X1 U22027 ( .B1(n19971), .B2(n19963), .A(n19962), .ZN(P1_U3481) );
  OAI22_X1 U22028 ( .A1(n22329), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22328), .ZN(n19964) );
  INV_X1 U22029 ( .A(n19964), .ZN(P1_U3460) );
  INV_X1 U22030 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19967) );
  NOR3_X1 U22031 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19965) );
  OAI21_X1 U22032 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19965), .A(n19971), .ZN(
        n19966) );
  OAI21_X1 U22033 ( .B1(n19971), .B2(n19967), .A(n19966), .ZN(P1_U2807) );
  OAI22_X1 U22034 ( .A1(n22329), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22328), .ZN(n19968) );
  INV_X1 U22035 ( .A(n19968), .ZN(P1_U3461) );
  OAI21_X1 U22036 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n19971), .ZN(n19969) );
  OAI21_X1 U22037 ( .B1(n19971), .B2(n19970), .A(n19969), .ZN(P1_U3482) );
  INV_X1 U22038 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n21398) );
  NAND2_X1 U22039 ( .A1(n19973), .A2(n19972), .ZN(n19974) );
  AND2_X1 U22040 ( .A1(n19975), .A2(n19974), .ZN(n21400) );
  AOI22_X1 U22041 ( .A1(n21405), .A2(n19986), .B1(n19985), .B2(n21400), .ZN(
        n19976) );
  OAI21_X1 U22042 ( .B1(n19989), .B2(n21398), .A(n19976), .ZN(P1_U2866) );
  INV_X1 U22043 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n19978) );
  INV_X1 U22044 ( .A(n21464), .ZN(n20023) );
  AOI22_X1 U22045 ( .A1(n20023), .A2(n19986), .B1(n19985), .B2(n21455), .ZN(
        n19977) );
  OAI21_X1 U22046 ( .B1(n19989), .B2(n19978), .A(n19977), .ZN(P1_U2860) );
  INV_X1 U22047 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n19983) );
  INV_X1 U22048 ( .A(n21438), .ZN(n19980) );
  OAI22_X1 U22049 ( .A1(n21440), .A2(n15965), .B1(n19980), .B2(n19979), .ZN(
        n19981) );
  INV_X1 U22050 ( .A(n19981), .ZN(n19982) );
  OAI21_X1 U22051 ( .B1(n19989), .B2(n19983), .A(n19982), .ZN(P1_U2862) );
  AOI22_X1 U22052 ( .A1(n20034), .A2(n19986), .B1(n19985), .B2(n19984), .ZN(
        n19987) );
  OAI21_X1 U22053 ( .B1(n19989), .B2(n19988), .A(n19987), .ZN(P1_U2855) );
  AOI22_X1 U22054 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20038), .B1(
        n21348), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19995) );
  OAI21_X1 U22055 ( .B1(n19990), .B2(n19992), .A(n19991), .ZN(n19993) );
  INV_X1 U22056 ( .A(n19993), .ZN(n21308) );
  AOI22_X1 U22057 ( .A1(n21308), .A2(n20039), .B1(n21732), .B2(n21379), .ZN(
        n19994) );
  OAI211_X1 U22058 ( .C1(n21382), .C2(n20043), .A(n19995), .B(n19994), .ZN(
        P1_U2995) );
  AOI22_X1 U22059 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20038), .B1(
        n21348), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n20001) );
  OAI21_X1 U22060 ( .B1(n19996), .B2(n19998), .A(n19997), .ZN(n19999) );
  INV_X1 U22061 ( .A(n19999), .ZN(n21326) );
  AOI22_X1 U22062 ( .A1(n21326), .A2(n20039), .B1(n21732), .B2(n21393), .ZN(
        n20000) );
  OAI211_X1 U22063 ( .C1(n21396), .C2(n20043), .A(n20001), .B(n20000), .ZN(
        P1_U2994) );
  AOI22_X1 U22064 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20038), .B1(
        n21348), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n20007) );
  NAND2_X1 U22065 ( .A1(n20003), .A2(n20004), .ZN(n20005) );
  NAND2_X1 U22066 ( .A1(n10999), .A2(n20005), .ZN(n21320) );
  AOI22_X1 U22067 ( .A1(n21320), .A2(n20039), .B1(n21732), .B2(n21405), .ZN(
        n20006) );
  OAI211_X1 U22068 ( .C1(n21408), .C2(n20043), .A(n20007), .B(n20006), .ZN(
        P1_U2993) );
  AOI22_X1 U22069 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20038), .B1(
        n21348), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n20013) );
  AOI21_X1 U22070 ( .B1(n20010), .B2(n20008), .A(n11007), .ZN(n21333) );
  AOI22_X1 U22071 ( .A1(n21333), .A2(n20039), .B1(n21732), .B2(n20011), .ZN(
        n20012) );
  OAI211_X1 U22072 ( .C1(n21420), .C2(n20043), .A(n20013), .B(n20012), .ZN(
        P1_U2992) );
  AOI22_X1 U22073 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20038), .B1(
        n21348), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n20016) );
  OAI22_X1 U22074 ( .A1(n21440), .A2(n20022), .B1(n21439), .B2(n20043), .ZN(
        n20014) );
  INV_X1 U22075 ( .A(n20014), .ZN(n20015) );
  OAI211_X1 U22076 ( .C1(n21574), .C2(n20017), .A(n20016), .B(n20015), .ZN(
        P1_U2989) );
  OAI22_X1 U22077 ( .A1(n20018), .A2(n21574), .B1(n21448), .B2(n20043), .ZN(
        n20019) );
  OAI21_X1 U22078 ( .B1(n20022), .B2(n21447), .A(n20021), .ZN(P1_U2988) );
  AOI22_X1 U22079 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20038), .B1(
        n21348), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n20025) );
  AOI22_X1 U22080 ( .A1(n21461), .A2(n20033), .B1(n21732), .B2(n20023), .ZN(
        n20024) );
  OAI211_X1 U22081 ( .C1(n20026), .C2(n21574), .A(n20025), .B(n20024), .ZN(
        P1_U2987) );
  XNOR2_X1 U22082 ( .A(n13755), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n20027) );
  XNOR2_X1 U22083 ( .A(n20028), .B(n20027), .ZN(n21340) );
  AOI22_X1 U22084 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20038), .B1(
        n21348), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n20031) );
  AOI22_X1 U22085 ( .A1(n21471), .A2(n21732), .B1(n20033), .B2(n20029), .ZN(
        n20030) );
  OAI211_X1 U22086 ( .C1(n21340), .C2(n21574), .A(n20031), .B(n20030), .ZN(
        P1_U2984) );
  AOI22_X1 U22087 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20038), .B1(
        n21348), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n20036) );
  AOI22_X1 U22088 ( .A1(n20034), .A2(n21732), .B1(n20033), .B2(n20032), .ZN(
        n20035) );
  OAI211_X1 U22089 ( .C1(n20037), .C2(n21574), .A(n20036), .B(n20035), .ZN(
        P1_U2982) );
  AOI22_X1 U22090 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n20038), .B1(
        n21348), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n20042) );
  AOI22_X1 U22091 ( .A1(n20040), .A2(n20039), .B1(n21732), .B2(n21499), .ZN(
        n20041) );
  OAI211_X1 U22092 ( .C1(n21491), .C2(n20043), .A(n20042), .B(n20041), .ZN(
        P1_U2980) );
  OAI21_X1 U22093 ( .B1(n20044), .B2(n21592), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20045) );
  OAI21_X1 U22094 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20046), .A(n20045), 
        .ZN(P1_U2803) );
  OAI21_X1 U22095 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21611), .A(n21614), 
        .ZN(n20047) );
  AOI22_X1 U22096 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n22328), .B1(n20048), 
        .B2(n20047), .ZN(P1_U2804) );
  AOI22_X1 U22097 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n20086), .ZN(n20050) );
  OAI21_X1 U22098 ( .B1(n14885), .B2(n20098), .A(n20050), .ZN(U247) );
  INV_X1 U22099 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20052) );
  AOI22_X1 U22100 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n20086), .ZN(n20051) );
  OAI21_X1 U22101 ( .B1(n20052), .B2(n20098), .A(n20051), .ZN(U246) );
  AOI22_X1 U22102 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n20086), .ZN(n20053) );
  OAI21_X1 U22103 ( .B1(n14891), .B2(n20098), .A(n20053), .ZN(U245) );
  INV_X1 U22104 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20055) );
  AOI22_X1 U22105 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n20086), .ZN(n20054) );
  OAI21_X1 U22106 ( .B1(n20055), .B2(n20098), .A(n20054), .ZN(U244) );
  INV_X1 U22107 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20057) );
  AOI22_X1 U22108 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n20086), .ZN(n20056) );
  OAI21_X1 U22109 ( .B1(n20057), .B2(n20098), .A(n20056), .ZN(U243) );
  INV_X1 U22110 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20059) );
  AOI22_X1 U22111 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n20086), .ZN(n20058) );
  OAI21_X1 U22112 ( .B1(n20059), .B2(n20098), .A(n20058), .ZN(U242) );
  INV_X1 U22113 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20061) );
  AOI22_X1 U22114 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n20086), .ZN(n20060) );
  OAI21_X1 U22115 ( .B1(n20061), .B2(n20098), .A(n20060), .ZN(U241) );
  INV_X1 U22116 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20063) );
  AOI22_X1 U22117 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n20086), .ZN(n20062) );
  OAI21_X1 U22118 ( .B1(n20063), .B2(n20098), .A(n20062), .ZN(U240) );
  INV_X1 U22119 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20065) );
  AOI22_X1 U22120 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n20086), .ZN(n20064) );
  OAI21_X1 U22121 ( .B1(n20065), .B2(n20098), .A(n20064), .ZN(U239) );
  AOI22_X1 U22122 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n20086), .ZN(n20066) );
  OAI21_X1 U22123 ( .B1(n20067), .B2(n20098), .A(n20066), .ZN(U238) );
  INV_X1 U22124 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20069) );
  AOI22_X1 U22125 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n20086), .ZN(n20068) );
  OAI21_X1 U22126 ( .B1(n20069), .B2(n20098), .A(n20068), .ZN(U237) );
  AOI22_X1 U22127 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n20086), .ZN(n20070) );
  OAI21_X1 U22128 ( .B1(n20071), .B2(n20098), .A(n20070), .ZN(U236) );
  INV_X1 U22129 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20073) );
  AOI22_X1 U22130 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n20086), .ZN(n20072) );
  OAI21_X1 U22131 ( .B1(n20073), .B2(n20098), .A(n20072), .ZN(U235) );
  AOI22_X1 U22132 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n20086), .ZN(n20074) );
  OAI21_X1 U22133 ( .B1(n20075), .B2(n20098), .A(n20074), .ZN(U234) );
  AOI22_X1 U22134 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n20095), .ZN(n20076) );
  OAI21_X1 U22135 ( .B1(n20077), .B2(n20098), .A(n20076), .ZN(U233) );
  AOI22_X1 U22136 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n20086), .ZN(n20078) );
  OAI21_X1 U22137 ( .B1(n16035), .B2(n20098), .A(n20078), .ZN(U232) );
  AOI22_X1 U22138 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n20095), .ZN(n20079) );
  OAI21_X1 U22139 ( .B1(n21747), .B2(n20098), .A(n20079), .ZN(U231) );
  INV_X1 U22140 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n21937) );
  AOI22_X1 U22141 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n20086), .ZN(n20080) );
  OAI21_X1 U22142 ( .B1(n21937), .B2(n20098), .A(n20080), .ZN(U230) );
  INV_X1 U22143 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n21979) );
  AOI22_X1 U22144 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n20086), .ZN(n20081) );
  OAI21_X1 U22145 ( .B1(n21979), .B2(n20098), .A(n20081), .ZN(U229) );
  INV_X1 U22146 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n22027) );
  AOI22_X1 U22147 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n20095), .ZN(n20082) );
  OAI21_X1 U22148 ( .B1(n22027), .B2(n20098), .A(n20082), .ZN(U228) );
  INV_X1 U22149 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n22072) );
  AOI22_X1 U22150 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n20086), .ZN(n20083) );
  OAI21_X1 U22151 ( .B1(n22072), .B2(n20098), .A(n20083), .ZN(U227) );
  AOI22_X1 U22152 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n20095), .ZN(n20084) );
  OAI21_X1 U22153 ( .B1(n22119), .B2(n20098), .A(n20084), .ZN(U226) );
  INV_X1 U22154 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n22169) );
  AOI22_X1 U22155 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n20086), .ZN(n20085) );
  OAI21_X1 U22156 ( .B1(n22169), .B2(n20098), .A(n20085), .ZN(U225) );
  INV_X1 U22157 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n22220) );
  AOI22_X1 U22158 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n20086), .ZN(n20087) );
  OAI21_X1 U22159 ( .B1(n22220), .B2(n20098), .A(n20087), .ZN(U224) );
  INV_X1 U22160 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n21734) );
  AOI22_X1 U22161 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n20095), .ZN(n20088) );
  OAI21_X1 U22162 ( .B1(n21734), .B2(n20098), .A(n20088), .ZN(U223) );
  AOI22_X1 U22163 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n20095), .ZN(n20089) );
  OAI21_X1 U22164 ( .B1(n16549), .B2(n20098), .A(n20089), .ZN(U222) );
  INV_X1 U22165 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n21978) );
  AOI22_X1 U22166 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n20095), .ZN(n20091) );
  OAI21_X1 U22167 ( .B1(n21978), .B2(n20098), .A(n20091), .ZN(U221) );
  INV_X1 U22168 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n22024) );
  AOI22_X1 U22169 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n20095), .ZN(n20092) );
  OAI21_X1 U22170 ( .B1(n22024), .B2(n20098), .A(n20092), .ZN(U220) );
  INV_X1 U22171 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n22070) );
  AOI22_X1 U22172 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n20095), .ZN(n20093) );
  OAI21_X1 U22173 ( .B1(n22070), .B2(n20098), .A(n20093), .ZN(U219) );
  INV_X1 U22174 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n22116) );
  AOI22_X1 U22175 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n20095), .ZN(n20094) );
  OAI21_X1 U22176 ( .B1(n22116), .B2(n20098), .A(n20094), .ZN(U218) );
  AOI22_X1 U22177 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20090), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n20095), .ZN(n20096) );
  OAI21_X1 U22178 ( .B1(n22166), .B2(n20098), .A(n20096), .ZN(U217) );
  OAI222_X1 U22179 ( .A1(U212), .A2(n20099), .B1(n20098), .B2(n22214), .C1(
        U214), .C2(n20097), .ZN(U216) );
  AOI22_X1 U22180 ( .A1(n22328), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20100), 
        .B2(n22329), .ZN(P1_U3483) );
  OAI21_X1 U22181 ( .B1(n21607), .B2(n20102), .A(n20101), .ZN(n20103) );
  AOI21_X1 U22182 ( .B1(n20104), .B2(n21256), .A(n20103), .ZN(n20112) );
  AOI21_X1 U22183 ( .B1(n20106), .B2(n21602), .A(n20105), .ZN(n20107) );
  OAI211_X1 U22184 ( .C1(n20108), .C2(n20107), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n21652), .ZN(n20109) );
  AOI21_X1 U22185 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20109), .A(n21248), 
        .ZN(n20111) );
  NAND2_X1 U22186 ( .A1(n20112), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20110) );
  OAI21_X1 U22187 ( .B1(n20112), .B2(n20111), .A(n20110), .ZN(P3_U3296) );
  AOI22_X1 U22188 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20130), .ZN(n20116) );
  OAI21_X1 U22189 ( .B1(n20749), .B2(n20166), .A(n20116), .ZN(P3_U2768) );
  AOI22_X1 U22190 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20130), .ZN(n20117) );
  OAI21_X1 U22191 ( .B1(n20118), .B2(n20166), .A(n20117), .ZN(P3_U2769) );
  AOI22_X1 U22192 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20130), .ZN(n20119) );
  OAI21_X1 U22193 ( .B1(n20120), .B2(n20166), .A(n20119), .ZN(P3_U2770) );
  AOI22_X1 U22194 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20130), .ZN(n20121) );
  OAI21_X1 U22195 ( .B1(n20676), .B2(n20166), .A(n20121), .ZN(P3_U2771) );
  AOI22_X1 U22196 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20130), .ZN(n20122) );
  OAI21_X1 U22197 ( .B1(n20123), .B2(n20166), .A(n20122), .ZN(P3_U2772) );
  AOI22_X1 U22198 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20130), .ZN(n20124) );
  OAI21_X1 U22199 ( .B1(n20125), .B2(n20166), .A(n20124), .ZN(P3_U2773) );
  AOI22_X1 U22200 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20130), .ZN(n20126) );
  OAI21_X1 U22201 ( .B1(n20671), .B2(n20166), .A(n20126), .ZN(P3_U2774) );
  AOI22_X1 U22202 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20130), .ZN(n20127) );
  OAI21_X1 U22203 ( .B1(n20736), .B2(n20166), .A(n20127), .ZN(P3_U2775) );
  AOI22_X1 U22204 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20130), .ZN(n20128) );
  OAI21_X1 U22205 ( .B1(n20729), .B2(n20166), .A(n20128), .ZN(P3_U2776) );
  AOI22_X1 U22206 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20130), .ZN(n20129) );
  OAI21_X1 U22207 ( .B1(n20691), .B2(n20166), .A(n20129), .ZN(P3_U2777) );
  AOI22_X1 U22208 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20163), .ZN(n20131) );
  OAI21_X1 U22209 ( .B1(n20132), .B2(n20166), .A(n20131), .ZN(P3_U2778) );
  AOI22_X1 U22210 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20163), .ZN(n20133) );
  OAI21_X1 U22211 ( .B1(n20134), .B2(n20166), .A(n20133), .ZN(P3_U2779) );
  AOI22_X1 U22212 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20164), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20163), .ZN(n20135) );
  OAI21_X1 U22213 ( .B1(n20717), .B2(n20166), .A(n20135), .ZN(P3_U2780) );
  AOI22_X1 U22214 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20149), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20163), .ZN(n20136) );
  OAI21_X1 U22215 ( .B1(n20137), .B2(n20166), .A(n20136), .ZN(P3_U2781) );
  AOI22_X1 U22216 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20149), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20163), .ZN(n20138) );
  OAI21_X1 U22217 ( .B1(n20711), .B2(n20166), .A(n20138), .ZN(P3_U2782) );
  AOI22_X1 U22218 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20149), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20163), .ZN(n20139) );
  OAI21_X1 U22219 ( .B1(n20785), .B2(n20166), .A(n20139), .ZN(P3_U2783) );
  AOI22_X1 U22220 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20149), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20163), .ZN(n20140) );
  OAI21_X1 U22221 ( .B1(n20141), .B2(n20166), .A(n20140), .ZN(P3_U2784) );
  AOI22_X1 U22222 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20149), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20163), .ZN(n20142) );
  OAI21_X1 U22223 ( .B1(n20648), .B2(n20166), .A(n20142), .ZN(P3_U2785) );
  AOI22_X1 U22224 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20149), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20163), .ZN(n20143) );
  OAI21_X1 U22225 ( .B1(n20144), .B2(n20166), .A(n20143), .ZN(P3_U2786) );
  AOI22_X1 U22226 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20149), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20163), .ZN(n20145) );
  OAI21_X1 U22227 ( .B1(n20623), .B2(n20166), .A(n20145), .ZN(P3_U2787) );
  AOI22_X1 U22228 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20149), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20163), .ZN(n20146) );
  OAI21_X1 U22229 ( .B1(n20147), .B2(n20166), .A(n20146), .ZN(P3_U2788) );
  AOI22_X1 U22230 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20149), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20163), .ZN(n20148) );
  OAI21_X1 U22231 ( .B1(n20624), .B2(n20166), .A(n20148), .ZN(P3_U2789) );
  AOI22_X1 U22232 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20149), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20163), .ZN(n20150) );
  OAI21_X1 U22233 ( .B1(n20151), .B2(n20166), .A(n20150), .ZN(P3_U2790) );
  AOI22_X1 U22234 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20164), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20163), .ZN(n20152) );
  OAI21_X1 U22235 ( .B1(n20772), .B2(n20166), .A(n20152), .ZN(P3_U2791) );
  AOI22_X1 U22236 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20164), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20163), .ZN(n20153) );
  OAI21_X1 U22237 ( .B1(n20154), .B2(n20166), .A(n20153), .ZN(P3_U2792) );
  AOI22_X1 U22238 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20164), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20163), .ZN(n20155) );
  OAI21_X1 U22239 ( .B1(n20156), .B2(n20166), .A(n20155), .ZN(P3_U2793) );
  AOI22_X1 U22240 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20164), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20163), .ZN(n20157) );
  OAI21_X1 U22241 ( .B1(n20611), .B2(n20166), .A(n20157), .ZN(P3_U2794) );
  AOI22_X1 U22242 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20164), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20163), .ZN(n20158) );
  OAI21_X1 U22243 ( .B1(n20159), .B2(n20166), .A(n20158), .ZN(P3_U2795) );
  AOI22_X1 U22244 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20164), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20163), .ZN(n20160) );
  OAI21_X1 U22245 ( .B1(n20161), .B2(n20166), .A(n20160), .ZN(P3_U2796) );
  AOI22_X1 U22246 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20164), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20163), .ZN(n20162) );
  OAI21_X1 U22247 ( .B1(n20758), .B2(n20166), .A(n20162), .ZN(P3_U2797) );
  AOI22_X1 U22248 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20164), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20163), .ZN(n20165) );
  OAI21_X1 U22249 ( .B1(n20167), .B2(n20166), .A(n20165), .ZN(P3_U2798) );
  INV_X1 U22250 ( .A(n14557), .ZN(n20816) );
  OAI21_X1 U22251 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20816), .A(
        n20822), .ZN(n20805) );
  OAI22_X1 U22252 ( .A1(n20168), .A2(n20586), .B1(n20805), .B2(n20197), .ZN(
        n20175) );
  NOR2_X1 U22253 ( .A1(n21243), .A2(n20523), .ZN(n20301) );
  INV_X1 U22254 ( .A(n20301), .ZN(n20352) );
  NOR2_X1 U22255 ( .A1(n20169), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20195) );
  AOI21_X1 U22256 ( .B1(n20229), .B2(n20170), .A(n20556), .ZN(n20182) );
  OAI211_X1 U22257 ( .C1(n20195), .C2(n20173), .A(n20561), .B(n20182), .ZN(
        n20172) );
  NAND2_X1 U22258 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20185) );
  OAI211_X1 U22259 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20445), .B(n20185), .ZN(n20171) );
  OAI211_X1 U22260 ( .C1(n20352), .C2(n20173), .A(n20172), .B(n20171), .ZN(
        n20174) );
  AOI211_X1 U22261 ( .C1(n20588), .C2(P3_EBX_REG_2__SCAN_IN), .A(n20175), .B(
        n20174), .ZN(n20179) );
  NOR3_X1 U22262 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20190) );
  AOI211_X1 U22263 ( .C1(n20176), .C2(P3_EBX_REG_2__SCAN_IN), .A(n20564), .B(
        n20190), .ZN(n20177) );
  INV_X1 U22264 ( .A(n20177), .ZN(n20178) );
  OAI211_X1 U22265 ( .C1(n20582), .C2(n20180), .A(n20179), .B(n20178), .ZN(
        P3_U2669) );
  AOI21_X1 U22266 ( .B1(n11427), .B2(n20822), .A(n17832), .ZN(n20830) );
  INV_X1 U22267 ( .A(n20830), .ZN(n20193) );
  NAND3_X1 U22268 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n20211) );
  NAND2_X1 U22269 ( .A1(n20445), .A2(n20211), .ZN(n20184) );
  NAND2_X1 U22270 ( .A1(n20586), .A2(n20184), .ZN(n20204) );
  OAI22_X1 U22271 ( .A1(n20181), .A2(n20582), .B1(n20516), .B2(n20189), .ZN(
        n20188) );
  XOR2_X1 U22272 ( .A(n20183), .B(n20182), .Z(n20186) );
  OAI22_X1 U22273 ( .A1(n21243), .A2(n20186), .B1(n20185), .B2(n20184), .ZN(
        n20187) );
  AOI211_X1 U22274 ( .C1(P3_REIP_REG_3__SCAN_IN), .C2(n20204), .A(n20188), .B(
        n20187), .ZN(n20192) );
  NAND2_X1 U22275 ( .A1(n20190), .A2(n20189), .ZN(n20194) );
  OAI211_X1 U22276 ( .C1(n20190), .C2(n20189), .A(n20587), .B(n20194), .ZN(
        n20191) );
  OAI211_X1 U22277 ( .C1(n20193), .C2(n20197), .A(n20192), .B(n20191), .ZN(
        P3_U2668) );
  NOR2_X1 U22278 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20194), .ZN(n20222) );
  AOI211_X1 U22279 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20194), .A(n20222), .B(
        n20564), .ZN(n20210) );
  INV_X1 U22280 ( .A(n20195), .ZN(n20429) );
  OAI21_X1 U22281 ( .B1(n20196), .B2(n20429), .A(n20523), .ZN(n20213) );
  NOR3_X1 U22282 ( .A1(n20199), .A2(n21243), .A3(n20213), .ZN(n20209) );
  AOI21_X1 U22283 ( .B1(n11506), .B2(n20198), .A(n20197), .ZN(n20203) );
  OAI21_X1 U22284 ( .B1(n20200), .B2(n20556), .A(n20199), .ZN(n20201) );
  OAI22_X1 U22285 ( .A1(n20324), .A2(n20201), .B1(n20200), .B2(n20582), .ZN(
        n20202) );
  AOI211_X1 U22286 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n20204), .A(n20203), .B(
        n20202), .ZN(n20206) );
  OR3_X1 U22287 ( .A1(n20450), .A2(n20211), .A3(P3_REIP_REG_4__SCAN_IN), .ZN(
        n20205) );
  OAI211_X1 U22288 ( .C1(n20207), .C2(n20516), .A(n20206), .B(n20205), .ZN(
        n20208) );
  OR4_X1 U22289 ( .A1(n10979), .A2(n20210), .A3(n20209), .A4(n20208), .ZN(
        P3_U2667) );
  NOR2_X1 U22290 ( .A1(n20890), .A2(n20211), .ZN(n20212) );
  NAND2_X1 U22291 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n20212), .ZN(n20252) );
  AOI21_X1 U22292 ( .B1(n20445), .B2(n20252), .A(n20461), .ZN(n20246) );
  NAND3_X1 U22293 ( .A1(n20212), .A2(n20445), .A3(n20252), .ZN(n20218) );
  INV_X1 U22294 ( .A(n20214), .ZN(n20216) );
  INV_X1 U22295 ( .A(n20213), .ZN(n20215) );
  OAI221_X1 U22296 ( .B1(n20216), .B2(n20215), .C1(n20214), .C2(n20213), .A(
        n20561), .ZN(n20217) );
  OAI211_X1 U22297 ( .C1(n20246), .C2(n20219), .A(n20218), .B(n20217), .ZN(
        n20220) );
  AOI211_X1 U22298 ( .C1(n20588), .C2(P3_EBX_REG_5__SCAN_IN), .A(n10979), .B(
        n20220), .ZN(n20224) );
  INV_X1 U22299 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20221) );
  NAND2_X1 U22300 ( .A1(n20222), .A2(n20221), .ZN(n20226) );
  OAI211_X1 U22301 ( .C1(n20222), .C2(n20221), .A(n20587), .B(n20226), .ZN(
        n20223) );
  OAI211_X1 U22302 ( .C1(n20582), .C2(n20225), .A(n20224), .B(n20223), .ZN(
        P3_U2666) );
  NOR2_X1 U22303 ( .A1(n20450), .A2(n20252), .ZN(n20239) );
  INV_X1 U22304 ( .A(n20239), .ZN(n20238) );
  AOI211_X1 U22305 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20226), .A(n20248), .B(
        n20564), .ZN(n20235) );
  NAND2_X1 U22306 ( .A1(n20227), .A2(n20229), .ZN(n20268) );
  NAND2_X1 U22307 ( .A1(n20228), .A2(n20268), .ZN(n20233) );
  NAND2_X1 U22308 ( .A1(n20561), .A2(n20229), .ZN(n20267) );
  OAI21_X1 U22309 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20267), .A(
        n20352), .ZN(n20230) );
  AOI22_X1 U22310 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20532), .B1(
        n20231), .B2(n20230), .ZN(n20232) );
  OAI211_X1 U22311 ( .C1(n20571), .C2(n20233), .A(n20232), .B(n11764), .ZN(
        n20234) );
  AOI211_X1 U22312 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20588), .A(n20235), .B(
        n20234), .ZN(n20236) );
  OAI221_X1 U22313 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n20238), .C1(n20237), 
        .C2(n20246), .A(n20236), .ZN(P3_U2665) );
  NAND2_X1 U22314 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n20253) );
  OAI211_X1 U22315 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n20239), .B(n20253), .ZN(n20244) );
  NAND2_X1 U22316 ( .A1(n11013), .A2(n20268), .ZN(n20241) );
  AOI21_X1 U22317 ( .B1(n20242), .B2(n20241), .A(n21243), .ZN(n20240) );
  OAI21_X1 U22318 ( .B1(n20242), .B2(n20241), .A(n20240), .ZN(n20243) );
  OAI211_X1 U22319 ( .C1(n20246), .C2(n20245), .A(n20244), .B(n20243), .ZN(
        n20247) );
  AOI211_X1 U22320 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n20532), .A(
        n10979), .B(n20247), .ZN(n20250) );
  NAND2_X1 U22321 ( .A1(n20248), .A2(n20251), .ZN(n20254) );
  OAI211_X1 U22322 ( .C1(n20248), .C2(n20251), .A(n20587), .B(n20254), .ZN(
        n20249) );
  OAI211_X1 U22323 ( .C1(n20251), .C2(n20516), .A(n20250), .B(n20249), .ZN(
        P3_U2664) );
  NOR2_X1 U22324 ( .A1(n20253), .A2(n20252), .ZN(n20259) );
  NAND2_X1 U22325 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n20259), .ZN(n20288) );
  AOI21_X1 U22326 ( .B1(n20445), .B2(n20288), .A(n20461), .ZN(n20284) );
  AOI211_X1 U22327 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n20254), .A(n20275), .B(
        n20564), .ZN(n20264) );
  OAI21_X1 U22328 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20255), .A(
        n20523), .ZN(n20256) );
  XNOR2_X1 U22329 ( .A(n20257), .B(n20256), .ZN(n20260) );
  INV_X1 U22330 ( .A(n20288), .ZN(n20273) );
  NOR2_X1 U22331 ( .A1(n20273), .A2(n20450), .ZN(n20258) );
  AOI22_X1 U22332 ( .A1(n20561), .A2(n20260), .B1(n20259), .B2(n20258), .ZN(
        n20261) );
  OAI211_X1 U22333 ( .C1(n20262), .C2(n20582), .A(n20261), .B(n11764), .ZN(
        n20263) );
  AOI211_X1 U22334 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n20588), .A(n20264), .B(
        n20263), .ZN(n20265) );
  OAI21_X1 U22335 ( .B1(n20284), .B2(n20266), .A(n20265), .ZN(P3_U2663) );
  AOI22_X1 U22336 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n20532), .B1(
        n20588), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n20279) );
  OAI21_X1 U22337 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n20267), .A(
        n20352), .ZN(n20271) );
  NOR2_X1 U22338 ( .A1(n20269), .A2(n20268), .ZN(n20297) );
  OAI21_X1 U22339 ( .B1(n20571), .B2(n20297), .A(n20272), .ZN(n20270) );
  OAI21_X1 U22340 ( .B1(n20272), .B2(n20271), .A(n20270), .ZN(n20277) );
  NAND3_X1 U22341 ( .A1(n20445), .A2(n20273), .A3(n20289), .ZN(n20283) );
  NAND2_X1 U22342 ( .A1(n20275), .A2(n20274), .ZN(n20285) );
  OAI211_X1 U22343 ( .C1(n20275), .C2(n20274), .A(n20587), .B(n20285), .ZN(
        n20276) );
  AND4_X1 U22344 ( .A1(n20277), .A2(n11764), .A3(n20283), .A4(n20276), .ZN(
        n20278) );
  OAI211_X1 U22345 ( .C1(n20284), .C2(n20289), .A(n20279), .B(n20278), .ZN(
        P3_U2662) );
  NOR2_X1 U22346 ( .A1(n20297), .A2(n20556), .ZN(n20280) );
  XOR2_X1 U22347 ( .A(n20281), .B(n20280), .Z(n20282) );
  AOI22_X1 U22348 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20532), .B1(
        n20561), .B2(n20282), .ZN(n20293) );
  AOI21_X1 U22349 ( .B1(n20284), .B2(n20283), .A(n20290), .ZN(n20287) );
  AOI211_X1 U22350 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20285), .A(n20306), .B(
        n20564), .ZN(n20286) );
  AOI211_X1 U22351 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20588), .A(n20287), .B(
        n20286), .ZN(n20292) );
  NOR2_X1 U22352 ( .A1(n20289), .A2(n20288), .ZN(n20294) );
  NAND3_X1 U22353 ( .A1(n20445), .A2(n20294), .A3(n20290), .ZN(n20291) );
  NAND4_X1 U22354 ( .A1(n20293), .A2(n20292), .A3(n11764), .A4(n20291), .ZN(
        P3_U2661) );
  NAND2_X1 U22355 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n20294), .ZN(n20296) );
  NOR2_X1 U22356 ( .A1(n20295), .A2(n20296), .ZN(n20382) );
  OAI21_X1 U22357 ( .B1(n20382), .B2(n20450), .A(n20586), .ZN(n20337) );
  NOR2_X1 U22358 ( .A1(n20450), .A2(n20296), .ZN(n20315) );
  NAND2_X1 U22359 ( .A1(n20298), .A2(n20297), .ZN(n20349) );
  NAND2_X1 U22360 ( .A1(n20349), .A2(n20523), .ZN(n20310) );
  INV_X1 U22361 ( .A(n20310), .ZN(n20312) );
  AOI221_X1 U22362 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20302), .C1(
        n20299), .C2(n20302), .A(n21243), .ZN(n20300) );
  OAI22_X1 U22363 ( .A1(n20302), .A2(n20312), .B1(n20301), .B2(n20300), .ZN(
        n20303) );
  OAI211_X1 U22364 ( .C1(n20516), .C2(n20305), .A(n11764), .B(n20303), .ZN(
        n20304) );
  AOI221_X1 U22365 ( .B1(P3_REIP_REG_11__SCAN_IN), .B2(n20337), .C1(n20315), 
        .C2(n20337), .A(n20304), .ZN(n20308) );
  NAND2_X1 U22366 ( .A1(n20306), .A2(n20305), .ZN(n20316) );
  OAI211_X1 U22367 ( .C1(n20306), .C2(n20305), .A(n20587), .B(n20316), .ZN(
        n20307) );
  OAI211_X1 U22368 ( .C1(n20582), .C2(n20309), .A(n20308), .B(n20307), .ZN(
        P3_U2660) );
  INV_X1 U22369 ( .A(n20337), .ZN(n20320) );
  INV_X1 U22370 ( .A(n20311), .ZN(n20313) );
  AOI221_X1 U22371 ( .B1(n20313), .B2(n20312), .C1(n20311), .C2(n20310), .A(
        n21243), .ZN(n20314) );
  AOI211_X1 U22372 ( .C1(n20588), .C2(P3_EBX_REG_12__SCAN_IN), .A(n10979), .B(
        n20314), .ZN(n20319) );
  NAND2_X1 U22373 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n20315), .ZN(n20372) );
  NOR2_X1 U22374 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n20372), .ZN(n20326) );
  AOI211_X1 U22375 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20316), .A(n20332), .B(
        n20564), .ZN(n20317) );
  AOI211_X1 U22376 ( .C1(n20532), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20326), .B(n20317), .ZN(n20318) );
  OAI211_X1 U22377 ( .C1(n20320), .C2(n20321), .A(n20319), .B(n20318), .ZN(
        P3_U2659) );
  NOR2_X1 U22378 ( .A1(n20321), .A2(n20372), .ZN(n20338) );
  OAI21_X1 U22379 ( .B1(n20322), .B2(n20349), .A(n20523), .ZN(n20339) );
  NAND2_X1 U22380 ( .A1(n20561), .A2(n20323), .ZN(n20329) );
  AOI211_X1 U22381 ( .C1(n11013), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20324), .B(n20323), .ZN(n20325) );
  AOI211_X1 U22382 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n20532), .A(
        n10979), .B(n20325), .ZN(n20328) );
  OAI21_X1 U22383 ( .B1(n20326), .B2(n20337), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n20327) );
  OAI211_X1 U22384 ( .C1(n20339), .C2(n20329), .A(n20328), .B(n20327), .ZN(
        n20330) );
  AOI21_X1 U22385 ( .B1(n20338), .B2(n20331), .A(n20330), .ZN(n20334) );
  NAND2_X1 U22386 ( .A1(n20332), .A2(n20335), .ZN(n20336) );
  OAI211_X1 U22387 ( .C1(n20332), .C2(n20335), .A(n20587), .B(n20336), .ZN(
        n20333) );
  OAI211_X1 U22388 ( .C1(n20335), .C2(n20516), .A(n20334), .B(n20333), .ZN(
        P3_U2658) );
  NOR2_X1 U22389 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20336), .ZN(n20354) );
  AOI211_X1 U22390 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20336), .A(n20354), .B(
        n20564), .ZN(n20344) );
  NAND3_X1 U22391 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_14__SCAN_IN), 
        .A3(P3_REIP_REG_12__SCAN_IN), .ZN(n20370) );
  NOR2_X1 U22392 ( .A1(n20445), .A2(n20461), .ZN(n20501) );
  INV_X1 U22393 ( .A(n20501), .ZN(n20585) );
  AOI21_X1 U22394 ( .B1(n20370), .B2(n20585), .A(n20337), .ZN(n20365) );
  AOI21_X1 U22395 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n20338), .A(
        P3_REIP_REG_14__SCAN_IN), .ZN(n20342) );
  XOR2_X1 U22396 ( .A(n20340), .B(n20339), .Z(n20341) );
  OAI22_X1 U22397 ( .A1(n20365), .A2(n20342), .B1(n21243), .B2(n20341), .ZN(
        n20343) );
  AOI211_X1 U22398 ( .C1(n20532), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20344), .B(n20343), .ZN(n20345) );
  OAI211_X1 U22399 ( .C1(n20516), .C2(n20346), .A(n20345), .B(n11764), .ZN(
        P3_U2657) );
  OAI21_X1 U22400 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20347), .A(
        n11013), .ZN(n20361) );
  INV_X1 U22401 ( .A(n20348), .ZN(n20350) );
  NOR2_X1 U22402 ( .A1(n20350), .A2(n20349), .ZN(n20392) );
  OAI21_X1 U22403 ( .B1(n20392), .B2(n20353), .A(n20561), .ZN(n20351) );
  AOI22_X1 U22404 ( .A1(n20353), .A2(n20361), .B1(n20352), .B2(n20351), .ZN(
        n20359) );
  INV_X1 U22405 ( .A(n20354), .ZN(n20355) );
  NOR2_X1 U22406 ( .A1(n20355), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n20366) );
  AOI211_X1 U22407 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n20355), .A(n20366), .B(
        n20564), .ZN(n20358) );
  AOI22_X1 U22408 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20532), .B1(
        n20588), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n20356) );
  INV_X1 U22409 ( .A(n20356), .ZN(n20357) );
  NOR4_X1 U22410 ( .A1(n10979), .A2(n20359), .A3(n20358), .A4(n20357), .ZN(
        n20360) );
  OAI211_X1 U22411 ( .C1(n20365), .C2(n20371), .A(n20360), .B(n20364), .ZN(
        P3_U2656) );
  XNOR2_X1 U22412 ( .A(n20362), .B(n20361), .ZN(n20363) );
  AOI22_X1 U22413 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n20532), .B1(
        n20561), .B2(n20363), .ZN(n20377) );
  AOI21_X1 U22414 ( .B1(n20365), .B2(n20364), .A(n20373), .ZN(n20369) );
  INV_X1 U22415 ( .A(n20366), .ZN(n20367) );
  AOI211_X1 U22416 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20367), .A(n20385), .B(
        n20564), .ZN(n20368) );
  AOI211_X1 U22417 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20588), .A(n20369), .B(
        n20368), .ZN(n20376) );
  NOR2_X1 U22418 ( .A1(n20371), .A2(n20370), .ZN(n20381) );
  INV_X1 U22419 ( .A(n20372), .ZN(n20374) );
  NAND3_X1 U22420 ( .A1(n20381), .A2(n20374), .A3(n20373), .ZN(n20375) );
  NAND4_X1 U22421 ( .A1(n20377), .A2(n20376), .A3(n11764), .A4(n20375), .ZN(
        P3_U2655) );
  INV_X1 U22422 ( .A(n20378), .ZN(n20393) );
  AOI21_X1 U22423 ( .B1(n20393), .B2(n20392), .A(n20556), .ZN(n20380) );
  XNOR2_X1 U22424 ( .A(n20380), .B(n20379), .ZN(n20390) );
  NAND3_X1 U22425 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n20382), .A3(n20381), 
        .ZN(n20383) );
  NOR2_X1 U22426 ( .A1(n20450), .A2(n20383), .ZN(n20391) );
  NOR2_X1 U22427 ( .A1(n21158), .A2(n20383), .ZN(n20422) );
  OAI21_X1 U22428 ( .B1(n20422), .B2(n20450), .A(n20586), .ZN(n20412) );
  OAI21_X1 U22429 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n20391), .A(n20412), 
        .ZN(n20387) );
  NAND2_X1 U22430 ( .A1(n20385), .A2(n20384), .ZN(n20399) );
  OAI211_X1 U22431 ( .C1(n20385), .C2(n20384), .A(n20587), .B(n20399), .ZN(
        n20386) );
  OAI211_X1 U22432 ( .C1(n20582), .C2(n20395), .A(n20387), .B(n20386), .ZN(
        n20388) );
  AOI211_X1 U22433 ( .C1(n20588), .C2(P3_EBX_REG_17__SCAN_IN), .A(n10979), .B(
        n20388), .ZN(n20389) );
  OAI21_X1 U22434 ( .B1(n21243), .B2(n20390), .A(n20389), .ZN(P3_U2654) );
  NAND2_X1 U22435 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n20391), .ZN(n20407) );
  INV_X1 U22436 ( .A(n20412), .ZN(n20406) );
  NAND2_X1 U22437 ( .A1(n20393), .A2(n20392), .ZN(n20394) );
  OAI21_X1 U22438 ( .B1(n20395), .B2(n20394), .A(n20523), .ZN(n20397) );
  OAI21_X1 U22439 ( .B1(n20398), .B2(n20397), .A(n20561), .ZN(n20396) );
  AOI21_X1 U22440 ( .B1(n20398), .B2(n20397), .A(n20396), .ZN(n20404) );
  AOI211_X1 U22441 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20399), .A(n20418), .B(
        n20564), .ZN(n20403) );
  OAI22_X1 U22442 ( .A1(n20401), .A2(n20582), .B1(n20516), .B2(n20400), .ZN(
        n20402) );
  NOR4_X1 U22443 ( .A1(n10979), .A2(n20404), .A3(n20403), .A4(n20402), .ZN(
        n20405) );
  OAI221_X1 U22444 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n20407), .C1(n21152), 
        .C2(n20406), .A(n20405), .ZN(P3_U2653) );
  AOI221_X1 U22445 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n20408), .C2(n21152), .A(n20407), .ZN(n20411) );
  INV_X1 U22446 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20417) );
  OAI22_X1 U22447 ( .A1(n20409), .A2(n20582), .B1(n20516), .B2(n20417), .ZN(
        n20410) );
  AOI211_X1 U22448 ( .C1(n20412), .C2(P3_REIP_REG_19__SCAN_IN), .A(n20411), 
        .B(n20410), .ZN(n20421) );
  OAI21_X1 U22449 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20413), .A(
        n11013), .ZN(n20415) );
  AOI21_X1 U22450 ( .B1(n20416), .B2(n20415), .A(n21243), .ZN(n20414) );
  OAI21_X1 U22451 ( .B1(n20416), .B2(n20415), .A(n20414), .ZN(n20420) );
  NAND2_X1 U22452 ( .A1(n20418), .A2(n20417), .ZN(n20426) );
  OAI211_X1 U22453 ( .C1(n20418), .C2(n20417), .A(n20587), .B(n20426), .ZN(
        n20419) );
  NAND4_X1 U22454 ( .A1(n20421), .A2(n11764), .A3(n20420), .A4(n20419), .ZN(
        P3_U2652) );
  NAND3_X1 U22455 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n20422), .ZN(n20424) );
  NOR2_X1 U22456 ( .A1(n20425), .A2(n20424), .ZN(n20449) );
  OAI21_X1 U22457 ( .B1(n20449), .B2(n20450), .A(n20586), .ZN(n20444) );
  INV_X1 U22458 ( .A(n20444), .ZN(n20423) );
  AOI221_X1 U22459 ( .B1(n20450), .B2(n20425), .C1(n20424), .C2(n20425), .A(
        n20423), .ZN(n20428) );
  AOI211_X1 U22460 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n20426), .A(n20439), .B(
        n20564), .ZN(n20427) );
  AOI211_X1 U22461 ( .C1(n20532), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n20428), .B(n20427), .ZN(n20434) );
  OAI21_X1 U22462 ( .B1(n20430), .B2(n20429), .A(n11012), .ZN(n20431) );
  NAND2_X1 U22463 ( .A1(n20432), .A2(n20431), .ZN(n20436) );
  OAI211_X1 U22464 ( .C1(n20432), .C2(n20431), .A(n20561), .B(n20436), .ZN(
        n20433) );
  OAI211_X1 U22465 ( .C1(n20435), .C2(n20516), .A(n20434), .B(n20433), .ZN(
        P3_U2651) );
  NAND2_X1 U22466 ( .A1(n11013), .A2(n20436), .ZN(n20437) );
  NAND2_X1 U22467 ( .A1(n20438), .A2(n20437), .ZN(n20454) );
  OAI211_X1 U22468 ( .C1(n20438), .C2(n20437), .A(n20561), .B(n20454), .ZN(
        n20441) );
  NAND2_X1 U22469 ( .A1(n20439), .A2(n20448), .ZN(n20451) );
  OAI211_X1 U22470 ( .C1(n20439), .C2(n20448), .A(n20587), .B(n20451), .ZN(
        n20440) );
  OAI211_X1 U22471 ( .C1(n20582), .C2(n20442), .A(n20441), .B(n20440), .ZN(
        n20443) );
  AOI21_X1 U22472 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n20444), .A(n20443), 
        .ZN(n20447) );
  NAND3_X1 U22473 ( .A1(n20445), .A2(n20449), .A3(n20846), .ZN(n20446) );
  OAI211_X1 U22474 ( .C1(n20448), .C2(n20516), .A(n20447), .B(n20446), .ZN(
        P3_U2650) );
  AOI22_X1 U22475 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20532), .B1(
        n20588), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n20459) );
  NAND2_X1 U22476 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n20449), .ZN(n20462) );
  OAI221_X1 U22477 ( .B1(n20450), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n20450), 
        .C2(n20449), .A(n20586), .ZN(n20453) );
  AOI211_X1 U22478 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n20451), .A(n20468), .B(
        n20564), .ZN(n20452) );
  AOI221_X1 U22479 ( .B1(n20460), .B2(n20463), .C1(n20453), .C2(
        P3_REIP_REG_22__SCAN_IN), .A(n20452), .ZN(n20458) );
  OAI211_X1 U22480 ( .C1(n20456), .C2(n20455), .A(n20561), .B(n20464), .ZN(
        n20457) );
  NAND3_X1 U22481 ( .A1(n20459), .A2(n20458), .A3(n20457), .ZN(P3_U2649) );
  NAND2_X1 U22482 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n20460), .ZN(n20473) );
  OR4_X1 U22483 ( .A1(n20463), .A2(n20474), .A3(n20462), .A4(n20461), .ZN(
        n20487) );
  NAND2_X1 U22484 ( .A1(n20585), .A2(n20487), .ZN(n20485) );
  AOI22_X1 U22485 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20532), .B1(
        n20588), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n20471) );
  OAI211_X1 U22486 ( .C1(n20466), .C2(n20465), .A(n20561), .B(n20480), .ZN(
        n20470) );
  INV_X1 U22487 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20467) );
  NAND2_X1 U22488 ( .A1(n20468), .A2(n20467), .ZN(n20475) );
  OAI211_X1 U22489 ( .C1(n20468), .C2(n20467), .A(n20587), .B(n20475), .ZN(
        n20469) );
  AND3_X1 U22490 ( .A1(n20471), .A2(n20470), .A3(n20469), .ZN(n20472) );
  OAI221_X1 U22491 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(n20473), .C1(n20474), 
        .C2(n20485), .A(n20472), .ZN(P3_U2648) );
  AOI211_X1 U22492 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n20475), .A(n20489), .B(
        n20564), .ZN(n20479) );
  OAI22_X1 U22493 ( .A1(n20477), .A2(n20582), .B1(n20516), .B2(n20476), .ZN(
        n20478) );
  AOI211_X1 U22494 ( .C1(n20486), .C2(n20488), .A(n20479), .B(n20478), .ZN(
        n20484) );
  NAND2_X1 U22495 ( .A1(n20523), .A2(n20480), .ZN(n20481) );
  NAND2_X1 U22496 ( .A1(n20482), .A2(n20481), .ZN(n20494) );
  OAI211_X1 U22497 ( .C1(n20482), .C2(n20481), .A(n20561), .B(n20494), .ZN(
        n20483) );
  OAI211_X1 U22498 ( .C1(n20485), .C2(n20488), .A(n20484), .B(n20483), .ZN(
        P3_U2647) );
  NAND2_X1 U22499 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20486), .ZN(n20514) );
  NOR2_X1 U22500 ( .A1(n20488), .A2(n20487), .ZN(n20502) );
  NOR3_X1 U22501 ( .A1(n20501), .A2(n20502), .A3(n20500), .ZN(n20493) );
  NAND2_X1 U22502 ( .A1(n20489), .A2(n20491), .ZN(n20503) );
  OAI211_X1 U22503 ( .C1(n20489), .C2(n20491), .A(n20587), .B(n20503), .ZN(
        n20490) );
  OAI21_X1 U22504 ( .B1(n20491), .B2(n20516), .A(n20490), .ZN(n20492) );
  AOI211_X1 U22505 ( .C1(n20532), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n20493), .B(n20492), .ZN(n20498) );
  NAND2_X1 U22506 ( .A1(n20523), .A2(n20494), .ZN(n20495) );
  NAND2_X1 U22507 ( .A1(n20496), .A2(n20495), .ZN(n20507) );
  OAI211_X1 U22508 ( .C1(n20496), .C2(n20495), .A(n20561), .B(n20507), .ZN(
        n20497) );
  OAI211_X1 U22509 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n20514), .A(n20498), 
        .B(n20497), .ZN(P3_U2646) );
  NAND2_X1 U22510 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n20499), .ZN(n20512) );
  NOR2_X1 U22511 ( .A1(n20500), .A2(n20499), .ZN(n20513) );
  AOI21_X1 U22512 ( .B1(n20513), .B2(n20502), .A(n20501), .ZN(n20547) );
  AOI211_X1 U22513 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20503), .A(n20520), .B(
        n20564), .ZN(n20506) );
  AOI22_X1 U22514 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20532), .B1(
        n20588), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n20504) );
  INV_X1 U22515 ( .A(n20504), .ZN(n20505) );
  AOI211_X1 U22516 ( .C1(n20547), .C2(P3_REIP_REG_26__SCAN_IN), .A(n20506), 
        .B(n20505), .ZN(n20511) );
  NAND2_X1 U22517 ( .A1(n20523), .A2(n20507), .ZN(n20508) );
  OAI211_X1 U22518 ( .C1(n20509), .C2(n20508), .A(n20561), .B(n20522), .ZN(
        n20510) );
  OAI211_X1 U22519 ( .C1(n20512), .C2(n20514), .A(n20511), .B(n20510), .ZN(
        P3_U2645) );
  INV_X1 U22520 ( .A(n20513), .ZN(n20515) );
  INV_X1 U22521 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n20519) );
  OAI22_X1 U22522 ( .A1(n20517), .A2(n20582), .B1(n20516), .B2(n20519), .ZN(
        n20518) );
  AOI221_X1 U22523 ( .B1(n20547), .B2(P3_REIP_REG_27__SCAN_IN), .C1(n20558), 
        .C2(n20529), .A(n20518), .ZN(n20528) );
  NAND2_X1 U22524 ( .A1(n20520), .A2(n20519), .ZN(n20531) );
  OAI211_X1 U22525 ( .C1(n20520), .C2(n20519), .A(n20587), .B(n20531), .ZN(
        n20527) );
  INV_X1 U22526 ( .A(n20521), .ZN(n20525) );
  OAI211_X1 U22527 ( .C1(n20525), .C2(n20524), .A(n20561), .B(n20530), .ZN(
        n20526) );
  NAND3_X1 U22528 ( .A1(n20528), .A2(n20527), .A3(n20526), .ZN(P3_U2644) );
  NAND2_X1 U22529 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n20558), .ZN(n20540) );
  AOI21_X1 U22530 ( .B1(n20558), .B2(n20529), .A(n20547), .ZN(n20538) );
  XOR2_X1 U22531 ( .A(n20544), .B(n20543), .Z(n20536) );
  NOR2_X1 U22532 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n20531), .ZN(n20542) );
  AOI211_X1 U22533 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n20531), .A(n20542), .B(
        n20564), .ZN(n20535) );
  AOI22_X1 U22534 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20532), .B1(
        n20588), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n20533) );
  INV_X1 U22535 ( .A(n20533), .ZN(n20534) );
  AOI211_X1 U22536 ( .C1(n20536), .C2(n20561), .A(n20535), .B(n20534), .ZN(
        n20537) );
  OAI221_X1 U22537 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(n20540), .C1(n20539), 
        .C2(n20538), .A(n20537), .ZN(P3_U2643) );
  INV_X1 U22538 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n20541) );
  NOR2_X1 U22539 ( .A1(n20542), .A2(n20541), .ZN(n20555) );
  NAND2_X1 U22540 ( .A1(n20542), .A2(n20541), .ZN(n20563) );
  NAND2_X1 U22541 ( .A1(n20587), .A2(n20563), .ZN(n20567) );
  OAI21_X1 U22542 ( .B1(n20544), .B2(n20556), .A(n20543), .ZN(n20545) );
  NOR2_X1 U22543 ( .A1(n20546), .A2(n20545), .ZN(n20557) );
  AOI211_X1 U22544 ( .C1(n20546), .C2(n20545), .A(n20557), .B(n21243), .ZN(
        n20551) );
  NAND3_X1 U22545 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n20548) );
  AOI21_X1 U22546 ( .B1(n20548), .B2(n20585), .A(n20547), .ZN(n20577) );
  OAI22_X1 U22547 ( .A1(n20577), .A2(n20552), .B1(n20549), .B2(n20582), .ZN(
        n20550) );
  AOI211_X1 U22548 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n20588), .A(n20551), .B(
        n20550), .ZN(n20554) );
  NAND4_X1 U22549 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n20558), .A4(n20552), .ZN(n20553) );
  OAI211_X1 U22550 ( .C1(n20555), .C2(n20567), .A(n20554), .B(n20553), .ZN(
        P3_U2642) );
  XOR2_X1 U22551 ( .A(n20573), .B(n20572), .Z(n20562) );
  NAND4_X1 U22552 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n20558), .ZN(n20568) );
  NOR2_X1 U22553 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n20568), .ZN(n20574) );
  OAI22_X1 U22554 ( .A1(n20577), .A2(n20569), .B1(n20559), .B2(n20582), .ZN(
        n20560) );
  NOR2_X1 U22555 ( .A1(n20564), .A2(n20563), .ZN(n20580) );
  OAI21_X1 U22556 ( .B1(n20588), .B2(n20580), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n20565) );
  OAI211_X1 U22557 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n20567), .A(n20566), .B(
        n20565), .ZN(P3_U2641) );
  NOR3_X1 U22558 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n20569), .A3(n20568), 
        .ZN(n20570) );
  AOI21_X1 U22559 ( .B1(n20588), .B2(P3_EBX_REG_31__SCAN_IN), .A(n20570), .ZN(
        n20581) );
  INV_X1 U22560 ( .A(n20574), .ZN(n20576) );
  AOI21_X1 U22561 ( .B1(n20577), .B2(n20576), .A(n20575), .ZN(n20578) );
  AOI22_X1 U22562 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n20585), .B1(n20584), 
        .B2(n11421), .ZN(n20591) );
  NAND3_X1 U22563 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20586), .A3(
        n20808), .ZN(n20590) );
  OAI21_X1 U22564 ( .B1(n20588), .B2(n20587), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n20589) );
  NAND3_X1 U22565 ( .A1(n20591), .A2(n20590), .A3(n20589), .ZN(P3_U2671) );
  NAND4_X1 U22566 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n20593) );
  NAND4_X1 U22567 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_7__SCAN_IN), .ZN(n20592) );
  NOR2_X1 U22568 ( .A1(n20593), .A2(n20592), .ZN(n20655) );
  INV_X1 U22569 ( .A(n20655), .ZN(n20767) );
  NAND2_X1 U22570 ( .A1(n20768), .A2(n20621), .ZN(n20784) );
  NAND2_X1 U22571 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20619), .ZN(n20612) );
  NOR2_X1 U22572 ( .A1(n20611), .A2(n20612), .ZN(n20605) );
  NAND2_X1 U22573 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n20605), .ZN(n20604) );
  NAND2_X1 U22574 ( .A1(n20604), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n20603) );
  NOR2_X2 U22575 ( .A1(n20788), .A2(n20775), .ZN(n20781) );
  AOI22_X1 U22576 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20782), .B1(n20781), .B2(
        n20601), .ZN(n20602) );
  OAI221_X1 U22577 ( .B1(n20604), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n20603), 
        .C2(n20757), .A(n20602), .ZN(P3_U2722) );
  INV_X1 U22578 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n20608) );
  INV_X1 U22579 ( .A(n20604), .ZN(n20755) );
  AOI21_X1 U22580 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n20777), .A(n20605), .ZN(
        n20607) );
  OAI222_X1 U22581 ( .A1(n20645), .A2(n20608), .B1(n20755), .B2(n20607), .C1(
        n20739), .C2(n20606), .ZN(P3_U2723) );
  NAND2_X1 U22582 ( .A1(n20777), .A2(n20612), .ZN(n20615) );
  AOI22_X1 U22583 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20782), .B1(n20781), .B2(
        n20609), .ZN(n20610) );
  OAI221_X1 U22584 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n20612), .C1(n20611), 
        .C2(n20615), .A(n20610), .ZN(P3_U2724) );
  NOR2_X1 U22585 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20619), .ZN(n20614) );
  OAI222_X1 U22586 ( .A1(n20645), .A2(n14607), .B1(n20615), .B2(n20614), .C1(
        n20739), .C2(n20613), .ZN(P3_U2725) );
  INV_X1 U22587 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n20620) );
  AOI21_X1 U22588 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n20777), .A(n20616), .ZN(
        n20618) );
  OAI222_X1 U22589 ( .A1(n20645), .A2(n20620), .B1(n20619), .B2(n20618), .C1(
        n20739), .C2(n20617), .ZN(P3_U2726) );
  NAND3_X1 U22590 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(n20621), .ZN(n20776) );
  NOR3_X1 U22591 ( .A1(n20622), .A2(n20648), .A3(n20776), .ZN(n20647) );
  NAND2_X1 U22592 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n20647), .ZN(n20637) );
  NOR2_X1 U22593 ( .A1(n20623), .A2(n20637), .ZN(n20640) );
  NAND2_X1 U22594 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n20640), .ZN(n20628) );
  NOR2_X1 U22595 ( .A1(n20624), .A2(n20628), .ZN(n20632) );
  AOI21_X1 U22596 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n20777), .A(n20632), .ZN(
        n20626) );
  OAI222_X1 U22597 ( .A1(n20741), .A2(n20645), .B1(n20627), .B2(n20626), .C1(
        n20739), .C2(n20625), .ZN(P3_U2728) );
  INV_X1 U22598 ( .A(n20628), .ZN(n20635) );
  AOI21_X1 U22599 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n20777), .A(n20635), .ZN(
        n20631) );
  INV_X1 U22600 ( .A(n20629), .ZN(n20630) );
  OAI222_X1 U22601 ( .A1(n20674), .A2(n20645), .B1(n20632), .B2(n20631), .C1(
        n20739), .C2(n20630), .ZN(P3_U2729) );
  AOI21_X1 U22602 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n20777), .A(n20640), .ZN(
        n20634) );
  OAI222_X1 U22603 ( .A1(n20636), .A2(n20645), .B1(n20635), .B2(n20634), .C1(
        n20739), .C2(n20633), .ZN(P3_U2730) );
  INV_X1 U22604 ( .A(n20637), .ZN(n20644) );
  AOI21_X1 U22605 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n20777), .A(n20644), .ZN(
        n20639) );
  OAI222_X1 U22606 ( .A1(n20641), .A2(n20645), .B1(n20640), .B2(n20639), .C1(
        n20739), .C2(n20638), .ZN(P3_U2731) );
  AOI21_X1 U22607 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n20777), .A(n20647), .ZN(
        n20643) );
  OAI222_X1 U22608 ( .A1(n20646), .A2(n20645), .B1(n20644), .B2(n20643), .C1(
        n20739), .C2(n20642), .ZN(P3_U2732) );
  AOI211_X1 U22609 ( .C1(n20648), .C2(n20776), .A(n20757), .B(n20647), .ZN(
        n20649) );
  AOI21_X1 U22610 ( .B1(n20782), .B2(BUF2_REG_2__SCAN_IN), .A(n20649), .ZN(
        n20650) );
  OAI21_X1 U22611 ( .B1(n20651), .B2(n20739), .A(n20650), .ZN(P3_U2733) );
  NOR2_X1 U22612 ( .A1(n20777), .A2(n20652), .ZN(n20744) );
  NAND2_X1 U22613 ( .A1(n20653), .A2(n20757), .ZN(n20740) );
  AOI22_X1 U22614 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20747), .B1(n20781), .B2(
        n20654), .ZN(n20659) );
  NAND4_X1 U22615 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_11__SCAN_IN), .ZN(n20657)
         );
  NAND4_X1 U22616 ( .A1(n20655), .A2(P3_EAX_REG_8__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .A4(P3_EAX_REG_14__SCAN_IN), .ZN(n20656) );
  NAND2_X1 U22617 ( .A1(n20764), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n20763) );
  NAND3_X1 U22618 ( .A1(n20768), .A2(n20748), .A3(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n20686) );
  NAND2_X1 U22619 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n20682), .ZN(n20681) );
  NAND2_X1 U22620 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20675), .ZN(n20661) );
  AND2_X1 U22621 ( .A1(n20777), .A2(n20661), .ZN(n20669) );
  NOR2_X1 U22622 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n20661), .ZN(n20668) );
  AOI21_X1 U22623 ( .B1(n20669), .B2(P3_EAX_REG_21__SCAN_IN), .A(n20668), .ZN(
        n20658) );
  OAI211_X1 U22624 ( .C1(n20660), .C2(n20754), .A(n20659), .B(n20658), .ZN(
        P3_U2714) );
  AOI22_X1 U22625 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20747), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20744), .ZN(n20663) );
  OAI211_X1 U22626 ( .C1(n20675), .C2(P3_EAX_REG_20__SCAN_IN), .A(n20777), .B(
        n20661), .ZN(n20662) );
  OAI211_X1 U22627 ( .C1(n20664), .C2(n20739), .A(n20663), .B(n20662), .ZN(
        P3_U2715) );
  OAI22_X1 U22628 ( .A1(n20666), .A2(n20739), .B1(n20665), .B2(n20754), .ZN(
        n20667) );
  AOI221_X1 U22629 ( .B1(n20669), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n20668), 
        .C2(P3_EAX_REG_22__SCAN_IN), .A(n20667), .ZN(n20673) );
  NAND4_X1 U22630 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_21__SCAN_IN), .A4(P3_EAX_REG_20__SCAN_IN), .ZN(n20670)
         );
  NOR2_X1 U22631 ( .A1(n20676), .A2(n20670), .ZN(n20690) );
  NAND4_X1 U22632 ( .A1(n20748), .A2(n20768), .A3(n20690), .A4(n20671), .ZN(
        n20672) );
  OAI211_X1 U22633 ( .C1(n20740), .C2(n20674), .A(n20673), .B(n20672), .ZN(
        P3_U2713) );
  AOI22_X1 U22634 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20747), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20744), .ZN(n20679) );
  AOI211_X1 U22635 ( .C1(n20676), .C2(n20681), .A(n20675), .B(n20757), .ZN(
        n20677) );
  INV_X1 U22636 ( .A(n20677), .ZN(n20678) );
  OAI211_X1 U22637 ( .C1(n20680), .C2(n20739), .A(n20679), .B(n20678), .ZN(
        P3_U2716) );
  AOI22_X1 U22638 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20747), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20744), .ZN(n20684) );
  OAI211_X1 U22639 ( .C1(n20682), .C2(P3_EAX_REG_18__SCAN_IN), .A(n20777), .B(
        n20681), .ZN(n20683) );
  OAI211_X1 U22640 ( .C1(n20685), .C2(n20739), .A(n20684), .B(n20683), .ZN(
        P3_U2717) );
  AOI22_X1 U22641 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20747), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20744), .ZN(n20688) );
  OAI211_X1 U22642 ( .C1(n20748), .C2(P3_EAX_REG_17__SCAN_IN), .A(n20777), .B(
        n20686), .ZN(n20687) );
  OAI211_X1 U22643 ( .C1(n20689), .C2(n20739), .A(n20688), .B(n20687), .ZN(
        P3_U2718) );
  AOI22_X1 U22644 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20747), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20744), .ZN(n20694) );
  NAND3_X1 U22645 ( .A1(n20748), .A2(n20690), .A3(P3_EAX_REG_22__SCAN_IN), 
        .ZN(n20737) );
  NAND2_X1 U22646 ( .A1(n20768), .A2(n20735), .ZN(n20728) );
  AOI211_X1 U22647 ( .C1(n20691), .C2(n20731), .A(n20697), .B(n20757), .ZN(
        n20692) );
  INV_X1 U22648 ( .A(n20692), .ZN(n20693) );
  OAI211_X1 U22649 ( .C1(n20695), .C2(n20739), .A(n20694), .B(n20693), .ZN(
        P3_U2710) );
  INV_X1 U22650 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n20700) );
  AOI22_X1 U22651 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20747), .B1(n20781), .B2(
        n20696), .ZN(n20699) );
  NAND2_X1 U22652 ( .A1(n20697), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n20701) );
  OAI211_X1 U22653 ( .C1(n20697), .C2(P3_EAX_REG_26__SCAN_IN), .A(n20777), .B(
        n20701), .ZN(n20698) );
  OAI211_X1 U22654 ( .C1(n20754), .C2(n20700), .A(n20699), .B(n20698), .ZN(
        P3_U2709) );
  NAND2_X1 U22655 ( .A1(n20716), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n20712) );
  NOR2_X1 U22656 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n20712), .ZN(n20703) );
  NAND2_X1 U22657 ( .A1(n20777), .A2(n20712), .ZN(n20710) );
  OAI21_X1 U22658 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n20784), .A(n20710), .ZN(
        n20702) );
  AOI22_X1 U22659 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n20703), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n20702), .ZN(n20704) );
  OAI21_X1 U22660 ( .B1(n20705), .B2(n20754), .A(n20704), .ZN(P3_U2704) );
  OAI22_X1 U22661 ( .A1(n20707), .A2(n20739), .B1(n20706), .B2(n20754), .ZN(
        n20708) );
  AOI21_X1 U22662 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n20747), .A(n20708), .ZN(
        n20709) );
  OAI221_X1 U22663 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n20712), .C1(n20711), 
        .C2(n20710), .A(n20709), .ZN(P3_U2705) );
  AOI22_X1 U22664 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20747), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20744), .ZN(n20714) );
  OAI211_X1 U22665 ( .C1(n20716), .C2(P3_EAX_REG_29__SCAN_IN), .A(n20777), .B(
        n20712), .ZN(n20713) );
  OAI211_X1 U22666 ( .C1(n20715), .C2(n20739), .A(n20714), .B(n20713), .ZN(
        P3_U2706) );
  INV_X1 U22667 ( .A(n20716), .ZN(n20719) );
  OAI21_X1 U22668 ( .B1(n20757), .B2(n20717), .A(n20723), .ZN(n20718) );
  AOI22_X1 U22669 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n20744), .B1(n20719), .B2(
        n20718), .ZN(n20722) );
  AOI22_X1 U22670 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20747), .B1(n20781), .B2(
        n20720), .ZN(n20721) );
  NAND2_X1 U22671 ( .A1(n20722), .A2(n20721), .ZN(P3_U2707) );
  AOI22_X1 U22672 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20747), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n20744), .ZN(n20726) );
  OAI211_X1 U22673 ( .C1(n20724), .C2(P3_EAX_REG_27__SCAN_IN), .A(n20777), .B(
        n20723), .ZN(n20725) );
  OAI211_X1 U22674 ( .C1(n20727), .C2(n20739), .A(n20726), .B(n20725), .ZN(
        P3_U2708) );
  OAI21_X1 U22675 ( .B1(n20757), .B2(n20729), .A(n20728), .ZN(n20730) );
  AOI22_X1 U22676 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n20744), .B1(n20731), .B2(
        n20730), .ZN(n20734) );
  AOI22_X1 U22677 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20747), .B1(n20781), .B2(
        n20732), .ZN(n20733) );
  NAND2_X1 U22678 ( .A1(n20734), .A2(n20733), .ZN(P3_U2711) );
  AOI211_X1 U22679 ( .C1(n20737), .C2(n20736), .A(n20757), .B(n20735), .ZN(
        n20743) );
  OAI22_X1 U22680 ( .A1(n20741), .A2(n20740), .B1(n20739), .B2(n20738), .ZN(
        n20742) );
  AOI211_X1 U22681 ( .C1(n20744), .C2(BUF2_REG_23__SCAN_IN), .A(n20743), .B(
        n20742), .ZN(n20745) );
  INV_X1 U22682 ( .A(n20745), .ZN(P3_U2712) );
  AOI22_X1 U22683 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20747), .B1(n20781), .B2(
        n20746), .ZN(n20752) );
  AOI211_X1 U22684 ( .C1(n20763), .C2(n20749), .A(n20757), .B(n20748), .ZN(
        n20750) );
  INV_X1 U22685 ( .A(n20750), .ZN(n20751) );
  OAI211_X1 U22686 ( .C1(n20754), .C2(n20753), .A(n20752), .B(n20751), .ZN(
        P3_U2719) );
  NAND2_X1 U22687 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n20755), .ZN(n20761) );
  AOI22_X1 U22688 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20782), .B1(n20781), .B2(
        n20756), .ZN(n20760) );
  OR3_X1 U22689 ( .A1(n20758), .A2(n20757), .A3(n20764), .ZN(n20759) );
  OAI211_X1 U22690 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n20761), .A(n20760), .B(
        n20759), .ZN(P3_U2721) );
  AOI22_X1 U22691 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20782), .B1(n20781), .B2(
        n20762), .ZN(n20766) );
  OAI211_X1 U22692 ( .C1(n20764), .C2(P3_EAX_REG_15__SCAN_IN), .A(n20777), .B(
        n20763), .ZN(n20765) );
  NAND2_X1 U22693 ( .A1(n20766), .A2(n20765), .ZN(P3_U2720) );
  AOI21_X1 U22694 ( .B1(n20768), .B2(n20767), .A(n20775), .ZN(n20771) );
  AOI22_X1 U22695 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20782), .B1(n20781), .B2(
        n20769), .ZN(n20770) );
  OAI221_X1 U22696 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n20773), .C1(n20772), 
        .C2(n20771), .A(n20770), .ZN(P3_U2727) );
  AOI22_X1 U22697 ( .A1(n20782), .A2(BUF2_REG_1__SCAN_IN), .B1(n20781), .B2(
        n20774), .ZN(n20779) );
  NOR2_X1 U22698 ( .A1(n20775), .A2(n20785), .ZN(n20786) );
  OAI211_X1 U22699 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n20786), .A(n20777), .B(
        n20776), .ZN(n20778) );
  NAND2_X1 U22700 ( .A1(n20779), .A2(n20778), .ZN(P3_U2734) );
  AOI22_X1 U22701 ( .A1(n20782), .A2(BUF2_REG_0__SCAN_IN), .B1(n20781), .B2(
        n20780), .ZN(n20783) );
  OAI221_X1 U22702 ( .B1(n20786), .B2(n20785), .C1(n20786), .C2(n20784), .A(
        n20783), .ZN(P3_U2735) );
  INV_X1 U22703 ( .A(n20787), .ZN(n21247) );
  NAND2_X1 U22704 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20809) );
  NAND2_X1 U22705 ( .A1(n20943), .A2(n20788), .ZN(n20793) );
  AOI22_X1 U22706 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21007), .B1(
        n20793), .B2(n11421), .ZN(n21212) );
  OAI21_X1 U22707 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n21212), .A(n20789), 
        .ZN(n20790) );
  AOI22_X1 U22708 ( .A1(n21247), .A2(n11421), .B1(n20809), .B2(n20790), .ZN(
        n20791) );
  INV_X1 U22709 ( .A(n20833), .ZN(n20831) );
  AOI22_X1 U22710 ( .A1(n20833), .A2(n11421), .B1(n20791), .B2(n20831), .ZN(
        P3_U3290) );
  INV_X1 U22711 ( .A(n20792), .ZN(n20795) );
  AOI22_X1 U22712 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n21071), .B2(n20864), .ZN(
        n20812) );
  AOI21_X1 U22713 ( .B1(n21192), .B2(n11421), .A(n21146), .ZN(n20797) );
  AOI22_X1 U22714 ( .A1(n20795), .A2(n20793), .B1(n20797), .B2(n11420), .ZN(
        n21214) );
  OAI22_X1 U22715 ( .A1(n20812), .A2(n20809), .B1(n21214), .B2(n20808), .ZN(
        n20794) );
  AOI21_X1 U22716 ( .B1(n21247), .B2(n20795), .A(n20794), .ZN(n20796) );
  AOI22_X1 U22717 ( .A1(n20833), .A2(n11420), .B1(n20796), .B2(n20831), .ZN(
        P3_U3289) );
  OAI22_X1 U22718 ( .A1(n20801), .A2(n20800), .B1(n20799), .B2(n20798), .ZN(
        n20821) );
  AOI211_X1 U22719 ( .C1(n11420), .C2(n20802), .A(n20820), .B(n20821), .ZN(
        n20804) );
  OAI22_X1 U22720 ( .A1(n20816), .A2(n20804), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n20803), .ZN(n20806) );
  AOI22_X1 U22721 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20806), .B1(
        n21204), .B2(n20805), .ZN(n20807) );
  INV_X1 U22722 ( .A(n20808), .ZN(n20829) );
  INV_X1 U22723 ( .A(n20809), .ZN(n20811) );
  AOI222_X1 U22724 ( .A1(n21218), .A2(n20829), .B1(n20812), .B2(n20811), .C1(
        n20810), .C2(n21247), .ZN(n20815) );
  AOI21_X1 U22725 ( .B1(n21247), .B2(n14557), .A(n20833), .ZN(n20814) );
  OAI22_X1 U22726 ( .A1(n20833), .A2(n20815), .B1(n20814), .B2(n20813), .ZN(
        P3_U3288) );
  NOR2_X1 U22727 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20816), .ZN(
        n20817) );
  XOR2_X1 U22728 ( .A(n11427), .B(n20817), .Z(n20827) );
  NAND2_X1 U22729 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20818) );
  AOI222_X1 U22730 ( .A1(n20822), .A2(n20821), .B1(n20820), .B2(n11421), .C1(
        n20819), .C2(n20818), .ZN(n20825) );
  OAI22_X1 U22731 ( .A1(n20825), .A2(n11427), .B1(n20824), .B2(n20823), .ZN(
        n20826) );
  AOI21_X1 U22732 ( .B1(n20827), .B2(n21204), .A(n20826), .ZN(n21211) );
  INV_X1 U22733 ( .A(n21211), .ZN(n20828) );
  AOI22_X1 U22734 ( .A1(n21247), .A2(n20830), .B1(n20829), .B2(n20828), .ZN(
        n20832) );
  AOI22_X1 U22735 ( .A1(n20833), .A2(n11427), .B1(n20832), .B2(n20831), .ZN(
        P3_U3285) );
  NOR2_X1 U22736 ( .A1(n21148), .A2(n20932), .ZN(n21133) );
  AOI21_X1 U22737 ( .B1(n21133), .B2(n20834), .A(n21192), .ZN(n20835) );
  AOI21_X1 U22738 ( .B1(n21204), .B2(n20836), .A(n20835), .ZN(n21117) );
  NOR2_X1 U22739 ( .A1(n21007), .A2(n21204), .ZN(n21181) );
  INV_X1 U22740 ( .A(n21181), .ZN(n20998) );
  AOI22_X1 U22741 ( .A1(n21203), .A2(n21091), .B1(n20837), .B2(n20998), .ZN(
        n20838) );
  OAI211_X1 U22742 ( .C1(n20839), .C2(n21137), .A(n21117), .B(n20838), .ZN(
        n20996) );
  AOI21_X1 U22743 ( .B1(n21188), .B2(n20840), .A(n21194), .ZN(n21115) );
  OAI21_X1 U22744 ( .B1(n20841), .B2(n20943), .A(n21115), .ZN(n20842) );
  OAI21_X1 U22745 ( .B1(n20996), .B2(n20842), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n20847) );
  NOR2_X1 U22746 ( .A1(n21089), .A2(n21194), .ZN(n21128) );
  AOI22_X1 U22747 ( .A1(n21196), .A2(n20844), .B1(n20843), .B2(n21128), .ZN(
        n20845) );
  OAI221_X1 U22748 ( .B1(n10979), .B2(n20847), .C1(n11764), .C2(n20846), .A(
        n20845), .ZN(P3_U2841) );
  NOR2_X1 U22749 ( .A1(n21204), .A2(n21188), .ZN(n21126) );
  AOI22_X1 U22750 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21192), .B1(
        n21126), .B2(n20994), .ZN(n20848) );
  AOI221_X1 U22751 ( .B1(n20856), .B2(n20850), .C1(n21203), .C2(n20849), .A(
        n20848), .ZN(n20852) );
  AOI22_X1 U22752 ( .A1(n10979), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21080), .ZN(n20851) );
  OAI21_X1 U22753 ( .B1(n20852), .B2(n21194), .A(n20851), .ZN(P3_U2862) );
  NAND2_X1 U22754 ( .A1(n21171), .A2(n21203), .ZN(n21015) );
  INV_X1 U22755 ( .A(n21162), .ZN(n21063) );
  NAND3_X1 U22756 ( .A1(n20864), .A2(n20853), .A3(n21063), .ZN(n20858) );
  NOR2_X1 U22757 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21126), .ZN(
        n20854) );
  AOI22_X1 U22758 ( .A1(n20856), .A2(n20855), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20854), .ZN(n20857) );
  NAND2_X1 U22759 ( .A1(n20858), .A2(n20857), .ZN(n20859) );
  AOI22_X1 U22760 ( .A1(n21171), .A2(n20859), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21080), .ZN(n20861) );
  NAND2_X1 U22761 ( .A1(n10979), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n20860) );
  OAI211_X1 U22762 ( .C1(n20862), .C2(n21015), .A(n20861), .B(n20860), .ZN(
        P3_U2861) );
  NAND2_X1 U22763 ( .A1(n10979), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n20871) );
  NOR3_X1 U22764 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n20864), .A3(
        n20872), .ZN(n20869) );
  NOR2_X1 U22765 ( .A1(n20864), .A2(n20994), .ZN(n20863) );
  AOI21_X1 U22766 ( .B1(n20863), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n20873), .ZN(n20867) );
  NAND2_X1 U22767 ( .A1(n20994), .A2(n21188), .ZN(n21134) );
  INV_X1 U22768 ( .A(n21134), .ZN(n21006) );
  OAI211_X1 U22769 ( .C1(n21006), .C2(n20864), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n21187), .ZN(n20865) );
  OAI211_X1 U22770 ( .C1(n20867), .C2(n21172), .A(n20866), .B(n20865), .ZN(
        n20868) );
  OAI21_X1 U22771 ( .B1(n20869), .B2(n20868), .A(n21171), .ZN(n20870) );
  OAI211_X1 U22772 ( .C1(n21094), .C2(n11522), .A(n20871), .B(n20870), .ZN(
        P3_U2860) );
  AOI22_X1 U22773 ( .A1(n10979), .A2(P3_REIP_REG_3__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21080), .ZN(n20881) );
  NAND2_X1 U22774 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20874) );
  OAI22_X1 U22775 ( .A1(n20873), .A2(n21172), .B1(n20872), .B2(n20874), .ZN(
        n20907) );
  INV_X1 U22776 ( .A(n20907), .ZN(n20877) );
  OAI21_X1 U22777 ( .B1(n21006), .B2(n20874), .A(n21187), .ZN(n20875) );
  OAI21_X1 U22778 ( .B1(n20876), .B2(n21172), .A(n20875), .ZN(n20893) );
  NOR2_X1 U22779 ( .A1(n11525), .A2(n20893), .ZN(n20887) );
  AOI211_X1 U22780 ( .C1(n20877), .C2(n11525), .A(n20887), .B(n21194), .ZN(
        n20878) );
  AOI21_X1 U22781 ( .B1(n20879), .B2(n20914), .A(n20878), .ZN(n20880) );
  OAI211_X1 U22782 ( .C1(n21015), .C2(n20882), .A(n20881), .B(n20880), .ZN(
        P3_U2859) );
  NAND2_X1 U22783 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21063), .ZN(
        n20886) );
  NAND3_X1 U22784 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n20883), .A3(
        n20907), .ZN(n20884) );
  OAI211_X1 U22785 ( .C1(n20887), .C2(n20886), .A(n20885), .B(n20884), .ZN(
        n20888) );
  AOI22_X1 U22786 ( .A1(n21171), .A2(n20888), .B1(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n21080), .ZN(n20889) );
  OAI21_X1 U22787 ( .B1(n11764), .B2(n20890), .A(n20889), .ZN(P3_U2858) );
  NAND2_X1 U22788 ( .A1(n21171), .A2(n20907), .ZN(n20900) );
  NAND3_X1 U22789 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n20891), .ZN(n20898) );
  INV_X1 U22790 ( .A(n21015), .ZN(n21081) );
  AOI22_X1 U22791 ( .A1(n10979), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n21081), 
        .B2(n20892), .ZN(n20897) );
  AOI21_X1 U22792 ( .B1(n21063), .B2(n20901), .A(n20893), .ZN(n20894) );
  OAI21_X1 U22793 ( .B1(n20894), .B2(n21194), .A(n21094), .ZN(n20899) );
  AOI22_X1 U22794 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20899), .B1(
        n20914), .B2(n20895), .ZN(n20896) );
  OAI211_X1 U22795 ( .C1(n20900), .C2(n20898), .A(n20897), .B(n20896), .ZN(
        P3_U2857) );
  AOI22_X1 U22796 ( .A1(n10979), .A2(P3_REIP_REG_6__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n20899), .ZN(n20905) );
  NOR3_X1 U22797 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n20901), .A3(
        n20900), .ZN(n20902) );
  AOI21_X1 U22798 ( .B1(n20903), .B2(n20914), .A(n20902), .ZN(n20904) );
  OAI211_X1 U22799 ( .C1(n21015), .C2(n20906), .A(n20905), .B(n20904), .ZN(
        P3_U2856) );
  AOI22_X1 U22800 ( .A1(n10979), .A2(P3_REIP_REG_7__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n21080), .ZN(n20916) );
  NAND2_X1 U22801 ( .A1(n20908), .A2(n20907), .ZN(n20927) );
  AOI21_X1 U22802 ( .B1(n20918), .B2(n20927), .A(n21194), .ZN(n20912) );
  AOI22_X1 U22803 ( .A1(n21204), .A2(n20910), .B1(n21187), .B2(n20909), .ZN(
        n20911) );
  NAND3_X1 U22804 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n20911), .A3(
        n21134), .ZN(n20919) );
  AOI22_X1 U22805 ( .A1(n20914), .A2(n20913), .B1(n20912), .B2(n20919), .ZN(
        n20915) );
  OAI211_X1 U22806 ( .C1(n21015), .C2(n20917), .A(n20916), .B(n20915), .ZN(
        P3_U2855) );
  AOI22_X1 U22807 ( .A1(n10979), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21080), .ZN(n20925) );
  OR3_X1 U22808 ( .A1(n20918), .A2(n20927), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20921) );
  NAND3_X1 U22809 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21063), .A3(
        n20919), .ZN(n20920) );
  OAI211_X1 U22810 ( .C1(n21137), .C2(n20922), .A(n20921), .B(n20920), .ZN(
        n20923) );
  AOI22_X1 U22811 ( .A1(n21171), .A2(n20923), .B1(n21196), .B2(n20922), .ZN(
        n20924) );
  OAI211_X1 U22812 ( .C1(n21015), .C2(n20926), .A(n20925), .B(n20924), .ZN(
        P3_U2854) );
  NAND2_X1 U22813 ( .A1(n20934), .A2(n20931), .ZN(n20942) );
  AOI22_X1 U22814 ( .A1(n10979), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n21196), 
        .B2(n20930), .ZN(n20941) );
  OAI21_X1 U22815 ( .B1(n20938), .B2(n20931), .A(n21204), .ZN(n20933) );
  NAND2_X1 U22816 ( .A1(n21007), .A2(n20932), .ZN(n21179) );
  OAI211_X1 U22817 ( .C1(n20934), .C2(n21192), .A(n20933), .B(n21179), .ZN(
        n20950) );
  NAND2_X1 U22818 ( .A1(n21137), .A2(n21050), .ZN(n21143) );
  NOR2_X1 U22819 ( .A1(n21138), .A2(n21137), .ZN(n20935) );
  NOR2_X1 U22820 ( .A1(n20978), .A2(n21172), .ZN(n20945) );
  AOI211_X1 U22821 ( .C1(n20936), .C2(n21203), .A(n20935), .B(n20945), .ZN(
        n21190) );
  OAI221_X1 U22822 ( .B1(n20943), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n20943), .C2(n20944), .A(n21190), .ZN(n20937) );
  AOI211_X1 U22823 ( .C1(n20938), .C2(n21143), .A(n21194), .B(n20937), .ZN(
        n21180) );
  OAI21_X1 U22824 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n20943), .A(
        n21180), .ZN(n20939) );
  OAI211_X1 U22825 ( .C1(n20950), .C2(n20939), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n11764), .ZN(n20940) );
  OAI211_X1 U22826 ( .C1(n20942), .C2(n21200), .A(n20941), .B(n20940), .ZN(
        P3_U2851) );
  AOI22_X1 U22827 ( .A1(n10979), .A2(P3_REIP_REG_12__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21080), .ZN(n20956) );
  NAND2_X1 U22828 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20946) );
  AOI21_X1 U22829 ( .B1(n20959), .B2(n20944), .A(n20943), .ZN(n20960) );
  AOI211_X1 U22830 ( .C1(n20946), .C2(n21007), .A(n20960), .B(n20945), .ZN(
        n20947) );
  OAI21_X1 U22831 ( .B1(n20948), .B2(n21050), .A(n20947), .ZN(n20949) );
  AOI211_X1 U22832 ( .C1(n21114), .C2(n20951), .A(n20950), .B(n20949), .ZN(
        n21170) );
  NOR3_X1 U22833 ( .A1(n21170), .A2(n20952), .A3(n21194), .ZN(n20953) );
  AOI21_X1 U22834 ( .B1(n21196), .B2(n20954), .A(n20953), .ZN(n20955) );
  OAI211_X1 U22835 ( .C1(n21200), .C2(n20957), .A(n20956), .B(n20955), .ZN(
        P3_U2850) );
  AOI22_X1 U22836 ( .A1(n10979), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21080), .ZN(n20971) );
  NAND2_X1 U22837 ( .A1(n20958), .A2(n20980), .ZN(n20967) );
  AOI21_X1 U22838 ( .B1(n20959), .B2(n20978), .A(n21172), .ZN(n20961) );
  AOI211_X1 U22839 ( .C1(n20962), .C2(n21007), .A(n20961), .B(n20960), .ZN(
        n20963) );
  OAI211_X1 U22840 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n21126), .A(
        n20963), .B(n21179), .ZN(n20964) );
  AOI22_X1 U22841 ( .A1(n21114), .A2(n20965), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n20964), .ZN(n20966) );
  OAI21_X1 U22842 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n20967), .A(
        n20966), .ZN(n20969) );
  AOI22_X1 U22843 ( .A1(n21171), .A2(n20969), .B1(n21081), .B2(n20968), .ZN(
        n20970) );
  OAI211_X1 U22844 ( .C1(n20972), .C2(n21168), .A(n20971), .B(n20970), .ZN(
        P3_U2848) );
  NOR2_X1 U22845 ( .A1(n20973), .A2(n21137), .ZN(n20975) );
  NOR2_X1 U22846 ( .A1(n21136), .A2(n21050), .ZN(n20983) );
  AOI22_X1 U22847 ( .A1(n20976), .A2(n20975), .B1(n20974), .B2(n20983), .ZN(
        n20991) );
  OAI22_X1 U22848 ( .A1(n20985), .A2(n21188), .B1(n21148), .B2(n21186), .ZN(
        n20977) );
  OAI211_X1 U22849 ( .C1(n20978), .C2(n21172), .A(n21179), .B(n20977), .ZN(
        n20981) );
  NAND3_X1 U22850 ( .A1(n20980), .A2(n20979), .A3(n20981), .ZN(n20990) );
  AOI21_X1 U22851 ( .B1(n20982), .B2(n20998), .A(n20981), .ZN(n21160) );
  AOI211_X1 U22852 ( .C1(n21114), .C2(n20984), .A(n20983), .B(n21194), .ZN(
        n21161) );
  AOI211_X1 U22853 ( .C1(n21160), .C2(n21161), .A(n10979), .B(n20985), .ZN(
        n20986) );
  AOI211_X1 U22854 ( .C1(n21196), .C2(n20988), .A(n20987), .B(n20986), .ZN(
        n20989) );
  OAI221_X1 U22855 ( .B1(n20992), .B2(n20991), .C1(n21194), .C2(n20990), .A(
        n20989), .ZN(P3_U2847) );
  NAND2_X1 U22856 ( .A1(n20993), .A2(n21133), .ZN(n21008) );
  OAI21_X1 U22857 ( .B1(n20994), .B2(n21008), .A(n21188), .ZN(n20995) );
  INV_X1 U22858 ( .A(n20995), .ZN(n20997) );
  AOI211_X1 U22859 ( .C1(n20999), .C2(n20998), .A(n20997), .B(n20996), .ZN(
        n21001) );
  OR2_X1 U22860 ( .A1(n21088), .A2(n21089), .ZN(n21000) );
  AOI221_X1 U22861 ( .B1(n21001), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), 
        .C1(n21000), .C2(n21087), .A(n21194), .ZN(n21002) );
  AOI21_X1 U22862 ( .B1(n21080), .B2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n21002), .ZN(n21004) );
  OAI211_X1 U22863 ( .C1(n21005), .C2(n21168), .A(n21004), .B(n21003), .ZN(
        P3_U2840) );
  AND2_X1 U22864 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21009) );
  AOI221_X1 U22865 ( .B1(n21188), .B2(n21008), .C1(n21007), .C2(n21008), .A(
        n21006), .ZN(n21095) );
  OAI211_X1 U22866 ( .C1(n21162), .C2(n21009), .A(n21099), .B(n21095), .ZN(
        n21023) );
  NOR2_X1 U22867 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21010), .ZN(
        n21011) );
  AOI22_X1 U22868 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21023), .B1(
        n21011), .B2(n21053), .ZN(n21012) );
  OAI21_X1 U22869 ( .B1(n21137), .B2(n21013), .A(n21012), .ZN(n21018) );
  OAI22_X1 U22870 ( .A1(n21168), .A2(n21016), .B1(n21015), .B2(n21014), .ZN(
        n21017) );
  AOI21_X1 U22871 ( .B1(n21171), .B2(n21018), .A(n21017), .ZN(n21020) );
  OAI211_X1 U22872 ( .C1(n21094), .C2(n21025), .A(n21020), .B(n21019), .ZN(
        P3_U2837) );
  INV_X1 U22873 ( .A(n21021), .ZN(n21033) );
  NOR2_X1 U22874 ( .A1(n21022), .A2(n21137), .ZN(n21024) );
  NAND2_X1 U22875 ( .A1(n21081), .A2(n21040), .ZN(n21026) );
  OAI221_X1 U22876 ( .B1(n21194), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), 
        .C1(n21194), .C2(n21027), .A(n21026), .ZN(n21030) );
  NOR4_X1 U22877 ( .A1(n21089), .A2(n21088), .A3(n21087), .A4(n21028), .ZN(
        n21029) );
  AOI222_X1 U22878 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21030), 
        .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n21080), .C1(n21030), 
        .C2(n21029), .ZN(n21031) );
  OAI211_X1 U22879 ( .C1(n21033), .C2(n21168), .A(n21032), .B(n21031), .ZN(
        P3_U2836) );
  NOR2_X1 U22880 ( .A1(n21034), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n21046) );
  AOI211_X1 U22881 ( .C1(n21114), .C2(n21037), .A(n21036), .B(n21035), .ZN(
        n21038) );
  OAI211_X1 U22882 ( .C1(n21146), .C2(n21039), .A(n21095), .B(n21038), .ZN(
        n21041) );
  AOI22_X1 U22883 ( .A1(n21171), .A2(n21041), .B1(n21081), .B2(n21040), .ZN(
        n21045) );
  AOI22_X1 U22884 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21080), .B1(
        n21196), .B2(n21042), .ZN(n21044) );
  OAI211_X1 U22885 ( .C1(n21046), .C2(n21045), .A(n21044), .B(n21043), .ZN(
        P3_U2835) );
  OAI221_X1 U22886 ( .B1(n21192), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), 
        .C1(n21192), .C2(n21048), .A(n21047), .ZN(n21061) );
  OAI22_X1 U22887 ( .A1(n21051), .A2(n21050), .B1(n21049), .B2(n21137), .ZN(
        n21066) );
  NAND3_X1 U22888 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n21054), .A3(
        n21053), .ZN(n21073) );
  OAI21_X1 U22889 ( .B1(n21055), .B2(n21137), .A(n21073), .ZN(n21056) );
  AOI21_X1 U22890 ( .B1(n21203), .B2(n21057), .A(n21056), .ZN(n21064) );
  NOR3_X1 U22891 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21064), .A3(
        n21194), .ZN(n21059) );
  AOI22_X1 U22892 ( .A1(n10979), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n21080), 
        .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21069) );
  AOI211_X1 U22893 ( .C1(n21063), .C2(n21062), .A(n21074), .B(n21061), .ZN(
        n21072) );
  INV_X1 U22894 ( .A(n21072), .ZN(n21067) );
  OAI21_X1 U22895 ( .B1(n21064), .B2(n21075), .A(n21074), .ZN(n21065) );
  OAI211_X1 U22896 ( .C1(n21067), .C2(n21066), .A(n21171), .B(n21065), .ZN(
        n21068) );
  OAI211_X1 U22897 ( .C1(n21070), .C2(n21168), .A(n21069), .B(n21068), .ZN(
        P3_U2832) );
  NOR3_X1 U22898 ( .A1(n21162), .A2(n21072), .A3(n21071), .ZN(n21077) );
  NOR4_X1 U22899 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21075), .A3(
        n21074), .A4(n21073), .ZN(n21076) );
  AOI211_X1 U22900 ( .C1(n21078), .C2(n21114), .A(n21077), .B(n21076), .ZN(
        n21086) );
  AOI21_X1 U22901 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21080), .A(
        n21079), .ZN(n21085) );
  AOI22_X1 U22902 ( .A1(n21196), .A2(n21083), .B1(n21082), .B2(n21081), .ZN(
        n21084) );
  OAI211_X1 U22903 ( .C1(n21086), .C2(n21194), .A(n21085), .B(n21084), .ZN(
        P3_U2831) );
  NOR3_X1 U22904 ( .A1(n21089), .A2(n21088), .A3(n21087), .ZN(n21090) );
  AOI21_X1 U22905 ( .B1(n21090), .B2(n21094), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21103) );
  OR2_X1 U22906 ( .A1(n21093), .A2(n21091), .ZN(n21098) );
  NOR2_X1 U22907 ( .A1(n21093), .A2(n21092), .ZN(n21096) );
  OAI211_X1 U22908 ( .C1(n21096), .C2(n21137), .A(n21095), .B(n21094), .ZN(
        n21097) );
  AOI21_X1 U22909 ( .B1(n21203), .B2(n21098), .A(n21097), .ZN(n21106) );
  NAND3_X1 U22910 ( .A1(n21099), .A2(n21106), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21100) );
  NAND2_X1 U22911 ( .A1(n21100), .A2(n11764), .ZN(n21104) );
  AOI22_X1 U22912 ( .A1(n10979), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n21196), 
        .B2(n21101), .ZN(n21102) );
  OAI21_X1 U22913 ( .B1(n21103), .B2(n21104), .A(n21102), .ZN(P3_U2839) );
  AOI211_X1 U22914 ( .C1(n21162), .C2(n21106), .A(n21105), .B(n21104), .ZN(
        n21107) );
  AOI21_X1 U22915 ( .B1(n21108), .B2(n21128), .A(n21107), .ZN(n21110) );
  OAI211_X1 U22916 ( .C1(n21111), .C2(n21168), .A(n21110), .B(n21109), .ZN(
        P3_U2838) );
  INV_X1 U22917 ( .A(n21128), .ZN(n21122) );
  AOI22_X1 U22918 ( .A1(n21114), .A2(n21113), .B1(n21203), .B2(n21112), .ZN(
        n21116) );
  NAND3_X1 U22919 ( .A1(n21117), .A2(n21116), .A3(n21115), .ZN(n21118) );
  NAND2_X1 U22920 ( .A1(n21118), .A2(n11764), .ZN(n21124) );
  AOI21_X1 U22921 ( .B1(n21196), .B2(n21120), .A(n21119), .ZN(n21121) );
  OAI221_X1 U22922 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21122), 
        .C1(n21123), .C2(n21124), .A(n21121), .ZN(P3_U2843) );
  NAND2_X1 U22923 ( .A1(n21123), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21125) );
  OAI21_X1 U22924 ( .B1(n21126), .B2(n21125), .A(n21124), .ZN(n21129) );
  AOI22_X1 U22925 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21129), .B1(
        n21128), .B2(n21127), .ZN(n21131) );
  OAI211_X1 U22926 ( .C1(n21168), .C2(n21132), .A(n21131), .B(n21130), .ZN(
        P3_U2842) );
  AND3_X1 U22927 ( .A1(n21134), .A2(n21133), .A3(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21145) );
  INV_X1 U22928 ( .A(n21135), .ZN(n21140) );
  OAI211_X1 U22929 ( .C1(n21138), .C2(n21137), .A(n21140), .B(n21136), .ZN(
        n21142) );
  AOI21_X1 U22930 ( .B1(n21140), .B2(n21139), .A(n21172), .ZN(n21141) );
  AOI211_X1 U22931 ( .C1(n21143), .C2(n21142), .A(n21141), .B(n21194), .ZN(
        n21144) );
  OAI21_X1 U22932 ( .B1(n21146), .B2(n21145), .A(n21144), .ZN(n21154) );
  OAI221_X1 U22933 ( .B1(n21154), .B2(n21187), .C1(n21154), .C2(n21147), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21153) );
  NOR2_X1 U22934 ( .A1(n21148), .A2(n21200), .ZN(n21163) );
  AOI22_X1 U22935 ( .A1(n21196), .A2(n21150), .B1(n21163), .B2(n21149), .ZN(
        n21151) );
  OAI221_X1 U22936 ( .B1(n10979), .B2(n21153), .C1(n11764), .C2(n21152), .A(
        n21151), .ZN(P3_U2844) );
  NAND2_X1 U22937 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21154), .ZN(
        n21159) );
  AOI22_X1 U22938 ( .A1(n21196), .A2(n21156), .B1(n21163), .B2(n21155), .ZN(
        n21157) );
  OAI221_X1 U22939 ( .B1(n10979), .B2(n21159), .C1(n11764), .C2(n21158), .A(
        n21157), .ZN(P3_U2845) );
  AOI221_X1 U22940 ( .B1(n21162), .B2(n21161), .C1(n21160), .C2(n21161), .A(
        n10979), .ZN(n21164) );
  AOI22_X1 U22941 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21164), .B1(
        n21163), .B2(n11551), .ZN(n21166) );
  OAI211_X1 U22942 ( .C1(n21168), .C2(n21167), .A(n21166), .B(n21165), .ZN(
        P3_U2846) );
  AOI22_X1 U22943 ( .A1(n10979), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21196), 
        .B2(n21169), .ZN(n21175) );
  OAI211_X1 U22944 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n21172), .A(
        n21171), .B(n21170), .ZN(n21173) );
  NAND3_X1 U22945 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11764), .A3(
        n21173), .ZN(n21174) );
  OAI211_X1 U22946 ( .C1(n21176), .C2(n21200), .A(n21175), .B(n21174), .ZN(
        P3_U2849) );
  NAND2_X1 U22947 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21177), .ZN(
        n21185) );
  AOI22_X1 U22948 ( .A1(n10979), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21196), 
        .B2(n21178), .ZN(n21184) );
  OAI211_X1 U22949 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n21181), .A(
        n21180), .B(n21179), .ZN(n21182) );
  NAND3_X1 U22950 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n11764), .A3(
        n21182), .ZN(n21183) );
  OAI211_X1 U22951 ( .C1(n21185), .C2(n21200), .A(n21184), .B(n21183), .ZN(
        P3_U2852) );
  OAI211_X1 U22952 ( .C1(n11543), .C2(n21188), .A(n21187), .B(n21186), .ZN(
        n21189) );
  OAI211_X1 U22953 ( .C1(n21192), .C2(n21191), .A(n21190), .B(n21189), .ZN(
        n21193) );
  OAI21_X1 U22954 ( .B1(n21194), .B2(n21193), .A(n11764), .ZN(n21198) );
  AOI22_X1 U22955 ( .A1(n10979), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n21196), 
        .B2(n21195), .ZN(n21197) );
  OAI221_X1 U22956 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21200), .C1(
        n21199), .C2(n21198), .A(n21197), .ZN(P3_U2853) );
  NAND2_X1 U22957 ( .A1(n21607), .A2(n18353), .ZN(n21242) );
  INV_X1 U22958 ( .A(n21201), .ZN(n21241) );
  INV_X1 U22959 ( .A(n21202), .ZN(n21238) );
  NOR2_X1 U22960 ( .A1(n21204), .A2(n21203), .ZN(n21206) );
  OAI222_X1 U22961 ( .A1(n21210), .A2(n21209), .B1(n21208), .B2(n21207), .C1(
        n21206), .C2(n21205), .ZN(n21258) );
  AOI22_X1 U22962 ( .A1(n21234), .A2(n11427), .B1(n21211), .B2(n21217), .ZN(
        n21225) );
  AND3_X1 U22963 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n21212), .ZN(n21213) );
  OAI22_X1 U22964 ( .A1(n21214), .A2(n21213), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n21212), .ZN(n21216) );
  AOI21_X1 U22965 ( .B1(n21216), .B2(n21217), .A(n21215), .ZN(n21220) );
  AOI221_X1 U22966 ( .B1(n21220), .B2(n21219), .C1(n21221), .C2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21224) );
  OAI21_X1 U22967 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n21221), .ZN(n21223) );
  AOI222_X1 U22968 ( .A1(n21225), .A2(n21224), .B1(n21225), .B2(n21223), .C1(
        n21224), .C2(n21222), .ZN(n21231) );
  AOI211_X1 U22969 ( .C1(n21228), .C2(n21652), .A(n21227), .B(n21226), .ZN(
        n21257) );
  OAI21_X1 U22970 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n21257), .ZN(n21229) );
  NAND4_X1 U22971 ( .A1(n21232), .A2(n21231), .A3(n21230), .A4(n21229), .ZN(
        n21233) );
  AOI211_X1 U22972 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n21234), .A(
        n21258), .B(n21233), .ZN(n21255) );
  OR3_X1 U22973 ( .A1(n21239), .A2(n21238), .A3(n21250), .ZN(n21240) );
  NAND4_X1 U22974 ( .A1(n21243), .A2(n21242), .A3(n21241), .A4(n21240), .ZN(
        P3_U2997) );
  OAI221_X1 U22975 ( .B1(n21246), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21246), 
        .C2(n21245), .A(n21244), .ZN(P3_U3282) );
  AOI22_X1 U22976 ( .A1(n21248), .A2(n21247), .B1(n21607), .B2(n18353), .ZN(
        n21249) );
  INV_X1 U22977 ( .A(n21249), .ZN(n21252) );
  OAI211_X1 U22978 ( .C1(n21255), .C2(n21256), .A(n21254), .B(n21253), .ZN(
        P3_U2996) );
  NOR2_X1 U22979 ( .A1(n21257), .A2(n21256), .ZN(n21261) );
  MUX2_X1 U22980 ( .A(P3_MORE_REG_SCAN_IN), .B(n21258), .S(n21261), .Z(
        P3_U3295) );
  OAI21_X1 U22981 ( .B1(n21261), .B2(n21260), .A(n21259), .ZN(P3_U2637) );
  AOI211_X1 U22982 ( .C1(n21264), .C2(n21667), .A(n21263), .B(n21262), .ZN(
        n21271) );
  INV_X1 U22983 ( .A(n21265), .ZN(n21267) );
  NAND4_X1 U22984 ( .A1(n21267), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n21266), 
        .A4(n21667), .ZN(n21268) );
  NAND2_X1 U22985 ( .A1(n21268), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n21270) );
  NOR2_X1 U22986 ( .A1(n21271), .A2(n21586), .ZN(n21269) );
  AOI22_X1 U22987 ( .A1(n21615), .A2(n21271), .B1(n21270), .B2(n21269), .ZN(
        P1_U3485) );
  INV_X1 U22988 ( .A(n21272), .ZN(n21274) );
  AOI22_X1 U22989 ( .A1(n21274), .A2(n21346), .B1(n21345), .B2(n21273), .ZN(
        n21282) );
  NAND2_X1 U22990 ( .A1(n21348), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n21281) );
  NAND4_X1 U22991 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21275), .A3(
        n16149), .A4(n21319), .ZN(n21280) );
  NOR2_X1 U22992 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21276), .ZN(
        n21278) );
  OAI21_X1 U22993 ( .B1(n21278), .B2(n21277), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21279) );
  NAND4_X1 U22994 ( .A1(n21282), .A2(n21281), .A3(n21280), .A4(n21279), .ZN(
        P1_U3017) );
  NOR2_X1 U22995 ( .A1(n21283), .A2(n21300), .ZN(n21286) );
  OAI21_X1 U22996 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21285), .A(
        n21284), .ZN(n21297) );
  AOI21_X1 U22997 ( .B1(n21305), .B2(n21286), .A(n21297), .ZN(n21296) );
  INV_X1 U22998 ( .A(n21287), .ZN(n21360) );
  NOR2_X1 U22999 ( .A1(n21288), .A2(n21369), .ZN(n21290) );
  NOR2_X1 U23000 ( .A1(n21289), .A2(n21304), .ZN(n21298) );
  AOI211_X1 U23001 ( .C1(n21360), .C2(n21345), .A(n21290), .B(n21298), .ZN(
        n21295) );
  INV_X1 U23002 ( .A(n21291), .ZN(n21293) );
  NOR2_X1 U23003 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21300), .ZN(
        n21292) );
  AOI22_X1 U23004 ( .A1(n21293), .A2(n21346), .B1(n21302), .B2(n21292), .ZN(
        n21294) );
  OAI211_X1 U23005 ( .C1(n21296), .C2(n21301), .A(n21295), .B(n21294), .ZN(
        P1_U3029) );
  AOI211_X1 U23006 ( .C1(n21301), .C2(n21299), .A(n21298), .B(n21297), .ZN(
        n21316) );
  AOI22_X1 U23007 ( .A1(n21371), .A2(n21345), .B1(n21348), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n21310) );
  NOR2_X1 U23008 ( .A1(n21301), .A2(n21300), .ZN(n21303) );
  AOI22_X1 U23009 ( .A1(n21305), .A2(n21304), .B1(n21303), .B2(n21302), .ZN(
        n21318) );
  AOI211_X1 U23010 ( .C1(n21311), .C2(n21317), .A(n21318), .B(n21306), .ZN(
        n21307) );
  AOI21_X1 U23011 ( .B1(n21308), .B2(n21346), .A(n21307), .ZN(n21309) );
  OAI211_X1 U23012 ( .C1(n21316), .C2(n21311), .A(n21310), .B(n21309), .ZN(
        P1_U3027) );
  INV_X1 U23013 ( .A(n21312), .ZN(n21313) );
  AOI222_X1 U23014 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n21348), .B1(n21345), 
        .B2(n21314), .C1(n21346), .C2(n21313), .ZN(n21315) );
  OAI221_X1 U23015 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21318), .C1(
        n21317), .C2(n21316), .A(n21315), .ZN(P1_U3028) );
  AOI22_X1 U23016 ( .A1(n21400), .A2(n21345), .B1(n21348), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n21322) );
  AOI22_X1 U23017 ( .A1(n21320), .A2(n21346), .B1(n21323), .B2(n21319), .ZN(
        n21321) );
  OAI211_X1 U23018 ( .C1(n21324), .C2(n21323), .A(n21322), .B(n21321), .ZN(
        P1_U3025) );
  AOI22_X1 U23019 ( .A1(n21326), .A2(n21346), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n21325), .ZN(n21332) );
  OAI22_X1 U23020 ( .A1(n21383), .A2(n21338), .B1(n21328), .B2(n21327), .ZN(
        n21329) );
  AOI211_X1 U23021 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n21348), .A(n21330), .B(
        n21329), .ZN(n21331) );
  NAND2_X1 U23022 ( .A1(n21332), .A2(n21331), .ZN(P1_U3026) );
  AOI222_X1 U23023 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n21348), .B1(n21345), 
        .B2(n21411), .C1(n21346), .C2(n21333), .ZN(n21335) );
  OAI211_X1 U23024 ( .C1(n21337), .C2(n21336), .A(n21335), .B(n21334), .ZN(
        P1_U3024) );
  NOR2_X1 U23025 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21352), .ZN(
        n21351) );
  OAI22_X1 U23026 ( .A1(n21340), .A2(n21339), .B1(n21338), .B2(n21469), .ZN(
        n21341) );
  AOI211_X1 U23027 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n21348), .A(n21351), 
        .B(n21341), .ZN(n21342) );
  OAI21_X1 U23028 ( .B1(n21349), .B2(n16138), .A(n21342), .ZN(P1_U3016) );
  INV_X1 U23029 ( .A(n21343), .ZN(n21347) );
  AOI22_X1 U23030 ( .A1(n21347), .A2(n21346), .B1(n21345), .B2(n21344), .ZN(
        n21358) );
  NAND2_X1 U23031 ( .A1(n21348), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n21357) );
  INV_X1 U23032 ( .A(n21349), .ZN(n21350) );
  OAI21_X1 U23033 ( .B1(n21351), .B2(n21350), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21356) );
  INV_X1 U23034 ( .A(n21352), .ZN(n21354) );
  NAND3_X1 U23035 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21354), .A3(
        n21353), .ZN(n21355) );
  NAND4_X1 U23036 ( .A1(n21358), .A2(n21357), .A3(n21356), .A4(n21355), .ZN(
        P1_U3015) );
  AOI21_X1 U23037 ( .B1(n21528), .B2(n15268), .A(n21359), .ZN(n21370) );
  AOI22_X1 U23038 ( .A1(n21519), .A2(n21360), .B1(n21551), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n21368) );
  INV_X1 U23039 ( .A(n21361), .ZN(n21362) );
  AOI22_X1 U23040 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n21564), .B1(
        n21521), .B2(n21362), .ZN(n21364) );
  NAND3_X1 U23041 ( .A1(n21528), .A2(P1_REIP_REG_1__SCAN_IN), .A3(n21369), 
        .ZN(n21363) );
  OAI211_X1 U23042 ( .C1(n21872), .C2(n21373), .A(n21364), .B(n21363), .ZN(
        n21365) );
  AOI21_X1 U23043 ( .B1(n21366), .B2(n21392), .A(n21365), .ZN(n21367) );
  OAI211_X1 U23044 ( .C1(n21370), .C2(n21369), .A(n21368), .B(n21367), .ZN(
        P1_U2838) );
  AOI22_X1 U23045 ( .A1(n21519), .A2(n21371), .B1(n21551), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n21372) );
  OAI21_X1 U23046 ( .B1(n21374), .B2(n21373), .A(n21372), .ZN(n21375) );
  AOI211_X1 U23047 ( .C1(n21564), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21492), .B(n21375), .ZN(n21381) );
  OAI21_X1 U23048 ( .B1(n21403), .B2(n21385), .A(n14514), .ZN(n21391) );
  OAI21_X1 U23049 ( .B1(n21403), .B2(n21377), .A(n21376), .ZN(n21378) );
  AOI22_X1 U23050 ( .A1(n21379), .A2(n21392), .B1(n21391), .B2(n21378), .ZN(
        n21380) );
  OAI211_X1 U23051 ( .C1(n21382), .C2(n21560), .A(n21381), .B(n21380), .ZN(
        P1_U2836) );
  INV_X1 U23052 ( .A(n21383), .ZN(n21384) );
  NAND2_X1 U23053 ( .A1(n21519), .A2(n21384), .ZN(n21390) );
  NAND2_X1 U23054 ( .A1(n21551), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n21389) );
  NAND2_X1 U23055 ( .A1(n21385), .A2(n21528), .ZN(n21386) );
  OAI21_X1 U23056 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n21386), .A(n21476), .ZN(
        n21387) );
  AOI21_X1 U23057 ( .B1(n21564), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n21387), .ZN(n21388) );
  AND3_X1 U23058 ( .A1(n21390), .A2(n21389), .A3(n21388), .ZN(n21395) );
  AOI22_X1 U23059 ( .A1(n21393), .A2(n21392), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n21391), .ZN(n21394) );
  OAI211_X1 U23060 ( .C1(n21396), .C2(n21560), .A(n21395), .B(n21394), .ZN(
        P1_U2835) );
  OAI22_X1 U23061 ( .A1(n21562), .A2(n21398), .B1(n21546), .B2(n21397), .ZN(
        n21399) );
  AOI211_X1 U23062 ( .C1(n21519), .C2(n21400), .A(n21492), .B(n21399), .ZN(
        n21407) );
  OAI21_X1 U23063 ( .B1(n21403), .B2(n21409), .A(n14514), .ZN(n21417) );
  OAI21_X1 U23064 ( .B1(n21403), .B2(n21402), .A(n21401), .ZN(n21404) );
  AOI22_X1 U23065 ( .A1(n21405), .A2(n21568), .B1(n21417), .B2(n21404), .ZN(
        n21406) );
  OAI211_X1 U23066 ( .C1(n21408), .C2(n21560), .A(n21407), .B(n21406), .ZN(
        P1_U2834) );
  AND2_X1 U23067 ( .A1(n21409), .A2(n21528), .ZN(n21421) );
  AOI22_X1 U23068 ( .A1(n21411), .A2(n21519), .B1(n21421), .B2(n21410), .ZN(
        n21419) );
  INV_X1 U23069 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21413) );
  NAND2_X1 U23070 ( .A1(n21551), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n21412) );
  OAI211_X1 U23071 ( .C1(n21413), .C2(n21546), .A(n21412), .B(n21476), .ZN(
        n21416) );
  NOR2_X1 U23072 ( .A1(n21414), .A2(n21553), .ZN(n21415) );
  AOI211_X1 U23073 ( .C1(P1_REIP_REG_7__SCAN_IN), .C2(n21417), .A(n21416), .B(
        n21415), .ZN(n21418) );
  OAI211_X1 U23074 ( .C1(n21420), .C2(n21560), .A(n21419), .B(n21418), .ZN(
        P1_U2833) );
  AOI21_X1 U23075 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n21421), .A(
        P1_REIP_REG_8__SCAN_IN), .ZN(n21430) );
  OAI22_X1 U23076 ( .A1(n21423), .A2(n21572), .B1(n21422), .B2(n21562), .ZN(
        n21424) );
  AOI211_X1 U23077 ( .C1(n21564), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n21492), .B(n21424), .ZN(n21428) );
  AOI22_X1 U23078 ( .A1(n21426), .A2(n21568), .B1(n21425), .B2(n21521), .ZN(
        n21427) );
  OAI211_X1 U23079 ( .C1(n21430), .C2(n21429), .A(n21428), .B(n21427), .ZN(
        P1_U2832) );
  NOR2_X1 U23080 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n21431), .ZN(n21432) );
  AOI22_X1 U23081 ( .A1(n21433), .A2(n21432), .B1(n21551), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n21444) );
  OR2_X1 U23082 ( .A1(n21534), .A2(n21434), .ZN(n21452) );
  OAI22_X1 U23083 ( .A1(n21436), .A2(n21546), .B1(n21435), .B2(n21452), .ZN(
        n21437) );
  AOI211_X1 U23084 ( .C1(n21438), .C2(n21519), .A(n21492), .B(n21437), .ZN(
        n21443) );
  OAI22_X1 U23085 ( .A1(n21440), .A2(n21553), .B1(n21439), .B2(n21560), .ZN(
        n21441) );
  INV_X1 U23086 ( .A(n21441), .ZN(n21442) );
  NAND3_X1 U23087 ( .A1(n21444), .A2(n21443), .A3(n21442), .ZN(P1_U2830) );
  AOI22_X1 U23088 ( .A1(n21551), .A2(P1_EBX_REG_11__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n21564), .ZN(n21445) );
  OAI211_X1 U23089 ( .C1(n21446), .C2(n21572), .A(n21445), .B(n21476), .ZN(
        n21450) );
  OAI22_X1 U23090 ( .A1(n21448), .A2(n21560), .B1(n21553), .B2(n21447), .ZN(
        n21449) );
  NOR2_X1 U23091 ( .A1(n21450), .A2(n21449), .ZN(n21451) );
  OAI221_X1 U23092 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n21454), .C1(n21453), 
        .C2(n21452), .A(n21451), .ZN(P1_U2829) );
  INV_X1 U23093 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21459) );
  AOI22_X1 U23094 ( .A1(n21455), .A2(n21519), .B1(n21551), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n21456) );
  OAI21_X1 U23095 ( .B1(n21459), .B2(n21457), .A(n21456), .ZN(n21458) );
  AOI211_X1 U23096 ( .C1(n21564), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n21492), .B(n21458), .ZN(n21463) );
  AOI22_X1 U23097 ( .A1(n21461), .A2(n21521), .B1(n21460), .B2(n21459), .ZN(
        n21462) );
  OAI211_X1 U23098 ( .C1(n21553), .C2(n21464), .A(n21463), .B(n21462), .ZN(
        P1_U2828) );
  AOI21_X1 U23099 ( .B1(n21564), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n21492), .ZN(n21465) );
  OAI21_X1 U23100 ( .B1(n21560), .B2(n21466), .A(n21465), .ZN(n21467) );
  AOI21_X1 U23101 ( .B1(n21551), .B2(P1_EBX_REG_15__SCAN_IN), .A(n21467), .ZN(
        n21468) );
  OAI21_X1 U23102 ( .B1(n21469), .B2(n21572), .A(n21468), .ZN(n21470) );
  AOI21_X1 U23103 ( .B1(n21471), .B2(n21568), .A(n21470), .ZN(n21472) );
  OAI221_X1 U23104 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n21475), .C1(n21474), 
        .C2(n21473), .A(n21472), .ZN(P1_U2825) );
  NAND2_X1 U23105 ( .A1(n21551), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n21477) );
  OAI211_X1 U23106 ( .C1(n21546), .C2(n21478), .A(n21477), .B(n21476), .ZN(
        n21481) );
  NOR2_X1 U23107 ( .A1(n21479), .A2(n21553), .ZN(n21480) );
  AOI211_X1 U23108 ( .C1(n21521), .C2(n21482), .A(n21481), .B(n21480), .ZN(
        n21485) );
  OAI211_X1 U23109 ( .C1(n21483), .C2(P1_REIP_REG_18__SCAN_IN), .A(n21567), 
        .B(n21488), .ZN(n21484) );
  OAI211_X1 U23110 ( .C1(n21486), .C2(n21572), .A(n21485), .B(n21484), .ZN(
        P1_U2822) );
  NAND2_X1 U23111 ( .A1(n21488), .A2(n21487), .ZN(n21490) );
  INV_X1 U23112 ( .A(n21506), .ZN(n21489) );
  NAND3_X1 U23113 ( .A1(n21490), .A2(n21567), .A3(n21489), .ZN(n21497) );
  INV_X1 U23114 ( .A(n21491), .ZN(n21493) );
  AOI21_X1 U23115 ( .B1(n21521), .B2(n21493), .A(n21492), .ZN(n21496) );
  NAND2_X1 U23116 ( .A1(n21551), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n21495) );
  NAND2_X1 U23117 ( .A1(n21564), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21494) );
  NAND4_X1 U23118 ( .A1(n21497), .A2(n21496), .A3(n21495), .A4(n21494), .ZN(
        n21498) );
  AOI21_X1 U23119 ( .B1(n21499), .B2(n21568), .A(n21498), .ZN(n21500) );
  OAI21_X1 U23120 ( .B1(n21572), .B2(n21501), .A(n21500), .ZN(P1_U2821) );
  AOI22_X1 U23121 ( .A1(n21551), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n21502), 
        .B2(n21521), .ZN(n21508) );
  NAND2_X1 U23122 ( .A1(n21518), .A2(n21567), .ZN(n21517) );
  OAI22_X1 U23123 ( .A1(n21504), .A2(n21553), .B1(n21503), .B2(n21572), .ZN(
        n21505) );
  AOI221_X1 U23124 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n21529), .C1(n21506), 
        .C2(n21529), .A(n21505), .ZN(n21507) );
  OAI211_X1 U23125 ( .C1(n21509), .C2(n21546), .A(n21508), .B(n21507), .ZN(
        P1_U2820) );
  AOI22_X1 U23126 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n21564), .B1(
        n21521), .B2(n21510), .ZN(n21512) );
  NAND2_X1 U23127 ( .A1(n21551), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n21511) );
  OAI211_X1 U23128 ( .C1(n21513), .C2(n21572), .A(n21512), .B(n21511), .ZN(
        n21514) );
  AOI21_X1 U23129 ( .B1(n21515), .B2(n21568), .A(n21514), .ZN(n21516) );
  OAI221_X1 U23130 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n21518), .C1(n21527), 
        .C2(n21517), .A(n21516), .ZN(P1_U2819) );
  AOI22_X1 U23131 ( .A1(n21551), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21564), .ZN(n21533) );
  AOI22_X1 U23132 ( .A1(n21522), .A2(n21521), .B1(n21520), .B2(n21519), .ZN(
        n21532) );
  INV_X1 U23133 ( .A(n21523), .ZN(n21526) );
  AOI22_X1 U23134 ( .A1(n21526), .A2(n21568), .B1(n21525), .B2(n21524), .ZN(
        n21531) );
  OAI221_X1 U23135 ( .B1(n21529), .B2(n21528), .C1(n21529), .C2(n21527), .A(
        P1_REIP_REG_22__SCAN_IN), .ZN(n21530) );
  NAND4_X1 U23136 ( .A1(n21533), .A2(n21532), .A3(n21531), .A4(n21530), .ZN(
        P1_U2818) );
  AOI22_X1 U23137 ( .A1(n21551), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n21564), .ZN(n21542) );
  NOR2_X1 U23138 ( .A1(n21556), .A2(n21534), .ZN(n21557) );
  NAND2_X1 U23139 ( .A1(n21536), .A2(n21535), .ZN(n21540) );
  OAI22_X1 U23140 ( .A1(n21538), .A2(n21553), .B1(n21537), .B2(n21572), .ZN(
        n21539) );
  AOI21_X1 U23141 ( .B1(n21557), .B2(n21540), .A(n21539), .ZN(n21541) );
  OAI211_X1 U23142 ( .C1(n21543), .C2(n21560), .A(n21542), .B(n21541), .ZN(
        P1_U2817) );
  INV_X1 U23143 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21547) );
  INV_X1 U23144 ( .A(n21544), .ZN(n21545) );
  OAI22_X1 U23145 ( .A1(n21547), .A2(n21546), .B1(n21560), .B2(n21545), .ZN(
        n21550) );
  NOR2_X1 U23146 ( .A1(n21548), .A2(n21572), .ZN(n21549) );
  AOI211_X1 U23147 ( .C1(n21551), .C2(P1_EBX_REG_24__SCAN_IN), .A(n21550), .B(
        n21549), .ZN(n21552) );
  OAI21_X1 U23148 ( .B1(n21554), .B2(n21553), .A(n21552), .ZN(n21555) );
  AOI221_X1 U23149 ( .B1(n21557), .B2(P1_REIP_REG_24__SCAN_IN), .C1(n21556), 
        .C2(n16096), .A(n21555), .ZN(n21558) );
  INV_X1 U23150 ( .A(n21558), .ZN(P1_U2816) );
  OAI22_X1 U23151 ( .A1(n21562), .A2(n21561), .B1(n21560), .B2(n21559), .ZN(
        n21563) );
  AOI21_X1 U23152 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n21564), .A(
        n21563), .ZN(n21571) );
  XNOR2_X1 U23153 ( .A(n21565), .B(P1_REIP_REG_25__SCAN_IN), .ZN(n21566) );
  AOI22_X1 U23154 ( .A1(n21569), .A2(n21568), .B1(n21567), .B2(n21566), .ZN(
        n21570) );
  OAI211_X1 U23155 ( .C1(n21573), .C2(n21572), .A(n21571), .B(n21570), .ZN(
        P1_U2815) );
  OAI21_X1 U23156 ( .B1(n21576), .B2(n21575), .A(n21574), .ZN(P1_U2806) );
  INV_X1 U23157 ( .A(n21586), .ZN(n21577) );
  OAI211_X1 U23158 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21667), .A(n21578), 
        .B(n21577), .ZN(n21580) );
  OAI21_X1 U23159 ( .B1(n21581), .B2(n21580), .A(n21579), .ZN(P1_U3163) );
  NOR2_X1 U23160 ( .A1(n21736), .A2(n21582), .ZN(n21583) );
  OAI21_X1 U23161 ( .B1(n21881), .B2(n21584), .A(n21583), .ZN(P1_U3466) );
  INV_X1 U23162 ( .A(n21584), .ZN(n21585) );
  AOI21_X1 U23163 ( .B1(n21587), .B2(n21586), .A(n21585), .ZN(n21588) );
  OAI22_X1 U23164 ( .A1(n21590), .A2(n21589), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n21588), .ZN(n21591) );
  OAI21_X1 U23165 ( .B1(n21593), .B2(n21592), .A(n21591), .ZN(P1_U3161) );
  AOI21_X1 U23166 ( .B1(n17151), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21595), 
        .ZN(n21594) );
  INV_X1 U23167 ( .A(n21594), .ZN(P1_U2805) );
  AOI21_X1 U23168 ( .B1(n17151), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n21595), 
        .ZN(n21596) );
  INV_X1 U23169 ( .A(n21596), .ZN(P1_U3465) );
  OAI21_X1 U23170 ( .B1(n21600), .B2(n21597), .A(n21598), .ZN(P2_U2818) );
  OAI21_X1 U23171 ( .B1(n21600), .B2(n21599), .A(n21598), .ZN(P2_U3592) );
  INV_X1 U23172 ( .A(n21601), .ZN(n21603) );
  OAI21_X1 U23173 ( .B1(n21605), .B2(n21602), .A(n21603), .ZN(P3_U2636) );
  OAI21_X1 U23174 ( .B1(n21605), .B2(n21604), .A(n21603), .ZN(P3_U3281) );
  INV_X1 U23175 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21644) );
  AOI21_X1 U23176 ( .B1(HOLD), .B2(n21606), .A(n21644), .ZN(n21608) );
  NAND2_X1 U23177 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n21607), .ZN(n21643) );
  INV_X1 U23178 ( .A(n21643), .ZN(n21656) );
  NOR2_X1 U23179 ( .A1(n21656), .A2(n21645), .ZN(n21660) );
  AOI21_X1 U23180 ( .B1(n21649), .B2(NA), .A(n21654), .ZN(n21658) );
  OAI22_X1 U23181 ( .A1(n18364), .A2(n21608), .B1(n21660), .B2(n21658), .ZN(
        P3_U3029) );
  AOI21_X1 U23182 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n21611), .A(n21653), .ZN(n21609) );
  AOI21_X1 U23183 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(
        P1_STATE_REG_1__SCAN_IN), .A(n21609), .ZN(n21613) );
  AOI22_X1 U23184 ( .A1(n21616), .A2(n21655), .B1(n21609), .B2(n21619), .ZN(
        n21612) );
  NOR2_X1 U23185 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21655), .ZN(n21610) );
  AOI21_X1 U23186 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21616), .A(n21614), 
        .ZN(n21623) );
  OAI33_X1 U23187 ( .A1(n21614), .A2(n21613), .A3(n21612), .B1(n21611), .B2(
        n21610), .B3(n21623), .ZN(P1_U3196) );
  AOI21_X1 U23188 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(HOLD), .A(n21615), .ZN(
        n21620) );
  AOI22_X1 U23189 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21616), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(n21620), .ZN(n21618) );
  OAI211_X1 U23190 ( .C1(n21619), .C2(n21653), .A(n21618), .B(n21617), .ZN(
        P1_U3195) );
  OAI21_X1 U23191 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21655), .A(n21620), 
        .ZN(n21621) );
  AOI21_X1 U23192 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(n21621), .ZN(
        n21622) );
  OAI22_X1 U23193 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21623), .B1(n22328), 
        .B2(n21622), .ZN(P1_U3194) );
  NAND2_X1 U23194 ( .A1(n21624), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21636) );
  NAND2_X1 U23195 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21636), .ZN(n21635) );
  NOR2_X1 U23196 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21655), .ZN(n21626) );
  AOI211_X1 U23197 ( .C1(n21640), .C2(n21635), .A(n21626), .B(n21625), .ZN(
        n21628) );
  AOI221_X1 U23198 ( .B1(n21629), .B2(n21628), .C1(n21653), .C2(n21628), .A(
        n21627), .ZN(P2_U3209) );
  INV_X1 U23199 ( .A(n21630), .ZN(n21634) );
  OAI211_X1 U23200 ( .C1(n21640), .C2(n21653), .A(P2_STATE_REG_0__SCAN_IN), 
        .B(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21633) );
  NAND2_X1 U23201 ( .A1(n21631), .A2(HOLD), .ZN(n21632) );
  NAND4_X1 U23202 ( .A1(n21634), .A2(n21633), .A3(n21636), .A4(n21632), .ZN(
        P2_U3210) );
  OAI22_X1 U23203 ( .A1(HOLD), .A2(n21635), .B1(P2_STATE_REG_0__SCAN_IN), .B2(
        n21655), .ZN(n21641) );
  OAI22_X1 U23204 ( .A1(NA), .A2(n21636), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21637) );
  OAI211_X1 U23205 ( .C1(HOLD), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n21637), .ZN(n21639) );
  OAI211_X1 U23206 ( .C1(n21641), .C2(n21640), .A(n21639), .B(n21638), .ZN(
        P2_U3211) );
  NOR2_X1 U23207 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21662)
         );
  NAND2_X1 U23208 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n21654), .ZN(n21642) );
  AOI221_X1 U23209 ( .B1(n21662), .B2(n21643), .C1(n21642), .C2(n21643), .A(
        n21648), .ZN(n21647) );
  AOI211_X1 U23210 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n21645), .B(
        n21644), .ZN(n21646) );
  AOI211_X1 U23211 ( .C1(n21649), .C2(n21648), .A(n21647), .B(n21646), .ZN(
        n21650) );
  OAI211_X1 U23212 ( .C1(n21652), .C2(n21651), .A(n21650), .B(n18365), .ZN(
        P3_U3030) );
  OAI22_X1 U23213 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n21654), .B2(n21653), .ZN(n21657)
         );
  OAI221_X1 U23214 ( .B1(n21657), .B2(n21656), .C1(n21657), .C2(n21655), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n21661) );
  INV_X1 U23215 ( .A(n21658), .ZN(n21659) );
  OAI22_X1 U23216 ( .A1(n21662), .A2(n21661), .B1(n21660), .B2(n21659), .ZN(
        P3_U3031) );
  INV_X1 U23217 ( .A(n21663), .ZN(n21664) );
  INV_X1 U23218 ( .A(n21665), .ZN(n21666) );
  OAI21_X2 U23219 ( .B1(n13547), .B2(n21667), .A(n21666), .ZN(n21718) );
  AOI22_X1 U23220 ( .A1(n21722), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n21721), .ZN(n21668) );
  OAI21_X1 U23221 ( .B1(n21729), .B2(n21724), .A(n21668), .ZN(P1_U2937) );
  AOI22_X1 U23222 ( .A1(n21718), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(
        P1_EAX_REG_0__SCAN_IN), .B2(n21721), .ZN(n21669) );
  OAI21_X1 U23223 ( .B1(n21729), .B2(n21724), .A(n21669), .ZN(P1_U2952) );
  AOI22_X1 U23224 ( .A1(n21718), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n21721), .ZN(n21670) );
  OAI21_X1 U23225 ( .B1(n21933), .B2(n21724), .A(n21670), .ZN(P1_U2938) );
  AOI22_X1 U23226 ( .A1(n21718), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(
        P1_EAX_REG_1__SCAN_IN), .B2(n21721), .ZN(n21671) );
  OAI21_X1 U23227 ( .B1(n21933), .B2(n21724), .A(n21671), .ZN(P1_U2953) );
  AOI22_X1 U23228 ( .A1(n21722), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n21721), .ZN(n21672) );
  OAI21_X1 U23229 ( .B1(n21976), .B2(n21724), .A(n21672), .ZN(P1_U2939) );
  AOI22_X1 U23230 ( .A1(n21722), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(
        P1_EAX_REG_2__SCAN_IN), .B2(n21721), .ZN(n21673) );
  OAI21_X1 U23231 ( .B1(n21976), .B2(n21724), .A(n21673), .ZN(P1_U2954) );
  AOI22_X1 U23232 ( .A1(n21722), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n21721), .ZN(n21674) );
  OAI21_X1 U23233 ( .B1(n22022), .B2(n21724), .A(n21674), .ZN(P1_U2940) );
  AOI22_X1 U23234 ( .A1(n21722), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(
        P1_EAX_REG_3__SCAN_IN), .B2(n21721), .ZN(n21675) );
  OAI21_X1 U23235 ( .B1(n22022), .B2(n21724), .A(n21675), .ZN(P1_U2955) );
  AOI22_X1 U23236 ( .A1(n21722), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n21721), .ZN(n21676) );
  OAI21_X1 U23237 ( .B1(n22068), .B2(n21724), .A(n21676), .ZN(P1_U2941) );
  AOI22_X1 U23238 ( .A1(n21722), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(
        P1_EAX_REG_4__SCAN_IN), .B2(n21721), .ZN(n21677) );
  OAI21_X1 U23239 ( .B1(n22068), .B2(n21724), .A(n21677), .ZN(P1_U2956) );
  AOI22_X1 U23240 ( .A1(n21722), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n21721), .ZN(n21678) );
  OAI21_X1 U23241 ( .B1(n22114), .B2(n21724), .A(n21678), .ZN(P1_U2942) );
  AOI22_X1 U23242 ( .A1(n21722), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(
        P1_EAX_REG_5__SCAN_IN), .B2(n21721), .ZN(n21679) );
  OAI21_X1 U23243 ( .B1(n22114), .B2(n21724), .A(n21679), .ZN(P1_U2957) );
  AOI22_X1 U23244 ( .A1(n21722), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n21721), .ZN(n21680) );
  OAI21_X1 U23245 ( .B1(n22164), .B2(n21724), .A(n21680), .ZN(P1_U2943) );
  AOI22_X1 U23246 ( .A1(n21722), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(
        P1_EAX_REG_6__SCAN_IN), .B2(n21721), .ZN(n21681) );
  OAI21_X1 U23247 ( .B1(n22164), .B2(n21724), .A(n21681), .ZN(P1_U2958) );
  AOI22_X1 U23248 ( .A1(n21722), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n21721), .ZN(n21682) );
  OAI21_X1 U23249 ( .B1(n22211), .B2(n21724), .A(n21682), .ZN(P1_U2944) );
  AOI22_X1 U23250 ( .A1(n21722), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(
        P1_EAX_REG_7__SCAN_IN), .B2(n21721), .ZN(n21683) );
  OAI21_X1 U23251 ( .B1(n22211), .B2(n21724), .A(n21683), .ZN(P1_U2959) );
  NOR2_X1 U23252 ( .A1(n21724), .A2(n21684), .ZN(n21687) );
  AOI21_X1 U23253 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n21722), .A(n21687), 
        .ZN(n21685) );
  OAI21_X1 U23254 ( .B1(n21686), .B2(n21720), .A(n21685), .ZN(P1_U2945) );
  AOI21_X1 U23255 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n21722), .A(n21687), 
        .ZN(n21688) );
  OAI21_X1 U23256 ( .B1(n15351), .B2(n21720), .A(n21688), .ZN(P1_U2960) );
  NOR2_X1 U23257 ( .A1(n21724), .A2(n21689), .ZN(n21692) );
  AOI21_X1 U23258 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n21722), .A(n21692), 
        .ZN(n21690) );
  OAI21_X1 U23259 ( .B1(n21691), .B2(n21720), .A(n21690), .ZN(P1_U2946) );
  AOI21_X1 U23260 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(n21722), .A(n21692), 
        .ZN(n21693) );
  OAI21_X1 U23261 ( .B1(n15449), .B2(n21720), .A(n21693), .ZN(P1_U2961) );
  NOR2_X1 U23262 ( .A1(n21724), .A2(n21694), .ZN(n21697) );
  AOI21_X1 U23263 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n21718), .A(n21697), 
        .ZN(n21695) );
  OAI21_X1 U23264 ( .B1(n21696), .B2(n21720), .A(n21695), .ZN(P1_U2947) );
  AOI21_X1 U23265 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n21722), .A(n21697), 
        .ZN(n21698) );
  OAI21_X1 U23266 ( .B1(n15462), .B2(n21720), .A(n21698), .ZN(P1_U2962) );
  NOR2_X1 U23267 ( .A1(n21724), .A2(n21699), .ZN(n21702) );
  AOI21_X1 U23268 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n21718), .A(n21702), 
        .ZN(n21700) );
  OAI21_X1 U23269 ( .B1(n21701), .B2(n21720), .A(n21700), .ZN(P1_U2948) );
  AOI21_X1 U23270 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(n21718), .A(n21702), 
        .ZN(n21703) );
  OAI21_X1 U23271 ( .B1(n15550), .B2(n21720), .A(n21703), .ZN(P1_U2963) );
  NOR2_X1 U23272 ( .A1(n21724), .A2(n21704), .ZN(n21707) );
  AOI21_X1 U23273 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n21718), .A(n21707), 
        .ZN(n21705) );
  OAI21_X1 U23274 ( .B1(n21706), .B2(n21720), .A(n21705), .ZN(P1_U2949) );
  AOI21_X1 U23275 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n21718), .A(n21707), 
        .ZN(n21708) );
  OAI21_X1 U23276 ( .B1(n15597), .B2(n21720), .A(n21708), .ZN(P1_U2964) );
  NOR2_X1 U23277 ( .A1(n21724), .A2(n21709), .ZN(n21712) );
  AOI21_X1 U23278 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n21718), .A(n21712), 
        .ZN(n21710) );
  OAI21_X1 U23279 ( .B1(n21711), .B2(n21720), .A(n21710), .ZN(P1_U2950) );
  AOI21_X1 U23280 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n21718), .A(n21712), 
        .ZN(n21713) );
  OAI21_X1 U23281 ( .B1(n15590), .B2(n21720), .A(n21713), .ZN(P1_U2965) );
  NOR2_X1 U23282 ( .A1(n21724), .A2(n21714), .ZN(n21717) );
  AOI21_X1 U23283 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n21718), .A(n21717), 
        .ZN(n21715) );
  OAI21_X1 U23284 ( .B1(n21716), .B2(n21720), .A(n21715), .ZN(P1_U2951) );
  AOI21_X1 U23285 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(n21718), .A(n21717), 
        .ZN(n21719) );
  OAI21_X1 U23286 ( .B1(n15621), .B2(n21720), .A(n21719), .ZN(P1_U2966) );
  AOI22_X1 U23287 ( .A1(n21722), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(
        P1_EAX_REG_15__SCAN_IN), .B2(n21721), .ZN(n21723) );
  OAI21_X1 U23288 ( .B1(n21725), .B2(n21724), .A(n21723), .ZN(P1_U2967) );
  INV_X1 U23289 ( .A(n22322), .ZN(n21726) );
  NAND2_X1 U23290 ( .A1(n21726), .A2(n21868), .ZN(n21727) );
  OAI21_X1 U23291 ( .B1(n21727), .B2(n22227), .A(n21869), .ZN(n21743) );
  INV_X1 U23292 ( .A(n21872), .ZN(n21728) );
  OR2_X1 U23293 ( .A1(n21823), .A2(n21728), .ZN(n21761) );
  NOR2_X1 U23294 ( .A1(n21761), .A2(n21903), .ZN(n21740) );
  NOR2_X1 U23295 ( .A1(n21738), .A2(n21917), .ZN(n21843) );
  INV_X1 U23296 ( .A(n21762), .ZN(n21841) );
  OR2_X1 U23297 ( .A1(n21824), .A2(n21841), .ZN(n21786) );
  INV_X1 U23298 ( .A(n21786), .ZN(n21745) );
  INV_X1 U23299 ( .A(n21922), .ZN(n21884) );
  INV_X1 U23300 ( .A(DATAI_24_), .ZN(n21733) );
  OAI22_X2 U23301 ( .A1(n21734), .A2(n22219), .B1(n21733), .B2(n22217), .ZN(
        n21909) );
  NOR2_X2 U23302 ( .A1(n22215), .A2(n21737), .ZN(n21921) );
  NOR3_X1 U23303 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21756) );
  INV_X1 U23304 ( .A(n21756), .ZN(n21753) );
  NOR2_X1 U23305 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21753), .ZN(
        n22216) );
  AOI22_X1 U23306 ( .A1(n22322), .A2(n21909), .B1(n21921), .B2(n22216), .ZN(
        n21749) );
  INV_X1 U23307 ( .A(n21738), .ZN(n21739) );
  NOR2_X1 U23308 ( .A1(n21739), .A2(n21917), .ZN(n21874) );
  NOR2_X1 U23309 ( .A1(n21874), .A2(n22212), .ZN(n21849) );
  INV_X1 U23310 ( .A(n21740), .ZN(n21742) );
  INV_X1 U23311 ( .A(n22216), .ZN(n21741) );
  AOI22_X1 U23312 ( .A1(n21743), .A2(n21742), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21741), .ZN(n21744) );
  OAI211_X1 U23313 ( .C1(n21745), .C2(n21917), .A(n21849), .B(n21744), .ZN(
        n22221) );
  AOI22_X1 U23314 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22221), .B1(
        n22227), .B2(n21929), .ZN(n21748) );
  OAI211_X1 U23315 ( .C1(n22224), .C2(n21884), .A(n21749), .B(n21748), .ZN(
        P1_U3033) );
  INV_X1 U23316 ( .A(n21929), .ZN(n21912) );
  INV_X1 U23317 ( .A(n21761), .ZN(n21774) );
  INV_X1 U23318 ( .A(n21752), .ZN(n21886) );
  NOR2_X1 U23319 ( .A1(n21885), .A2(n21753), .ZN(n22225) );
  AOI21_X1 U23320 ( .B1(n21774), .B2(n21886), .A(n22225), .ZN(n21754) );
  OAI22_X1 U23321 ( .A1(n21754), .A2(n21923), .B1(n21753), .B2(n21917), .ZN(
        n22226) );
  AOI22_X1 U23322 ( .A1(n22226), .A2(n21922), .B1(n21921), .B2(n22225), .ZN(
        n21758) );
  OAI211_X1 U23323 ( .C1(n21781), .C2(n21900), .A(n21896), .B(n21754), .ZN(
        n21755) );
  OAI211_X1 U23324 ( .C1(n21868), .C2(n21756), .A(n21926), .B(n21755), .ZN(
        n22228) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22228), .B1(
        n22227), .B2(n21909), .ZN(n21757) );
  OAI211_X1 U23326 ( .C1(n21912), .C2(n22231), .A(n21758), .B(n21757), .ZN(
        P1_U3041) );
  NAND2_X1 U23327 ( .A1(n22231), .A2(n21896), .ZN(n21760) );
  OAI21_X1 U23328 ( .B1(n22239), .B2(n21760), .A(n21869), .ZN(n21764) );
  NOR2_X1 U23329 ( .A1(n21761), .A2(n15264), .ZN(n21766) );
  NOR2_X1 U23330 ( .A1(n21762), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21801) );
  NOR3_X1 U23331 ( .A1(n21763), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21770) );
  NAND2_X1 U23332 ( .A1(n21885), .A2(n21770), .ZN(n22125) );
  INV_X1 U23333 ( .A(n22125), .ZN(n22232) );
  AOI22_X1 U23334 ( .A1(n22239), .A2(n21929), .B1(n21921), .B2(n22232), .ZN(
        n21769) );
  INV_X1 U23335 ( .A(n21764), .ZN(n21767) );
  NOR2_X1 U23336 ( .A1(n21801), .A2(n21917), .ZN(n21803) );
  AOI21_X1 U23337 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22125), .A(n21803), 
        .ZN(n21765) );
  OAI211_X1 U23338 ( .C1(n21767), .C2(n21766), .A(n21765), .B(n21849), .ZN(
        n22234) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22234), .B1(
        n22233), .B2(n21909), .ZN(n21768) );
  OAI211_X1 U23340 ( .C1(n22237), .C2(n21884), .A(n21769), .B(n21768), .ZN(
        P1_U3049) );
  INV_X1 U23341 ( .A(n21770), .ZN(n21777) );
  INV_X1 U23342 ( .A(n21771), .ZN(n21773) );
  NAND2_X1 U23343 ( .A1(n21773), .A2(n21772), .ZN(n21914) );
  INV_X1 U23344 ( .A(n21914), .ZN(n21812) );
  NOR2_X1 U23345 ( .A1(n21885), .A2(n21777), .ZN(n22238) );
  AOI21_X1 U23346 ( .B1(n21774), .B2(n21812), .A(n22238), .ZN(n21776) );
  AOI21_X1 U23347 ( .B1(n21781), .B2(n21868), .A(n21858), .ZN(n21780) );
  OAI22_X1 U23348 ( .A1(n21917), .A2(n21777), .B1(n21776), .B2(n21780), .ZN(
        n21775) );
  AOI22_X1 U23349 ( .A1(n22239), .A2(n21909), .B1(n22238), .B2(n21921), .ZN(
        n21783) );
  INV_X1 U23350 ( .A(n21776), .ZN(n21779) );
  INV_X1 U23351 ( .A(n21926), .ZN(n21860) );
  AOI21_X1 U23352 ( .B1(n21923), .B2(n21777), .A(n21860), .ZN(n21778) );
  OAI21_X1 U23353 ( .B1(n21780), .B2(n21779), .A(n21778), .ZN(n22240) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n22240), .B1(
        n22246), .B2(n21929), .ZN(n21782) );
  OAI211_X1 U23355 ( .C1(n22243), .C2(n21884), .A(n21783), .B(n21782), .ZN(
        P1_U3057) );
  NOR3_X1 U23356 ( .A1(n21875), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21796) );
  INV_X1 U23357 ( .A(n21796), .ZN(n21793) );
  NOR2_X1 U23358 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21793), .ZN(
        n22245) );
  INV_X1 U23359 ( .A(n21874), .ZN(n21899) );
  NOR2_X1 U23360 ( .A1(n21872), .A2(n21784), .ZN(n21813) );
  NAND3_X1 U23361 ( .A1(n21813), .A2(n21896), .A3(n15264), .ZN(n21785) );
  OAI21_X1 U23362 ( .B1(n21899), .B2(n21786), .A(n21785), .ZN(n22244) );
  AOI22_X1 U23363 ( .A1(n21921), .A2(n22245), .B1(n22244), .B2(n21922), .ZN(
        n21792) );
  INV_X1 U23364 ( .A(n22246), .ZN(n21787) );
  AOI21_X1 U23365 ( .B1(n21787), .B2(n22255), .A(n21900), .ZN(n21788) );
  AOI21_X1 U23366 ( .B1(n21813), .B2(n15264), .A(n21788), .ZN(n21789) );
  NOR2_X1 U23367 ( .A1(n21789), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21790) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n22247), .B1(
        n22246), .B2(n21909), .ZN(n21791) );
  OAI211_X1 U23369 ( .C1(n21912), .C2(n22255), .A(n21792), .B(n21791), .ZN(
        P1_U3065) );
  INV_X1 U23370 ( .A(n21909), .ZN(n21932) );
  NOR2_X1 U23371 ( .A1(n21885), .A2(n21793), .ZN(n22250) );
  AOI21_X1 U23372 ( .B1(n21813), .B2(n21886), .A(n22250), .ZN(n21794) );
  OAI22_X1 U23373 ( .A1(n21794), .A2(n21923), .B1(n21793), .B2(n21917), .ZN(
        n22251) );
  AOI22_X1 U23374 ( .A1(n22251), .A2(n21922), .B1(n21921), .B2(n22250), .ZN(
        n21798) );
  OAI21_X1 U23375 ( .B1(n21810), .B2(n21900), .A(n21794), .ZN(n21795) );
  OAI221_X1 U23376 ( .B1(n21868), .B2(n21796), .C1(n21923), .C2(n21795), .A(
        n21926), .ZN(n22252) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n22252), .B1(
        n22257), .B2(n21929), .ZN(n21797) );
  OAI211_X1 U23378 ( .C1(n21932), .C2(n22255), .A(n21798), .B(n21797), .ZN(
        P1_U3073) );
  INV_X1 U23379 ( .A(n22257), .ZN(n21799) );
  NAND2_X1 U23380 ( .A1(n21799), .A2(n21896), .ZN(n21800) );
  OAI21_X1 U23381 ( .B1(n21800), .B2(n22264), .A(n21869), .ZN(n21805) );
  AND2_X1 U23382 ( .A1(n21813), .A2(n21903), .ZN(n21802) );
  INV_X1 U23383 ( .A(n21916), .ZN(n21924) );
  NOR3_X2 U23384 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n21924), .ZN(n22256) );
  AOI22_X1 U23385 ( .A1(n22257), .A2(n21909), .B1(n21921), .B2(n22256), .ZN(
        n21808) );
  INV_X1 U23386 ( .A(n21802), .ZN(n21804) );
  AOI21_X1 U23387 ( .B1(n21805), .B2(n21804), .A(n21803), .ZN(n21806) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n22258), .B1(
        n22264), .B2(n21929), .ZN(n21807) );
  OAI211_X1 U23389 ( .C1(n22261), .C2(n21884), .A(n21808), .B(n21807), .ZN(
        P1_U3081) );
  INV_X1 U23390 ( .A(n21811), .ZN(n22262) );
  AOI21_X1 U23391 ( .B1(n21813), .B2(n21812), .A(n22262), .ZN(n21815) );
  NOR2_X1 U23392 ( .A1(n21924), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21817) );
  INV_X1 U23393 ( .A(n21817), .ZN(n21814) );
  OAI22_X1 U23394 ( .A1(n21815), .A2(n21923), .B1(n21814), .B2(n21917), .ZN(
        n22263) );
  AOI22_X1 U23395 ( .A1(n22263), .A2(n21922), .B1(n22262), .B2(n21921), .ZN(
        n21819) );
  OAI21_X1 U23396 ( .B1(n21817), .B2(n21816), .A(n21926), .ZN(n22265) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n21909), .ZN(n21818) );
  OAI211_X1 U23398 ( .C1(n21912), .C2(n22268), .A(n21819), .B(n21818), .ZN(
        P1_U3089) );
  INV_X1 U23399 ( .A(n21867), .ZN(n21822) );
  AND2_X1 U23400 ( .A1(n21823), .A2(n21872), .ZN(n21854) );
  NOR3_X1 U23401 ( .A1(n13778), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21836) );
  INV_X1 U23402 ( .A(n21836), .ZN(n21833) );
  NOR2_X1 U23403 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21833), .ZN(
        n22269) );
  AOI21_X1 U23404 ( .B1(n21854), .B2(n15264), .A(n22269), .ZN(n21828) );
  INV_X1 U23405 ( .A(n21843), .ZN(n21826) );
  INV_X1 U23406 ( .A(n21824), .ZN(n21825) );
  NOR2_X1 U23407 ( .A1(n21825), .A2(n21841), .ZN(n21873) );
  INV_X1 U23408 ( .A(n21873), .ZN(n21877) );
  OAI22_X1 U23409 ( .A1(n21828), .A2(n21923), .B1(n21826), .B2(n21877), .ZN(
        n22270) );
  AOI22_X1 U23410 ( .A1(n22270), .A2(n21922), .B1(n21921), .B2(n22269), .ZN(
        n21832) );
  INV_X1 U23411 ( .A(n22280), .ZN(n21827) );
  OAI21_X1 U23412 ( .B1(n21827), .B2(n22271), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21829) );
  NAND2_X1 U23413 ( .A1(n21829), .A2(n21828), .ZN(n21830) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n22272), .B1(
        n22271), .B2(n21909), .ZN(n21831) );
  OAI211_X1 U23415 ( .C1(n21912), .C2(n22280), .A(n21832), .B(n21831), .ZN(
        P1_U3097) );
  NOR2_X1 U23416 ( .A1(n21885), .A2(n21833), .ZN(n22275) );
  AOI21_X1 U23417 ( .B1(n21854), .B2(n21886), .A(n22275), .ZN(n21834) );
  OAI22_X1 U23418 ( .A1(n21834), .A2(n21923), .B1(n21833), .B2(n21917), .ZN(
        n22276) );
  AOI22_X1 U23419 ( .A1(n22276), .A2(n21922), .B1(n21921), .B2(n22275), .ZN(
        n21838) );
  OAI211_X1 U23420 ( .C1(n21859), .C2(n21900), .A(n21896), .B(n21834), .ZN(
        n21835) );
  OAI211_X1 U23421 ( .C1(n21896), .C2(n21836), .A(n21926), .B(n21835), .ZN(
        n22277) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22277), .B1(
        n22282), .B2(n21929), .ZN(n21837) );
  OAI211_X1 U23423 ( .C1(n21932), .C2(n22280), .A(n21838), .B(n21837), .ZN(
        P1_U3105) );
  INV_X1 U23424 ( .A(n22282), .ZN(n21839) );
  NAND2_X1 U23425 ( .A1(n21839), .A2(n21868), .ZN(n21840) );
  OAI21_X1 U23426 ( .B1(n21840), .B2(n22289), .A(n21869), .ZN(n21847) );
  AND2_X1 U23427 ( .A1(n21854), .A2(n21903), .ZN(n21844) );
  NAND2_X1 U23428 ( .A1(n21841), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21898) );
  INV_X1 U23429 ( .A(n21898), .ZN(n21842) );
  NAND3_X1 U23430 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n21875), .ZN(n21861) );
  NOR2_X1 U23431 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21861), .ZN(
        n22281) );
  AOI22_X1 U23432 ( .A1(n22282), .A2(n21909), .B1(n21921), .B2(n22281), .ZN(
        n21851) );
  INV_X1 U23433 ( .A(n21844), .ZN(n21846) );
  INV_X1 U23434 ( .A(n22281), .ZN(n21845) );
  AOI22_X1 U23435 ( .A1(n21847), .A2(n21846), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21845), .ZN(n21848) );
  NAND2_X1 U23436 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21898), .ZN(n21906) );
  NAND3_X1 U23437 ( .A1(n21849), .A2(n21848), .A3(n21906), .ZN(n22283) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n21929), .ZN(n21850) );
  OAI211_X1 U23439 ( .C1(n22286), .C2(n21884), .A(n21851), .B(n21850), .ZN(
        P1_U3113) );
  INV_X1 U23440 ( .A(n21854), .ZN(n21856) );
  NOR2_X1 U23441 ( .A1(n21885), .A2(n21861), .ZN(n22287) );
  INV_X1 U23442 ( .A(n22287), .ZN(n21855) );
  OAI21_X1 U23443 ( .B1(n21856), .B2(n21914), .A(n21855), .ZN(n21863) );
  INV_X1 U23444 ( .A(n21863), .ZN(n21857) );
  OAI22_X1 U23445 ( .A1(n21857), .A2(n21923), .B1(n21861), .B2(n21917), .ZN(
        n22288) );
  AOI22_X1 U23446 ( .A1(n22288), .A2(n21922), .B1(n21921), .B2(n22287), .ZN(
        n21866) );
  AOI21_X1 U23447 ( .B1(n21859), .B2(n21896), .A(n21858), .ZN(n21864) );
  AOI21_X1 U23448 ( .B1(n21861), .B2(n21923), .A(n21860), .ZN(n21862) );
  OAI21_X1 U23449 ( .B1(n21864), .B2(n21863), .A(n21862), .ZN(n22290) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n21909), .ZN(n21865) );
  OAI211_X1 U23451 ( .C1(n21912), .C2(n22293), .A(n21866), .B(n21865), .ZN(
        P1_U3121) );
  NAND3_X1 U23452 ( .A1(n22293), .A2(n21868), .A3(n22308), .ZN(n21870) );
  NAND2_X1 U23453 ( .A1(n21870), .A2(n21869), .ZN(n21879) );
  NOR2_X1 U23454 ( .A1(n21915), .A2(n21903), .ZN(n21876) );
  INV_X1 U23455 ( .A(n22308), .ZN(n22148) );
  NOR3_X1 U23456 ( .A1(n21875), .A2(n13778), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21890) );
  INV_X1 U23457 ( .A(n21890), .ZN(n21887) );
  NOR2_X1 U23458 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21887), .ZN(
        n22147) );
  AOI22_X1 U23459 ( .A1(n22148), .A2(n21929), .B1(n21921), .B2(n22147), .ZN(
        n21883) );
  INV_X1 U23460 ( .A(n21876), .ZN(n21878) );
  AOI22_X1 U23461 ( .A1(n21879), .A2(n21878), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21877), .ZN(n21880) );
  OAI211_X1 U23462 ( .C1(n22147), .C2(n21881), .A(n21907), .B(n21880), .ZN(
        n22298) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n22298), .B1(
        n22297), .B2(n21909), .ZN(n21882) );
  OAI211_X1 U23464 ( .C1(n22302), .C2(n21884), .A(n21883), .B(n21882), .ZN(
        P1_U3129) );
  NOR2_X1 U23465 ( .A1(n21885), .A2(n21887), .ZN(n22303) );
  AOI21_X1 U23466 ( .B1(n21904), .B2(n21886), .A(n22303), .ZN(n21888) );
  OAI22_X1 U23467 ( .A1(n21888), .A2(n21923), .B1(n21887), .B2(n21917), .ZN(
        n22304) );
  AOI22_X1 U23468 ( .A1(n22304), .A2(n21922), .B1(n21921), .B2(n22303), .ZN(
        n21893) );
  OAI211_X1 U23469 ( .C1(n21895), .C2(n21900), .A(n21896), .B(n21888), .ZN(
        n21889) );
  OAI211_X1 U23470 ( .C1(n21896), .C2(n21890), .A(n21926), .B(n21889), .ZN(
        n22305) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22305), .B1(
        n22312), .B2(n21929), .ZN(n21892) );
  OAI211_X1 U23472 ( .C1(n21932), .C2(n22308), .A(n21893), .B(n21892), .ZN(
        P1_U3137) );
  NOR3_X2 U23473 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13778), .A3(
        n21924), .ZN(n22310) );
  NAND3_X1 U23474 ( .A1(n21904), .A2(n21903), .A3(n21896), .ZN(n21897) );
  OAI21_X1 U23475 ( .B1(n21899), .B2(n21898), .A(n21897), .ZN(n22309) );
  AOI22_X1 U23476 ( .A1(n21921), .A2(n22310), .B1(n22309), .B2(n21922), .ZN(
        n21911) );
  INV_X1 U23477 ( .A(n22312), .ZN(n21901) );
  AOI21_X1 U23478 ( .B1(n21901), .B2(n22326), .A(n21900), .ZN(n21902) );
  AOI21_X1 U23479 ( .B1(n21904), .B2(n21903), .A(n21902), .ZN(n21905) );
  NOR2_X1 U23480 ( .A1(n21905), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21908) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n21909), .ZN(n21910) );
  OAI211_X1 U23482 ( .C1(n21912), .C2(n22326), .A(n21911), .B(n21910), .ZN(
        P1_U3145) );
  NAND2_X1 U23483 ( .A1(n21913), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21920) );
  OAI21_X1 U23484 ( .B1(n21915), .B2(n21914), .A(n21920), .ZN(n21927) );
  INV_X1 U23485 ( .A(n21927), .ZN(n21919) );
  NAND2_X1 U23486 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21916), .ZN(
        n21918) );
  OAI22_X1 U23487 ( .A1(n21919), .A2(n21923), .B1(n21918), .B2(n21917), .ZN(
        n22320) );
  INV_X1 U23488 ( .A(n21920), .ZN(n22317) );
  AOI22_X1 U23489 ( .A1(n22320), .A2(n21922), .B1(n21921), .B2(n22317), .ZN(
        n21931) );
  OAI21_X1 U23490 ( .B1(n21924), .B2(n13778), .A(n21923), .ZN(n21925) );
  OAI211_X1 U23491 ( .C1(n21928), .C2(n21927), .A(n21926), .B(n21925), .ZN(
        n22323) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n22323), .B1(
        n22322), .B2(n21929), .ZN(n21930) );
  OAI211_X1 U23493 ( .C1(n21932), .C2(n22326), .A(n21931), .B(n21930), .ZN(
        P1_U3153) );
  INV_X1 U23494 ( .A(DATAI_25_), .ZN(n21934) );
  OAI22_X2 U23495 ( .A1(n16549), .A2(n22219), .B1(n21934), .B2(n22217), .ZN(
        n21967) );
  NOR2_X2 U23496 ( .A1(n22215), .A2(n21935), .ZN(n21970) );
  AOI22_X1 U23497 ( .A1(n22322), .A2(n21967), .B1(n21970), .B2(n22216), .ZN(
        n21939) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22221), .B1(
        n22227), .B2(n21972), .ZN(n21938) );
  OAI211_X1 U23499 ( .C1(n22224), .C2(n21964), .A(n21939), .B(n21938), .ZN(
        P1_U3034) );
  AOI22_X1 U23500 ( .A1(n22226), .A2(n21971), .B1(n21970), .B2(n22225), .ZN(
        n21941) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22228), .B1(
        n22227), .B2(n21967), .ZN(n21940) );
  OAI211_X1 U23502 ( .C1(n11106), .C2(n22231), .A(n21941), .B(n21940), .ZN(
        P1_U3042) );
  AOI22_X1 U23503 ( .A1(n22239), .A2(n21972), .B1(n21970), .B2(n22232), .ZN(
        n21943) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n22234), .B1(
        n22233), .B2(n21967), .ZN(n21942) );
  OAI211_X1 U23505 ( .C1(n22237), .C2(n21964), .A(n21943), .B(n21942), .ZN(
        P1_U3050) );
  AOI22_X1 U23506 ( .A1(n22246), .A2(n21972), .B1(n21970), .B2(n22238), .ZN(
        n21945) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n21967), .ZN(n21944) );
  OAI211_X1 U23508 ( .C1(n22243), .C2(n21964), .A(n21945), .B(n21944), .ZN(
        P1_U3058) );
  AOI22_X1 U23509 ( .A1(n21970), .A2(n22245), .B1(n22244), .B2(n21971), .ZN(
        n21947) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n22247), .B1(
        n22246), .B2(n21967), .ZN(n21946) );
  OAI211_X1 U23511 ( .C1(n11106), .C2(n22255), .A(n21947), .B(n21946), .ZN(
        P1_U3066) );
  INV_X1 U23512 ( .A(n21967), .ZN(n21975) );
  AOI22_X1 U23513 ( .A1(n22251), .A2(n21971), .B1(n21970), .B2(n22250), .ZN(
        n21949) );
  AOI22_X1 U23514 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n22252), .B1(
        n22257), .B2(n21972), .ZN(n21948) );
  OAI211_X1 U23515 ( .C1(n21975), .C2(n22255), .A(n21949), .B(n21948), .ZN(
        P1_U3074) );
  AOI22_X1 U23516 ( .A1(n22257), .A2(n21967), .B1(n21970), .B2(n22256), .ZN(
        n21951) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n22258), .B1(
        n22264), .B2(n21972), .ZN(n21950) );
  OAI211_X1 U23518 ( .C1(n22261), .C2(n21964), .A(n21951), .B(n21950), .ZN(
        P1_U3082) );
  AOI22_X1 U23519 ( .A1(n22263), .A2(n21971), .B1(n22262), .B2(n21970), .ZN(
        n21953) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n21967), .ZN(n21952) );
  OAI211_X1 U23521 ( .C1(n11106), .C2(n22268), .A(n21953), .B(n21952), .ZN(
        P1_U3090) );
  AOI22_X1 U23522 ( .A1(n22270), .A2(n21971), .B1(n21970), .B2(n22269), .ZN(
        n21955) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n22272), .B1(
        n22271), .B2(n21967), .ZN(n21954) );
  OAI211_X1 U23524 ( .C1(n11106), .C2(n22280), .A(n21955), .B(n21954), .ZN(
        P1_U3098) );
  AOI22_X1 U23525 ( .A1(n22276), .A2(n21971), .B1(n21970), .B2(n22275), .ZN(
        n21957) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22277), .B1(
        n22282), .B2(n21972), .ZN(n21956) );
  OAI211_X1 U23527 ( .C1(n21975), .C2(n22280), .A(n21957), .B(n21956), .ZN(
        P1_U3106) );
  AOI22_X1 U23528 ( .A1(n22282), .A2(n21967), .B1(n21970), .B2(n22281), .ZN(
        n21959) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n21972), .ZN(n21958) );
  OAI211_X1 U23530 ( .C1(n22286), .C2(n21964), .A(n21959), .B(n21958), .ZN(
        P1_U3114) );
  AOI22_X1 U23531 ( .A1(n22288), .A2(n21971), .B1(n21970), .B2(n22287), .ZN(
        n21961) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n21967), .ZN(n21960) );
  OAI211_X1 U23533 ( .C1(n11106), .C2(n22293), .A(n21961), .B(n21960), .ZN(
        P1_U3122) );
  AOI22_X1 U23534 ( .A1(n22148), .A2(n21972), .B1(n21970), .B2(n22147), .ZN(
        n21963) );
  AOI22_X1 U23535 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n22298), .B1(
        n22297), .B2(n21967), .ZN(n21962) );
  OAI211_X1 U23536 ( .C1(n22302), .C2(n21964), .A(n21963), .B(n21962), .ZN(
        P1_U3130) );
  AOI22_X1 U23537 ( .A1(n22304), .A2(n21971), .B1(n21970), .B2(n22303), .ZN(
        n21966) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22305), .B1(
        n22312), .B2(n21972), .ZN(n21965) );
  OAI211_X1 U23539 ( .C1(n21975), .C2(n22308), .A(n21966), .B(n21965), .ZN(
        P1_U3138) );
  AOI22_X1 U23540 ( .A1(n21970), .A2(n22310), .B1(n22309), .B2(n21971), .ZN(
        n21969) );
  AOI22_X1 U23541 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n21967), .ZN(n21968) );
  OAI211_X1 U23542 ( .C1(n11106), .C2(n22326), .A(n21969), .B(n21968), .ZN(
        P1_U3146) );
  AOI22_X1 U23543 ( .A1(n22320), .A2(n21971), .B1(n21970), .B2(n22317), .ZN(
        n21974) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n22323), .B1(
        n22322), .B2(n21972), .ZN(n21973) );
  OAI211_X1 U23545 ( .C1(n21975), .C2(n22326), .A(n21974), .B(n21973), .ZN(
        P1_U3154) );
  INV_X1 U23546 ( .A(n22017), .ZN(n22009) );
  OAI22_X2 U23547 ( .A1(n21978), .A2(n22219), .B1(n21977), .B2(n22217), .ZN(
        n22012) );
  NOR2_X2 U23548 ( .A1(n22215), .A2(n13844), .ZN(n22016) );
  AOI22_X1 U23549 ( .A1(n22322), .A2(n22012), .B1(n22016), .B2(n22216), .ZN(
        n21982) );
  OAI22_X1 U23550 ( .A1(n21980), .A2(n22217), .B1(n21979), .B2(n22219), .ZN(
        n22018) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22221), .B1(
        n22227), .B2(n22018), .ZN(n21981) );
  OAI211_X1 U23552 ( .C1(n22224), .C2(n22009), .A(n21982), .B(n21981), .ZN(
        P1_U3035) );
  INV_X1 U23553 ( .A(n22018), .ZN(n22015) );
  AOI22_X1 U23554 ( .A1(n22226), .A2(n22017), .B1(n22016), .B2(n22225), .ZN(
        n21984) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22228), .B1(
        n22227), .B2(n22012), .ZN(n21983) );
  OAI211_X1 U23556 ( .C1(n22015), .C2(n22231), .A(n21984), .B(n21983), .ZN(
        P1_U3043) );
  AOI22_X1 U23557 ( .A1(n22239), .A2(n22018), .B1(n22016), .B2(n22232), .ZN(
        n21986) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22234), .B1(
        n22233), .B2(n22012), .ZN(n21985) );
  OAI211_X1 U23559 ( .C1(n22237), .C2(n22009), .A(n21986), .B(n21985), .ZN(
        P1_U3051) );
  AOI22_X1 U23560 ( .A1(n22246), .A2(n22018), .B1(n22238), .B2(n22016), .ZN(
        n21988) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n22012), .ZN(n21987) );
  OAI211_X1 U23562 ( .C1(n22243), .C2(n22009), .A(n21988), .B(n21987), .ZN(
        P1_U3059) );
  AOI22_X1 U23563 ( .A1(n22016), .A2(n22245), .B1(n22244), .B2(n22017), .ZN(
        n21990) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n22247), .B1(
        n22246), .B2(n22012), .ZN(n21989) );
  OAI211_X1 U23565 ( .C1(n22015), .C2(n22255), .A(n21990), .B(n21989), .ZN(
        P1_U3067) );
  INV_X1 U23566 ( .A(n22012), .ZN(n22021) );
  AOI22_X1 U23567 ( .A1(n22251), .A2(n22017), .B1(n22016), .B2(n22250), .ZN(
        n21992) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n22252), .B1(
        n22257), .B2(n22018), .ZN(n21991) );
  OAI211_X1 U23569 ( .C1(n22021), .C2(n22255), .A(n21992), .B(n21991), .ZN(
        P1_U3075) );
  AOI22_X1 U23570 ( .A1(n22257), .A2(n22012), .B1(n22016), .B2(n22256), .ZN(
        n21994) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n22258), .B1(
        n22264), .B2(n22018), .ZN(n21993) );
  OAI211_X1 U23572 ( .C1(n22261), .C2(n22009), .A(n21994), .B(n21993), .ZN(
        P1_U3083) );
  AOI22_X1 U23573 ( .A1(n22263), .A2(n22017), .B1(n22262), .B2(n22016), .ZN(
        n21996) );
  AOI22_X1 U23574 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n22012), .ZN(n21995) );
  OAI211_X1 U23575 ( .C1(n22015), .C2(n22268), .A(n21996), .B(n21995), .ZN(
        P1_U3091) );
  AOI22_X1 U23576 ( .A1(n22270), .A2(n22017), .B1(n22016), .B2(n22269), .ZN(
        n21998) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n22272), .B1(
        n22271), .B2(n22012), .ZN(n21997) );
  OAI211_X1 U23578 ( .C1(n22015), .C2(n22280), .A(n21998), .B(n21997), .ZN(
        P1_U3099) );
  AOI22_X1 U23579 ( .A1(n22276), .A2(n22017), .B1(n22016), .B2(n22275), .ZN(
        n22000) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22277), .B1(
        n22282), .B2(n22018), .ZN(n21999) );
  OAI211_X1 U23581 ( .C1(n22021), .C2(n22280), .A(n22000), .B(n21999), .ZN(
        P1_U3107) );
  AOI22_X1 U23582 ( .A1(n22289), .A2(n22018), .B1(n22016), .B2(n22281), .ZN(
        n22002) );
  AOI22_X1 U23583 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22283), .B1(
        n22282), .B2(n22012), .ZN(n22001) );
  OAI211_X1 U23584 ( .C1(n22286), .C2(n22009), .A(n22002), .B(n22001), .ZN(
        P1_U3115) );
  AOI22_X1 U23585 ( .A1(n22288), .A2(n22017), .B1(n22016), .B2(n22287), .ZN(
        n22004) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n22012), .ZN(n22003) );
  OAI211_X1 U23587 ( .C1(n22015), .C2(n22293), .A(n22004), .B(n22003), .ZN(
        P1_U3123) );
  INV_X1 U23588 ( .A(n22016), .ZN(n22005) );
  INV_X1 U23589 ( .A(n22147), .ZN(n22294) );
  OAI22_X1 U23590 ( .A1(n22308), .A2(n22015), .B1(n22005), .B2(n22294), .ZN(
        n22006) );
  INV_X1 U23591 ( .A(n22006), .ZN(n22008) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n22298), .B1(
        n22297), .B2(n22012), .ZN(n22007) );
  OAI211_X1 U23593 ( .C1(n22302), .C2(n22009), .A(n22008), .B(n22007), .ZN(
        P1_U3131) );
  AOI22_X1 U23594 ( .A1(n22304), .A2(n22017), .B1(n22016), .B2(n22303), .ZN(
        n22011) );
  AOI22_X1 U23595 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22305), .B1(
        n22312), .B2(n22018), .ZN(n22010) );
  OAI211_X1 U23596 ( .C1(n22021), .C2(n22308), .A(n22011), .B(n22010), .ZN(
        P1_U3139) );
  AOI22_X1 U23597 ( .A1(n22016), .A2(n22310), .B1(n22309), .B2(n22017), .ZN(
        n22014) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22012), .ZN(n22013) );
  OAI211_X1 U23599 ( .C1(n22015), .C2(n22326), .A(n22014), .B(n22013), .ZN(
        P1_U3147) );
  AOI22_X1 U23600 ( .A1(n22320), .A2(n22017), .B1(n22016), .B2(n22317), .ZN(
        n22020) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n22323), .B1(
        n22322), .B2(n22018), .ZN(n22019) );
  OAI211_X1 U23602 ( .C1(n22021), .C2(n22326), .A(n22020), .B(n22019), .ZN(
        P1_U3155) );
  INV_X1 U23603 ( .A(n22063), .ZN(n22056) );
  OAI22_X2 U23604 ( .A1(n22024), .A2(n22219), .B1(n22023), .B2(n22217), .ZN(
        n22059) );
  NOR2_X2 U23605 ( .A1(n22215), .A2(n22025), .ZN(n22062) );
  AOI22_X1 U23606 ( .A1(n22322), .A2(n22059), .B1(n22062), .B2(n22216), .ZN(
        n22029) );
  OAI22_X1 U23607 ( .A1(n22027), .A2(n22219), .B1(n22026), .B2(n22217), .ZN(
        n22064) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22221), .B1(
        n22227), .B2(n11105), .ZN(n22028) );
  OAI211_X1 U23609 ( .C1(n22224), .C2(n22056), .A(n22029), .B(n22028), .ZN(
        P1_U3036) );
  AOI22_X1 U23610 ( .A1(n22226), .A2(n22063), .B1(n22062), .B2(n22225), .ZN(
        n22031) );
  AOI22_X1 U23611 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n22228), .B1(
        n22227), .B2(n22059), .ZN(n22030) );
  OAI211_X1 U23612 ( .C1(n11104), .C2(n22231), .A(n22031), .B(n22030), .ZN(
        P1_U3044) );
  INV_X1 U23613 ( .A(n22059), .ZN(n22067) );
  INV_X1 U23614 ( .A(n22062), .ZN(n22032) );
  OAI22_X1 U23615 ( .A1(n22231), .A2(n22067), .B1(n22032), .B2(n22125), .ZN(
        n22033) );
  INV_X1 U23616 ( .A(n22033), .ZN(n22035) );
  AOI22_X1 U23617 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22234), .B1(
        n22239), .B2(n11105), .ZN(n22034) );
  OAI211_X1 U23618 ( .C1(n22237), .C2(n22056), .A(n22035), .B(n22034), .ZN(
        P1_U3052) );
  AOI22_X1 U23619 ( .A1(n22246), .A2(n11105), .B1(n22238), .B2(n22062), .ZN(
        n22037) );
  AOI22_X1 U23620 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n22059), .ZN(n22036) );
  OAI211_X1 U23621 ( .C1(n22243), .C2(n22056), .A(n22037), .B(n22036), .ZN(
        P1_U3060) );
  AOI22_X1 U23622 ( .A1(n22062), .A2(n22245), .B1(n22244), .B2(n22063), .ZN(
        n22039) );
  AOI22_X1 U23623 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n22247), .B1(
        n22246), .B2(n22059), .ZN(n22038) );
  OAI211_X1 U23624 ( .C1(n11104), .C2(n22255), .A(n22039), .B(n22038), .ZN(
        P1_U3068) );
  AOI22_X1 U23625 ( .A1(n22251), .A2(n22063), .B1(n22062), .B2(n22250), .ZN(
        n22041) );
  AOI22_X1 U23626 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n22252), .B1(
        n22257), .B2(n11105), .ZN(n22040) );
  OAI211_X1 U23627 ( .C1(n22067), .C2(n22255), .A(n22041), .B(n22040), .ZN(
        P1_U3076) );
  AOI22_X1 U23628 ( .A1(n22257), .A2(n22059), .B1(n22062), .B2(n22256), .ZN(
        n22043) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n22258), .B1(
        n22264), .B2(n11105), .ZN(n22042) );
  OAI211_X1 U23630 ( .C1(n22261), .C2(n22056), .A(n22043), .B(n22042), .ZN(
        P1_U3084) );
  AOI22_X1 U23631 ( .A1(n22263), .A2(n22063), .B1(n22262), .B2(n22062), .ZN(
        n22045) );
  AOI22_X1 U23632 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n22059), .ZN(n22044) );
  OAI211_X1 U23633 ( .C1(n11104), .C2(n22268), .A(n22045), .B(n22044), .ZN(
        P1_U3092) );
  AOI22_X1 U23634 ( .A1(n22270), .A2(n22063), .B1(n22062), .B2(n22269), .ZN(
        n22047) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n22272), .B1(
        n22271), .B2(n22059), .ZN(n22046) );
  OAI211_X1 U23636 ( .C1(n11104), .C2(n22280), .A(n22047), .B(n22046), .ZN(
        P1_U3100) );
  AOI22_X1 U23637 ( .A1(n22276), .A2(n22063), .B1(n22062), .B2(n22275), .ZN(
        n22049) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n22277), .B1(
        n22282), .B2(n11105), .ZN(n22048) );
  OAI211_X1 U23639 ( .C1(n22067), .C2(n22280), .A(n22049), .B(n22048), .ZN(
        P1_U3108) );
  AOI22_X1 U23640 ( .A1(n22282), .A2(n22059), .B1(n22062), .B2(n22281), .ZN(
        n22051) );
  AOI22_X1 U23641 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n11105), .ZN(n22050) );
  OAI211_X1 U23642 ( .C1(n22286), .C2(n22056), .A(n22051), .B(n22050), .ZN(
        P1_U3116) );
  AOI22_X1 U23643 ( .A1(n22288), .A2(n22063), .B1(n22062), .B2(n22287), .ZN(
        n22053) );
  AOI22_X1 U23644 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n22059), .ZN(n22052) );
  OAI211_X1 U23645 ( .C1(n11104), .C2(n22293), .A(n22053), .B(n22052), .ZN(
        P1_U3124) );
  AOI22_X1 U23646 ( .A1(n22148), .A2(n11105), .B1(n22062), .B2(n22147), .ZN(
        n22055) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n22298), .B1(
        n22297), .B2(n22059), .ZN(n22054) );
  OAI211_X1 U23648 ( .C1(n22302), .C2(n22056), .A(n22055), .B(n22054), .ZN(
        P1_U3132) );
  AOI22_X1 U23649 ( .A1(n22304), .A2(n22063), .B1(n22062), .B2(n22303), .ZN(
        n22058) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n22305), .B1(
        n22312), .B2(n11105), .ZN(n22057) );
  OAI211_X1 U23651 ( .C1(n22067), .C2(n22308), .A(n22058), .B(n22057), .ZN(
        P1_U3140) );
  AOI22_X1 U23652 ( .A1(n22062), .A2(n22310), .B1(n22309), .B2(n22063), .ZN(
        n22061) );
  AOI22_X1 U23653 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22059), .ZN(n22060) );
  OAI211_X1 U23654 ( .C1(n11104), .C2(n22326), .A(n22061), .B(n22060), .ZN(
        P1_U3148) );
  AOI22_X1 U23655 ( .A1(n22320), .A2(n22063), .B1(n22062), .B2(n22317), .ZN(
        n22066) );
  AOI22_X1 U23656 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n22323), .B1(
        n22322), .B2(n11105), .ZN(n22065) );
  OAI211_X1 U23657 ( .C1(n22067), .C2(n22326), .A(n22066), .B(n22065), .ZN(
        P1_U3156) );
  INV_X1 U23658 ( .A(n22109), .ZN(n22101) );
  OAI22_X2 U23659 ( .A1(n22070), .A2(n22219), .B1(n22069), .B2(n22217), .ZN(
        n22104) );
  NOR2_X2 U23660 ( .A1(n22215), .A2(n13474), .ZN(n22108) );
  AOI22_X1 U23661 ( .A1(n22322), .A2(n22104), .B1(n22108), .B2(n22216), .ZN(
        n22074) );
  OAI22_X1 U23662 ( .A1(n22072), .A2(n22219), .B1(n22071), .B2(n22217), .ZN(
        n22110) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22221), .B1(
        n22227), .B2(n22110), .ZN(n22073) );
  OAI211_X1 U23664 ( .C1(n22224), .C2(n22101), .A(n22074), .B(n22073), .ZN(
        P1_U3037) );
  INV_X1 U23665 ( .A(n22110), .ZN(n22107) );
  AOI22_X1 U23666 ( .A1(n22226), .A2(n22109), .B1(n22108), .B2(n22225), .ZN(
        n22076) );
  AOI22_X1 U23667 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22228), .B1(
        n22227), .B2(n22104), .ZN(n22075) );
  OAI211_X1 U23668 ( .C1(n22107), .C2(n22231), .A(n22076), .B(n22075), .ZN(
        P1_U3045) );
  AOI22_X1 U23669 ( .A1(n22233), .A2(n22104), .B1(n22108), .B2(n22232), .ZN(
        n22078) );
  AOI22_X1 U23670 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22234), .B1(
        n22239), .B2(n22110), .ZN(n22077) );
  OAI211_X1 U23671 ( .C1(n22237), .C2(n22101), .A(n22078), .B(n22077), .ZN(
        P1_U3053) );
  AOI22_X1 U23672 ( .A1(n22246), .A2(n22110), .B1(n22238), .B2(n22108), .ZN(
        n22080) );
  AOI22_X1 U23673 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n22104), .ZN(n22079) );
  OAI211_X1 U23674 ( .C1(n22243), .C2(n22101), .A(n22080), .B(n22079), .ZN(
        P1_U3061) );
  AOI22_X1 U23675 ( .A1(n22108), .A2(n22245), .B1(n22244), .B2(n22109), .ZN(
        n22082) );
  AOI22_X1 U23676 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n22247), .B1(
        n22246), .B2(n22104), .ZN(n22081) );
  OAI211_X1 U23677 ( .C1(n22107), .C2(n22255), .A(n22082), .B(n22081), .ZN(
        P1_U3069) );
  INV_X1 U23678 ( .A(n22104), .ZN(n22113) );
  AOI22_X1 U23679 ( .A1(n22251), .A2(n22109), .B1(n22108), .B2(n22250), .ZN(
        n22084) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n22252), .B1(
        n22257), .B2(n22110), .ZN(n22083) );
  OAI211_X1 U23681 ( .C1(n22113), .C2(n22255), .A(n22084), .B(n22083), .ZN(
        P1_U3077) );
  AOI22_X1 U23682 ( .A1(n22264), .A2(n22110), .B1(n22108), .B2(n22256), .ZN(
        n22086) );
  AOI22_X1 U23683 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n22258), .B1(
        n22257), .B2(n22104), .ZN(n22085) );
  OAI211_X1 U23684 ( .C1(n22261), .C2(n22101), .A(n22086), .B(n22085), .ZN(
        P1_U3085) );
  AOI22_X1 U23685 ( .A1(n22263), .A2(n22109), .B1(n22262), .B2(n22108), .ZN(
        n22088) );
  AOI22_X1 U23686 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n22104), .ZN(n22087) );
  OAI211_X1 U23687 ( .C1(n22107), .C2(n22268), .A(n22088), .B(n22087), .ZN(
        P1_U3093) );
  AOI22_X1 U23688 ( .A1(n22270), .A2(n22109), .B1(n22108), .B2(n22269), .ZN(
        n22090) );
  AOI22_X1 U23689 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n22272), .B1(
        n22271), .B2(n22104), .ZN(n22089) );
  OAI211_X1 U23690 ( .C1(n22107), .C2(n22280), .A(n22090), .B(n22089), .ZN(
        P1_U3101) );
  AOI22_X1 U23691 ( .A1(n22276), .A2(n22109), .B1(n22108), .B2(n22275), .ZN(
        n22092) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22277), .B1(
        n22282), .B2(n22110), .ZN(n22091) );
  OAI211_X1 U23693 ( .C1(n22113), .C2(n22280), .A(n22092), .B(n22091), .ZN(
        P1_U3109) );
  AOI22_X1 U23694 ( .A1(n22289), .A2(n22110), .B1(n22108), .B2(n22281), .ZN(
        n22094) );
  AOI22_X1 U23695 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22283), .B1(
        n22282), .B2(n22104), .ZN(n22093) );
  OAI211_X1 U23696 ( .C1(n22286), .C2(n22101), .A(n22094), .B(n22093), .ZN(
        P1_U3117) );
  AOI22_X1 U23697 ( .A1(n22288), .A2(n22109), .B1(n22108), .B2(n22287), .ZN(
        n22096) );
  AOI22_X1 U23698 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n22104), .ZN(n22095) );
  OAI211_X1 U23699 ( .C1(n22107), .C2(n22293), .A(n22096), .B(n22095), .ZN(
        P1_U3125) );
  INV_X1 U23700 ( .A(n22108), .ZN(n22097) );
  OAI22_X1 U23701 ( .A1(n22308), .A2(n22107), .B1(n22097), .B2(n22294), .ZN(
        n22098) );
  INV_X1 U23702 ( .A(n22098), .ZN(n22100) );
  AOI22_X1 U23703 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n22298), .B1(
        n22297), .B2(n22104), .ZN(n22099) );
  OAI211_X1 U23704 ( .C1(n22302), .C2(n22101), .A(n22100), .B(n22099), .ZN(
        P1_U3133) );
  AOI22_X1 U23705 ( .A1(n22304), .A2(n22109), .B1(n22108), .B2(n22303), .ZN(
        n22103) );
  AOI22_X1 U23706 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22305), .B1(
        n22312), .B2(n22110), .ZN(n22102) );
  OAI211_X1 U23707 ( .C1(n22113), .C2(n22308), .A(n22103), .B(n22102), .ZN(
        P1_U3141) );
  AOI22_X1 U23708 ( .A1(n22108), .A2(n22310), .B1(n22309), .B2(n22109), .ZN(
        n22106) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22104), .ZN(n22105) );
  OAI211_X1 U23710 ( .C1(n22107), .C2(n22326), .A(n22106), .B(n22105), .ZN(
        P1_U3149) );
  AOI22_X1 U23711 ( .A1(n22320), .A2(n22109), .B1(n22108), .B2(n22317), .ZN(
        n22112) );
  AOI22_X1 U23712 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n22323), .B1(
        n22322), .B2(n22110), .ZN(n22111) );
  OAI211_X1 U23713 ( .C1(n22113), .C2(n22326), .A(n22112), .B(n22111), .ZN(
        P1_U3157) );
  INV_X1 U23714 ( .A(n22159), .ZN(n22151) );
  OAI22_X2 U23715 ( .A1(n22116), .A2(n22219), .B1(n22115), .B2(n22217), .ZN(
        n22154) );
  NOR2_X2 U23716 ( .A1(n22215), .A2(n22117), .ZN(n22158) );
  AOI22_X1 U23717 ( .A1(n22322), .A2(n22154), .B1(n22158), .B2(n22216), .ZN(
        n22121) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22221), .B1(
        n22227), .B2(n22160), .ZN(n22120) );
  OAI211_X1 U23719 ( .C1(n22224), .C2(n22151), .A(n22121), .B(n22120), .ZN(
        P1_U3038) );
  INV_X1 U23720 ( .A(n22160), .ZN(n22157) );
  AOI22_X1 U23721 ( .A1(n22226), .A2(n22159), .B1(n22158), .B2(n22225), .ZN(
        n22123) );
  AOI22_X1 U23722 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22228), .B1(
        n22227), .B2(n22154), .ZN(n22122) );
  OAI211_X1 U23723 ( .C1(n22157), .C2(n22231), .A(n22123), .B(n22122), .ZN(
        P1_U3046) );
  INV_X1 U23724 ( .A(n22154), .ZN(n22163) );
  INV_X1 U23725 ( .A(n22158), .ZN(n22124) );
  OAI22_X1 U23726 ( .A1(n22231), .A2(n22163), .B1(n22125), .B2(n22124), .ZN(
        n22126) );
  INV_X1 U23727 ( .A(n22126), .ZN(n22128) );
  AOI22_X1 U23728 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22234), .B1(
        n22239), .B2(n22160), .ZN(n22127) );
  OAI211_X1 U23729 ( .C1(n22237), .C2(n22151), .A(n22128), .B(n22127), .ZN(
        P1_U3054) );
  AOI22_X1 U23730 ( .A1(n22239), .A2(n22154), .B1(n22238), .B2(n22158), .ZN(
        n22130) );
  AOI22_X1 U23731 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n22240), .B1(
        n22246), .B2(n22160), .ZN(n22129) );
  OAI211_X1 U23732 ( .C1(n22243), .C2(n22151), .A(n22130), .B(n22129), .ZN(
        P1_U3062) );
  AOI22_X1 U23733 ( .A1(n22158), .A2(n22245), .B1(n22244), .B2(n22159), .ZN(
        n22132) );
  AOI22_X1 U23734 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n22247), .B1(
        n22246), .B2(n22154), .ZN(n22131) );
  OAI211_X1 U23735 ( .C1(n22157), .C2(n22255), .A(n22132), .B(n22131), .ZN(
        P1_U3070) );
  AOI22_X1 U23736 ( .A1(n22251), .A2(n22159), .B1(n22158), .B2(n22250), .ZN(
        n22134) );
  AOI22_X1 U23737 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n22252), .B1(
        n22257), .B2(n22160), .ZN(n22133) );
  OAI211_X1 U23738 ( .C1(n22163), .C2(n22255), .A(n22134), .B(n22133), .ZN(
        P1_U3078) );
  AOI22_X1 U23739 ( .A1(n22264), .A2(n22160), .B1(n22158), .B2(n22256), .ZN(
        n22136) );
  AOI22_X1 U23740 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n22258), .B1(
        n22257), .B2(n22154), .ZN(n22135) );
  OAI211_X1 U23741 ( .C1(n22261), .C2(n22151), .A(n22136), .B(n22135), .ZN(
        P1_U3086) );
  AOI22_X1 U23742 ( .A1(n22263), .A2(n22159), .B1(n22262), .B2(n22158), .ZN(
        n22138) );
  AOI22_X1 U23743 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n22154), .ZN(n22137) );
  OAI211_X1 U23744 ( .C1(n22157), .C2(n22268), .A(n22138), .B(n22137), .ZN(
        P1_U3094) );
  AOI22_X1 U23745 ( .A1(n22270), .A2(n22159), .B1(n22158), .B2(n22269), .ZN(
        n22140) );
  AOI22_X1 U23746 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n22272), .B1(
        n22271), .B2(n22154), .ZN(n22139) );
  OAI211_X1 U23747 ( .C1(n22157), .C2(n22280), .A(n22140), .B(n22139), .ZN(
        P1_U3102) );
  AOI22_X1 U23748 ( .A1(n22276), .A2(n22159), .B1(n22158), .B2(n22275), .ZN(
        n22142) );
  AOI22_X1 U23749 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22277), .B1(
        n22282), .B2(n22160), .ZN(n22141) );
  OAI211_X1 U23750 ( .C1(n22163), .C2(n22280), .A(n22142), .B(n22141), .ZN(
        P1_U3110) );
  AOI22_X1 U23751 ( .A1(n22282), .A2(n22154), .B1(n22158), .B2(n22281), .ZN(
        n22144) );
  AOI22_X1 U23752 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n22160), .ZN(n22143) );
  OAI211_X1 U23753 ( .C1(n22286), .C2(n22151), .A(n22144), .B(n22143), .ZN(
        P1_U3118) );
  AOI22_X1 U23754 ( .A1(n22288), .A2(n22159), .B1(n22158), .B2(n22287), .ZN(
        n22146) );
  AOI22_X1 U23755 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n22154), .ZN(n22145) );
  OAI211_X1 U23756 ( .C1(n22157), .C2(n22293), .A(n22146), .B(n22145), .ZN(
        P1_U3126) );
  AOI22_X1 U23757 ( .A1(n22148), .A2(n22160), .B1(n22158), .B2(n22147), .ZN(
        n22150) );
  AOI22_X1 U23758 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n22298), .B1(
        n22297), .B2(n22154), .ZN(n22149) );
  OAI211_X1 U23759 ( .C1(n22302), .C2(n22151), .A(n22150), .B(n22149), .ZN(
        P1_U3134) );
  AOI22_X1 U23760 ( .A1(n22304), .A2(n22159), .B1(n22158), .B2(n22303), .ZN(
        n22153) );
  AOI22_X1 U23761 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22305), .B1(
        n22312), .B2(n22160), .ZN(n22152) );
  OAI211_X1 U23762 ( .C1(n22163), .C2(n22308), .A(n22153), .B(n22152), .ZN(
        P1_U3142) );
  AOI22_X1 U23763 ( .A1(n22158), .A2(n22310), .B1(n22309), .B2(n22159), .ZN(
        n22156) );
  AOI22_X1 U23764 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22154), .ZN(n22155) );
  OAI211_X1 U23765 ( .C1(n22157), .C2(n22326), .A(n22156), .B(n22155), .ZN(
        P1_U3150) );
  AOI22_X1 U23766 ( .A1(n22320), .A2(n22159), .B1(n22158), .B2(n22317), .ZN(
        n22162) );
  AOI22_X1 U23767 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n22323), .B1(
        n22322), .B2(n22160), .ZN(n22161) );
  OAI211_X1 U23768 ( .C1(n22163), .C2(n22326), .A(n22162), .B(n22161), .ZN(
        P1_U3158) );
  OAI22_X2 U23769 ( .A1(n22166), .A2(n22219), .B1(n22165), .B2(n22217), .ZN(
        n22201) );
  NOR2_X2 U23770 ( .A1(n22215), .A2(n22167), .ZN(n22205) );
  AOI22_X1 U23771 ( .A1(n22322), .A2(n22201), .B1(n22205), .B2(n22216), .ZN(
        n22171) );
  OAI22_X1 U23772 ( .A1(n22169), .A2(n22219), .B1(n22168), .B2(n22217), .ZN(
        n22207) );
  AOI22_X1 U23773 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22221), .B1(
        n22227), .B2(n22207), .ZN(n22170) );
  OAI211_X1 U23774 ( .C1(n22224), .C2(n22198), .A(n22171), .B(n22170), .ZN(
        P1_U3039) );
  INV_X1 U23775 ( .A(n22207), .ZN(n22204) );
  AOI22_X1 U23776 ( .A1(n22226), .A2(n22206), .B1(n22205), .B2(n22225), .ZN(
        n22173) );
  AOI22_X1 U23777 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n22228), .B1(
        n22227), .B2(n22201), .ZN(n22172) );
  OAI211_X1 U23778 ( .C1(n22204), .C2(n22231), .A(n22173), .B(n22172), .ZN(
        P1_U3047) );
  AOI22_X1 U23779 ( .A1(n22239), .A2(n22207), .B1(n22205), .B2(n22232), .ZN(
        n22175) );
  AOI22_X1 U23780 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22234), .B1(
        n22233), .B2(n22201), .ZN(n22174) );
  OAI211_X1 U23781 ( .C1(n22237), .C2(n22198), .A(n22175), .B(n22174), .ZN(
        P1_U3055) );
  AOI22_X1 U23782 ( .A1(n22246), .A2(n22207), .B1(n22238), .B2(n22205), .ZN(
        n22177) );
  AOI22_X1 U23783 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n22201), .ZN(n22176) );
  OAI211_X1 U23784 ( .C1(n22243), .C2(n22198), .A(n22177), .B(n22176), .ZN(
        P1_U3063) );
  AOI22_X1 U23785 ( .A1(n22205), .A2(n22245), .B1(n22244), .B2(n22206), .ZN(
        n22179) );
  AOI22_X1 U23786 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n22247), .B1(
        n22246), .B2(n22201), .ZN(n22178) );
  OAI211_X1 U23787 ( .C1(n22204), .C2(n22255), .A(n22179), .B(n22178), .ZN(
        P1_U3071) );
  INV_X1 U23788 ( .A(n22201), .ZN(n22210) );
  AOI22_X1 U23789 ( .A1(n22251), .A2(n22206), .B1(n22205), .B2(n22250), .ZN(
        n22181) );
  AOI22_X1 U23790 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n22252), .B1(
        n22257), .B2(n22207), .ZN(n22180) );
  OAI211_X1 U23791 ( .C1(n22210), .C2(n22255), .A(n22181), .B(n22180), .ZN(
        P1_U3079) );
  AOI22_X1 U23792 ( .A1(n22264), .A2(n22207), .B1(n22205), .B2(n22256), .ZN(
        n22183) );
  AOI22_X1 U23793 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n22258), .B1(
        n22257), .B2(n22201), .ZN(n22182) );
  OAI211_X1 U23794 ( .C1(n22261), .C2(n22198), .A(n22183), .B(n22182), .ZN(
        P1_U3087) );
  AOI22_X1 U23795 ( .A1(n22263), .A2(n22206), .B1(n22262), .B2(n22205), .ZN(
        n22185) );
  AOI22_X1 U23796 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n22201), .ZN(n22184) );
  OAI211_X1 U23797 ( .C1(n22204), .C2(n22268), .A(n22185), .B(n22184), .ZN(
        P1_U3095) );
  AOI22_X1 U23798 ( .A1(n22270), .A2(n22206), .B1(n22205), .B2(n22269), .ZN(
        n22187) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n22272), .B1(
        n22271), .B2(n22201), .ZN(n22186) );
  OAI211_X1 U23800 ( .C1(n22204), .C2(n22280), .A(n22187), .B(n22186), .ZN(
        P1_U3103) );
  AOI22_X1 U23801 ( .A1(n22276), .A2(n22206), .B1(n22205), .B2(n22275), .ZN(
        n22189) );
  AOI22_X1 U23802 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n22277), .B1(
        n22282), .B2(n22207), .ZN(n22188) );
  OAI211_X1 U23803 ( .C1(n22210), .C2(n22280), .A(n22189), .B(n22188), .ZN(
        P1_U3111) );
  AOI22_X1 U23804 ( .A1(n22282), .A2(n22201), .B1(n22205), .B2(n22281), .ZN(
        n22191) );
  AOI22_X1 U23805 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22283), .B1(
        n22289), .B2(n22207), .ZN(n22190) );
  OAI211_X1 U23806 ( .C1(n22286), .C2(n22198), .A(n22191), .B(n22190), .ZN(
        P1_U3119) );
  AOI22_X1 U23807 ( .A1(n22288), .A2(n22206), .B1(n22205), .B2(n22287), .ZN(
        n22193) );
  AOI22_X1 U23808 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n22201), .ZN(n22192) );
  OAI211_X1 U23809 ( .C1(n22204), .C2(n22293), .A(n22193), .B(n22192), .ZN(
        P1_U3127) );
  INV_X1 U23810 ( .A(n22205), .ZN(n22194) );
  OAI22_X1 U23811 ( .A1(n22308), .A2(n22204), .B1(n22194), .B2(n22294), .ZN(
        n22195) );
  INV_X1 U23812 ( .A(n22195), .ZN(n22197) );
  AOI22_X1 U23813 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n22298), .B1(
        n22297), .B2(n22201), .ZN(n22196) );
  OAI211_X1 U23814 ( .C1(n22302), .C2(n22198), .A(n22197), .B(n22196), .ZN(
        P1_U3135) );
  AOI22_X1 U23815 ( .A1(n22304), .A2(n22206), .B1(n22205), .B2(n22303), .ZN(
        n22200) );
  AOI22_X1 U23816 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n22305), .B1(
        n22312), .B2(n22207), .ZN(n22199) );
  OAI211_X1 U23817 ( .C1(n22210), .C2(n22308), .A(n22200), .B(n22199), .ZN(
        P1_U3143) );
  AOI22_X1 U23818 ( .A1(n22205), .A2(n22310), .B1(n22309), .B2(n22206), .ZN(
        n22203) );
  AOI22_X1 U23819 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22201), .ZN(n22202) );
  OAI211_X1 U23820 ( .C1(n22204), .C2(n22326), .A(n22203), .B(n22202), .ZN(
        P1_U3151) );
  AOI22_X1 U23821 ( .A1(n22320), .A2(n22206), .B1(n22205), .B2(n22317), .ZN(
        n22209) );
  AOI22_X1 U23822 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n22323), .B1(
        n22322), .B2(n22207), .ZN(n22208) );
  OAI211_X1 U23823 ( .C1(n22210), .C2(n22326), .A(n22209), .B(n22208), .ZN(
        P1_U3159) );
  INV_X1 U23824 ( .A(n22319), .ZN(n22301) );
  OAI22_X2 U23825 ( .A1(n22214), .A2(n22219), .B1(n22213), .B2(n22217), .ZN(
        n22311) );
  NOR2_X2 U23826 ( .A1(n22215), .A2(n13429), .ZN(n22318) );
  AOI22_X1 U23827 ( .A1(n22322), .A2(n22311), .B1(n22318), .B2(n22216), .ZN(
        n22223) );
  OAI22_X1 U23828 ( .A1(n22220), .A2(n22219), .B1(n22218), .B2(n22217), .ZN(
        n22321) );
  AOI22_X1 U23829 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22221), .B1(
        n22227), .B2(n22321), .ZN(n22222) );
  OAI211_X1 U23830 ( .C1(n22224), .C2(n22301), .A(n22223), .B(n22222), .ZN(
        P1_U3040) );
  INV_X1 U23831 ( .A(n22321), .ZN(n22316) );
  AOI22_X1 U23832 ( .A1(n22226), .A2(n22319), .B1(n22318), .B2(n22225), .ZN(
        n22230) );
  AOI22_X1 U23833 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22228), .B1(
        n22227), .B2(n22311), .ZN(n22229) );
  OAI211_X1 U23834 ( .C1(n22316), .C2(n22231), .A(n22230), .B(n22229), .ZN(
        P1_U3048) );
  AOI22_X1 U23835 ( .A1(n22239), .A2(n22321), .B1(n22232), .B2(n22318), .ZN(
        n22236) );
  AOI22_X1 U23836 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22234), .B1(
        n22233), .B2(n22311), .ZN(n22235) );
  OAI211_X1 U23837 ( .C1(n22237), .C2(n22301), .A(n22236), .B(n22235), .ZN(
        P1_U3056) );
  AOI22_X1 U23838 ( .A1(n22239), .A2(n22311), .B1(n22238), .B2(n22318), .ZN(
        n22242) );
  AOI22_X1 U23839 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22240), .B1(
        n22246), .B2(n22321), .ZN(n22241) );
  OAI211_X1 U23840 ( .C1(n22243), .C2(n22301), .A(n22242), .B(n22241), .ZN(
        P1_U3064) );
  AOI22_X1 U23841 ( .A1(n22318), .A2(n22245), .B1(n22244), .B2(n22319), .ZN(
        n22249) );
  AOI22_X1 U23842 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n22247), .B1(
        n22246), .B2(n22311), .ZN(n22248) );
  OAI211_X1 U23843 ( .C1(n22316), .C2(n22255), .A(n22249), .B(n22248), .ZN(
        P1_U3072) );
  INV_X1 U23844 ( .A(n22311), .ZN(n22327) );
  AOI22_X1 U23845 ( .A1(n22251), .A2(n22319), .B1(n22318), .B2(n22250), .ZN(
        n22254) );
  AOI22_X1 U23846 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n22252), .B1(
        n22257), .B2(n22321), .ZN(n22253) );
  OAI211_X1 U23847 ( .C1(n22327), .C2(n22255), .A(n22254), .B(n22253), .ZN(
        P1_U3080) );
  AOI22_X1 U23848 ( .A1(n22257), .A2(n22311), .B1(n22318), .B2(n22256), .ZN(
        n22260) );
  AOI22_X1 U23849 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n22258), .B1(
        n22264), .B2(n22321), .ZN(n22259) );
  OAI211_X1 U23850 ( .C1(n22261), .C2(n22301), .A(n22260), .B(n22259), .ZN(
        P1_U3088) );
  AOI22_X1 U23851 ( .A1(n22263), .A2(n22319), .B1(n22262), .B2(n22318), .ZN(
        n22267) );
  AOI22_X1 U23852 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n22265), .B1(
        n22264), .B2(n22311), .ZN(n22266) );
  OAI211_X1 U23853 ( .C1(n22316), .C2(n22268), .A(n22267), .B(n22266), .ZN(
        P1_U3096) );
  AOI22_X1 U23854 ( .A1(n22270), .A2(n22319), .B1(n22318), .B2(n22269), .ZN(
        n22274) );
  AOI22_X1 U23855 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n22272), .B1(
        n22271), .B2(n22311), .ZN(n22273) );
  OAI211_X1 U23856 ( .C1(n22316), .C2(n22280), .A(n22274), .B(n22273), .ZN(
        P1_U3104) );
  AOI22_X1 U23857 ( .A1(n22276), .A2(n22319), .B1(n22318), .B2(n22275), .ZN(
        n22279) );
  AOI22_X1 U23858 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22277), .B1(
        n22282), .B2(n22321), .ZN(n22278) );
  OAI211_X1 U23859 ( .C1(n22327), .C2(n22280), .A(n22279), .B(n22278), .ZN(
        P1_U3112) );
  AOI22_X1 U23860 ( .A1(n22289), .A2(n22321), .B1(n22318), .B2(n22281), .ZN(
        n22285) );
  AOI22_X1 U23861 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22283), .B1(
        n22282), .B2(n22311), .ZN(n22284) );
  OAI211_X1 U23862 ( .C1(n22286), .C2(n22301), .A(n22285), .B(n22284), .ZN(
        P1_U3120) );
  AOI22_X1 U23863 ( .A1(n22288), .A2(n22319), .B1(n22318), .B2(n22287), .ZN(
        n22292) );
  AOI22_X1 U23864 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n22290), .B1(
        n22289), .B2(n22311), .ZN(n22291) );
  OAI211_X1 U23865 ( .C1(n22316), .C2(n22293), .A(n22292), .B(n22291), .ZN(
        P1_U3128) );
  INV_X1 U23866 ( .A(n22318), .ZN(n22295) );
  OAI22_X1 U23867 ( .A1(n22308), .A2(n22316), .B1(n22295), .B2(n22294), .ZN(
        n22296) );
  INV_X1 U23868 ( .A(n22296), .ZN(n22300) );
  AOI22_X1 U23869 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22298), .B1(
        n22297), .B2(n22311), .ZN(n22299) );
  OAI211_X1 U23870 ( .C1(n22302), .C2(n22301), .A(n22300), .B(n22299), .ZN(
        P1_U3136) );
  AOI22_X1 U23871 ( .A1(n22304), .A2(n22319), .B1(n22318), .B2(n22303), .ZN(
        n22307) );
  AOI22_X1 U23872 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22305), .B1(
        n22312), .B2(n22321), .ZN(n22306) );
  OAI211_X1 U23873 ( .C1(n22327), .C2(n22308), .A(n22307), .B(n22306), .ZN(
        P1_U3144) );
  AOI22_X1 U23874 ( .A1(n22318), .A2(n22310), .B1(n22309), .B2(n22319), .ZN(
        n22315) );
  AOI22_X1 U23875 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22313), .B1(
        n22312), .B2(n22311), .ZN(n22314) );
  OAI211_X1 U23876 ( .C1(n22316), .C2(n22326), .A(n22315), .B(n22314), .ZN(
        P1_U3152) );
  AOI22_X1 U23877 ( .A1(n22320), .A2(n22319), .B1(n22318), .B2(n22317), .ZN(
        n22325) );
  AOI22_X1 U23878 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n22323), .B1(
        n22322), .B2(n22321), .ZN(n22324) );
  OAI211_X1 U23879 ( .C1(n22327), .C2(n22326), .A(n22325), .B(n22324), .ZN(
        P1_U3160) );
  OAI22_X1 U23880 ( .A1(n22329), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n22328), .ZN(n22330) );
  INV_X1 U23881 ( .A(n22330), .ZN(P1_U3486) );
  AND2_X2 U15237 ( .A1(n14764), .A2(n14915), .ZN(n13445) );
  INV_X2 U11097 ( .A(n11093), .ZN(n17823) );
  CLKBUF_X3 U13143 ( .A(n11508), .Z(n17848) );
  BUF_X2 U11372 ( .A(n11469), .Z(n17852) );
  BUF_X2 U11134 ( .A(n11437), .Z(n17833) );
  CLKBUF_X2 U11118 ( .A(n13476), .Z(n13831) );
  CLKBUF_X2 U11136 ( .A(n11560), .Z(n17725) );
  INV_X2 U11197 ( .A(n17747), .ZN(n17861) );
  CLKBUF_X1 U11365 ( .A(n15508), .Z(n10984) );
  CLKBUF_X1 U11391 ( .A(n13489), .Z(n13490) );
  CLKBUF_X1 U11392 ( .A(n13470), .Z(n22167) );
  CLKBUF_X1 U11414 ( .A(n15933), .Z(n15934) );
  CLKBUF_X1 U11436 ( .A(n15844), .Z(n15845) );
  CLKBUF_X1 U11457 ( .A(n12944), .Z(n15331) );
  CLKBUF_X1 U12052 ( .A(n17465), .Z(n17473) );
  CLKBUF_X1 U12228 ( .A(n12633), .Z(n19642) );
  CLKBUF_X1 U12248 ( .A(n15564), .Z(n11002) );
  CLKBUF_X1 U12343 ( .A(n16705), .Z(n16727) );
  CLKBUF_X1 U12384 ( .A(n20149), .Z(n20164) );
  INV_X2 U12487 ( .A(n18195), .ZN(n18141) );
  INV_X1 U13040 ( .A(n19882), .ZN(n19907) );
  AOI211_X1 U13145 ( .C1(n20033), .C2(n16069), .A(n16068), .B(n16067), .ZN(
        n16070) );
  CLKBUF_X1 U15325 ( .A(n18745), .Z(n19080) );
endmodule

