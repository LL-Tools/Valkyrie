

module b20_C_AntiSAT_k_256_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, ADD_1068_U4, ADD_1068_U55, 
        ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, 
        ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, 
        ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, 
        ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, 
        P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, 
        P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, 
        P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, 
        P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, 
        P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, 
        P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, 
        P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, 
        P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, 
        P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, 
        P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, 
        P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, 
        P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502;

  NAND2_X1 U5001 ( .A1(n8441), .A2(n6617), .ZN(n8440) );
  INV_X1 U5002 ( .A(n6279), .ZN(n8048) );
  CLKBUF_X1 U5003 ( .A(n6297), .Z(n6451) );
  CLKBUF_X3 U5004 ( .A(n6120), .Z(n7352) );
  NAND2_X1 U5005 ( .A1(n8648), .A2(n7865), .ZN(n6120) );
  XNOR2_X1 U5007 ( .A(n5135), .B(n5144), .ZN(n5664) );
  AND2_X1 U5009 ( .A1(n6629), .A2(n6628), .ZN(n4496) );
  OAI21_X1 U5010 ( .B1(n6626), .B2(n5023), .A(n5019), .ZN(n4497) );
  XNOR2_X2 U5011 ( .A(n6082), .B(n6081), .ZN(n4498) );
  OAI21_X1 U5012 ( .B1(n6626), .B2(n5023), .A(n5019), .ZN(n8294) );
  XNOR2_X1 U5013 ( .A(n6082), .B(n6081), .ZN(n6084) );
  NAND2_X1 U5014 ( .A1(n8067), .A2(n8063), .ZN(n7186) );
  AND2_X1 U5015 ( .A1(n4910), .A2(n4909), .ZN(n5003) );
  INV_X2 U5016 ( .A(n5967), .ZN(n5991) );
  NAND3_X1 U5017 ( .A1(n4752), .A2(n4750), .A3(n4753), .ZN(n6074) );
  CLKBUF_X2 U5018 ( .A(n6157), .Z(n6410) );
  OR2_X1 U5019 ( .A1(n7603), .A2(n7602), .ZN(n4926) );
  OR2_X1 U5020 ( .A1(n6441), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6456) );
  INV_X1 U5021 ( .A(n8070), .ZN(n9990) );
  INV_X1 U5022 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8644) );
  INV_X1 U5023 ( .A(n8890), .ZN(n5485) );
  INV_X1 U5024 ( .A(n9171), .ZN(n9349) );
  INV_X1 U5025 ( .A(n6680), .ZN(n7856) );
  NAND4_X1 U5027 ( .A1(n5245), .A2(n5244), .A3(n5243), .A4(n5242), .ZN(n9050)
         );
  NAND2_X2 U5028 ( .A1(n6568), .A2(n6567), .ZN(n8494) );
  OAI21_X2 U5029 ( .B1(n10058), .B2(n8496), .A(n7744), .ZN(n6568) );
  XNOR2_X2 U5030 ( .A(n7875), .B(n7874), .ZN(n7882) );
  NOR2_X1 U5031 ( .A1(n6074), .A2(n6680), .ZN(n4499) );
  NOR2_X1 U5032 ( .A1(n6074), .A2(n6680), .ZN(n6297) );
  NAND2_X4 U5033 ( .A1(n6110), .A2(n4914), .ZN(n6846) );
  NAND2_X4 U5034 ( .A1(n5757), .A2(n6007), .ZN(n5988) );
  NAND2_X2 U5035 ( .A1(n5756), .A2(n9032), .ZN(n5757) );
  XNOR2_X2 U5036 ( .A(n6078), .B(P2_IR_REG_29__SCAN_IN), .ZN(n6083) );
  NAND2_X2 U5037 ( .A1(n8643), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6082) );
  OAI22_X2 U5038 ( .A1(n7590), .A2(n6565), .B1(n7682), .B2(n10045), .ZN(n7680)
         );
  OAI22_X2 U5039 ( .A1(n7547), .A2(n8036), .B1(n8226), .B2(n7552), .ZN(n7590)
         );
  INV_X4 U5040 ( .A(n6726), .ZN(n5665) );
  AOI21_X2 U5041 ( .B1(n9661), .B2(n5678), .A(n5677), .ZN(n6980) );
  OAI21_X2 U5042 ( .B1(n6883), .B2(n5240), .A(n8903), .ZN(n9661) );
  INV_X2 U5043 ( .A(n5003), .ZN(n5100) );
  NAND2_X2 U5044 ( .A1(n5664), .A2(n5669), .ZN(n6707) );
  XNOR2_X2 U5045 ( .A(n5272), .B(n5249), .ZN(n7072) );
  NAND2_X1 U5046 ( .A1(n5318), .A2(n5317), .ZN(n9751) );
  NAND2_X1 U5047 ( .A1(n9986), .A2(n9990), .ZN(n9985) );
  AND3_X1 U5048 ( .A1(n5238), .A2(n5237), .A3(n5236), .ZN(n9691) );
  BUF_X2 U5049 ( .A(n5792), .Z(n5948) );
  CLKBUF_X2 U5050 ( .A(n6147), .Z(n6344) );
  NAND4_X2 U5051 ( .A1(n5202), .A2(n5201), .A3(n5203), .A4(n5200), .ZN(n6884)
         );
  CLKBUF_X2 U5052 ( .A(n5241), .Z(n5647) );
  CLKBUF_X1 U5053 ( .A(n5664), .Z(n4502) );
  OR2_X1 U5054 ( .A1(n6065), .A2(n4872), .ZN(n4752) );
  AND2_X1 U5055 ( .A1(n4987), .A2(n4674), .ZN(n4673) );
  OAI21_X1 U5056 ( .B1(n8336), .B2(n10000), .A(n8335), .ZN(n8570) );
  AND2_X1 U5057 ( .A1(n8314), .A2(n8313), .ZN(n8316) );
  NAND2_X1 U5058 ( .A1(n4898), .A2(n4901), .ZN(n8345) );
  NAND2_X1 U5059 ( .A1(n8206), .A2(n8193), .ZN(n8185) );
  NAND2_X1 U5060 ( .A1(n5706), .A2(n9148), .ZN(n8900) );
  NAND2_X1 U5061 ( .A1(n9174), .A2(n9183), .ZN(n8974) );
  NAND2_X1 U5062 ( .A1(n8425), .A2(n8151), .ZN(n8412) );
  NAND2_X1 U5063 ( .A1(n6453), .A2(n6452), .ZN(n8511) );
  XNOR2_X1 U5064 ( .A(n5615), .B(n5614), .ZN(n7787) );
  NAND2_X1 U5065 ( .A1(n5582), .A2(n5581), .ZN(n9370) );
  NAND2_X1 U5066 ( .A1(n8436), .A2(n8435), .ZN(n8434) );
  NAND2_X1 U5067 ( .A1(n5568), .A2(n5567), .ZN(n9375) );
  NAND2_X1 U5068 ( .A1(n5552), .A2(n5551), .ZN(n9384) );
  NAND2_X1 U5069 ( .A1(n6385), .A2(n6384), .ZN(n8594) );
  NAND2_X1 U5070 ( .A1(n5534), .A2(n5533), .ZN(n9248) );
  OR2_X1 U5071 ( .A1(n5850), .A2(n5849), .ZN(n5035) );
  NAND2_X1 U5072 ( .A1(n5850), .A2(n5849), .ZN(n7698) );
  NAND2_X1 U5073 ( .A1(n6375), .A2(n6374), .ZN(n8600) );
  NAND2_X1 U5074 ( .A1(n5562), .A2(n5561), .ZN(n5575) );
  NAND2_X1 U5075 ( .A1(n6355), .A2(n6354), .ZN(n8612) );
  NAND2_X1 U5076 ( .A1(n6366), .A2(n6365), .ZN(n8606) );
  OR2_X1 U5077 ( .A1(n7601), .A2(n4911), .ZN(n7481) );
  NAND2_X1 U5078 ( .A1(n5424), .A2(n5423), .ZN(n9431) );
  INV_X1 U5079 ( .A(n8823), .ZN(n8820) );
  NAND2_X1 U5080 ( .A1(n5376), .A2(n5375), .ZN(n9616) );
  NOR2_X1 U5081 ( .A1(n7411), .A2(n4949), .ZN(n4948) );
  NAND2_X1 U5082 ( .A1(n7219), .A2(n6559), .ZN(n4889) );
  AND2_X1 U5083 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n5584), .ZN(n5600) );
  NAND2_X1 U5084 ( .A1(n5309), .A2(n5308), .ZN(n5326) );
  INV_X2 U5085 ( .A(n10005), .ZN(n4500) );
  AND2_X1 U5086 ( .A1(n6162), .A2(n6161), .ZN(n10032) );
  NAND2_X1 U5087 ( .A1(n9883), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9882) );
  NOR2_X2 U5088 ( .A1(n6009), .A2(P1_U3086), .ZN(n6010) );
  AOI21_X1 U5089 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7087), .A(n9493), .ZN(
        n9510) );
  AND2_X1 U5090 ( .A1(n6855), .A2(n6858), .ZN(n9883) );
  INV_X1 U5091 ( .A(n9664), .ZN(n9651) );
  AOI21_X1 U5092 ( .B1(n5263), .B2(n5109), .A(n5108), .ZN(n5290) );
  NAND2_X1 U5093 ( .A1(n6133), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6106) );
  INV_X1 U5094 ( .A(n5971), .ZN(n5990) );
  NAND4_X1 U5095 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .ZN(n7187)
         );
  NAND4_X1 U5096 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n9049)
         );
  BUF_X2 U5097 ( .A(n6117), .Z(n7347) );
  AND2_X1 U5098 ( .A1(n6056), .A2(n6055), .ZN(n6467) );
  OR2_X1 U5099 ( .A1(n5425), .A2(n7723), .ZN(n5447) );
  NAND2_X1 U5100 ( .A1(n8648), .A2(n6083), .ZN(n6147) );
  NAND2_X1 U5101 ( .A1(n9842), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9868) );
  AND2_X1 U5102 ( .A1(n5749), .A2(n6007), .ZN(n5754) );
  AOI21_X1 U5103 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9549), .A(n9539), .ZN(
        n9557) );
  CLKBUF_X3 U5104 ( .A(n5226), .Z(n6722) );
  INV_X1 U5105 ( .A(n6084), .ZN(n8648) );
  OR2_X1 U5106 ( .A1(n5704), .A2(n5703), .ZN(n5755) );
  AND2_X1 U5107 ( .A1(n5122), .A2(n5121), .ZN(n5168) );
  INV_X1 U5108 ( .A(n6083), .ZN(n7865) );
  NAND2_X2 U5109 ( .A1(n4529), .A2(n6512), .ZN(n8273) );
  AND2_X1 U5110 ( .A1(n7862), .A2(n7849), .ZN(n5226) );
  NAND2_X1 U5111 ( .A1(n6707), .A2(n8014), .ZN(n5209) );
  AND2_X1 U5112 ( .A1(n5702), .A2(n6001), .ZN(n5750) );
  AND2_X1 U5113 ( .A1(n5151), .A2(n7849), .ZN(n5223) );
  NAND2_X1 U5114 ( .A1(n5151), .A2(n5149), .ZN(n5199) );
  NAND3_X1 U5115 ( .A1(n5728), .A2(n5745), .A3(n7751), .ZN(n6007) );
  NAND2_X1 U5116 ( .A1(n5660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5712) );
  OR2_X1 U5117 ( .A1(n6080), .A2(n8644), .ZN(n6078) );
  INV_X1 U5118 ( .A(n6001), .ZN(n5701) );
  OR2_X1 U5119 ( .A1(n9451), .A2(n9452), .ZN(n5145) );
  XNOR2_X1 U5120 ( .A(n4760), .B(n4759), .ZN(n6001) );
  NAND2_X2 U5121 ( .A1(n6680), .A2(P2_U3151), .ZN(n8650) );
  NAND2_X1 U5122 ( .A1(n6042), .A2(n6041), .ZN(n6063) );
  AND2_X1 U5123 ( .A1(n5657), .A2(n5075), .ZN(n5082) );
  INV_X1 U5124 ( .A(n5420), .ZN(n4501) );
  NAND4_X1 U5125 ( .A1(n4761), .A2(n4510), .A3(n4654), .A4(n4505), .ZN(n5456)
         );
  NOR2_X1 U5126 ( .A1(n6029), .A2(n6028), .ZN(n5074) );
  AND3_X1 U5127 ( .A1(n5130), .A2(n5270), .A3(n5235), .ZN(n5195) );
  OR2_X1 U5128 ( .A1(n5235), .A2(n9452), .ZN(n5272) );
  INV_X1 U5130 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5351) );
  INV_X1 U5131 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n10274) );
  NOR2_X1 U5132 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5270) );
  NOR2_X1 U5133 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5235) );
  INV_X4 U5134 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5135 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n10333) );
  NOR2_X2 U5136 ( .A1(n9300), .A2(n5468), .ZN(n9287) );
  OAI211_X1 U5137 ( .C1(n6675), .C2(n6846), .A(n6101), .B(n4754), .ZN(n6553)
         );
  NOR2_X1 U5138 ( .A1(n4508), .A2(n8500), .ZN(n4870) );
  INV_X1 U5139 ( .A(n5433), .ZN(n5434) );
  INV_X1 U5140 ( .A(n8745), .ZN(n4647) );
  NAND2_X1 U5141 ( .A1(n9225), .A2(n4799), .ZN(n4795) );
  NOR2_X1 U5142 ( .A1(n5693), .A2(n4802), .ZN(n4799) );
  OAI21_X1 U5143 ( .B1(n8072), .B2(n8182), .A(n8073), .ZN(n4757) );
  AND2_X1 U5144 ( .A1(n8129), .A2(n8482), .ZN(n4749) );
  NAND2_X1 U5145 ( .A1(n4728), .A2(n4729), .ZN(n8177) );
  OR2_X1 U5146 ( .A1(n8162), .A2(n4733), .ZN(n4728) );
  NOR2_X1 U5147 ( .A1(n7289), .A2(n7288), .ZN(n5043) );
  NAND2_X1 U5148 ( .A1(n4723), .A2(n4722), .ZN(n4721) );
  NOR2_X1 U5149 ( .A1(n9740), .A2(n4892), .ZN(n5680) );
  NOR2_X1 U5150 ( .A1(n5680), .A2(n7390), .ZN(n4780) );
  INV_X1 U5151 ( .A(n4970), .ZN(n4969) );
  OAI21_X1 U5152 ( .B1(n5574), .B2(n4971), .A(n5591), .ZN(n4970) );
  AND2_X1 U5153 ( .A1(n5470), .A2(SI_18_), .ZN(n5475) );
  INV_X1 U5154 ( .A(n6410), .ZN(n7829) );
  OR2_X1 U5155 ( .A1(n8284), .A2(n8287), .ZN(n8207) );
  NAND2_X1 U5156 ( .A1(n4755), .A2(n6553), .ZN(n6602) );
  OR2_X1 U5157 ( .A1(n7352), .A2(n6121), .ZN(n6122) );
  OR2_X1 U5158 ( .A1(n8588), .A2(n7966), .ZN(n8175) );
  OR2_X1 U5159 ( .A1(n8600), .A2(n6574), .ZN(n8165) );
  OR2_X1 U5160 ( .A1(n6618), .A2(n7907), .ZN(n8151) );
  INV_X1 U5161 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4998) );
  OR2_X1 U5162 ( .A1(n8625), .A2(n8001), .ZN(n8146) );
  NAND2_X1 U5163 ( .A1(n8687), .A2(n5947), .ZN(n5953) );
  INV_X1 U5164 ( .A(n5752), .ZN(n5749) );
  AOI21_X1 U5165 ( .B1(n7630), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7629), .ZN(
        n7717) );
  INV_X1 U5166 ( .A(n9179), .ZN(n4873) );
  NOR2_X1 U5167 ( .A1(n9256), .A2(n9262), .ZN(n9240) );
  NAND2_X1 U5168 ( .A1(n9782), .A2(n9788), .ZN(n4818) );
  NOR2_X1 U5169 ( .A1(n7469), .A2(n9616), .ZN(n4666) );
  INV_X1 U5170 ( .A(n5680), .ZN(n4781) );
  OR2_X1 U5171 ( .A1(n9050), .A2(n9698), .ZN(n5678) );
  NAND2_X1 U5172 ( .A1(n7855), .A2(n7854), .ZN(n8013) );
  OR2_X1 U5173 ( .A1(n7853), .A2(n7852), .ZN(n7854) );
  OR2_X1 U5174 ( .A1(n7851), .A2(n7850), .ZN(n7855) );
  NAND2_X1 U5175 ( .A1(n5081), .A2(n5053), .ZN(n5055) );
  AND2_X1 U5176 ( .A1(n5056), .A2(n5058), .ZN(n5053) );
  NOR2_X1 U5177 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5056) );
  OAI21_X1 U5178 ( .B1(n5511), .B2(n5510), .A(n5509), .ZN(n5513) );
  NOR2_X1 U5179 ( .A1(n5418), .A2(n4985), .ZN(n4984) );
  INV_X1 U5180 ( .A(SI_15_), .ZN(n4985) );
  NAND2_X1 U5181 ( .A1(n4857), .A2(n4855), .ZN(n5303) );
  AND2_X1 U5182 ( .A1(n4856), .A2(n5126), .ZN(n4855) );
  XNOR2_X1 U5183 ( .A(n5299), .B(SI_9_), .ZN(n5302) );
  NOR2_X1 U5184 ( .A1(n4521), .A2(n4556), .ZN(n4753) );
  NAND2_X1 U5185 ( .A1(n6065), .A2(n4751), .ZN(n4750) );
  INV_X1 U5186 ( .A(n6344), .ZN(n6591) );
  INV_X1 U5187 ( .A(n7349), .ZN(n6593) );
  OR2_X1 U5188 ( .A1(n6262), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6263) );
  INV_X1 U5189 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U5190 ( .A1(n6077), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6511) );
  INV_X1 U5191 ( .A(n8185), .ZN(n8188) );
  INV_X1 U5192 ( .A(n6427), .ZN(n6426) );
  OR2_X1 U5193 ( .A1(n6386), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6401) );
  AND4_X1 U5194 ( .A1(n6141), .A2(n6140), .A3(n6139), .A4(n6138), .ZN(n8096)
         );
  NAND2_X1 U5195 ( .A1(n4886), .A2(n8484), .ZN(n6643) );
  XNOR2_X1 U5196 ( .A(n6600), .B(n8185), .ZN(n4886) );
  AND2_X1 U5197 ( .A1(n8304), .A2(n8320), .ZN(n6587) );
  OR2_X1 U5198 ( .A1(n8172), .A2(n8332), .ZN(n6625) );
  INV_X1 U5199 ( .A(n8319), .ZN(n8348) );
  OR2_X1 U5200 ( .A1(n6575), .A2(n7966), .ZN(n5071) );
  NAND2_X1 U5201 ( .A1(n5009), .A2(n5013), .ZN(n5010) );
  INV_X1 U5202 ( .A(n8375), .ZN(n5009) );
  OR2_X1 U5203 ( .A1(n8621), .A2(n7907), .ZN(n5077) );
  OR2_X1 U5204 ( .A1(n4866), .A2(n4536), .ZN(n4863) );
  AOI21_X1 U5205 ( .B1(n4869), .B2(n4867), .A(n4522), .ZN(n4865) );
  AND2_X1 U5206 ( .A1(n6030), .A2(n6031), .ZN(n4957) );
  INV_X1 U5207 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6031) );
  OAI21_X1 U5208 ( .B1(n5064), .B2(n5066), .A(n5068), .ZN(n5063) );
  INV_X1 U5209 ( .A(n6531), .ZN(n5068) );
  NAND2_X1 U5210 ( .A1(n5887), .A2(n8655), .ZN(n8656) );
  NAND2_X1 U5211 ( .A1(n4650), .A2(n5886), .ZN(n5887) );
  OAI21_X1 U5212 ( .B1(n7758), .B2(n5038), .A(n4648), .ZN(n4650) );
  INV_X1 U5213 ( .A(n5064), .ZN(n4612) );
  NAND2_X1 U5214 ( .A1(n8722), .A2(n5066), .ZN(n4613) );
  NAND2_X1 U5215 ( .A1(n5241), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5216) );
  OAI22_X1 U5216 ( .A1(n9252), .A2(n5691), .B1(n9401), .B2(n9277), .ZN(n9239)
         );
  INV_X1 U5217 ( .A(n4807), .ZN(n4806) );
  OAI21_X1 U5218 ( .B1(n4504), .B2(n9004), .A(n5685), .ZN(n4807) );
  OR2_X1 U5219 ( .A1(n9616), .A2(n9788), .ZN(n9609) );
  AOI22_X1 U5220 ( .A1(n9625), .A2(n9627), .B1(n9748), .B2(n9759), .ZN(n7464)
         );
  INV_X1 U5221 ( .A(n6707), .ZN(n5484) );
  AOI21_X1 U5223 ( .B1(n4974), .B2(n4976), .A(n4973), .ZN(n4972) );
  INV_X1 U5224 ( .A(n4976), .ZN(n4975) );
  INV_X1 U5225 ( .A(n5363), .ZN(n4973) );
  NAND2_X1 U5226 ( .A1(n5370), .A2(n5369), .ZN(n5384) );
  NAND2_X1 U5227 ( .A1(n5326), .A2(n4982), .ZN(n4978) );
  NAND2_X1 U5228 ( .A1(n5326), .A2(n5325), .ZN(n5339) );
  INV_X1 U5229 ( .A(n8297), .ZN(n8333) );
  INV_X1 U5230 ( .A(n8251), .ZN(n8279) );
  OR2_X1 U5231 ( .A1(n9876), .A2(n4627), .ZN(n4624) );
  NAND2_X1 U5232 ( .A1(n4629), .A2(n4628), .ZN(n4627) );
  INV_X1 U5233 ( .A(n9877), .ZN(n4628) );
  INV_X1 U5234 ( .A(n9893), .ZN(n4629) );
  INV_X1 U5235 ( .A(n4626), .ZN(n4625) );
  OAI22_X1 U5236 ( .A1(n9893), .A2(n4630), .B1(n6830), .B2(n9888), .ZN(n4626)
         );
  AND2_X1 U5237 ( .A1(n6000), .A2(n8777), .ZN(n4652) );
  INV_X1 U5238 ( .A(n9149), .ZN(n4826) );
  NAND2_X1 U5239 ( .A1(n4827), .A2(n9777), .ZN(n4823) );
  OAI22_X1 U5240 ( .A1(n9359), .A2(n9787), .B1(n9789), .B2(n9148), .ZN(n9149)
         );
  OAI21_X1 U5241 ( .B1(n8805), .B2(n8909), .A(n8804), .ZN(n4677) );
  INV_X1 U5242 ( .A(n8836), .ZN(n4692) );
  AND2_X1 U5243 ( .A1(n9317), .A2(n4695), .ZN(n4694) );
  NAND2_X1 U5244 ( .A1(n8929), .A2(n4696), .ZN(n4695) );
  OR2_X1 U5245 ( .A1(n8930), .A2(n4697), .ZN(n4696) );
  INV_X1 U5246 ( .A(n8926), .ZN(n4697) );
  NOR2_X1 U5247 ( .A1(n8930), .A2(n4699), .ZN(n4698) );
  INV_X1 U5248 ( .A(n8847), .ZN(n4699) );
  NAND2_X1 U5249 ( .A1(n4709), .A2(n4708), .ZN(n8161) );
  AOI21_X1 U5250 ( .B1(n4732), .B2(n4730), .A(n4550), .ZN(n4729) );
  INV_X1 U5251 ( .A(n8163), .ZN(n4730) );
  NAND2_X1 U5252 ( .A1(n8187), .A2(n4514), .ZN(n4715) );
  AND2_X1 U5253 ( .A1(n4688), .A2(n4689), .ZN(n4685) );
  NOR2_X1 U5254 ( .A1(n8792), .A2(n4511), .ZN(n4689) );
  INV_X1 U5255 ( .A(n5576), .ZN(n4971) );
  OR2_X1 U5256 ( .A1(n6654), .A2(n6599), .ZN(n8206) );
  OR2_X1 U5257 ( .A1(n8557), .A2(n8051), .ZN(n8212) );
  NOR2_X1 U5258 ( .A1(n4714), .A2(n4721), .ZN(n4713) );
  NAND2_X1 U5259 ( .A1(n6848), .A2(n6847), .ZN(n6850) );
  INV_X1 U5260 ( .A(n7430), .ZN(n4929) );
  AOI21_X1 U5261 ( .B1(n7430), .B2(n7551), .A(n7433), .ZN(n4928) );
  NAND2_X1 U5262 ( .A1(n4926), .A2(n4925), .ZN(n4924) );
  NAND2_X1 U5263 ( .A1(n8236), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4925) );
  INV_X1 U5264 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6233) );
  NOR2_X1 U5265 ( .A1(n6367), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U5266 ( .A1(n4607), .A2(n6300), .ZN(n6314) );
  NOR2_X1 U5267 ( .A1(n6287), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n4607) );
  INV_X1 U5268 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7619) );
  NOR2_X1 U5269 ( .A1(n6245), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n4606) );
  INV_X1 U5270 ( .A(n4890), .ZN(n4888) );
  NAND2_X1 U5271 ( .A1(n10032), .A2(n4891), .ZN(n4890) );
  OR2_X1 U5272 ( .A1(n4891), .A2(n10032), .ZN(n6559) );
  NAND2_X1 U5273 ( .A1(n6602), .A2(n8069), .ZN(n8070) );
  NAND2_X1 U5274 ( .A1(n6548), .A2(n6549), .ZN(n8067) );
  NAND3_X1 U5275 ( .A1(n6467), .A2(n6466), .A3(n10318), .ZN(n6471) );
  OR2_X1 U5276 ( .A1(n8511), .A2(n8333), .ZN(n8020) );
  NAND2_X1 U5277 ( .A1(n5022), .A2(n8021), .ZN(n5021) );
  INV_X1 U5278 ( .A(n5024), .ZN(n5022) );
  AND2_X1 U5279 ( .A1(n8511), .A2(n8333), .ZN(n8184) );
  AND2_X1 U5280 ( .A1(n6576), .A2(n4540), .ZN(n4899) );
  OR2_X1 U5281 ( .A1(n6623), .A2(n8347), .ZN(n8176) );
  AOI21_X1 U5282 ( .B1(n4851), .B2(n8413), .A(n4849), .ZN(n4848) );
  INV_X1 U5283 ( .A(n8391), .ZN(n4849) );
  INV_X1 U5284 ( .A(n4851), .ZN(n4850) );
  NOR2_X1 U5285 ( .A1(n6572), .A2(n4852), .ZN(n4851) );
  INV_X1 U5286 ( .A(n8403), .ZN(n4852) );
  OR2_X1 U5287 ( .A1(n8606), .A2(n7915), .ZN(n8058) );
  AND2_X1 U5288 ( .A1(n5034), .A2(n8130), .ZN(n5033) );
  NAND2_X1 U5289 ( .A1(n6613), .A2(n6614), .ZN(n5034) );
  INV_X1 U5290 ( .A(n8131), .ZN(n5030) );
  INV_X2 U5291 ( .A(n6063), .ZN(n6065) );
  AOI21_X1 U5292 ( .B1(n4617), .B2(n4615), .A(n4525), .ZN(n4614) );
  INV_X1 U5293 ( .A(n4617), .ZN(n4616) );
  NOR2_X1 U5294 ( .A1(n5052), .A2(n5049), .ZN(n5048) );
  INV_X1 U5295 ( .A(n5903), .ZN(n5049) );
  AND2_X1 U5296 ( .A1(n5923), .A2(n5051), .ZN(n5050) );
  OR2_X1 U5297 ( .A1(n8715), .A2(n5052), .ZN(n5051) );
  INV_X1 U5298 ( .A(n5963), .ZN(n4767) );
  NAND2_X1 U5299 ( .A1(n4568), .A2(n5040), .ZN(n5039) );
  OR2_X1 U5300 ( .A1(n9691), .A2(n5798), .ZN(n5780) );
  AND2_X1 U5301 ( .A1(n5784), .A2(n5783), .ZN(n5787) );
  NAND2_X1 U5302 ( .A1(n5892), .A2(n5891), .ZN(n5895) );
  NAND2_X1 U5303 ( .A1(n8656), .A2(n8654), .ZN(n5892) );
  NAND2_X1 U5304 ( .A1(n8984), .A2(n4991), .ZN(n9012) );
  NOR2_X1 U5305 ( .A1(n9156), .A2(n4992), .ZN(n4991) );
  NAND2_X1 U5306 ( .A1(n4997), .A2(n4993), .ZN(n4992) );
  AND2_X1 U5307 ( .A1(n8896), .A2(n9128), .ZN(n9018) );
  NAND2_X1 U5308 ( .A1(n4687), .A2(n4686), .ZN(n8895) );
  OR2_X1 U5309 ( .A1(n8979), .A2(n9031), .ZN(n4686) );
  NAND2_X1 U5310 ( .A1(n8894), .A2(n8979), .ZN(n4687) );
  OR2_X1 U5311 ( .A1(n9413), .A2(n9417), .ZN(n8844) );
  NAND2_X1 U5312 ( .A1(n8665), .A2(n9612), .ZN(n4817) );
  INV_X1 U5313 ( .A(n8830), .ZN(n9606) );
  NAND2_X1 U5314 ( .A1(n4774), .A2(n4773), .ZN(n4772) );
  NOR2_X1 U5315 ( .A1(n4780), .A2(n7264), .ZN(n4773) );
  OR2_X1 U5316 ( .A1(n4573), .A2(n4780), .ZN(n4775) );
  INV_X1 U5317 ( .A(n7397), .ZN(n4787) );
  INV_X1 U5318 ( .A(n7263), .ZN(n4774) );
  NAND2_X1 U5319 ( .A1(n4893), .A2(n4892), .ZN(n8824) );
  NAND2_X1 U5320 ( .A1(n7293), .A2(n4789), .ZN(n4788) );
  NAND2_X1 U5321 ( .A1(n7262), .A2(n7163), .ZN(n8803) );
  INV_X1 U5322 ( .A(n5677), .ZN(n8908) );
  AND2_X1 U5323 ( .A1(n9723), .A2(n9729), .ZN(n4792) );
  XNOR2_X1 U5324 ( .A(n7853), .B(n7852), .ZN(n7851) );
  AOI21_X1 U5325 ( .B1(n5630), .B2(n5629), .A(n4598), .ZN(n5641) );
  INV_X1 U5326 ( .A(n5631), .ZN(n4598) );
  NAND2_X1 U5327 ( .A1(n5081), .A2(n5058), .ZN(n5057) );
  OAI21_X1 U5328 ( .B1(n5420), .B2(n5057), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5716) );
  AND2_X1 U5329 ( .A1(n5576), .A2(n5566), .ZN(n5574) );
  OR2_X1 U5330 ( .A1(n5475), .A2(n5474), .ZN(n5494) );
  OR2_X1 U5331 ( .A1(n5471), .A2(n5475), .ZN(n5493) );
  NOR2_X1 U5332 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5128) );
  NOR2_X1 U5333 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5127) );
  AND4_X1 U5334 ( .A1(n5130), .A2(n5270), .A3(n5235), .A4(n5058), .ZN(n4761)
         );
  AND4_X1 U5335 ( .A1(n5351), .A2(n5345), .A3(n5129), .A4(n5405), .ZN(n4505)
         );
  OAI21_X1 U5336 ( .B1(n5400), .B2(SI_14_), .A(n5399), .ZN(n5402) );
  NAND2_X1 U5337 ( .A1(n5384), .A2(n5383), .ZN(n5400) );
  NAND2_X1 U5338 ( .A1(n5365), .A2(SI_13_), .ZN(n5383) );
  NAND2_X1 U5339 ( .A1(n5340), .A2(SI_12_), .ZN(n5363) );
  NOR2_X1 U5340 ( .A1(n5338), .A2(n4983), .ZN(n4982) );
  INV_X1 U5341 ( .A(n5325), .ZN(n4983) );
  INV_X1 U5342 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5345) );
  XNOR2_X1 U5343 ( .A(n5337), .B(SI_11_), .ZN(n5338) );
  XNOR2_X1 U5344 ( .A(n5123), .B(SI_8_), .ZN(n5156) );
  AOI21_X1 U5345 ( .B1(n5168), .B2(n4861), .A(n4860), .ZN(n4859) );
  INV_X1 U5346 ( .A(n5122), .ZN(n4860) );
  INV_X1 U5347 ( .A(n5118), .ZN(n4861) );
  INV_X1 U5348 ( .A(n5168), .ZN(n4862) );
  NAND2_X1 U5349 ( .A1(n5119), .A2(SI_7_), .ZN(n5122) );
  INV_X1 U5350 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5344) );
  INV_X1 U5351 ( .A(SI_5_), .ZN(n10364) );
  NOR2_X1 U5352 ( .A1(n4554), .A2(n4952), .ZN(n4951) );
  INV_X1 U5353 ( .A(n4954), .ZN(n4952) );
  OAI21_X1 U5354 ( .B1(n7231), .B2(n4947), .A(n4945), .ZN(n6230) );
  INV_X1 U5355 ( .A(n4948), .ZN(n4947) );
  AOI21_X1 U5356 ( .B1(n4946), .B2(n4948), .A(n4543), .ZN(n4945) );
  NOR2_X1 U5357 ( .A1(n6498), .A2(n4935), .ZN(n4934) );
  INV_X1 U5358 ( .A(n6450), .ZN(n4935) );
  INV_X1 U5359 ( .A(n8228), .ZN(n6609) );
  NOR2_X1 U5360 ( .A1(n7939), .A2(n4938), .ZN(n4937) );
  INV_X1 U5361 ( .A(n6322), .ZN(n4938) );
  NAND2_X1 U5362 ( .A1(n4941), .A2(n7946), .ZN(n7919) );
  OR2_X1 U5363 ( .A1(n7973), .A2(n4933), .ZN(n4932) );
  INV_X1 U5364 ( .A(n6353), .ZN(n4933) );
  OR2_X1 U5365 ( .A1(n7652), .A2(n8223), .ZN(n4955) );
  OR2_X1 U5366 ( .A1(n7020), .A2(n7019), .ZN(n7334) );
  NAND2_X1 U5367 ( .A1(n6474), .A2(n6473), .ZN(n6776) );
  INV_X1 U5368 ( .A(n7732), .ZN(n6474) );
  AND2_X1 U5369 ( .A1(n7480), .A2(n7604), .ZN(n7601) );
  XNOR2_X1 U5370 ( .A(n4924), .B(n4923), .ZN(n9908) );
  NOR2_X1 U5371 ( .A1(n9908), .A2(n6266), .ZN(n9907) );
  INV_X1 U5372 ( .A(n8259), .ZN(n4640) );
  AND2_X1 U5373 ( .A1(n7486), .A2(n7485), .ZN(n7611) );
  OR2_X1 U5374 ( .A1(n4641), .A2(n4594), .ZN(n4639) );
  OR2_X1 U5375 ( .A1(n9941), .A2(n9940), .ZN(n4918) );
  OR2_X1 U5376 ( .A1(n9978), .A2(n9977), .ZN(n4922) );
  OR2_X1 U5377 ( .A1(n9978), .A2(n4921), .ZN(n4919) );
  OR2_X1 U5378 ( .A1(n4535), .A2(n9475), .ZN(n4920) );
  OR2_X1 U5379 ( .A1(n9475), .A2(n9977), .ZN(n4921) );
  NAND2_X1 U5380 ( .A1(n4605), .A2(n6411), .ZN(n6427) );
  OR2_X1 U5381 ( .A1(n6345), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U5382 ( .A1(n8440), .A2(n4547), .ZN(n8425) );
  OR2_X1 U5383 ( .A1(n6314), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6330) );
  AOI21_X1 U5384 ( .B1(n8449), .B2(n8144), .A(n6616), .ZN(n8441) );
  NAND2_X1 U5385 ( .A1(n8451), .A2(n5076), .ZN(n8436) );
  OR2_X1 U5386 ( .A1(n7936), .A2(n8001), .ZN(n5076) );
  AND2_X1 U5387 ( .A1(n10054), .A2(n8224), .ZN(n6566) );
  INV_X1 U5388 ( .A(n8482), .ZN(n8127) );
  INV_X1 U5389 ( .A(n8227), .ZN(n7549) );
  NAND2_X1 U5390 ( .A1(n7375), .A2(n8082), .ZN(n5017) );
  NAND2_X1 U5391 ( .A1(n5017), .A2(n5016), .ZN(n7587) );
  AND2_X1 U5392 ( .A1(n8036), .A2(n8104), .ZN(n5016) );
  OR2_X1 U5393 ( .A1(n6198), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6212) );
  NOR2_X1 U5394 ( .A1(n6555), .A2(n4838), .ZN(n4837) );
  INV_X1 U5395 ( .A(n6554), .ZN(n4838) );
  NAND2_X1 U5396 ( .A1(n4841), .A2(n7194), .ZN(n4840) );
  NAND2_X1 U5397 ( .A1(n8070), .A2(n9991), .ZN(n4839) );
  NAND2_X1 U5398 ( .A1(n6297), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4754) );
  INV_X1 U5399 ( .A(n8026), .ZN(n8064) );
  INV_X1 U5400 ( .A(n6642), .ZN(n5006) );
  NAND2_X1 U5401 ( .A1(n4569), .A2(n4900), .ZN(n4895) );
  NOR2_X1 U5402 ( .A1(n8053), .A2(n5025), .ZN(n5024) );
  INV_X1 U5403 ( .A(n6625), .ZN(n5025) );
  OR2_X1 U5404 ( .A1(n8183), .A2(n8184), .ZN(n8307) );
  NAND2_X1 U5405 ( .A1(n6424), .A2(n6423), .ZN(n8172) );
  OR2_X1 U5406 ( .A1(n6637), .A2(n8182), .ZN(n9993) );
  OR2_X1 U5407 ( .A1(n8182), .A2(n6632), .ZN(n9995) );
  AOI21_X1 U5408 ( .B1(n5013), .B2(n5012), .A(n4731), .ZN(n5011) );
  INV_X1 U5409 ( .A(n8056), .ZN(n5012) );
  AND2_X1 U5410 ( .A1(n5015), .A2(n8176), .ZN(n8359) );
  NAND2_X1 U5411 ( .A1(n6622), .A2(n8165), .ZN(n8375) );
  NAND2_X1 U5412 ( .A1(n4853), .A2(n4851), .ZN(n8402) );
  NAND2_X1 U5413 ( .A1(n8414), .A2(n6620), .ZN(n4853) );
  NAND2_X1 U5414 ( .A1(n6343), .A2(n6342), .ZN(n6618) );
  NAND2_X1 U5415 ( .A1(n8453), .A2(n8452), .ZN(n8451) );
  AOI21_X1 U5416 ( .B1(n4868), .B2(n4508), .A(n4559), .ZN(n4867) );
  INV_X1 U5417 ( .A(n9993), .ZN(n8479) );
  NAND2_X1 U5418 ( .A1(n6601), .A2(n8209), .ZN(n8484) );
  INV_X1 U5419 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6464) );
  OAI21_X1 U5420 ( .B1(n6032), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6033) );
  INV_X1 U5421 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n10184) );
  AND2_X1 U5422 ( .A1(n4957), .A2(n6037), .ZN(n4956) );
  NAND2_X1 U5423 ( .A1(n6098), .A2(n8644), .ZN(n4916) );
  XNOR2_X1 U5424 ( .A(n5760), .B(n5981), .ZN(n5766) );
  AOI21_X1 U5425 ( .B1(n6884), .B2(n5990), .A(n5762), .ZN(n5765) );
  NAND2_X1 U5426 ( .A1(n5939), .A2(n4549), .ZN(n8687) );
  NOR2_X1 U5427 ( .A1(n4771), .A2(n4767), .ZN(n4766) );
  AOI21_X1 U5428 ( .B1(n4770), .B2(n4585), .A(n8723), .ZN(n4769) );
  INV_X1 U5429 ( .A(n8666), .ZN(n4770) );
  XNOR2_X1 U5430 ( .A(n4653), .B(n5981), .ZN(n5806) );
  OAI21_X1 U5431 ( .B1(n5798), .B2(n9705), .A(n5799), .ZN(n4653) );
  NAND2_X1 U5432 ( .A1(n4619), .A2(n7756), .ZN(n7758) );
  NOR2_X1 U5433 ( .A1(n5953), .A2(n5952), .ZN(n8745) );
  NAND2_X1 U5434 ( .A1(n5953), .A2(n5952), .ZN(n8743) );
  AND2_X1 U5435 ( .A1(n5751), .A2(n6007), .ZN(n5753) );
  INV_X1 U5436 ( .A(n9018), .ZN(n9030) );
  AND2_X1 U5437 ( .A1(n9338), .A2(n8983), .ZN(n9015) );
  AND2_X1 U5438 ( .A1(n5272), .A2(n5271), .ZN(n5275) );
  NOR2_X1 U5439 ( .A1(n9544), .A2(n7080), .ZN(n9562) );
  XNOR2_X1 U5440 ( .A(n4603), .B(n4602), .ZN(n7881) );
  INV_X1 U5441 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n4602) );
  NAND2_X1 U5442 ( .A1(n9119), .A2(n7878), .ZN(n4603) );
  INV_X1 U5443 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7887) );
  OAI21_X1 U5444 ( .B1(n9178), .B2(n5698), .A(n5697), .ZN(n9161) );
  NAND2_X1 U5445 ( .A1(n5696), .A2(n9367), .ZN(n5697) );
  NAND2_X1 U5446 ( .A1(n4876), .A2(n8949), .ZN(n4875) );
  INV_X1 U5447 ( .A(n4878), .ZN(n4876) );
  OR2_X1 U5448 ( .A1(n9213), .A2(n4877), .ZN(n4874) );
  OR2_X1 U5449 ( .A1(n4880), .A2(n5590), .ZN(n4877) );
  INV_X1 U5450 ( .A(n4797), .ZN(n4796) );
  OAI21_X1 U5451 ( .B1(n5693), .B2(n4798), .A(n4800), .ZN(n4797) );
  NAND2_X1 U5452 ( .A1(n4801), .A2(n4533), .ZN(n4798) );
  OR2_X1 U5453 ( .A1(n9375), .A2(n9380), .ZN(n9191) );
  OAI22_X1 U5454 ( .A1(n9239), .A2(n5692), .B1(n9397), .B2(n9248), .ZN(n9225)
         );
  AOI21_X1 U5455 ( .B1(n9237), .B2(n9238), .A(n5542), .ZN(n9223) );
  NAND2_X1 U5456 ( .A1(n4905), .A2(n4903), .ZN(n9237) );
  AOI21_X1 U5457 ( .B1(n4906), .B2(n9275), .A(n4904), .ZN(n4903) );
  NAND2_X1 U5458 ( .A1(n9276), .A2(n4906), .ZN(n4905) );
  INV_X1 U5459 ( .A(n8865), .ZN(n4904) );
  AND2_X1 U5460 ( .A1(n9254), .A2(n8863), .ZN(n4906) );
  OR2_X1 U5461 ( .A1(n9276), .A2(n9275), .ZN(n4907) );
  AND2_X1 U5462 ( .A1(n9285), .A2(n8844), .ZN(n9276) );
  NAND2_X1 U5463 ( .A1(n5462), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5488) );
  OR2_X1 U5464 ( .A1(n5684), .A2(n4538), .ZN(n4504) );
  OR2_X1 U5465 ( .A1(n9426), .A2(n9418), .ZN(n9298) );
  AND2_X1 U5466 ( .A1(n9298), .A2(n8857), .ZN(n9317) );
  NAND2_X1 U5467 ( .A1(n5683), .A2(n5682), .ZN(n7811) );
  NAND2_X1 U5468 ( .A1(n9605), .A2(n4908), .ZN(n7693) );
  AND2_X1 U5469 ( .A1(n5398), .A2(n9609), .ZN(n4908) );
  NAND2_X1 U5470 ( .A1(n4814), .A2(n4818), .ZN(n4813) );
  INV_X1 U5471 ( .A(n4815), .ZN(n4814) );
  AOI21_X1 U5472 ( .B1(n8999), .B2(n4819), .A(n4816), .ZN(n4815) );
  NAND2_X1 U5473 ( .A1(n9607), .A2(n8928), .ZN(n9605) );
  NAND2_X1 U5474 ( .A1(n4820), .A2(n9611), .ZN(n4819) );
  AOI21_X1 U5475 ( .B1(n4830), .B2(n4832), .A(n4829), .ZN(n4828) );
  INV_X1 U5476 ( .A(n8827), .ZN(n4829) );
  NAND2_X1 U5477 ( .A1(n7465), .A2(n8999), .ZN(n9607) );
  NOR2_X1 U5478 ( .A1(n7363), .A2(n9636), .ZN(n9637) );
  AND2_X1 U5479 ( .A1(n5319), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5331) );
  OAI22_X1 U5480 ( .A1(n7362), .A2(n7361), .B1(n9629), .B2(n9751), .ZN(n9625)
         );
  NOR2_X1 U5481 ( .A1(n4792), .A2(n4783), .ZN(n4782) );
  NAND2_X1 U5482 ( .A1(n4788), .A2(n4793), .ZN(n4783) );
  INV_X1 U5483 ( .A(n4786), .ZN(n4785) );
  NAND2_X1 U5484 ( .A1(n4790), .A2(n4788), .ZN(n9643) );
  NAND2_X1 U5485 ( .A1(n7140), .A2(n8803), .ZN(n7387) );
  AOI22_X1 U5486 ( .A1(n7146), .A2(n8986), .B1(n7262), .B2(n9713), .ZN(n7263)
         );
  OR2_X1 U5487 ( .A1(n9662), .A2(n9705), .ZN(n8802) );
  OAI22_X1 U5488 ( .A1(n6984), .A2(n4528), .B1(n6988), .B2(n9662), .ZN(n7146)
         );
  NAND2_X1 U5489 ( .A1(n5461), .A2(n5460), .ZN(n9421) );
  OR2_X1 U5490 ( .A1(n5997), .A2(n4502), .ZN(n9787) );
  XNOR2_X1 U5491 ( .A(n8017), .B(n8016), .ZN(n8889) );
  OAI21_X1 U5492 ( .B1(n8013), .B2(n8012), .A(n8011), .ZN(n8017) );
  XNOR2_X1 U5493 ( .A(n8013), .B(n8012), .ZN(n8885) );
  NOR2_X1 U5494 ( .A1(n5055), .A2(n4679), .ZN(n4678) );
  NAND2_X1 U5495 ( .A1(n4821), .A2(n5134), .ZN(n4679) );
  NOR2_X1 U5496 ( .A1(n5055), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n4680) );
  NAND2_X1 U5497 ( .A1(n4586), .A2(n5543), .ZN(n4961) );
  INV_X1 U5498 ( .A(n5526), .ZN(n4962) );
  NOR2_X1 U5499 ( .A1(n5527), .A2(n4960), .ZN(n4959) );
  INV_X1 U5500 ( .A(n5543), .ZN(n4960) );
  XNOR2_X1 U5501 ( .A(n5662), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8988) );
  XNOR2_X1 U5502 ( .A(n5483), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U5503 ( .A1(n5482), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5483) );
  INV_X1 U5504 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5405) );
  AND2_X1 U5505 ( .A1(n5404), .A2(n5389), .ZN(n7630) );
  AND2_X1 U5506 ( .A1(n5374), .A2(n5386), .ZN(n7312) );
  OAI21_X1 U5507 ( .B1(n5340), .B2(SI_12_), .A(n5363), .ZN(n5341) );
  NOR2_X1 U5508 ( .A1(n4977), .A2(n5341), .ZN(n4976) );
  INV_X1 U5509 ( .A(n4979), .ZN(n4977) );
  NAND2_X1 U5510 ( .A1(n4981), .A2(n4980), .ZN(n4979) );
  INV_X1 U5511 ( .A(SI_11_), .ZN(n4980) );
  INV_X1 U5512 ( .A(n5337), .ZN(n4981) );
  INV_X1 U5513 ( .A(n5310), .ZN(n5308) );
  NAND2_X1 U5514 ( .A1(n5292), .A2(n5113), .ZN(n5192) );
  AND2_X1 U5515 ( .A1(n5118), .A2(n5117), .ZN(n5191) );
  NAND2_X1 U5516 ( .A1(n5192), .A2(n5191), .ZN(n5194) );
  AND2_X1 U5517 ( .A1(n6392), .A2(n6391), .ZN(n7960) );
  AND2_X1 U5518 ( .A1(n7989), .A2(n4934), .ZN(n7840) );
  NAND2_X1 U5519 ( .A1(n6993), .A2(n4548), .ZN(n7127) );
  NAND2_X1 U5520 ( .A1(n6326), .A2(n6325), .ZN(n8538) );
  OR2_X1 U5521 ( .A1(n6995), .A2(n6996), .ZN(n6993) );
  INV_X1 U5522 ( .A(n8405), .ZN(n8424) );
  NAND2_X1 U5523 ( .A1(n6265), .A2(n6264), .ZN(n8129) );
  OR2_X1 U5524 ( .A1(n6781), .A2(n6279), .ZN(n6265) );
  NAND2_X1 U5525 ( .A1(n6500), .A2(n9989), .ZN(n7968) );
  INV_X1 U5526 ( .A(n8454), .ZN(n8423) );
  OR2_X1 U5527 ( .A1(n6931), .A2(n8214), .ZN(n7994) );
  AOI21_X1 U5528 ( .B1(n4736), .B2(n4735), .A(n4734), .ZN(n8213) );
  AND2_X1 U5529 ( .A1(n8284), .A2(n8287), .ZN(n4734) );
  AOI21_X1 U5530 ( .B1(n8211), .B2(n4596), .A(n4518), .ZN(n4735) );
  NAND2_X1 U5531 ( .A1(n6462), .A2(n6461), .ZN(n8297) );
  NAND2_X1 U5532 ( .A1(n6447), .A2(n6446), .ZN(n8319) );
  NAND4_X2 U5533 ( .A1(n6156), .A2(n6155), .A3(n6154), .A4(n6153), .ZN(n8230)
         );
  XNOR2_X1 U5534 ( .A(n6796), .B(n6805), .ZN(n9838) );
  NOR2_X1 U5535 ( .A1(n6772), .A2(n6806), .ZN(n9837) );
  AND2_X1 U5536 ( .A1(n4624), .A2(n4587), .ZN(n6908) );
  INV_X1 U5537 ( .A(n6832), .ZN(n4623) );
  NAND2_X1 U5538 ( .A1(n6914), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7030) );
  NOR2_X1 U5539 ( .A1(n6910), .A2(n6909), .ZN(n7014) );
  AND2_X1 U5540 ( .A1(n6284), .A2(n6295), .ZN(n9914) );
  OR2_X1 U5541 ( .A1(n6178), .A2(n5008), .ZN(n6310) );
  INV_X1 U5542 ( .A(n5074), .ZN(n5008) );
  XNOR2_X1 U5543 ( .A(n8277), .B(n8276), .ZN(n4644) );
  AOI21_X1 U5544 ( .B1(n9964), .B2(n8279), .A(n4643), .ZN(n4642) );
  OAI21_X1 U5545 ( .B1(n9897), .B2(n5000), .A(n8278), .ZN(n4643) );
  AOI21_X1 U5546 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n9468), .A(n9473), .ZN(
        n8242) );
  OR2_X1 U5547 ( .A1(n8233), .A2(n8215), .ZN(n9875) );
  NAND2_X1 U5548 ( .A1(n6440), .A2(n6439), .ZN(n8340) );
  NAND2_X1 U5549 ( .A1(n6261), .A2(n6260), .ZN(n7748) );
  OR2_X1 U5550 ( .A1(n6743), .A2(n6279), .ZN(n6261) );
  INV_X1 U5551 ( .A(n6553), .ZN(n10013) );
  OR2_X1 U5552 ( .A1(n6668), .A2(n10079), .ZN(n6671) );
  NAND2_X1 U5553 ( .A1(n6397), .A2(n6396), .ZN(n8588) );
  NAND2_X1 U5554 ( .A1(n6472), .A2(n7767), .ZN(n6735) );
  XNOR2_X1 U5555 ( .A(n6061), .B(n6060), .ZN(n8251) );
  XNOR2_X1 U5556 ( .A(n6160), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6917) );
  OR2_X1 U5557 ( .A1(n6159), .A2(n8644), .ZN(n6160) );
  NAND2_X1 U5558 ( .A1(n5061), .A2(n6532), .ZN(n5060) );
  NAND2_X1 U5559 ( .A1(n5062), .A2(n5064), .ZN(n5061) );
  INV_X1 U5560 ( .A(n5063), .ZN(n5062) );
  AND4_X1 U5561 ( .A1(n5508), .A2(n5507), .A3(n5506), .A4(n5505), .ZN(n9288)
         );
  AND2_X1 U5562 ( .A1(n5069), .A2(n4574), .ZN(n6533) );
  AND4_X1 U5563 ( .A1(n5382), .A2(n5381), .A3(n5380), .A4(n5379), .ZN(n9788)
         );
  AND4_X1 U5564 ( .A1(n5336), .A2(n5335), .A3(n5334), .A4(n5333), .ZN(n9748)
         );
  INV_X1 U5565 ( .A(n8697), .ZN(n5067) );
  INV_X1 U5566 ( .A(n6010), .ZN(n8750) );
  AND2_X1 U5567 ( .A1(n6011), .A2(n5998), .ZN(n8777) );
  INV_X1 U5568 ( .A(n4986), .ZN(n4674) );
  NAND2_X1 U5569 ( .A1(n4988), .A2(n5701), .ZN(n4987) );
  OAI21_X1 U5570 ( .B1(n9023), .B2(n5701), .A(n9024), .ZN(n4986) );
  AOI21_X1 U5571 ( .B1(n9028), .B2(n9021), .A(n8899), .ZN(n4675) );
  NAND2_X1 U5572 ( .A1(n5226), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U5573 ( .A1(n5537), .A2(n6957), .ZN(n5242) );
  NAND2_X1 U5574 ( .A1(n5226), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4672) );
  AND3_X1 U5575 ( .A1(n5217), .A2(n5216), .A3(n5215), .ZN(n5218) );
  CLKBUF_X1 U5576 ( .A(n5703), .Z(n9021) );
  NAND2_X1 U5577 ( .A1(n5517), .A2(n5516), .ZN(n9262) );
  NAND2_X1 U5578 ( .A1(n5355), .A2(n5354), .ZN(n7469) );
  OR2_X1 U5579 ( .A1(n6743), .A2(n5209), .ZN(n5355) );
  NAND2_X1 U5580 ( .A1(n9348), .A2(n4604), .ZN(n9437) );
  AND2_X1 U5581 ( .A1(n4822), .A2(n9347), .ZN(n4604) );
  CLKBUF_X1 U5582 ( .A(n5704), .Z(n7542) );
  OAI21_X1 U5583 ( .B1(n4758), .B2(n8061), .A(n4756), .ZN(n8093) );
  NAND2_X1 U5584 ( .A1(n8065), .A2(n4544), .ZN(n4758) );
  INV_X1 U5585 ( .A(n4757), .ZN(n4756) );
  OAI21_X1 U5586 ( .B1(n8807), .B2(n9031), .A(n4676), .ZN(n8813) );
  AOI21_X1 U5587 ( .B1(n4677), .B2(n4516), .A(n4561), .ZN(n4676) );
  AOI21_X1 U5588 ( .B1(n4565), .B2(n8128), .A(n4746), .ZN(n4745) );
  NOR2_X1 U5589 ( .A1(n8125), .A2(n4747), .ZN(n4746) );
  INV_X1 U5590 ( .A(n4749), .ZN(n4747) );
  AOI21_X1 U5591 ( .B1(n4745), .B2(n4748), .A(n4744), .ZN(n4743) );
  NOR2_X1 U5592 ( .A1(n8128), .A2(n4749), .ZN(n4748) );
  NAND2_X1 U5593 ( .A1(n4712), .A2(n8142), .ZN(n8149) );
  NAND2_X1 U5594 ( .A1(n8138), .A2(n6617), .ZN(n4712) );
  NAND2_X1 U5595 ( .A1(n4710), .A2(n8199), .ZN(n4709) );
  NAND2_X1 U5596 ( .A1(n8149), .A2(n4711), .ZN(n4710) );
  AND2_X1 U5597 ( .A1(n8154), .A2(n8151), .ZN(n4711) );
  NAND2_X1 U5598 ( .A1(n8143), .A2(n8182), .ZN(n4708) );
  OR2_X1 U5599 ( .A1(n8836), .A2(n4581), .ZN(n4693) );
  OAI21_X1 U5600 ( .B1(n4700), .B2(n4694), .A(n4692), .ZN(n4691) );
  NOR3_X1 U5601 ( .A1(n8869), .A2(n4506), .A3(n4706), .ZN(n4705) );
  INV_X1 U5602 ( .A(n8954), .ZN(n4706) );
  AOI21_X1 U5603 ( .B1(n4704), .B2(n4703), .A(n4707), .ZN(n4702) );
  NAND2_X1 U5604 ( .A1(n8867), .A2(n8868), .ZN(n4707) );
  NOR2_X1 U5605 ( .A1(n4506), .A2(n4553), .ZN(n4704) );
  INV_X1 U5606 ( .A(n8869), .ZN(n4703) );
  AOI21_X1 U5607 ( .B1(n4727), .B2(n4733), .A(n4567), .ZN(n4726) );
  AND2_X1 U5608 ( .A1(n4729), .A2(n5013), .ZN(n4727) );
  INV_X1 U5609 ( .A(n5183), .ZN(n8815) );
  AND2_X1 U5610 ( .A1(n8814), .A2(n7388), .ZN(n8810) );
  NAND2_X1 U5611 ( .A1(n8809), .A2(n8824), .ZN(n5183) );
  INV_X1 U5612 ( .A(n5156), .ZN(n4858) );
  NAND2_X1 U5613 ( .A1(n4723), .A2(n4724), .ZN(n4720) );
  NOR2_X1 U5614 ( .A1(n8192), .A2(n8191), .ZN(n8198) );
  INV_X1 U5615 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4999) );
  NAND2_X1 U5616 ( .A1(n7792), .A2(n5037), .ZN(n5036) );
  NOR2_X1 U5617 ( .A1(n5038), .A2(n4618), .ZN(n4617) );
  INV_X1 U5618 ( .A(n7756), .ZN(n4618) );
  INV_X1 U5619 ( .A(n5911), .ZN(n5052) );
  NAND2_X1 U5620 ( .A1(n7289), .A2(n7288), .ZN(n5044) );
  NOR2_X1 U5621 ( .A1(n5042), .A2(n5043), .ZN(n5041) );
  INV_X1 U5622 ( .A(n5043), .ZN(n5040) );
  NOR2_X1 U5623 ( .A1(n9179), .A2(n4994), .ZN(n4993) );
  NAND2_X1 U5624 ( .A1(n4996), .A2(n4995), .ZN(n4994) );
  INV_X1 U5625 ( .A(n9193), .ZN(n4995) );
  NOR2_X1 U5626 ( .A1(n9214), .A2(n9011), .ZN(n4996) );
  INV_X1 U5627 ( .A(n9276), .ZN(n8970) );
  AND2_X1 U5628 ( .A1(n7469), .A2(n9611), .ZN(n8830) );
  NAND2_X1 U5629 ( .A1(n5645), .A2(n5644), .ZN(n7853) );
  OAI21_X1 U5630 ( .B1(n5003), .B2(n5002), .A(n5001), .ZN(n5091) );
  NOR2_X1 U5631 ( .A1(n6067), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4751) );
  INV_X1 U5632 ( .A(n7230), .ZN(n4946) );
  AND2_X1 U5633 ( .A1(n4912), .A2(n9866), .ZN(n9842) );
  NAND2_X1 U5634 ( .A1(n4913), .A2(n9847), .ZN(n4912) );
  INV_X1 U5635 ( .A(n6850), .ZN(n4913) );
  OAI21_X1 U5636 ( .B1(n7030), .B2(n7032), .A(n4562), .ZN(n7428) );
  OR2_X1 U5637 ( .A1(n7029), .A2(n7032), .ZN(n4927) );
  NOR2_X1 U5638 ( .A1(n7480), .A2(n7604), .ZN(n4911) );
  AND2_X1 U5639 ( .A1(n7612), .A2(n7613), .ZN(n4641) );
  NOR2_X1 U5640 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6026) );
  INV_X1 U5641 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6024) );
  INV_X1 U5642 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6025) );
  INV_X1 U5643 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6238) );
  INV_X1 U5644 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6280) );
  AND2_X1 U5645 ( .A1(n6022), .A2(n6158), .ZN(n6023) );
  INV_X1 U5646 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U5647 ( .A1(n6065), .A2(n6064), .ZN(n6077) );
  NOR2_X1 U5648 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(n6401), .ZN(n4605) );
  INV_X1 U5649 ( .A(n8428), .ZN(n6619) );
  NAND4_X1 U5650 ( .A1(n6547), .A2(n6544), .A3(n6545), .A4(n6546), .ZN(n6550)
         );
  NOR2_X1 U5651 ( .A1(n6584), .A2(n4897), .ZN(n4896) );
  INV_X1 U5652 ( .A(n4899), .ZN(n4897) );
  INV_X1 U5653 ( .A(n4867), .ZN(n4866) );
  NOR2_X1 U5654 ( .A1(n6733), .A2(n6488), .ZN(n6658) );
  INV_X1 U5655 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6338) );
  NOR2_X1 U5656 ( .A1(n6236), .A2(n6235), .ZN(n6239) );
  OR2_X1 U5657 ( .A1(n6178), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6206) );
  NOR2_X1 U5658 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n6021) );
  AND2_X1 U5659 ( .A1(n5884), .A2(n4649), .ZN(n4648) );
  NAND2_X1 U5660 ( .A1(n7792), .A2(n5037), .ZN(n4649) );
  NAND2_X1 U5661 ( .A1(n7578), .A2(n5845), .ZN(n5850) );
  NAND2_X1 U5662 ( .A1(n8713), .A2(n5911), .ZN(n8677) );
  XNOR2_X1 U5663 ( .A(n4762), .B(n5988), .ZN(n5819) );
  NOR2_X1 U5664 ( .A1(n4537), .A2(n4763), .ZN(n4762) );
  NOR2_X1 U5665 ( .A1(n7293), .A2(n5967), .ZN(n4763) );
  NAND2_X1 U5666 ( .A1(n4688), .A2(n4684), .ZN(n4683) );
  INV_X1 U5667 ( .A(n8984), .ZN(n4684) );
  AOI21_X1 U5668 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n7084), .A(n9570), .ZN(
        n9494) );
  INV_X1 U5669 ( .A(n8882), .ZN(n8962) );
  NOR2_X1 U5670 ( .A1(n9152), .A2(n4670), .ZN(n4669) );
  INV_X1 U5671 ( .A(n4671), .ZN(n4670) );
  NOR2_X1 U5672 ( .A1(n9352), .A2(n9362), .ZN(n4671) );
  OR2_X1 U5673 ( .A1(n9152), .A2(n9349), .ZN(n8961) );
  NAND2_X1 U5674 ( .A1(n8868), .A2(n8936), .ZN(n4880) );
  AND2_X1 U5675 ( .A1(n5535), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5553) );
  AND2_X1 U5676 ( .A1(n8866), .A2(n8936), .ZN(n9010) );
  INV_X1 U5677 ( .A(n5518), .ZN(n5519) );
  AND2_X1 U5678 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(n5519), .ZN(n5535) );
  AND2_X1 U5679 ( .A1(n4520), .A2(n9273), .ZN(n4656) );
  NOR2_X1 U5680 ( .A1(n9421), .A2(n9426), .ZN(n4658) );
  NAND2_X1 U5681 ( .A1(n8993), .A2(n8820), .ZN(n4832) );
  AND2_X1 U5682 ( .A1(n8998), .A2(n8823), .ZN(n4830) );
  AND2_X1 U5683 ( .A1(n8826), .A2(n8827), .ZN(n8998) );
  NAND2_X1 U5684 ( .A1(n4662), .A2(n4660), .ZN(n7363) );
  AND2_X1 U5685 ( .A1(n4664), .A2(n4661), .ZN(n4660) );
  NOR2_X1 U5686 ( .A1(n4663), .A2(n9740), .ZN(n4661) );
  NAND2_X1 U5687 ( .A1(n9723), .A2(n4794), .ZN(n4663) );
  AND2_X1 U5688 ( .A1(n9050), .A2(n9698), .ZN(n5677) );
  NOR2_X1 U5689 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4821) );
  NAND2_X1 U5690 ( .A1(n4967), .A2(n4965), .ZN(n5609) );
  AOI21_X1 U5691 ( .B1(n4969), .B2(n4971), .A(n4966), .ZN(n4965) );
  INV_X1 U5692 ( .A(n5593), .ZN(n4966) );
  AND2_X1 U5693 ( .A1(n5628), .A2(n5597), .ZN(n5608) );
  AND2_X1 U5694 ( .A1(n5593), .A2(n5580), .ZN(n5591) );
  INV_X1 U5695 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5711) );
  OR2_X1 U5696 ( .A1(n5082), .A2(n9452), .ZN(n4760) );
  INV_X1 U5697 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5656) );
  INV_X1 U5698 ( .A(n4982), .ZN(n4974) );
  NAND2_X1 U5699 ( .A1(n5304), .A2(SI_10_), .ZN(n5325) );
  NAND2_X1 U5700 ( .A1(n6400), .A2(n7966), .ZN(n4943) );
  AND2_X1 U5701 ( .A1(n7985), .A2(n6437), .ZN(n7921) );
  AND2_X1 U5702 ( .A1(n7920), .A2(n6422), .ZN(n7946) );
  INV_X1 U5703 ( .A(n6205), .ZN(n4949) );
  NAND2_X1 U5704 ( .A1(n7231), .A2(n7230), .ZN(n4950) );
  NAND2_X1 U5705 ( .A1(n7652), .A2(n8223), .ZN(n4954) );
  AND2_X1 U5706 ( .A1(n6232), .A2(n6251), .ZN(n4939) );
  NAND2_X1 U5707 ( .A1(n7453), .A2(n7454), .ZN(n4940) );
  NAND2_X1 U5708 ( .A1(n6351), .A2(n7973), .ZN(n7976) );
  INV_X1 U5709 ( .A(n4597), .ZN(n4596) );
  OAI21_X1 U5710 ( .B1(n8556), .B2(n8212), .A(n8210), .ZN(n4597) );
  INV_X1 U5711 ( .A(n8201), .ZN(n4740) );
  NAND2_X1 U5712 ( .A1(n6046), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6490) );
  OR2_X1 U5713 ( .A1(n7352), .A2(n6829), .ZN(n6155) );
  OR2_X1 U5714 ( .A1(n6854), .A2(n6853), .ZN(n6855) );
  OR2_X1 U5715 ( .A1(n9876), .A2(n9877), .ZN(n4631) );
  NAND2_X1 U5716 ( .A1(n7327), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7431) );
  AND2_X1 U5717 ( .A1(n7431), .A2(n7430), .ZN(n7432) );
  NOR2_X1 U5718 ( .A1(n7611), .A2(n4641), .ZN(n8260) );
  NAND2_X1 U5719 ( .A1(n4637), .A2(n4636), .ZN(n9919) );
  AOI21_X1 U5720 ( .B1(n4527), .B2(n4639), .A(n4593), .ZN(n4636) );
  NOR2_X1 U5721 ( .A1(n8238), .A2(n9907), .ZN(n9925) );
  INV_X1 U5722 ( .A(n4924), .ZN(n8237) );
  AND2_X1 U5723 ( .A1(n4918), .A2(n4539), .ZN(n9958) );
  OR2_X1 U5724 ( .A1(n6501), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7822) );
  INV_X1 U5725 ( .A(n4605), .ZN(n6412) );
  NAND2_X1 U5726 ( .A1(n4608), .A2(n6376), .ZN(n6386) );
  INV_X1 U5727 ( .A(n4608), .ZN(n6377) );
  NAND2_X1 U5728 ( .A1(n6357), .A2(n6356), .ZN(n6367) );
  INV_X1 U5729 ( .A(n6358), .ZN(n6357) );
  OR2_X1 U5730 ( .A1(n8443), .A2(n8423), .ZN(n5072) );
  INV_X1 U5731 ( .A(n6330), .ZN(n6329) );
  INV_X1 U5732 ( .A(n4607), .ZN(n6301) );
  NAND2_X1 U5733 ( .A1(n6269), .A2(n6268), .ZN(n6287) );
  INV_X1 U5734 ( .A(n8467), .ZN(n8497) );
  NAND2_X1 U5735 ( .A1(n4606), .A2(n7619), .ZN(n6270) );
  INV_X1 U5736 ( .A(n4606), .ZN(n6253) );
  INV_X1 U5737 ( .A(n8223), .ZN(n8496) );
  INV_X1 U5738 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6210) );
  INV_X1 U5739 ( .A(n6212), .ZN(n6211) );
  OR2_X1 U5740 ( .A1(n6219), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U5741 ( .A1(n6561), .A2(n6560), .ZN(n7371) );
  NOR2_X1 U5742 ( .A1(n4555), .A2(n4888), .ZN(n4887) );
  NAND2_X1 U5743 ( .A1(n6184), .A2(n6183), .ZN(n6198) );
  INV_X1 U5744 ( .A(n6185), .ZN(n6184) );
  NAND2_X1 U5745 ( .A1(n4889), .A2(n4890), .ZN(n7277) );
  OR2_X1 U5746 ( .A1(n6163), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U5747 ( .A1(n6149), .A2(n6148), .ZN(n6163) );
  INV_X1 U5748 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6148) );
  INV_X1 U5749 ( .A(n6150), .ZN(n6149) );
  NAND2_X1 U5750 ( .A1(n7201), .A2(n8076), .ZN(n7106) );
  INV_X1 U5751 ( .A(n4840), .ZN(n4835) );
  AND4_X1 U5752 ( .A1(n6547), .A2(n6545), .A3(n6546), .A4(n6544), .ZN(n9996)
         );
  NOR2_X1 U5753 ( .A1(n7187), .A2(n6932), .ZN(n7179) );
  NAND2_X1 U5754 ( .A1(n6590), .A2(n6589), .ZN(n6654) );
  OR2_X1 U5755 ( .A1(n8184), .A2(n8054), .ZN(n5023) );
  INV_X1 U5756 ( .A(n5020), .ZN(n5019) );
  OAI21_X1 U5757 ( .B1(n8184), .B2(n5021), .A(n8020), .ZN(n5020) );
  AND2_X1 U5758 ( .A1(n6625), .A2(n8179), .ZN(n8352) );
  NAND2_X1 U5759 ( .A1(n6409), .A2(n6408), .ZN(n6623) );
  NAND2_X1 U5760 ( .A1(n4843), .A2(n4842), .ZN(n8379) );
  AOI21_X1 U5761 ( .B1(n4844), .B2(n4512), .A(n8167), .ZN(n4842) );
  NOR2_X1 U5762 ( .A1(n4847), .A2(n8377), .ZN(n4844) );
  NAND2_X1 U5763 ( .A1(n4845), .A2(n4846), .ZN(n8390) );
  OR2_X1 U5764 ( .A1(n8414), .A2(n4512), .ZN(n4845) );
  NOR2_X1 U5765 ( .A1(n8155), .A2(n5005), .ZN(n5004) );
  INV_X1 U5766 ( .A(n8058), .ZN(n5005) );
  NAND2_X1 U5767 ( .A1(n8412), .A2(n8413), .ZN(n6621) );
  AOI21_X1 U5768 ( .B1(n5033), .B2(n5031), .A(n5030), .ZN(n5029) );
  INV_X1 U5769 ( .A(n5033), .ZN(n5032) );
  INV_X1 U5770 ( .A(n6614), .ZN(n5031) );
  AND2_X1 U5771 ( .A1(n6467), .A2(n6466), .ZN(n6477) );
  INV_X1 U5772 ( .A(n6477), .ZN(n6733) );
  NOR2_X1 U5773 ( .A1(n5027), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U5774 ( .A1(n6064), .A2(n5028), .ZN(n5027) );
  INV_X1 U5775 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U5776 ( .A1(n4563), .A2(n5065), .ZN(n5064) );
  OR2_X1 U5777 ( .A1(n8696), .A2(n5963), .ZN(n5065) );
  NAND2_X1 U5778 ( .A1(n5792), .A2(n9683), .ZN(n5768) );
  NAND2_X1 U5779 ( .A1(n5933), .A2(n5083), .ZN(n5939) );
  INV_X1 U5780 ( .A(n5583), .ZN(n5584) );
  INV_X1 U5781 ( .A(n8696), .ZN(n5066) );
  INV_X1 U5782 ( .A(n4610), .ZN(n4609) );
  INV_X1 U5783 ( .A(n5809), .ZN(n4611) );
  NAND2_X1 U5784 ( .A1(n8703), .A2(n5903), .ZN(n8714) );
  NAND2_X1 U5785 ( .A1(n8714), .A2(n8715), .ZN(n8713) );
  AND2_X1 U5786 ( .A1(n5553), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5569) );
  OR2_X1 U5787 ( .A1(n5178), .A2(n5161), .ZN(n5163) );
  NOR2_X1 U5788 ( .A1(n5163), .A2(n7581), .ZN(n5319) );
  AND2_X1 U5789 ( .A1(n5789), .A2(n5791), .ZN(n6897) );
  NOR2_X1 U5790 ( .A1(n5447), .A2(n7780), .ZN(n5462) );
  NAND2_X2 U5791 ( .A1(n4531), .A2(n5815), .ZN(n7160) );
  INV_X1 U5792 ( .A(n5814), .ZN(n5815) );
  NAND2_X1 U5793 ( .A1(n7159), .A2(n7161), .ZN(n5816) );
  INV_X1 U5794 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5184) );
  INV_X1 U5795 ( .A(n5891), .ZN(n4621) );
  NOR2_X1 U5796 ( .A1(n5392), .A2(n7316), .ZN(n5410) );
  NAND2_X1 U5797 ( .A1(n4990), .A2(n4989), .ZN(n4988) );
  OR2_X1 U5798 ( .A1(n9022), .A2(n9021), .ZN(n4990) );
  AOI21_X1 U5799 ( .B1(n7084), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9574), .ZN(
        n9498) );
  AOI21_X1 U5800 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7090), .A(n9513), .ZN(
        n9105) );
  AOI21_X1 U5801 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9489), .A(n9484), .ZN(
        n9587) );
  AOI21_X1 U5802 ( .B1(n9489), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9481), .ZN(
        n9592) );
  NOR2_X1 U5803 ( .A1(n7718), .A2(n7719), .ZN(n7720) );
  NAND2_X1 U5804 ( .A1(n7720), .A2(n7721), .ZN(n7775) );
  NAND2_X1 U5805 ( .A1(n8887), .A2(n8886), .ZN(n8979) );
  AND2_X1 U5806 ( .A1(n9180), .A2(n4667), .ZN(n9132) );
  AND2_X1 U5807 ( .A1(n4669), .A2(n9142), .ZN(n4667) );
  AND2_X1 U5809 ( .A1(n8962), .A2(n8900), .ZN(n8984) );
  NAND2_X1 U5810 ( .A1(n9180), .A2(n4669), .ZN(n9150) );
  AND2_X1 U5811 ( .A1(n5649), .A2(n5621), .ZN(n9168) );
  OAI21_X1 U5812 ( .B1(n9162), .B2(n5626), .A(n4997), .ZN(n9165) );
  NAND2_X1 U5813 ( .A1(n5695), .A2(n5694), .ZN(n9178) );
  NAND2_X1 U5814 ( .A1(n4795), .A2(n4524), .ZN(n5695) );
  NOR2_X1 U5815 ( .A1(n9206), .A2(n9370), .ZN(n9180) );
  NOR2_X1 U5816 ( .A1(n9193), .A2(n5589), .ZN(n4878) );
  AND4_X1 U5817 ( .A1(n5558), .A2(n5557), .A3(n5556), .A4(n5555), .ZN(n9216)
         );
  NOR2_X1 U5818 ( .A1(n9384), .A2(n9241), .ZN(n9226) );
  INV_X1 U5819 ( .A(n9010), .ZN(n9224) );
  NAND2_X1 U5820 ( .A1(n9240), .A2(n9392), .ZN(n9241) );
  OR2_X1 U5821 ( .A1(n9406), .A2(n9398), .ZN(n5689) );
  NOR2_X1 U5822 ( .A1(n9273), .A2(n9288), .ZN(n5690) );
  NOR2_X1 U5823 ( .A1(n5488), .A2(n7885), .ZN(n5504) );
  AND2_X1 U5824 ( .A1(n8844), .A2(n8902), .ZN(n9286) );
  NAND2_X1 U5825 ( .A1(n4804), .A2(n4803), .ZN(n9284) );
  AOI21_X1 U5826 ( .B1(n4515), .B2(n4504), .A(n4558), .ZN(n4803) );
  NAND2_X1 U5827 ( .A1(n7812), .A2(n4658), .ZN(n9303) );
  NOR3_X1 U5828 ( .A1(n9326), .A2(n5467), .A3(n9302), .ZN(n9300) );
  OR2_X1 U5829 ( .A1(n7798), .A2(n4885), .ZN(n4883) );
  NAND2_X1 U5830 ( .A1(n8929), .A2(n8849), .ZN(n4885) );
  NAND2_X1 U5831 ( .A1(n8929), .A2(n9004), .ZN(n4884) );
  AND2_X2 U5832 ( .A1(n4883), .A2(n4881), .ZN(n9326) );
  NOR2_X1 U5833 ( .A1(n9327), .A2(n4882), .ZN(n4881) );
  INV_X1 U5834 ( .A(n4884), .ZN(n4882) );
  NAND2_X1 U5835 ( .A1(n7812), .A2(n9325), .ZN(n9319) );
  NOR2_X1 U5836 ( .A1(n7798), .A2(n5431), .ZN(n7815) );
  NAND2_X1 U5837 ( .A1(n9637), .A2(n4665), .ZN(n7813) );
  AND2_X1 U5838 ( .A1(n4507), .A2(n9532), .ZN(n4665) );
  NOR2_X1 U5839 ( .A1(n7799), .A2(n9002), .ZN(n7798) );
  NAND2_X1 U5840 ( .A1(n4526), .A2(n4817), .ZN(n4811) );
  NAND2_X1 U5841 ( .A1(n9637), .A2(n4666), .ZN(n9620) );
  OR2_X1 U5842 ( .A1(n5377), .A2(n7250), .ZN(n5392) );
  OR2_X1 U5843 ( .A1(n5357), .A2(n5356), .ZN(n5377) );
  NAND2_X1 U5844 ( .A1(n9637), .A2(n4820), .ZN(n9619) );
  NAND2_X1 U5845 ( .A1(n7358), .A2(n8820), .ZN(n9628) );
  NAND2_X1 U5846 ( .A1(n5331), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U5847 ( .A1(n4833), .A2(n7361), .ZN(n7358) );
  NAND2_X1 U5848 ( .A1(n4779), .A2(n4778), .ZN(n7362) );
  NAND2_X1 U5849 ( .A1(n4786), .A2(n4523), .ZN(n4778) );
  NAND2_X1 U5850 ( .A1(n4775), .A2(n4772), .ZN(n4779) );
  NAND2_X1 U5851 ( .A1(n4662), .A2(n4661), .ZN(n7383) );
  NOR2_X1 U5852 ( .A1(n9654), .A2(n4663), .ZN(n7404) );
  NOR2_X1 U5853 ( .A1(n9654), .A2(n9653), .ZN(n9655) );
  NOR2_X1 U5854 ( .A1(n5280), .A2(n5184), .ZN(n5186) );
  NAND2_X1 U5855 ( .A1(n5281), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U5856 ( .A1(n5296), .A2(n5295), .ZN(n7140) );
  NAND2_X1 U5857 ( .A1(n8803), .A2(n8913), .ZN(n8986) );
  AND2_X1 U5858 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5281) );
  NAND2_X1 U5859 ( .A1(n9674), .A2(n9698), .ZN(n9672) );
  NOR2_X1 U5860 ( .A1(n9672), .A2(n6988), .ZN(n7143) );
  AOI21_X1 U5861 ( .B1(n9671), .B2(n9670), .A(n5679), .ZN(n6984) );
  NAND2_X1 U5862 ( .A1(n5678), .A2(n8908), .ZN(n9670) );
  AND3_X1 U5863 ( .A1(n9691), .A2(n8905), .A3(n6889), .ZN(n9674) );
  OAI21_X1 U5864 ( .B1(n6872), .B2(n6873), .A(n5673), .ZN(n6888) );
  NAND2_X1 U5865 ( .A1(n5674), .A2(n8903), .ZN(n8987) );
  NAND2_X1 U5866 ( .A1(n6872), .A2(n6876), .ZN(n6875) );
  NOR2_X1 U5867 ( .A1(n6712), .A2(n6889), .ZN(n6876) );
  AND4_X1 U5868 ( .A1(n5573), .A2(n5572), .A3(n5571), .A4(n5570), .ZN(n9380)
         );
  AOI21_X1 U5869 ( .B1(n9643), .B2(n4561), .A(n4792), .ZN(n7395) );
  AND2_X1 U5870 ( .A1(n5294), .A2(n5293), .ZN(n9713) );
  AND3_X1 U5871 ( .A1(n5279), .A2(n5278), .A3(n5277), .ZN(n9705) );
  INV_X1 U5872 ( .A(n9784), .ZN(n9772) );
  XNOR2_X1 U5873 ( .A(n5641), .B(n5640), .ZN(n7808) );
  XNOR2_X1 U5874 ( .A(n5138), .B(n5137), .ZN(n5669) );
  NAND2_X1 U5875 ( .A1(n5136), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5138) );
  XNOR2_X1 U5876 ( .A(n5715), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5728) );
  XNOR2_X1 U5877 ( .A(n5609), .B(n5608), .ZN(n7766) );
  XNOR2_X1 U5878 ( .A(n5592), .B(n5591), .ZN(n7730) );
  NAND2_X1 U5879 ( .A1(n4968), .A2(n5576), .ZN(n5592) );
  NAND2_X1 U5880 ( .A1(n5575), .A2(n5574), .ZN(n4968) );
  NOR2_X1 U5881 ( .A1(n5720), .A2(n5719), .ZN(n5745) );
  NAND2_X1 U5882 ( .A1(n4963), .A2(n5526), .ZN(n5545) );
  OAI21_X1 U5883 ( .B1(n5500), .B2(n5499), .A(n5498), .ZN(n5511) );
  OR2_X1 U5884 ( .A1(n5493), .A2(n5495), .ZN(n5499) );
  AND2_X1 U5885 ( .A1(n5497), .A2(n5496), .ZN(n5498) );
  OR2_X1 U5886 ( .A1(n5495), .A2(n5494), .ZN(n5497) );
  XNOR2_X1 U5887 ( .A(n5481), .B(n5495), .ZN(n7304) );
  AND2_X1 U5888 ( .A1(n5476), .A2(n5494), .ZN(n5481) );
  XNOR2_X1 U5889 ( .A(n5455), .B(n5473), .ZN(n7285) );
  INV_X1 U5890 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4654) );
  AND2_X1 U5891 ( .A1(n5383), .A2(n5368), .ZN(n5369) );
  NOR2_X1 U5892 ( .A1(n5300), .A2(SI_9_), .ZN(n5301) );
  OAI21_X1 U5893 ( .B1(n5194), .B2(n4862), .A(n4859), .ZN(n5157) );
  AND2_X1 U5894 ( .A1(n5174), .A2(n5173), .ZN(n7087) );
  INV_X1 U5895 ( .A(n5264), .ZN(n5108) );
  AND2_X1 U5896 ( .A1(n5113), .A2(n5112), .ZN(n5289) );
  NAND2_X1 U5897 ( .A1(n7151), .A2(n7150), .ZN(n7149) );
  NAND2_X1 U5898 ( .A1(n6278), .A2(n6277), .ZN(n7890) );
  NAND2_X1 U5899 ( .A1(n4953), .A2(n4951), .ZN(n6278) );
  NAND2_X1 U5900 ( .A1(n7976), .A2(n6353), .ZN(n7903) );
  AND2_X1 U5901 ( .A1(n6419), .A2(n6418), .ZN(n8347) );
  NAND2_X1 U5902 ( .A1(n7931), .A2(n7930), .ZN(n7929) );
  NAND2_X1 U5903 ( .A1(n7929), .A2(n6322), .ZN(n7938) );
  NAND2_X1 U5904 ( .A1(n4950), .A2(n6205), .ZN(n7410) );
  NAND2_X1 U5905 ( .A1(n4931), .A2(n4930), .ZN(n7954) );
  AOI21_X1 U5906 ( .B1(n4513), .B2(n4933), .A(n4545), .ZN(n4930) );
  NAND2_X1 U5907 ( .A1(n4953), .A2(n4954), .ZN(n7735) );
  NAND2_X1 U5908 ( .A1(n4940), .A2(n6232), .ZN(n7665) );
  INV_X1 U5909 ( .A(n7981), .ZN(n8006) );
  XNOR2_X1 U5910 ( .A(n6490), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8218) );
  AND2_X1 U5911 ( .A1(n7355), .A2(n7354), .ZN(n8287) );
  INV_X1 U5912 ( .A(n8332), .ZN(n8360) );
  INV_X1 U5913 ( .A(n8347), .ZN(n8369) );
  INV_X1 U5914 ( .A(n7960), .ZN(n8395) );
  OR2_X1 U5915 ( .A1(n6797), .A2(n9832), .ZN(n4635) );
  NOR2_X1 U5916 ( .A1(n7014), .A2(n4622), .ZN(n7020) );
  AND2_X1 U5917 ( .A1(n7015), .A2(n7016), .ZN(n4622) );
  INV_X1 U5918 ( .A(n7334), .ZN(n7333) );
  NOR2_X1 U5919 ( .A1(n7033), .A2(n7032), .ZN(n7325) );
  AND2_X1 U5920 ( .A1(n7030), .A2(n7029), .ZN(n7033) );
  AND2_X1 U5921 ( .A1(n4638), .A2(n4640), .ZN(n9903) );
  NAND2_X1 U5922 ( .A1(n4638), .A2(n4527), .ZN(n9902) );
  OR2_X1 U5923 ( .A1(n7611), .A2(n4639), .ZN(n4638) );
  INV_X1 U5924 ( .A(n4918), .ZN(n9939) );
  NAND2_X1 U5925 ( .A1(n6770), .A2(n6769), .ZN(n9964) );
  INV_X1 U5926 ( .A(n4922), .ZN(n9976) );
  AND2_X1 U5927 ( .A1(n4922), .A2(n4535), .ZN(n9474) );
  NAND2_X1 U5928 ( .A1(n8019), .A2(n8018), .ZN(n8284) );
  NAND2_X1 U5929 ( .A1(n5006), .A2(n6643), .ZN(n7821) );
  NAND2_X1 U5930 ( .A1(n6456), .A2(n6442), .ZN(n8339) );
  NAND2_X1 U5931 ( .A1(n8440), .A2(n8139), .ZN(n8427) );
  NAND2_X1 U5932 ( .A1(n6243), .A2(n6242), .ZN(n10054) );
  NAND2_X1 U5933 ( .A1(n5017), .A2(n8104), .ZN(n7544) );
  NAND2_X1 U5934 ( .A1(n4836), .A2(n4840), .ZN(n7198) );
  NAND2_X1 U5935 ( .A1(n4839), .A2(n4837), .ZN(n4836) );
  AND2_X1 U5936 ( .A1(n7121), .A2(n9989), .ZN(n10005) );
  OR2_X1 U5937 ( .A1(n7121), .A2(n9987), .ZN(n8442) );
  OR2_X1 U5938 ( .A1(n6718), .A2(n6663), .ZN(n9989) );
  INV_X1 U5939 ( .A(n8442), .ZN(n8473) );
  INV_X1 U5940 ( .A(n8284), .ZN(n8556) );
  NAND2_X1 U5941 ( .A1(n8050), .A2(n8049), .ZN(n8557) );
  NAND2_X1 U5942 ( .A1(n4566), .A2(n5006), .ZN(n6668) );
  INV_X1 U5943 ( .A(n6654), .ZN(n7823) );
  OAI21_X1 U5944 ( .B1(n8300), .B2(n10000), .A(n8299), .ZN(n8560) );
  NAND2_X1 U5945 ( .A1(n5018), .A2(n8021), .ZN(n8308) );
  NAND2_X1 U5946 ( .A1(n6626), .A2(n5024), .ZN(n5018) );
  INV_X1 U5947 ( .A(n8340), .ZN(n8571) );
  XNOR2_X1 U5948 ( .A(n8331), .B(n4722), .ZN(n8336) );
  OAI22_X1 U5949 ( .A1(n8333), .A2(n9993), .B1(n9995), .B2(n8332), .ZN(n8334)
         );
  NAND2_X1 U5950 ( .A1(n6626), .A2(n6625), .ZN(n8328) );
  INV_X1 U5951 ( .A(n8172), .ZN(n8576) );
  NAND2_X1 U5952 ( .A1(n5010), .A2(n5011), .ZN(n8357) );
  NAND2_X1 U5953 ( .A1(n8375), .A2(n8056), .ZN(n5014) );
  AND2_X1 U5954 ( .A1(n4853), .A2(n4854), .ZN(n8404) );
  INV_X1 U5955 ( .A(n6618), .ZN(n8621) );
  NAND2_X1 U5956 ( .A1(n6313), .A2(n6312), .ZN(n8625) );
  AND2_X1 U5957 ( .A1(n8456), .A2(n8455), .ZN(n8623) );
  NAND2_X1 U5958 ( .A1(n6299), .A2(n6298), .ZN(n8631) );
  NAND2_X1 U5959 ( .A1(n4864), .A2(n4867), .ZN(n8466) );
  NAND2_X1 U5960 ( .A1(n8494), .A2(n4868), .ZN(n4864) );
  NAND2_X1 U5961 ( .A1(n6286), .A2(n6285), .ZN(n8637) );
  AOI21_X1 U5962 ( .B1(n8494), .B2(n8500), .A(n4508), .ZN(n8478) );
  INV_X1 U5963 ( .A(n8620), .ZN(n8638) );
  AND2_X1 U5964 ( .A1(n6673), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6737) );
  XNOR2_X1 U5965 ( .A(n6043), .B(n6064), .ZN(n7767) );
  XNOR2_X1 U5966 ( .A(n6465), .B(n6464), .ZN(n7732) );
  INV_X1 U5967 ( .A(n8218), .ZN(n7540) );
  NAND2_X1 U5968 ( .A1(n6058), .A2(n4957), .ZN(n6044) );
  INV_X1 U5969 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7305) );
  INV_X1 U5970 ( .A(n4915), .ZN(n4914) );
  OAI21_X1 U5971 ( .B1(n6070), .B2(n4917), .A(n4916), .ZN(n4915) );
  NAND2_X1 U5972 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4917) );
  NAND2_X1 U5973 ( .A1(n6072), .A2(n6071), .ZN(n6805) );
  INV_X1 U5974 ( .A(n4768), .ZN(n8668) );
  NAND2_X1 U5975 ( .A1(n5035), .A2(n7698), .ZN(n7639) );
  AND4_X1 U5976 ( .A1(n5182), .A2(n5181), .A3(n5180), .A4(n5179), .ZN(n9729)
         );
  NAND2_X1 U5977 ( .A1(n5939), .A2(n5938), .ZN(n8689) );
  NAND2_X1 U5978 ( .A1(n4765), .A2(n4764), .ZN(n8697) );
  AOI21_X1 U5979 ( .B1(n8743), .B2(n4519), .A(n4557), .ZN(n4764) );
  AND3_X1 U5980 ( .A1(n5466), .A2(n5465), .A3(n5464), .ZN(n9330) );
  INV_X1 U5981 ( .A(n4769), .ZN(n4646) );
  AOI21_X1 U5982 ( .B1(n8668), .B2(n8666), .A(n4771), .ZN(n8724) );
  XNOR2_X1 U5983 ( .A(n5806), .B(n5807), .ZN(n6965) );
  AND4_X1 U5984 ( .A1(n5324), .A2(n5323), .A3(n5322), .A4(n5321), .ZN(n7704)
         );
  AND4_X1 U5985 ( .A1(n5524), .A2(n5523), .A3(n5522), .A4(n5521), .ZN(n9277)
         );
  NAND2_X1 U5986 ( .A1(n7791), .A2(n7792), .ZN(n7790) );
  NAND2_X1 U5987 ( .A1(n7758), .A2(n5869), .ZN(n7791) );
  INV_X1 U5988 ( .A(n9044), .ZN(n9418) );
  AND4_X1 U5989 ( .A1(n5492), .A2(n5491), .A3(n5490), .A4(n5489), .ZN(n9417)
         );
  AND2_X1 U5990 ( .A1(n6013), .A2(n7068), .ZN(n8767) );
  AND2_X1 U5991 ( .A1(n5620), .A2(n5603), .ZN(n9184) );
  AND4_X1 U5992 ( .A1(n5430), .A2(n5429), .A3(n5428), .A4(n5427), .ZN(n9329)
         );
  INV_X1 U5993 ( .A(n8767), .ZN(n8779) );
  NAND4_X1 U5994 ( .A1(n5261), .A2(n5260), .A3(n5259), .A4(n5258), .ZN(n9662)
         );
  OR2_X1 U5995 ( .A1(n5199), .A2(n5257), .ZN(n5261) );
  NAND2_X1 U5996 ( .A1(n4530), .A2(n5229), .ZN(n5779) );
  AND2_X1 U5997 ( .A1(n5228), .A2(n5227), .ZN(n5229) );
  NAND2_X1 U5998 ( .A1(n5226), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5203) );
  OR2_X1 U5999 ( .A1(n6679), .A2(n6678), .ZN(n9051) );
  AND2_X1 U6000 ( .A1(n5276), .A2(n5287), .ZN(n9549) );
  AOI21_X1 U6001 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7312), .A(n7311), .ZN(
        n7315) );
  AOI21_X1 U6002 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7312), .A(n7308), .ZN(
        n7310) );
  NOR2_X1 U6003 ( .A1(n7711), .A2(n7710), .ZN(n7714) );
  AOI21_X1 U6004 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n7776), .A(n7771), .ZN(
        n7772) );
  OAI21_X1 U6005 ( .B1(n9604), .B2(n7887), .A(n7886), .ZN(n4601) );
  AND2_X1 U6006 ( .A1(n8892), .A2(n8891), .ZN(n9338) );
  INV_X1 U6007 ( .A(n8979), .ZN(n9341) );
  OR2_X1 U6008 ( .A1(n9157), .A2(n9156), .ZN(n9342) );
  NAND2_X1 U6009 ( .A1(n4874), .A2(n4875), .ZN(n9177) );
  NAND2_X1 U6010 ( .A1(n4795), .A2(n4796), .ZN(n9194) );
  OAI21_X1 U6011 ( .B1(n9225), .B2(n4533), .A(n4801), .ZN(n9205) );
  AND4_X1 U6012 ( .A1(n5541), .A2(n5540), .A3(n5539), .A4(n5538), .ZN(n9381)
         );
  NAND2_X1 U6013 ( .A1(n4907), .A2(n4906), .ZN(n9253) );
  AND2_X1 U6014 ( .A1(n4907), .A2(n8863), .ZN(n9255) );
  INV_X1 U6015 ( .A(n9268), .ZN(n9269) );
  OR2_X1 U6016 ( .A1(n7811), .A2(n4504), .ZN(n4805) );
  AND2_X1 U6017 ( .A1(n4808), .A2(n4809), .ZN(n9318) );
  NAND2_X1 U6018 ( .A1(n7811), .A2(n9004), .ZN(n4808) );
  NAND2_X1 U6019 ( .A1(n9605), .A2(n9609), .ZN(n7691) );
  NAND2_X1 U6020 ( .A1(n4812), .A2(n4813), .ZN(n7687) );
  NAND2_X1 U6021 ( .A1(n7464), .A2(n4534), .ZN(n4812) );
  OR2_X1 U6022 ( .A1(n6781), .A2(n5209), .ZN(n5376) );
  OAI21_X1 U6023 ( .B1(n7464), .B2(n8999), .A(n4819), .ZN(n9618) );
  NAND2_X1 U6024 ( .A1(n5330), .A2(n5329), .ZN(n9636) );
  AND2_X1 U6025 ( .A1(n4777), .A2(n4776), .ZN(n7380) );
  OR2_X1 U6026 ( .A1(n4785), .A2(n4784), .ZN(n4777) );
  NAND2_X1 U6027 ( .A1(n4790), .A2(n4782), .ZN(n4776) );
  NAND2_X1 U6028 ( .A1(n6003), .A2(n9026), .ZN(n9664) );
  OR2_X1 U6029 ( .A1(n9634), .A2(n6791), .ZN(n9668) );
  NAND2_X1 U6030 ( .A1(n6945), .A2(n6887), .ZN(n9677) );
  OR2_X1 U6031 ( .A1(n6540), .A2(n6783), .ZN(n9823) );
  INV_X2 U6032 ( .A(n9823), .ZN(n9825) );
  AND2_X1 U6033 ( .A1(n6699), .A2(n9026), .ZN(n9681) );
  XNOR2_X1 U6034 ( .A(n5148), .B(n5147), .ZN(n7849) );
  NAND2_X1 U6035 ( .A1(n5146), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6036 ( .A1(n4655), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5135) );
  CLKBUF_X1 U6037 ( .A(n5669), .Z(n7867) );
  INV_X1 U6038 ( .A(n5728), .ZN(n7770) );
  AND2_X1 U6039 ( .A1(n5722), .A2(n4532), .ZN(n7751) );
  AND2_X1 U6040 ( .A1(n4958), .A2(n4961), .ZN(n5560) );
  INV_X1 U6041 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10379) );
  INV_X1 U6042 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7307) );
  INV_X1 U6043 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7104) );
  NAND2_X1 U6044 ( .A1(n4978), .A2(n4976), .ZN(n5364) );
  NAND2_X1 U6045 ( .A1(n4978), .A2(n4979), .ZN(n5342) );
  NAND2_X1 U6046 ( .A1(n5169), .A2(n5168), .ZN(n5171) );
  NAND2_X1 U6047 ( .A1(n5194), .A2(n5118), .ZN(n5169) );
  NAND2_X1 U6048 ( .A1(n7989), .A2(n4583), .ZN(n4936) );
  NAND2_X1 U6049 ( .A1(n6993), .A2(n6128), .ZN(n7002) );
  NAND2_X1 U6050 ( .A1(n4624), .A2(n4625), .ZN(n6833) );
  INV_X1 U6051 ( .A(n4926), .ZN(n8235) );
  OAI21_X1 U6052 ( .B1(n4644), .B2(n9875), .A(n4642), .ZN(n8280) );
  OAI211_X1 U6053 ( .C1(n6533), .C2(n5999), .A(n4651), .B(n6020), .ZN(P1_U3220) );
  NAND2_X1 U6054 ( .A1(n6533), .A2(n4652), .ZN(n4651) );
  OAI21_X1 U6055 ( .B1(n4675), .B2(n9032), .A(n4673), .ZN(n9040) );
  OAI211_X1 U6056 ( .C1(n7884), .C2(n5702), .A(n4600), .B(n4599), .ZN(P1_U3262) );
  INV_X1 U6057 ( .A(n4601), .ZN(n4600) );
  OR2_X1 U6058 ( .A1(n7883), .A2(n9021), .ZN(n4599) );
  NAND2_X1 U6059 ( .A1(n4825), .A2(n4592), .ZN(P1_U3550) );
  NAND2_X1 U6060 ( .A1(n9437), .A2(n9825), .ZN(n4825) );
  INV_X1 U6061 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n4824) );
  AND2_X1 U6062 ( .A1(n9238), .A2(n4541), .ZN(n4506) );
  AND2_X1 U6063 ( .A1(n4666), .A2(n8665), .ZN(n4507) );
  NOR2_X1 U6064 ( .A1(n8129), .A2(n8482), .ZN(n4508) );
  INV_X1 U6065 ( .A(n8229), .ZN(n4891) );
  INV_X1 U6066 ( .A(n4585), .ZN(n4771) );
  NOR2_X1 U6067 ( .A1(n4942), .A2(n4943), .ZN(n4509) );
  AND4_X2 U6068 ( .A1(n5128), .A2(n5127), .A3(n5344), .A4(n10274), .ZN(n4510)
         );
  INV_X1 U6069 ( .A(n5223), .ZN(n6726) );
  AND2_X1 U6070 ( .A1(n9431), .A2(n9045), .ZN(n5684) );
  AND2_X1 U6071 ( .A1(n8612), .A2(n8405), .ZN(n6572) );
  AND4_X1 U6072 ( .A1(n8876), .A2(n9174), .A3(n9183), .A4(n9031), .ZN(n4511)
         );
  NAND2_X1 U6073 ( .A1(n4647), .A2(n4551), .ZN(n4768) );
  OR2_X1 U6074 ( .A1(n4850), .A2(n8392), .ZN(n4512) );
  INV_X1 U6075 ( .A(n4733), .ZN(n4732) );
  AND2_X1 U6076 ( .A1(n7904), .A2(n4932), .ZN(n4513) );
  OR2_X1 U6077 ( .A1(n8179), .A2(n8199), .ZN(n4514) );
  AND2_X1 U6078 ( .A1(n4806), .A2(n4546), .ZN(n4515) );
  AND2_X1 U6079 ( .A1(n8806), .A2(n9031), .ZN(n4516) );
  INV_X1 U6080 ( .A(n9183), .ZN(n9359) );
  AND4_X1 U6081 ( .A1(n8207), .A2(n8052), .A3(n8195), .A4(n8212), .ZN(n4517)
         );
  AND2_X1 U6082 ( .A1(n4517), .A2(n6661), .ZN(n4518) );
  AND2_X1 U6083 ( .A1(n9191), .A2(n8939), .ZN(n8868) );
  AND2_X1 U6084 ( .A1(n4766), .A2(n8746), .ZN(n4519) );
  AND2_X1 U6085 ( .A1(n4658), .A2(n4657), .ZN(n4520) );
  AND2_X1 U6086 ( .A1(n6066), .A2(n8644), .ZN(n4521) );
  AND2_X1 U6087 ( .A1(n8631), .A2(n8480), .ZN(n4522) );
  AND2_X1 U6088 ( .A1(n4793), .A2(n4781), .ZN(n4523) );
  AND2_X1 U6089 ( .A1(n4796), .A2(n4552), .ZN(n4524) );
  NAND2_X1 U6090 ( .A1(n5160), .A2(n5159), .ZN(n9732) );
  INV_X1 U6091 ( .A(n9732), .ZN(n4794) );
  AND4_X1 U6092 ( .A1(n5190), .A2(n5189), .A3(n5188), .A4(n5187), .ZN(n7293)
         );
  NAND2_X1 U6093 ( .A1(n5036), .A2(n5883), .ZN(n4525) );
  INV_X1 U6094 ( .A(n8169), .ZN(n4731) );
  NAND2_X1 U6095 ( .A1(n4813), .A2(n4577), .ZN(n4526) );
  OR2_X1 U6096 ( .A1(n8594), .A2(n7960), .ZN(n8168) );
  AND2_X1 U6097 ( .A1(n5409), .A2(n5408), .ZN(n9532) );
  INV_X1 U6098 ( .A(n8022), .ZN(n5015) );
  INV_X1 U6099 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5137) );
  INV_X1 U6100 ( .A(n7469), .ZN(n4820) );
  AND2_X1 U6101 ( .A1(n4640), .A2(n9904), .ZN(n4527) );
  NAND2_X1 U6102 ( .A1(n5143), .A2(n5142), .ZN(n9740) );
  INV_X1 U6103 ( .A(n9740), .ZN(n4893) );
  AND2_X1 U6104 ( .A1(n8802), .A2(n8904), .ZN(n4528) );
  OR2_X1 U6105 ( .A1(n6077), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4529) );
  INV_X1 U6106 ( .A(n7792), .ZN(n5038) );
  AND2_X1 U6107 ( .A1(n5225), .A2(n5224), .ZN(n4530) );
  AND2_X1 U6108 ( .A1(n6964), .A2(n5809), .ZN(n4531) );
  NAND2_X1 U6109 ( .A1(n5218), .A2(n4672), .ZN(n6712) );
  NAND2_X1 U6110 ( .A1(n6143), .A2(n6023), .ZN(n6178) );
  XNOR2_X1 U6111 ( .A(n6884), .B(n5761), .ZN(n6872) );
  NAND2_X1 U6112 ( .A1(n4501), .A2(n5054), .ZN(n5718) );
  OR2_X1 U6113 ( .A1(n5055), .A2(n5420), .ZN(n4532) );
  NOR2_X1 U6114 ( .A1(n9384), .A2(n9388), .ZN(n4533) );
  AND2_X1 U6115 ( .A1(n8165), .A2(n8164), .ZN(n8392) );
  AND2_X1 U6116 ( .A1(n4818), .A2(n4819), .ZN(n4534) );
  XNOR2_X1 U6117 ( .A(n5712), .B(n5711), .ZN(n5704) );
  OR2_X1 U6118 ( .A1(n9965), .A2(n8240), .ZN(n4535) );
  AND2_X1 U6119 ( .A1(n8010), .A2(n6615), .ZN(n4536) );
  INV_X1 U6120 ( .A(n8232), .ZN(n4755) );
  INV_X1 U6121 ( .A(n5869), .ZN(n5037) );
  NAND2_X1 U6122 ( .A1(n5487), .A2(n5486), .ZN(n9413) );
  INV_X1 U6123 ( .A(n9413), .ZN(n4657) );
  NAND2_X1 U6124 ( .A1(n5391), .A2(n5390), .ZN(n9793) );
  AND2_X1 U6125 ( .A1(n7268), .A2(n5948), .ZN(n4537) );
  NAND2_X1 U6126 ( .A1(n5446), .A2(n5445), .ZN(n9426) );
  NAND2_X1 U6127 ( .A1(n5599), .A2(n5598), .ZN(n9362) );
  NAND2_X1 U6128 ( .A1(n5617), .A2(n5616), .ZN(n9352) );
  AND2_X1 U6129 ( .A1(n9426), .A2(n9044), .ZN(n4538) );
  OR2_X1 U6130 ( .A1(n9931), .A2(n8239), .ZN(n4539) );
  AND4_X1 U6131 ( .A1(n5155), .A2(n5154), .A3(n5153), .A4(n5152), .ZN(n9747)
         );
  INV_X1 U6132 ( .A(n9747), .ZN(n4892) );
  OR2_X1 U6133 ( .A1(n9406), .A2(n9288), .ZN(n8863) );
  OR2_X1 U6134 ( .A1(n8612), .A2(n8424), .ZN(n8154) );
  OR2_X1 U6135 ( .A1(n6623), .A2(n8369), .ZN(n4540) );
  NOR2_X1 U6136 ( .A1(n8865), .A2(n8899), .ZN(n4541) );
  AND2_X1 U6137 ( .A1(n5067), .A2(n5066), .ZN(n4542) );
  AND2_X1 U6138 ( .A1(n6218), .A2(n8226), .ZN(n4543) );
  AND2_X1 U6139 ( .A1(n8098), .A2(n8182), .ZN(n4544) );
  AND2_X1 U6140 ( .A1(n6364), .A2(n8424), .ZN(n4545) );
  OR2_X1 U6141 ( .A1(n9421), .A2(n9043), .ZN(n4546) );
  INV_X1 U6142 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9452) );
  AND2_X1 U6143 ( .A1(n6619), .A2(n8139), .ZN(n4547) );
  INV_X1 U6144 ( .A(n6584), .ZN(n4900) );
  INV_X1 U6145 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4759) );
  AND2_X1 U6146 ( .A1(n4944), .A2(n6128), .ZN(n4548) );
  AND2_X1 U6147 ( .A1(n5944), .A2(n5938), .ZN(n4549) );
  INV_X1 U6148 ( .A(n4902), .ZN(n4901) );
  AND2_X1 U6149 ( .A1(n8057), .A2(n8182), .ZN(n4550) );
  INV_X1 U6150 ( .A(n4847), .ZN(n4846) );
  NOR2_X1 U6151 ( .A1(n4848), .A2(n8392), .ZN(n4847) );
  NAND2_X1 U6152 ( .A1(n8743), .A2(n8746), .ZN(n4551) );
  NAND2_X1 U6153 ( .A1(n9145), .A2(n8974), .ZN(n9164) );
  INV_X1 U6154 ( .A(n9164), .ZN(n4997) );
  OR2_X1 U6155 ( .A1(n9370), .A2(n9042), .ZN(n4552) );
  AND2_X1 U6156 ( .A1(n9238), .A2(n8864), .ZN(n4553) );
  AND2_X1 U6157 ( .A1(n7733), .A2(n8482), .ZN(n4554) );
  AND2_X1 U6158 ( .A1(n6609), .A2(n10036), .ZN(n4555) );
  INV_X1 U6159 ( .A(n4802), .ZN(n4801) );
  NOR2_X1 U6160 ( .A1(n9227), .A2(n9216), .ZN(n4802) );
  AND2_X1 U6161 ( .A1(n4871), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4556) );
  INV_X1 U6162 ( .A(n7264), .ZN(n4791) );
  AND2_X1 U6163 ( .A1(n8799), .A2(n8806), .ZN(n7264) );
  NOR2_X1 U6164 ( .A1(n4769), .A2(n4767), .ZN(n4557) );
  NOR2_X1 U6165 ( .A1(n9312), .A2(n9330), .ZN(n4558) );
  AND4_X1 U6166 ( .A1(n5167), .A2(n5166), .A3(n5165), .A4(n5164), .ZN(n7582)
         );
  NOR2_X1 U6167 ( .A1(n8637), .A2(n8467), .ZN(n4559) );
  NAND2_X1 U6168 ( .A1(n6058), .A2(n6030), .ZN(n4560) );
  INV_X1 U6169 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5144) );
  OR2_X1 U6170 ( .A1(n9213), .A2(n4880), .ZN(n4879) );
  NAND2_X1 U6171 ( .A1(n8808), .A2(n7388), .ZN(n4561) );
  AOI21_X1 U6172 ( .B1(n8722), .B2(n5062), .A(n5060), .ZN(n5059) );
  AND2_X1 U6173 ( .A1(n4927), .A2(n7326), .ZN(n4562) );
  NOR2_X1 U6174 ( .A1(n8764), .A2(n8765), .ZN(n4563) );
  AND4_X2 U6175 ( .A1(n6125), .A2(n6124), .A3(n6123), .A4(n6122), .ZN(n9994)
         );
  INV_X1 U6176 ( .A(n9994), .ZN(n4841) );
  AND3_X1 U6177 ( .A1(n8961), .A2(n8974), .A3(n8899), .ZN(n4564) );
  INV_X2 U6178 ( .A(n5199), .ZN(n5537) );
  INV_X1 U6179 ( .A(n4869), .ZN(n4868) );
  OR2_X1 U6180 ( .A1(n4870), .A2(n6570), .ZN(n4869) );
  NAND2_X1 U6181 ( .A1(n4613), .A2(n4612), .ZN(n5069) );
  AND2_X1 U6182 ( .A1(n4823), .A2(n4826), .ZN(n9348) );
  NAND2_X1 U6183 ( .A1(n8125), .A2(n4508), .ZN(n4565) );
  AND2_X1 U6184 ( .A1(n5073), .A2(n6643), .ZN(n4566) );
  OR2_X1 U6185 ( .A1(n8022), .A2(n4731), .ZN(n4567) );
  NAND2_X1 U6186 ( .A1(n7170), .A2(n5044), .ZN(n4568) );
  INV_X1 U6187 ( .A(n4793), .ZN(n4784) );
  NAND2_X1 U6188 ( .A1(n7582), .A2(n4794), .ZN(n4793) );
  OR2_X1 U6189 ( .A1(n6578), .A2(n4902), .ZN(n4569) );
  INV_X1 U6190 ( .A(n8884), .ZN(n4688) );
  AND2_X1 U6191 ( .A1(n4859), .A2(n4858), .ZN(n4570) );
  OR2_X1 U6192 ( .A1(n6399), .A2(n6398), .ZN(n7945) );
  INV_X1 U6193 ( .A(n7945), .ZN(n4942) );
  NAND2_X1 U6194 ( .A1(n8340), .A2(n8348), .ZN(n8021) );
  AND2_X1 U6195 ( .A1(n5014), .A2(n8168), .ZN(n4571) );
  AND2_X1 U6196 ( .A1(n5011), .A2(n5015), .ZN(n4572) );
  AND2_X1 U6197 ( .A1(n4782), .A2(n4781), .ZN(n4573) );
  AND2_X1 U6198 ( .A1(n8130), .A2(n8131), .ZN(n8487) );
  INV_X1 U6199 ( .A(n8487), .ZN(n4744) );
  NOR2_X1 U6200 ( .A1(n6532), .A2(n6531), .ZN(n4574) );
  AND2_X1 U6201 ( .A1(n8175), .A2(n8168), .ZN(n5013) );
  NAND2_X1 U6202 ( .A1(n5503), .A2(n5502), .ZN(n9406) );
  AND2_X1 U6203 ( .A1(n4875), .A2(n4873), .ZN(n4575) );
  AND2_X1 U6204 ( .A1(n9751), .A2(n7704), .ZN(n8823) );
  AND2_X1 U6205 ( .A1(n4879), .A2(n4878), .ZN(n4576) );
  NAND2_X1 U6206 ( .A1(n9793), .A2(n9047), .ZN(n4577) );
  OR2_X1 U6207 ( .A1(n8180), .A2(n4715), .ZN(n4578) );
  INV_X1 U6208 ( .A(n4872), .ZN(n4871) );
  AND2_X1 U6209 ( .A1(n6023), .A2(n5007), .ZN(n4579) );
  AND2_X1 U6210 ( .A1(n4534), .A2(n4817), .ZN(n4580) );
  INV_X1 U6211 ( .A(n8036), .ZN(n7546) );
  AND2_X1 U6212 ( .A1(n8086), .A2(n8110), .ZN(n8036) );
  NAND2_X1 U6213 ( .A1(n9317), .A2(n4698), .ZN(n4581) );
  INV_X1 U6214 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6215 ( .A1(n5634), .A2(n5633), .ZN(n9152) );
  INV_X1 U6216 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5002) );
  NAND2_X1 U6217 ( .A1(n6621), .A2(n8154), .ZN(n8401) );
  AND2_X1 U6218 ( .A1(n4805), .A2(n4806), .ZN(n4582) );
  OR2_X1 U6219 ( .A1(n8053), .A2(n8054), .ZN(n8330) );
  INV_X1 U6220 ( .A(n8330), .ZN(n4722) );
  AND3_X1 U6221 ( .A1(n7831), .A2(n4934), .A3(n7997), .ZN(n4583) );
  INV_X1 U6222 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5028) );
  INV_X1 U6223 ( .A(n9046), .ZN(n9790) );
  NOR2_X1 U6224 ( .A1(n7813), .A2(n9431), .ZN(n7812) );
  NOR2_X1 U6225 ( .A1(n7815), .A2(n9004), .ZN(n4584) );
  AND4_X1 U6226 ( .A1(n5362), .A2(n5361), .A3(n5360), .A4(n5359), .ZN(n9611)
         );
  INV_X1 U6227 ( .A(n9698), .ZN(n6958) );
  AND3_X1 U6228 ( .A1(n5255), .A2(n5254), .A3(n5253), .ZN(n9698) );
  NAND2_X1 U6229 ( .A1(n7812), .A2(n4520), .ZN(n4659) );
  NAND2_X1 U6230 ( .A1(n5959), .A2(n5958), .ZN(n4585) );
  INV_X1 U6231 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6475) );
  OR2_X1 U6232 ( .A1(n5544), .A2(n4962), .ZN(n4586) );
  NAND2_X1 U6233 ( .A1(n6407), .A2(n6406), .ZN(n8380) );
  INV_X1 U6234 ( .A(n8380), .ZN(n7966) );
  NAND2_X1 U6235 ( .A1(n6586), .A2(n6585), .ZN(n8304) );
  AND2_X1 U6236 ( .A1(n4625), .A2(n4623), .ZN(n4587) );
  AND2_X1 U6237 ( .A1(n4961), .A2(n5559), .ZN(n4588) );
  INV_X1 U6238 ( .A(n6572), .ZN(n4854) );
  INV_X1 U6239 ( .A(n9899), .ZN(n4923) );
  NAND2_X1 U6240 ( .A1(n4774), .A2(n4791), .ZN(n4790) );
  INV_X1 U6241 ( .A(n8182), .ZN(n8199) );
  NAND2_X1 U6242 ( .A1(n8218), .A2(n8064), .ZN(n8182) );
  AND2_X1 U6243 ( .A1(n9637), .A2(n4507), .ZN(n4589) );
  NAND2_X1 U6244 ( .A1(n4839), .A2(n6554), .ZN(n7192) );
  XNOR2_X1 U6245 ( .A(n6230), .B(n7682), .ZN(n7453) );
  NAND2_X1 U6246 ( .A1(n5045), .A2(n7170), .ZN(n7287) );
  INV_X2 U6247 ( .A(n9801), .ZN(n9802) );
  OR2_X1 U6248 ( .A1(n6540), .A2(n6539), .ZN(n9801) );
  INV_X1 U6249 ( .A(n7755), .ZN(n4615) );
  INV_X1 U6250 ( .A(n9617), .ZN(n4816) );
  OAI21_X1 U6251 ( .B1(n6954), .B2(n4611), .A(n4609), .ZN(n7159) );
  NAND2_X1 U6252 ( .A1(n5841), .A2(n5840), .ZN(n7578) );
  NAND2_X1 U6253 ( .A1(n4940), .A2(n4939), .ZN(n7663) );
  AND2_X1 U6254 ( .A1(n4950), .A2(n4948), .ZN(n4590) );
  AND2_X1 U6255 ( .A1(n8257), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4591) );
  OR2_X1 U6256 ( .A1(n7265), .A2(n7268), .ZN(n9654) );
  INV_X1 U6257 ( .A(n9654), .ZN(n4662) );
  OR2_X1 U6258 ( .A1(n9825), .A2(n4824), .ZN(n4592) );
  NOR2_X1 U6259 ( .A1(n8261), .A2(n4923), .ZN(n4593) );
  INV_X1 U6260 ( .A(n5684), .ZN(n4809) );
  INV_X1 U6261 ( .A(n7268), .ZN(n4789) );
  AND2_X1 U6262 ( .A1(n7616), .A2(n8244), .ZN(n4594) );
  INV_X1 U6263 ( .A(n9751), .ZN(n4664) );
  NAND2_X1 U6264 ( .A1(n5774), .A2(n5085), .ZN(n6760) );
  NAND2_X1 U6265 ( .A1(n5776), .A2(n5775), .ZN(n7841) );
  NAND2_X1 U6266 ( .A1(n6954), .A2(n5805), .ZN(n6964) );
  NAND2_X1 U6267 ( .A1(n5819), .A2(n5820), .ZN(n5046) );
  INV_X1 U6268 ( .A(n5046), .ZN(n5042) );
  AND2_X1 U6269 ( .A1(n4631), .A2(n4630), .ZN(n4595) );
  NAND2_X1 U6270 ( .A1(n6080), .A2(n6079), .ZN(n8643) );
  INV_X1 U6271 ( .A(n6661), .ZN(n8203) );
  XNOR2_X1 U6272 ( .A(n6048), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6661) );
  NOR2_X1 U6273 ( .A1(n5146), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n9451) );
  INV_X1 U6274 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6135) );
  INV_X1 U6275 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5000) );
  AND3_X2 U6276 ( .A1(n5074), .A2(n4579), .A3(n6143), .ZN(n6042) );
  NAND2_X1 U6277 ( .A1(n8464), .A2(n8135), .ZN(n8449) );
  NAND2_X1 U6278 ( .A1(n6624), .A2(n8176), .ZN(n8353) );
  AOI21_X1 U6279 ( .B1(n8061), .B2(n8023), .A(n6603), .ZN(n6604) );
  OAI21_X1 U6280 ( .B1(n5326), .B2(n4975), .A(n4972), .ZN(n5370) );
  NAND2_X1 U6281 ( .A1(n5194), .A2(n4570), .ZN(n4857) );
  INV_X1 U6282 ( .A(n8202), .ZN(n4741) );
  INV_X1 U6283 ( .A(n4719), .ZN(n4718) );
  NOR2_X2 U6284 ( .A1(n8185), .A2(n8186), .ZN(n4723) );
  INV_X2 U6285 ( .A(n5100), .ZN(n6680) );
  NAND2_X1 U6286 ( .A1(n4958), .A2(n4588), .ZN(n5562) );
  OR2_X1 U6287 ( .A1(n9994), .A2(n7194), .ZN(n8074) );
  OAI21_X1 U6288 ( .B1(n4741), .B2(n4740), .A(n4738), .ZN(n4737) );
  OAI21_X1 U6289 ( .B1(n4724), .B2(n4722), .A(n4723), .ZN(n4719) );
  AND4_X1 U6290 ( .A1(n8200), .A2(n8199), .A3(n8212), .A4(n8206), .ZN(n4739)
         );
  OAI211_X1 U6291 ( .C1(n8181), .C2(n4715), .A(n4718), .B(n4578), .ZN(n8192)
         );
  NAND2_X1 U6292 ( .A1(n4737), .A2(n8203), .ZN(n4736) );
  OAI21_X1 U6293 ( .B1(n8197), .B2(n8304), .A(n4739), .ZN(n4738) );
  OAI21_X1 U6294 ( .B1(n4721), .B2(n4514), .A(n4720), .ZN(n4717) );
  INV_X1 U6295 ( .A(n4716), .ZN(n8189) );
  NAND2_X2 U6296 ( .A1(n8353), .A2(n8179), .ZN(n6626) );
  NAND2_X1 U6297 ( .A1(n9985), .A2(n6602), .ZN(n8061) );
  OAI21_X1 U6298 ( .B1(n6668), .B2(n10065), .A(n6653), .ZN(n6655) );
  NAND2_X1 U6299 ( .A1(n6801), .A2(n6802), .ZN(n6848) );
  XNOR2_X1 U6300 ( .A(n8239), .B(n9931), .ZN(n9941) );
  AOI21_X2 U6301 ( .B1(n7630), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7627), .ZN(
        n7709) );
  OAI21_X1 U6302 ( .B1(n5805), .B2(n4611), .A(n5814), .ZN(n4610) );
  NAND2_X2 U6303 ( .A1(n6953), .A2(n6955), .ZN(n6954) );
  AOI21_X2 U6304 ( .B1(n4768), .B2(n4585), .A(n4646), .ZN(n8722) );
  NAND2_X1 U6305 ( .A1(n7702), .A2(n7755), .ZN(n4619) );
  OAI21_X1 U6306 ( .B1(n7702), .B2(n4616), .A(n4614), .ZN(n5888) );
  INV_X1 U6307 ( .A(n5888), .ZN(n5881) );
  AND2_X2 U6308 ( .A1(n5895), .A2(n4620), .ZN(n8776) );
  NAND3_X1 U6309 ( .A1(n8656), .A2(n4621), .A3(n8654), .ZN(n4620) );
  NAND2_X2 U6310 ( .A1(n8776), .A2(n8775), .ZN(n8774) );
  INV_X1 U6311 ( .A(n4631), .ZN(n9874) );
  NAND2_X1 U6312 ( .A1(n6827), .A2(n9863), .ZN(n4630) );
  NAND2_X1 U6313 ( .A1(n4635), .A2(n4632), .ZN(n6825) );
  NAND2_X1 U6314 ( .A1(n4634), .A2(n4633), .ZN(n4632) );
  INV_X1 U6315 ( .A(n9837), .ZN(n4633) );
  MUX2_X1 U6316 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n8273), .Z(n6772) );
  INV_X1 U6317 ( .A(n9838), .ZN(n4634) );
  MUX2_X1 U6318 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8273), .Z(n6796) );
  NAND2_X1 U6319 ( .A1(n7611), .A2(n4527), .ZN(n4637) );
  NAND2_X1 U6320 ( .A1(n4645), .A2(n5039), .ZN(n7558) );
  NAND3_X1 U6321 ( .A1(n5816), .A2(n7160), .A3(n5041), .ZN(n4645) );
  INV_X1 U6322 ( .A(n5456), .ZN(n5657) );
  NAND3_X1 U6323 ( .A1(n4761), .A2(n4510), .A3(n4505), .ZN(n5443) );
  NAND2_X1 U6324 ( .A1(n5456), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6325 ( .A1(n4501), .A2(n4680), .ZN(n5136) );
  NAND3_X1 U6326 ( .A1(n4501), .A2(n4680), .A3(n5137), .ZN(n4655) );
  NAND2_X1 U6327 ( .A1(n7812), .A2(n4656), .ZN(n9256) );
  INV_X1 U6328 ( .A(n4659), .ZN(n9291) );
  AND2_X1 U6329 ( .A1(n9180), .A2(n4671), .ZN(n9167) );
  NAND2_X1 U6330 ( .A1(n9180), .A2(n5696), .ZN(n9181) );
  NAND2_X1 U6331 ( .A1(n4678), .A2(n4501), .ZN(n5146) );
  NAND2_X1 U6332 ( .A1(n8880), .A2(n4564), .ZN(n4682) );
  NAND2_X1 U6333 ( .A1(n4681), .A2(n4683), .ZN(n8894) );
  NAND3_X1 U6334 ( .A1(n4682), .A2(n8881), .A3(n4685), .ZN(n4681) );
  INV_X1 U6335 ( .A(n8845), .ZN(n4690) );
  OAI21_X1 U6336 ( .B1(n4690), .B2(n4693), .A(n4691), .ZN(n8837) );
  INV_X1 U6337 ( .A(n9007), .ZN(n4700) );
  NAND2_X1 U6338 ( .A1(n4701), .A2(n4702), .ZN(n8871) );
  NAND3_X1 U6339 ( .A1(n8862), .A2(n4705), .A3(n8861), .ZN(n4701) );
  AOI21_X1 U6340 ( .B1(n4713), .B2(n8181), .A(n4717), .ZN(n4716) );
  INV_X1 U6341 ( .A(n8180), .ZN(n4714) );
  INV_X1 U6342 ( .A(n8187), .ZN(n4724) );
  NAND2_X1 U6343 ( .A1(n4725), .A2(n4726), .ZN(n8170) );
  NAND2_X1 U6344 ( .A1(n8162), .A2(n4727), .ZN(n4725) );
  NAND2_X1 U6345 ( .A1(n8167), .A2(n8166), .ZN(n4733) );
  NAND2_X1 U6346 ( .A1(n4742), .A2(n4743), .ZN(n8133) );
  NAND2_X1 U6347 ( .A1(n8126), .A2(n4745), .ZN(n4742) );
  NAND3_X1 U6348 ( .A1(n5195), .A2(n4510), .A3(n4505), .ZN(n5420) );
  NAND2_X1 U6349 ( .A1(n8745), .A2(n4766), .ZN(n4765) );
  OAI21_X1 U6350 ( .B1(n4561), .B2(n4792), .A(n4787), .ZN(n4786) );
  OR2_X1 U6351 ( .A1(n9375), .A2(n9228), .ZN(n4800) );
  NAND2_X1 U6352 ( .A1(n7811), .A2(n4515), .ZN(n4804) );
  NAND2_X1 U6353 ( .A1(n5754), .A2(n6884), .ZN(n5759) );
  NAND2_X1 U6354 ( .A1(n7464), .A2(n4580), .ZN(n4810) );
  NAND2_X1 U6355 ( .A1(n4810), .A2(n4811), .ZN(n7802) );
  NAND3_X1 U6356 ( .A1(n9158), .A2(n9784), .A3(n9342), .ZN(n4822) );
  NAND2_X1 U6357 ( .A1(n5676), .A2(n5675), .ZN(n9671) );
  OAI21_X1 U6358 ( .B1(n9268), .B2(n5690), .A(n5689), .ZN(n9252) );
  AOI22_X1 U6359 ( .A1(n9161), .A2(n9164), .B1(n9174), .B2(n9359), .ZN(n9157)
         );
  MUX2_X1 U6360 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9437), .S(n9802), .Z(
        P1_U3518) );
  XNOR2_X1 U6361 ( .A(n9147), .B(n9146), .ZN(n4827) );
  NAND2_X1 U6362 ( .A1(n4831), .A2(n4828), .ZN(n7465) );
  NAND3_X1 U6363 ( .A1(n4833), .A2(n8998), .A3(n4832), .ZN(n4831) );
  INV_X1 U6364 ( .A(n7360), .ZN(n4833) );
  NAND3_X1 U6365 ( .A1(n8070), .A2(n4840), .A3(n9991), .ZN(n4834) );
  OAI211_X1 U6366 ( .C1(n4837), .C2(n4835), .A(n6605), .B(n4834), .ZN(n6556)
         );
  NAND2_X1 U6367 ( .A1(n8414), .A2(n4844), .ZN(n4843) );
  NAND3_X1 U6368 ( .A1(n4859), .A2(n4862), .A3(n4858), .ZN(n4856) );
  OAI22_X2 U6369 ( .A1(n8494), .A2(n4863), .B1(n4865), .B2(n4536), .ZN(n8453)
         );
  NAND3_X1 U6370 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .A3(P2_IR_REG_31__SCAN_IN), .ZN(n4872) );
  NOR2_X2 U6371 ( .A1(n6112), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6143) );
  AND2_X2 U6372 ( .A1(n4874), .A2(n4575), .ZN(n9162) );
  INV_X1 U6373 ( .A(n4879), .ZN(n9212) );
  NAND2_X1 U6374 ( .A1(n4883), .A2(n4884), .ZN(n9328) );
  NAND2_X1 U6375 ( .A1(n4889), .A2(n4887), .ZN(n6561) );
  NAND2_X1 U6376 ( .A1(n6577), .A2(n4896), .ZN(n4894) );
  NAND2_X1 U6377 ( .A1(n6577), .A2(n4899), .ZN(n4898) );
  NAND2_X1 U6378 ( .A1(n4894), .A2(n4895), .ZN(n8295) );
  NAND2_X1 U6379 ( .A1(n6577), .A2(n6576), .ZN(n8358) );
  NOR2_X1 U6380 ( .A1(n8585), .A2(n8347), .ZN(n4902) );
  INV_X1 U6381 ( .A(n4907), .ZN(n9274) );
  MUX2_X1 U6382 ( .A(n5219), .B(n6086), .S(n5003), .Z(n5094) );
  NAND3_X1 U6383 ( .A1(n4998), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4909) );
  NAND3_X1 U6384 ( .A1(n5000), .A2(n7887), .A3(n4999), .ZN(n4910) );
  NOR2_X2 U6385 ( .A1(n7481), .A2(n6244), .ZN(n7600) );
  NOR2_X2 U6386 ( .A1(n9923), .A2(n4591), .ZN(n8239) );
  NAND2_X1 U6387 ( .A1(n4920), .A2(n4919), .ZN(n9473) );
  XNOR2_X1 U6388 ( .A(n8240), .B(n9965), .ZN(n9978) );
  OAI21_X1 U6389 ( .B1(n4929), .B2(n7327), .A(n4928), .ZN(n7478) );
  INV_X1 U6390 ( .A(n7478), .ZN(n7477) );
  NAND2_X1 U6391 ( .A1(n6351), .A2(n4513), .ZN(n4931) );
  NAND2_X1 U6392 ( .A1(n7989), .A2(n6450), .ZN(n6499) );
  OAI211_X1 U6393 ( .C1(n7840), .C2(n7839), .A(n4936), .B(n7838), .ZN(P2_U3160) );
  NAND2_X1 U6394 ( .A1(n7929), .A2(n4937), .ZN(n7937) );
  NAND2_X1 U6395 ( .A1(n7945), .A2(n4943), .ZN(n4941) );
  NAND2_X1 U6396 ( .A1(n7945), .A2(n6400), .ZN(n7897) );
  NAND2_X1 U6397 ( .A1(n7127), .A2(n6171), .ZN(n7131) );
  AND2_X1 U6398 ( .A1(n7131), .A2(n6177), .ZN(n7151) );
  INV_X1 U6399 ( .A(n7003), .ZN(n4944) );
  NAND2_X1 U6400 ( .A1(n7654), .A2(n4955), .ZN(n4953) );
  NAND2_X1 U6401 ( .A1(n6058), .A2(n4956), .ZN(n6046) );
  NAND2_X1 U6402 ( .A1(n6032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U6403 ( .A1(n6476), .A2(n6475), .ZN(n6054) );
  NAND2_X1 U6404 ( .A1(n6033), .A2(n10184), .ZN(n6463) );
  NAND3_X1 U6405 ( .A1(n5513), .A2(n5512), .A3(n4959), .ZN(n4958) );
  NAND3_X1 U6406 ( .A1(n5513), .A2(n5512), .A3(n4964), .ZN(n4963) );
  NAND2_X1 U6407 ( .A1(n5513), .A2(n5512), .ZN(n5528) );
  INV_X1 U6408 ( .A(n5527), .ZN(n4964) );
  NAND2_X1 U6409 ( .A1(n5575), .A2(n4969), .ZN(n4967) );
  OAI22_X2 U6410 ( .A1(n5416), .A2(n4984), .B1(SI_15_), .B2(n5417), .ZN(n5437)
         );
  OAI21_X2 U6411 ( .B1(n5437), .B2(n5436), .A(n5435), .ZN(n5500) );
  NAND3_X1 U6412 ( .A1(n9020), .A2(n9021), .A3(n9030), .ZN(n4989) );
  NAND2_X1 U6413 ( .A1(n5003), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U6414 ( .A1(n6621), .A2(n5004), .ZN(n8388) );
  NAND2_X1 U6415 ( .A1(n8388), .A2(n8059), .ZN(n6622) );
  NAND2_X1 U6416 ( .A1(n5010), .A2(n4572), .ZN(n6624) );
  AND2_X2 U6417 ( .A1(n6065), .A2(n5026), .ZN(n6080) );
  OAI21_X1 U6418 ( .B1(n8501), .B2(n5032), .A(n5029), .ZN(n8464) );
  OAI21_X1 U6419 ( .B1(n8501), .B2(n6613), .A(n6614), .ZN(n8488) );
  NAND3_X1 U6420 ( .A1(n5035), .A2(n7698), .A3(n5853), .ZN(n7638) );
  NAND3_X1 U6421 ( .A1(n5816), .A2(n7160), .A3(n5046), .ZN(n5045) );
  NAND2_X1 U6422 ( .A1(n5816), .A2(n7160), .ZN(n7169) );
  NAND2_X1 U6423 ( .A1(n5047), .A2(n5050), .ZN(n5933) );
  NAND2_X1 U6424 ( .A1(n8703), .A2(n5048), .ZN(n5047) );
  NOR2_X1 U6425 ( .A1(n5057), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5054) );
  AND2_X1 U6426 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  AOI21_X2 U6427 ( .B1(n7117), .B2(n6558), .A(n6557), .ZN(n7219) );
  NAND2_X1 U6428 ( .A1(n6497), .A2(n7997), .ZN(n6530) );
  XNOR2_X1 U6429 ( .A(n5700), .B(n8984), .ZN(n9137) );
  INV_X1 U6430 ( .A(n5091), .ZN(n5090) );
  NAND2_X1 U6431 ( .A1(n5609), .A2(n5608), .ZN(n5630) );
  NAND2_X1 U6432 ( .A1(n5641), .A2(n5640), .ZN(n5645) );
  NAND2_X1 U6433 ( .A1(n6052), .A2(n6051), .ZN(n6056) );
  NAND2_X1 U6434 ( .A1(n6034), .A2(n6463), .ZN(n6472) );
  OR2_X1 U6435 ( .A1(n6033), .A2(n10184), .ZN(n6034) );
  NAND2_X1 U6436 ( .A1(n7149), .A2(n6193), .ZN(n7231) );
  INV_X1 U6437 ( .A(n5230), .ZN(n5232) );
  INV_X1 U6438 ( .A(n6120), .ZN(n6133) );
  XNOR2_X1 U6439 ( .A(n5303), .B(n5302), .ZN(n6721) );
  NAND2_X1 U6440 ( .A1(n6499), .A2(n6498), .ZN(n6497) );
  INV_X1 U6441 ( .A(n7186), .ZN(n8024) );
  AOI21_X2 U6442 ( .B1(n5303), .B2(n5302), .A(n5301), .ZN(n5309) );
  OAI21_X1 U6443 ( .B1(n6530), .B2(n7840), .A(n5087), .ZN(P2_U3154) );
  NAND2_X1 U6444 ( .A1(n6550), .A2(n10007), .ZN(n8063) );
  INV_X1 U6445 ( .A(n6550), .ZN(n6548) );
  AND2_X1 U6446 ( .A1(n6042), .A2(n6035), .ZN(n6058) );
  AOI21_X1 U6447 ( .B1(n6563), .B2(n7549), .A(n6562), .ZN(n7547) );
  NAND4_X2 U6448 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n8232)
         );
  NAND2_X1 U6449 ( .A1(n4498), .A2(n7865), .ZN(n6118) );
  NAND2_X1 U6450 ( .A1(n6496), .A2(n6495), .ZN(n7997) );
  INV_X2 U6451 ( .A(n10065), .ZN(n10063) );
  OR2_X1 U6452 ( .A1(n7823), .A2(n8537), .ZN(n5070) );
  OR2_X1 U6453 ( .A1(n6644), .A2(n10046), .ZN(n5073) );
  AND2_X1 U6454 ( .A1(n5656), .A2(n5655), .ZN(n5075) );
  INV_X4 U6455 ( .A(n6680), .ZN(n8014) );
  OR2_X1 U6456 ( .A1(n7823), .A2(n8620), .ZN(n5078) );
  OR2_X1 U6457 ( .A1(n9825), .A2(n5747), .ZN(n5079) );
  NOR2_X1 U6458 ( .A1(n5331), .A2(n5320), .ZN(n5080) );
  INV_X1 U6459 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5088) );
  INV_X1 U6460 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5161) );
  AND2_X1 U6461 ( .A1(n9346), .A2(n9345), .ZN(n9347) );
  AND4_X1 U6462 ( .A1(n5133), .A2(n5132), .A3(n5131), .A4(n5656), .ZN(n5081)
         );
  AND2_X1 U6463 ( .A1(n5978), .A2(n5977), .ZN(n6531) );
  INV_X1 U6464 ( .A(n9152), .ZN(n9343) );
  NAND2_X1 U6465 ( .A1(n6792), .A2(n9664), .ZN(n9296) );
  OR2_X1 U6466 ( .A1(n6002), .A2(n5750), .ZN(n9781) );
  AND2_X1 U6467 ( .A1(n8732), .A2(n5932), .ZN(n5083) );
  OR2_X1 U6468 ( .A1(n6707), .A2(n7073), .ZN(n5084) );
  OR2_X1 U6469 ( .A1(n6007), .A2(n5770), .ZN(n5085) );
  INV_X1 U6470 ( .A(n5703), .ZN(n5702) );
  INV_X1 U6471 ( .A(n8435), .ZN(n6617) );
  INV_X1 U6472 ( .A(n9362), .ZN(n5696) );
  AND2_X1 U6473 ( .A1(n8511), .A2(n8297), .ZN(n5086) );
  AND2_X1 U6474 ( .A1(n6529), .A2(n6528), .ZN(n5087) );
  INV_X1 U6475 ( .A(n8797), .ZN(n8915) );
  INV_X1 U6476 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5129) );
  INV_X1 U6477 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6027) );
  INV_X1 U6478 ( .A(n8900), .ZN(n8883) );
  INV_X1 U6479 ( .A(n9781), .ZN(n9344) );
  INV_X1 U6480 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6064) );
  INV_X1 U6481 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6035) );
  INV_X1 U6482 ( .A(n7640), .ZN(n5853) );
  INV_X1 U6483 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6134) );
  INV_X1 U6484 ( .A(n6270), .ZN(n6269) );
  INV_X1 U6485 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6183) );
  OR2_X1 U6486 ( .A1(n8588), .A2(n8380), .ZN(n6576) );
  OR2_X1 U6487 ( .A1(n7748), .A2(n8223), .ZN(n6567) );
  INV_X1 U6488 ( .A(n8098), .ZN(n6603) );
  INV_X1 U6489 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U6490 ( .A1(n9152), .A2(n9171), .ZN(n5699) );
  AND2_X1 U6491 ( .A1(n5473), .A2(n5472), .ZN(n5474) );
  NOR2_X1 U6492 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5130) );
  NAND2_X1 U6493 ( .A1(n6135), .A2(n6134), .ZN(n6150) );
  INV_X1 U6494 ( .A(n6429), .ZN(n6117) );
  INV_X1 U6495 ( .A(n6456), .ZN(n6455) );
  NAND2_X1 U6496 ( .A1(n6329), .A2(n6328), .ZN(n6345) );
  NAND2_X1 U6497 ( .A1(n6211), .A2(n6210), .ZN(n6219) );
  NAND2_X1 U6498 ( .A1(n7153), .A2(n8228), .ZN(n6560) );
  NAND2_X1 U6499 ( .A1(n7187), .A2(n7215), .ZN(n7185) );
  NAND2_X1 U6500 ( .A1(n6571), .A2(n5077), .ZN(n8414) );
  OR2_X1 U6501 ( .A1(n6206), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U6502 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n5569), .ZN(n5583) );
  AND2_X1 U6503 ( .A1(n5600), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5618) );
  INV_X1 U6504 ( .A(n7849), .ZN(n5149) );
  INV_X1 U6505 ( .A(n9240), .ZN(n9257) );
  NOR2_X1 U6506 ( .A1(n9321), .A2(n5702), .ZN(n6003) );
  NAND2_X1 U6507 ( .A1(n5400), .A2(SI_14_), .ZN(n5401) );
  AND2_X1 U6508 ( .A1(n5262), .A2(n5104), .ZN(n5246) );
  INV_X1 U6509 ( .A(n8437), .ZN(n7907) );
  AND2_X1 U6510 ( .A1(n6095), .A2(n7185), .ZN(n6940) );
  NAND2_X1 U6511 ( .A1(n6426), .A2(n6425), .ZN(n6441) );
  INV_X1 U6512 ( .A(n8468), .ZN(n8001) );
  OR2_X1 U6513 ( .A1(n6118), .A2(n6088), .ZN(n6094) );
  AND2_X1 U6514 ( .A1(n6771), .A2(n7809), .ZN(n6803) );
  NAND2_X1 U6515 ( .A1(n6455), .A2(n6454), .ZN(n6501) );
  AND2_X1 U6516 ( .A1(n7374), .A2(n8105), .ZN(n8101) );
  OR2_X1 U6517 ( .A1(n10057), .A2(n7116), .ZN(n9987) );
  NOR2_X1 U6518 ( .A1(n7109), .A2(n7111), .ZN(n6659) );
  INV_X1 U6519 ( .A(n8334), .ZN(n8335) );
  AND2_X1 U6520 ( .A1(n8135), .A2(n8448), .ZN(n8463) );
  INV_X1 U6521 ( .A(n8484), .ZN(n10000) );
  NAND2_X1 U6522 ( .A1(n6470), .A2(n6469), .ZN(n7109) );
  INV_X1 U6523 ( .A(n8733), .ZN(n5938) );
  INV_X1 U6524 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7581) );
  INV_X1 U6525 ( .A(n4502), .ZN(n7068) );
  INV_X1 U6526 ( .A(n9142), .ZN(n5706) );
  INV_X1 U6527 ( .A(n9180), .ZN(n9195) );
  AND2_X1 U6528 ( .A1(n8809), .A2(n8814), .ZN(n7397) );
  OR2_X1 U6529 ( .A1(n6002), .A2(n5701), .ZN(n9321) );
  INV_X1 U6530 ( .A(n8998), .ZN(n9627) );
  AND2_X1 U6531 ( .A1(n5724), .A2(n9026), .ZN(n6784) );
  NOR2_X1 U6532 ( .A1(n5727), .A2(n7770), .ZN(n6698) );
  AND2_X1 U6533 ( .A1(n5561), .A2(n5550), .ZN(n5559) );
  NAND2_X1 U6534 ( .A1(n5496), .A2(n5480), .ZN(n5495) );
  NAND2_X1 U6535 ( .A1(n6109), .A2(n6108), .ZN(n6995) );
  INV_X1 U6536 ( .A(n7994), .ZN(n8003) );
  AOI21_X1 U6537 ( .B1(n7890), .B2(n7891), .A(n6294), .ZN(n8000) );
  AND2_X1 U6538 ( .A1(n6434), .A2(n6433), .ZN(n8332) );
  AND4_X1 U6539 ( .A1(n6250), .A2(n6249), .A3(n6248), .A4(n6247), .ZN(n8116)
         );
  AND4_X1 U6540 ( .A1(n6224), .A2(n6223), .A3(n6222), .A4(n6221), .ZN(n7682)
         );
  INV_X1 U6541 ( .A(n9875), .ZN(n9973) );
  AND2_X1 U6542 ( .A1(n6803), .A2(n8273), .ZN(n9974) );
  XNOR2_X1 U6543 ( .A(n8304), .B(n8320), .ZN(n8296) );
  INV_X1 U6544 ( .A(n9989), .ZN(n8472) );
  NAND2_X1 U6545 ( .A1(n6610), .A2(n8101), .ZN(n7375) );
  INV_X1 U6546 ( .A(n9995), .ZN(n8481) );
  INV_X1 U6547 ( .A(n8476), .ZN(n8502) );
  INV_X1 U6548 ( .A(n8537), .ZN(n8549) );
  OR3_X1 U6549 ( .A1(n6660), .A2(n6659), .A3(n6718), .ZN(n7107) );
  INV_X1 U6550 ( .A(n6620), .ZN(n8413) );
  OR2_X1 U6551 ( .A1(n6649), .A2(n6648), .ZN(n6650) );
  NAND2_X1 U6552 ( .A1(n6776), .A2(n6737), .ZN(n6718) );
  NOR2_X1 U6553 ( .A1(n6241), .A2(n6240), .ZN(n7613) );
  INV_X1 U6554 ( .A(n9705), .ZN(n6988) );
  AND4_X1 U6555 ( .A1(n5607), .A2(n5606), .A3(n5605), .A4(n5604), .ZN(n9367)
         );
  AND4_X1 U6556 ( .A1(n5588), .A2(n5587), .A3(n5586), .A4(n5585), .ZN(n9358)
         );
  AND4_X1 U6557 ( .A1(n5397), .A2(n5396), .A3(n5395), .A4(n5394), .ZN(n9612)
         );
  AND2_X1 U6558 ( .A1(n6751), .A2(n6750), .ZN(n7067) );
  OR2_X1 U6559 ( .A1(n7069), .A2(n7068), .ZN(n9599) );
  AND2_X1 U6560 ( .A1(n7067), .A2(n9064), .ZN(n9590) );
  INV_X1 U6561 ( .A(n9321), .ZN(n9673) );
  INV_X1 U6562 ( .A(n8868), .ZN(n9214) );
  AND2_X1 U6563 ( .A1(n8831), .A2(n9606), .ZN(n8999) );
  INV_X1 U6564 ( .A(n9264), .ZN(n9676) );
  INV_X1 U6565 ( .A(n9668), .ZN(n9652) );
  INV_X1 U6566 ( .A(n9777), .ZN(n9754) );
  NAND2_X1 U6567 ( .A1(n9626), .A2(n9796), .ZN(n9784) );
  AND2_X1 U6568 ( .A1(n6706), .A2(n5723), .ZN(n9026) );
  AND2_X1 U6569 ( .A1(n5327), .A2(n5316), .ZN(n9489) );
  INV_X1 U6570 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10367) );
  INV_X1 U6571 ( .A(n7997), .ZN(n7970) );
  NAND2_X1 U6572 ( .A1(n6507), .A2(n6506), .ZN(n8320) );
  OR2_X1 U6573 ( .A1(P2_U3150), .A2(n6777), .ZN(n9897) );
  OR2_X1 U6574 ( .A1(n6798), .A2(n8273), .ZN(n9980) );
  AND2_X1 U6575 ( .A1(n8439), .A2(n8438), .ZN(n8541) );
  NAND2_X1 U6576 ( .A1(n4500), .A2(n7178), .ZN(n8476) );
  NAND2_X1 U6577 ( .A1(n10081), .A2(n10055), .ZN(n8537) );
  INV_X1 U6578 ( .A(n10081), .ZN(n10079) );
  INV_X1 U6579 ( .A(n6623), .ZN(n8585) );
  OR2_X1 U6580 ( .A1(n10065), .A2(n10059), .ZN(n8615) );
  OR2_X1 U6581 ( .A1(n10065), .A2(n10057), .ZN(n8620) );
  AND2_X1 U6582 ( .A1(n6651), .A2(n6650), .ZN(n10065) );
  INV_X1 U6583 ( .A(n10105), .ZN(n6748) );
  NAND2_X1 U6584 ( .A1(n6734), .A2(n6733), .ZN(n10105) );
  INV_X1 U6585 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7102) );
  INV_X1 U6586 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6731) );
  INV_X1 U6587 ( .A(n8768), .ZN(n8780) );
  INV_X1 U6588 ( .A(n8777), .ZN(n8754) );
  INV_X1 U6589 ( .A(n8769), .ZN(n8786) );
  INV_X1 U6590 ( .A(n9380), .ZN(n9228) );
  OR2_X1 U6591 ( .A1(n6792), .A2(n9021), .ZN(n9264) );
  INV_X1 U6592 ( .A(n9677), .ZN(n9336) );
  INV_X1 U6593 ( .A(n9296), .ZN(n9666) );
  NAND2_X1 U6594 ( .A1(n9801), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6542) );
  INV_X1 U6595 ( .A(n9681), .ZN(n9680) );
  INV_X1 U6596 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10251) );
  INV_X1 U6597 ( .A(n8233), .ZN(P2_U3893) );
  INV_X1 U6598 ( .A(SI_1_), .ZN(n5089) );
  NAND2_X1 U6599 ( .A1(n5090), .A2(n5089), .ZN(n5092) );
  NAND2_X1 U6600 ( .A1(n5091), .A2(SI_1_), .ZN(n5096) );
  NAND2_X1 U6601 ( .A1(n5092), .A2(n5096), .ZN(n5206) );
  INV_X1 U6602 ( .A(n5206), .ZN(n5095) );
  INV_X1 U6603 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6086) );
  INV_X1 U6604 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5219) );
  INV_X1 U6605 ( .A(SI_0_), .ZN(n5093) );
  NOR2_X1 U6606 ( .A1(n5094), .A2(n5093), .ZN(n5204) );
  NAND2_X1 U6607 ( .A1(n5095), .A2(n5204), .ZN(n5208) );
  NAND2_X1 U6608 ( .A1(n5208), .A2(n5096), .ZN(n5230) );
  MUX2_X1 U6609 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5100), .Z(n5097) );
  NAND2_X1 U6610 ( .A1(n5097), .A2(SI_2_), .ZN(n5099) );
  OAI21_X1 U6611 ( .B1(n5097), .B2(SI_2_), .A(n5099), .ZN(n5231) );
  INV_X1 U6612 ( .A(n5231), .ZN(n5098) );
  NAND2_X1 U6613 ( .A1(n5230), .A2(n5098), .ZN(n5233) );
  NAND2_X1 U6614 ( .A1(n5233), .A2(n5099), .ZN(n5247) );
  MUX2_X1 U6615 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5100), .Z(n5101) );
  NAND2_X1 U6616 ( .A1(n5101), .A2(SI_3_), .ZN(n5262) );
  INV_X1 U6617 ( .A(n5101), .ZN(n5103) );
  INV_X1 U6618 ( .A(SI_3_), .ZN(n5102) );
  NAND2_X1 U6619 ( .A1(n5103), .A2(n5102), .ZN(n5104) );
  NAND2_X1 U6620 ( .A1(n5247), .A2(n5246), .ZN(n5263) );
  MUX2_X1 U6621 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n8014), .Z(n5105) );
  NAND2_X1 U6622 ( .A1(n5105), .A2(SI_4_), .ZN(n5265) );
  AND2_X1 U6623 ( .A1(n5262), .A2(n5265), .ZN(n5109) );
  INV_X1 U6624 ( .A(n5105), .ZN(n5107) );
  INV_X1 U6625 ( .A(SI_4_), .ZN(n5106) );
  NAND2_X1 U6626 ( .A1(n5107), .A2(n5106), .ZN(n5264) );
  MUX2_X1 U6627 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8014), .Z(n5110) );
  NAND2_X1 U6628 ( .A1(n5110), .A2(SI_5_), .ZN(n5113) );
  INV_X1 U6629 ( .A(n5110), .ZN(n5111) );
  NAND2_X1 U6630 ( .A1(n5111), .A2(n10364), .ZN(n5112) );
  NAND2_X1 U6631 ( .A1(n5290), .A2(n5289), .ZN(n5292) );
  MUX2_X1 U6632 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n8014), .Z(n5114) );
  NAND2_X1 U6633 ( .A1(n5114), .A2(SI_6_), .ZN(n5118) );
  INV_X1 U6634 ( .A(n5114), .ZN(n5116) );
  INV_X1 U6635 ( .A(SI_6_), .ZN(n5115) );
  NAND2_X1 U6636 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  MUX2_X1 U6637 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8014), .Z(n5119) );
  INV_X1 U6638 ( .A(n5119), .ZN(n5120) );
  INV_X1 U6639 ( .A(SI_7_), .ZN(n10320) );
  NAND2_X1 U6640 ( .A1(n5120), .A2(n10320), .ZN(n5121) );
  MUX2_X1 U6641 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n8014), .Z(n5123) );
  INV_X1 U6642 ( .A(n5123), .ZN(n5125) );
  INV_X1 U6643 ( .A(SI_8_), .ZN(n5124) );
  NAND2_X1 U6644 ( .A1(n5125), .A2(n5124), .ZN(n5126) );
  MUX2_X1 U6645 ( .A(n6731), .B(n10251), .S(n8014), .Z(n5299) );
  NOR2_X1 U6646 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5133) );
  NOR2_X1 U6647 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5132) );
  NOR2_X1 U6648 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5131) );
  INV_X1 U6649 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5134) );
  INV_X2 U6650 ( .A(n5209), .ZN(n8888) );
  NAND2_X1 U6651 ( .A1(n6721), .A2(n8888), .ZN(n5143) );
  INV_X1 U6652 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6653 ( .A1(n5195), .A2(n5139), .ZN(n5348) );
  NAND2_X1 U6654 ( .A1(n5348), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5172) );
  OAI21_X1 U6655 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6656 ( .A1(n5172), .A2(n5140), .ZN(n5313) );
  INV_X1 U6657 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5141) );
  XNOR2_X1 U6658 ( .A(n5313), .B(n5141), .ZN(n9108) );
  AOI22_X1 U6659 ( .A1(n5485), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5484), .B2(
        n9108), .ZN(n5142) );
  XNOR2_X2 U6660 ( .A(n5145), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5151) );
  INV_X1 U6661 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6662 ( .A1(n5665), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5155) );
  NOR2_X2 U6663 ( .A1(n5151), .A2(n7849), .ZN(n5241) );
  NAND2_X1 U6664 ( .A1(n5241), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6665 ( .A1(n5186), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5178) );
  AND2_X1 U6666 ( .A1(n5163), .A2(n7581), .ZN(n5150) );
  NOR2_X1 U6667 ( .A1(n5319), .A2(n5150), .ZN(n7584) );
  NAND2_X1 U6668 ( .A1(n5537), .A2(n7584), .ZN(n5153) );
  INV_X1 U6669 ( .A(n5151), .ZN(n7862) );
  NAND2_X1 U6670 ( .A1(n6722), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5152) );
  XNOR2_X1 U6671 ( .A(n5157), .B(n5156), .ZN(n6709) );
  NAND2_X1 U6672 ( .A1(n6709), .A2(n8888), .ZN(n5160) );
  NAND2_X1 U6673 ( .A1(n5172), .A2(n5344), .ZN(n5174) );
  NAND2_X1 U6674 ( .A1(n5174), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5158) );
  XNOR2_X1 U6675 ( .A(n5158), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7090) );
  AOI22_X1 U6676 ( .A1(n5485), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5484), .B2(
        n7090), .ZN(n5159) );
  NAND2_X1 U6677 ( .A1(n5665), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6678 ( .A1(n6722), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6679 ( .A1(n5178), .A2(n5161), .ZN(n5162) );
  AND2_X1 U6680 ( .A1(n5163), .A2(n5162), .ZN(n7399) );
  NAND2_X1 U6681 ( .A1(n5537), .A2(n7399), .ZN(n5165) );
  NAND2_X1 U6682 ( .A1(n5241), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5164) );
  OR2_X1 U6683 ( .A1(n9732), .A2(n7582), .ZN(n8809) );
  NAND2_X1 U6684 ( .A1(n9732), .A2(n7582), .ZN(n8814) );
  OR2_X1 U6685 ( .A1(n5169), .A2(n5168), .ZN(n5170) );
  NAND2_X1 U6686 ( .A1(n5171), .A2(n5170), .ZN(n6703) );
  OR2_X1 U6687 ( .A1(n6703), .A2(n5209), .ZN(n5176) );
  OR2_X1 U6688 ( .A1(n5172), .A2(n5344), .ZN(n5173) );
  AOI22_X1 U6689 ( .A1(n5485), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5484), .B2(
        n7087), .ZN(n5175) );
  NAND2_X1 U6690 ( .A1(n5176), .A2(n5175), .ZN(n9653) );
  NAND2_X1 U6691 ( .A1(n5665), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6692 ( .A1(n5647), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5181) );
  OR2_X1 U6693 ( .A1(n5186), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5177) );
  AND2_X1 U6694 ( .A1(n5178), .A2(n5177), .ZN(n9650) );
  NAND2_X1 U6695 ( .A1(n5537), .A2(n9650), .ZN(n5180) );
  NAND2_X1 U6696 ( .A1(n6722), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6697 ( .A1(n9653), .A2(n9729), .ZN(n7388) );
  NAND2_X1 U6698 ( .A1(n9740), .A2(n9747), .ZN(n8819) );
  OAI21_X1 U6699 ( .B1(n5183), .B2(n8810), .A(n8819), .ZN(n5297) );
  NAND2_X1 U6700 ( .A1(n5647), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6701 ( .A1(n5665), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5189) );
  AND2_X1 U6702 ( .A1(n5280), .A2(n5184), .ZN(n5185) );
  NOR2_X1 U6703 ( .A1(n5186), .A2(n5185), .ZN(n7267) );
  NAND2_X1 U6704 ( .A1(n5537), .A2(n7267), .ZN(n5188) );
  NAND2_X1 U6705 ( .A1(n6722), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5187) );
  OR2_X1 U6706 ( .A1(n5192), .A2(n5191), .ZN(n5193) );
  NAND2_X1 U6707 ( .A1(n5194), .A2(n5193), .ZN(n6697) );
  OR2_X1 U6708 ( .A1(n6697), .A2(n5209), .ZN(n5198) );
  OR2_X1 U6709 ( .A1(n5195), .A2(n9452), .ZN(n5196) );
  XNOR2_X1 U6710 ( .A(n5196), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7084) );
  AOI22_X1 U6711 ( .A1(n5485), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5484), .B2(
        n7084), .ZN(n5197) );
  NAND2_X1 U6712 ( .A1(n5198), .A2(n5197), .ZN(n7268) );
  NAND2_X1 U6713 ( .A1(n7293), .A2(n7268), .ZN(n8806) );
  INV_X1 U6714 ( .A(n8806), .ZN(n8800) );
  OR2_X1 U6715 ( .A1(n5297), .A2(n8800), .ZN(n8996) );
  INV_X1 U6716 ( .A(n5199), .ZN(n5222) );
  NAND2_X1 U6717 ( .A1(n5222), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U6718 ( .A1(n5223), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6719 ( .A1(n5241), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5200) );
  OR2_X1 U6720 ( .A1(n8890), .A2(n5002), .ZN(n5214) );
  INV_X1 U6721 ( .A(n5204), .ZN(n5205) );
  NAND2_X1 U6722 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  AND2_X1 U6723 ( .A1(n5208), .A2(n5207), .ZN(n6073) );
  INV_X1 U6724 ( .A(n6073), .ZN(n6684) );
  OR2_X1 U6725 ( .A1(n5209), .A2(n6684), .ZN(n5212) );
  INV_X1 U6726 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6727 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5210) );
  XNOR2_X1 U6728 ( .A(n5211), .B(n5210), .ZN(n7073) );
  AND2_X1 U6729 ( .A1(n5212), .A2(n5084), .ZN(n5213) );
  NAND2_X2 U6730 ( .A1(n5214), .A2(n5213), .ZN(n5761) );
  NAND2_X1 U6731 ( .A1(n5222), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6732 ( .A1(n5223), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5215) );
  INV_X1 U6733 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U6734 ( .A1(n8014), .A2(SI_0_), .ZN(n5220) );
  XNOR2_X1 U6735 ( .A(n5220), .B(n5219), .ZN(n9459) );
  MUX2_X1 U6736 ( .A(n9072), .B(n9459), .S(n6707), .Z(n6889) );
  INV_X1 U6737 ( .A(n6884), .ZN(n6795) );
  NAND2_X1 U6738 ( .A1(n6795), .A2(n5761), .ZN(n5221) );
  NAND2_X1 U6739 ( .A1(n6875), .A2(n5221), .ZN(n6883) );
  NAND2_X1 U6740 ( .A1(n5222), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6741 ( .A1(n5223), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6742 ( .A1(n5226), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6743 ( .A1(n5241), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5227) );
  INV_X1 U6744 ( .A(n5779), .ZN(n5239) );
  NAND2_X1 U6745 ( .A1(n5232), .A2(n5231), .ZN(n5234) );
  AND2_X1 U6746 ( .A1(n5234), .A2(n5233), .ZN(n6100) );
  INV_X1 U6747 ( .A(n6100), .ZN(n6682) );
  OR2_X1 U6748 ( .A1(n5209), .A2(n6682), .ZN(n5238) );
  INV_X1 U6749 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6683) );
  OR2_X1 U6750 ( .A1(n8890), .A2(n6683), .ZN(n5237) );
  INV_X1 U6751 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5249) );
  OR2_X1 U6752 ( .A1(n6707), .A2(n7072), .ZN(n5236) );
  NAND2_X1 U6753 ( .A1(n5239), .A2(n6902), .ZN(n5674) );
  INV_X1 U6754 ( .A(n5674), .ZN(n5240) );
  NAND2_X1 U6755 ( .A1(n5779), .A2(n9691), .ZN(n8903) );
  NAND2_X1 U6756 ( .A1(n5665), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6757 ( .A1(n5241), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5243) );
  INV_X1 U6758 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6957) );
  OR2_X1 U6759 ( .A1(n5247), .A2(n5246), .ZN(n5248) );
  AND2_X1 U6760 ( .A1(n5263), .A2(n5248), .ZN(n6114) );
  INV_X1 U6761 ( .A(n6114), .ZN(n6686) );
  OR2_X1 U6762 ( .A1(n6686), .A2(n5209), .ZN(n5255) );
  INV_X1 U6763 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6687) );
  OR2_X1 U6764 ( .A1(n8890), .A2(n6687), .ZN(n5254) );
  NAND2_X1 U6765 ( .A1(n5272), .A2(n5249), .ZN(n5250) );
  NAND2_X1 U6766 ( .A1(n5250), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5252) );
  INV_X1 U6767 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5251) );
  XNOR2_X1 U6768 ( .A(n5252), .B(n5251), .ZN(n7076) );
  OR2_X1 U6769 ( .A1(n6707), .A2(n7076), .ZN(n5253) );
  NOR2_X1 U6770 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5256) );
  NOR2_X1 U6771 ( .A1(n5281), .A2(n5256), .ZN(n6987) );
  INV_X1 U6772 ( .A(n6987), .ZN(n5257) );
  NAND2_X1 U6773 ( .A1(n5226), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U6774 ( .A1(n5223), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6775 ( .A1(n5241), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6776 ( .A1(n5263), .A2(n5262), .ZN(n5267) );
  AND2_X1 U6777 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  NAND2_X1 U6778 ( .A1(n5267), .A2(n5266), .ZN(n5269) );
  OR2_X1 U6779 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  AND2_X1 U6780 ( .A1(n5269), .A2(n5268), .ZN(n6688) );
  NAND2_X1 U6781 ( .A1(n8888), .A2(n6688), .ZN(n5279) );
  OR2_X1 U6782 ( .A1(n5270), .A2(n9452), .ZN(n5271) );
  INV_X1 U6783 ( .A(n5275), .ZN(n5273) );
  NAND2_X1 U6784 ( .A1(n5273), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5276) );
  INV_X1 U6785 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6786 ( .A1(n5275), .A2(n5274), .ZN(n5287) );
  INV_X1 U6787 ( .A(n9549), .ZN(n6690) );
  OR2_X1 U6788 ( .A1(n6707), .A2(n6690), .ZN(n5278) );
  INV_X1 U6789 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6692) );
  OR2_X1 U6790 ( .A1(n8890), .A2(n6692), .ZN(n5277) );
  NAND2_X1 U6791 ( .A1(n9662), .A2(n9705), .ZN(n8904) );
  NAND2_X1 U6792 ( .A1(n6980), .A2(n8904), .ZN(n8797) );
  NAND2_X1 U6793 ( .A1(n8797), .A2(n8802), .ZN(n5296) );
  NAND2_X1 U6794 ( .A1(n5241), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6795 ( .A1(n5665), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5285) );
  OAI21_X1 U6796 ( .B1(n5281), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5280), .ZN(
        n7164) );
  INV_X1 U6797 ( .A(n7164), .ZN(n5282) );
  NAND2_X1 U6798 ( .A1(n5537), .A2(n5282), .ZN(n5284) );
  NAND2_X1 U6799 ( .A1(n6722), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5283) );
  INV_X1 U6800 ( .A(n9049), .ZN(n7262) );
  NAND2_X1 U6801 ( .A1(n5287), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5288) );
  XNOR2_X1 U6802 ( .A(n5288), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7082) );
  AOI22_X1 U6803 ( .A1(n5485), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5484), .B2(
        n7082), .ZN(n5294) );
  OR2_X1 U6804 ( .A1(n5290), .A2(n5289), .ZN(n5291) );
  NAND2_X1 U6805 ( .A1(n5292), .A2(n5291), .ZN(n6694) );
  OR2_X1 U6806 ( .A1(n6694), .A2(n5209), .ZN(n5293) );
  INV_X1 U6807 ( .A(n9713), .ZN(n7163) );
  NAND2_X1 U6808 ( .A1(n9049), .A2(n9713), .ZN(n8913) );
  INV_X1 U6809 ( .A(n8986), .ZN(n5295) );
  OR2_X1 U6810 ( .A1(n9653), .A2(n9729), .ZN(n8808) );
  OR2_X1 U6811 ( .A1(n7268), .A2(n7293), .ZN(n8799) );
  NAND3_X1 U6812 ( .A1(n8808), .A2(n8815), .A3(n8799), .ZN(n8994) );
  INV_X1 U6813 ( .A(n8994), .ZN(n5298) );
  OR2_X1 U6814 ( .A1(n5298), .A2(n5297), .ZN(n8917) );
  OAI21_X1 U6815 ( .B1(n8996), .B2(n7387), .A(n8917), .ZN(n7360) );
  INV_X1 U6816 ( .A(n5299), .ZN(n5300) );
  MUX2_X1 U6817 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n8014), .Z(n5304) );
  INV_X1 U6818 ( .A(n5304), .ZN(n5306) );
  INV_X1 U6819 ( .A(SI_10_), .ZN(n5305) );
  NAND2_X1 U6820 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  NAND2_X1 U6821 ( .A1(n5325), .A2(n5307), .ZN(n5310) );
  INV_X1 U6822 ( .A(n5309), .ZN(n5311) );
  NAND2_X1 U6823 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  NAND2_X1 U6824 ( .A1(n5326), .A2(n5312), .ZN(n6717) );
  OR2_X1 U6825 ( .A1(n6717), .A2(n5209), .ZN(n5318) );
  OR2_X1 U6826 ( .A1(n5313), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6827 ( .A1(n5314), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6828 ( .A1(n5315), .A2(n10274), .ZN(n5327) );
  OR2_X1 U6829 ( .A1(n5315), .A2(n10274), .ZN(n5316) );
  AOI22_X1 U6830 ( .A1(n5485), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5484), .B2(
        n9489), .ZN(n5317) );
  NAND2_X1 U6831 ( .A1(n5665), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6832 ( .A1(n5647), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5323) );
  NOR2_X1 U6833 ( .A1(n5319), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6834 ( .A1(n5537), .A2(n5080), .ZN(n5322) );
  NAND2_X1 U6835 ( .A1(n6722), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5321) );
  OR2_X1 U6836 ( .A1(n9751), .A2(n7704), .ZN(n8916) );
  NAND2_X1 U6837 ( .A1(n8916), .A2(n8820), .ZN(n8993) );
  MUX2_X1 U6838 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n8014), .Z(n5337) );
  XNOR2_X1 U6839 ( .A(n5339), .B(n5338), .ZN(n6738) );
  NAND2_X1 U6840 ( .A1(n6738), .A2(n8888), .ZN(n5330) );
  NAND2_X1 U6841 ( .A1(n5327), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5328) );
  XNOR2_X1 U6842 ( .A(n5328), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9585) );
  AOI22_X1 U6843 ( .A1(n5485), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5484), .B2(
        n9585), .ZN(n5329) );
  NAND2_X1 U6844 ( .A1(n5665), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6845 ( .A1(n6722), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5335) );
  OR2_X1 U6846 ( .A1(n5331), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5332) );
  AND2_X1 U6847 ( .A1(n5357), .A2(n5332), .ZN(n9635) );
  NAND2_X1 U6848 ( .A1(n5537), .A2(n9635), .ZN(n5334) );
  NAND2_X1 U6849 ( .A1(n5647), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5333) );
  OR2_X1 U6850 ( .A1(n9636), .A2(n9748), .ZN(n8826) );
  NAND2_X1 U6851 ( .A1(n9636), .A2(n9748), .ZN(n8827) );
  MUX2_X1 U6852 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n8014), .Z(n5340) );
  NAND2_X1 U6853 ( .A1(n5342), .A2(n5341), .ZN(n5343) );
  NAND2_X1 U6854 ( .A1(n5343), .A2(n5364), .ZN(n6743) );
  NOR2_X1 U6855 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5346) );
  NAND4_X1 U6856 ( .A1(n5346), .A2(n5345), .A3(n10274), .A4(n5344), .ZN(n5347)
         );
  OR2_X1 U6857 ( .A1(n5348), .A2(n5347), .ZN(n5350) );
  NAND2_X1 U6858 ( .A1(n5350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5349) );
  MUX2_X1 U6859 ( .A(n5349), .B(P1_IR_REG_31__SCAN_IN), .S(n5351), .Z(n5353)
         );
  INV_X1 U6860 ( .A(n5350), .ZN(n5352) );
  NAND2_X1 U6861 ( .A1(n5352), .A2(n5351), .ZN(n5373) );
  NAND2_X1 U6862 ( .A1(n5353), .A2(n5373), .ZN(n7097) );
  INV_X1 U6863 ( .A(n7097), .ZN(n7246) );
  AOI22_X1 U6864 ( .A1(n5485), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5484), .B2(
        n7246), .ZN(n5354) );
  NAND2_X1 U6865 ( .A1(n5665), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6866 ( .A1(n6722), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5361) );
  INV_X1 U6867 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6868 ( .A1(n5357), .A2(n5356), .ZN(n5358) );
  AND2_X1 U6869 ( .A1(n5377), .A2(n5358), .ZN(n7763) );
  NAND2_X1 U6870 ( .A1(n5537), .A2(n7763), .ZN(n5360) );
  NAND2_X1 U6871 ( .A1(n5647), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5359) );
  OR2_X1 U6872 ( .A1(n7469), .A2(n9611), .ZN(n8831) );
  MUX2_X1 U6873 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n8014), .Z(n5365) );
  INV_X1 U6874 ( .A(n5365), .ZN(n5367) );
  INV_X1 U6875 ( .A(SI_13_), .ZN(n5366) );
  NAND2_X1 U6876 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  OR2_X1 U6877 ( .A1(n5370), .A2(n5369), .ZN(n5371) );
  NAND2_X1 U6878 ( .A1(n5384), .A2(n5371), .ZN(n6781) );
  NAND2_X1 U6879 ( .A1(n5373), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5372) );
  MUX2_X1 U6880 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5372), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n5374) );
  OR2_X1 U6881 ( .A1(n5373), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5386) );
  AOI22_X1 U6882 ( .A1(n5485), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5484), .B2(
        n7312), .ZN(n5375) );
  NAND2_X1 U6883 ( .A1(n5665), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6884 ( .A1(n6722), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5381) );
  INV_X1 U6885 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7250) );
  NAND2_X1 U6886 ( .A1(n5377), .A2(n7250), .ZN(n5378) );
  AND2_X1 U6887 ( .A1(n5392), .A2(n5378), .ZN(n9615) );
  NAND2_X1 U6888 ( .A1(n5537), .A2(n9615), .ZN(n5380) );
  NAND2_X1 U6889 ( .A1(n5647), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6890 ( .A1(n9616), .A2(n9788), .ZN(n8847) );
  AND2_X1 U6891 ( .A1(n8847), .A2(n9606), .ZN(n8928) );
  MUX2_X1 U6892 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7856), .Z(n5399) );
  XNOR2_X1 U6893 ( .A(n5399), .B(SI_14_), .ZN(n5385) );
  XNOR2_X1 U6894 ( .A(n5400), .B(n5385), .ZN(n6927) );
  NAND2_X1 U6895 ( .A1(n6927), .A2(n8888), .ZN(n5391) );
  NAND2_X1 U6896 ( .A1(n5386), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5388) );
  INV_X1 U6897 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6898 ( .A1(n5388), .A2(n5387), .ZN(n5404) );
  OR2_X1 U6899 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  AOI22_X1 U6900 ( .A1(n5485), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5484), .B2(
        n7630), .ZN(n5390) );
  NAND2_X1 U6901 ( .A1(n5647), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6902 ( .A1(n5665), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5396) );
  INV_X1 U6903 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7316) );
  AND2_X1 U6904 ( .A1(n5392), .A2(n7316), .ZN(n5393) );
  NOR2_X1 U6905 ( .A1(n5410), .A2(n5393), .ZN(n8662) );
  NAND2_X1 U6906 ( .A1(n5537), .A2(n8662), .ZN(n5395) );
  NAND2_X1 U6907 ( .A1(n6722), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5394) );
  OR2_X1 U6908 ( .A1(n9793), .A2(n9612), .ZN(n8850) );
  NAND2_X1 U6909 ( .A1(n9793), .A2(n9612), .ZN(n8846) );
  NAND2_X1 U6910 ( .A1(n8850), .A2(n8846), .ZN(n9001) );
  INV_X1 U6911 ( .A(n9001), .ZN(n5398) );
  NAND2_X1 U6912 ( .A1(n7693), .A2(n8846), .ZN(n7799) );
  NAND2_X1 U6913 ( .A1(n5402), .A2(n5401), .ZN(n5416) );
  MUX2_X1 U6914 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7856), .Z(n5417) );
  XNOR2_X1 U6915 ( .A(n5417), .B(SI_15_), .ZN(n5403) );
  XNOR2_X1 U6916 ( .A(n5416), .B(n5403), .ZN(n7009) );
  NAND2_X1 U6917 ( .A1(n7009), .A2(n8888), .ZN(n5409) );
  NAND2_X1 U6918 ( .A1(n5404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5406) );
  XNOR2_X1 U6919 ( .A(n5406), .B(n5405), .ZN(n7716) );
  INV_X1 U6920 ( .A(n7716), .ZN(n5407) );
  AOI22_X1 U6921 ( .A1(n5485), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5484), .B2(
        n5407), .ZN(n5408) );
  NAND2_X1 U6922 ( .A1(n5665), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6923 ( .A1(n5647), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5414) );
  OR2_X1 U6924 ( .A1(n5410), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6925 ( .A1(n5410), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5425) );
  AND2_X1 U6926 ( .A1(n5411), .A2(n5425), .ZN(n8783) );
  NAND2_X1 U6927 ( .A1(n5537), .A2(n8783), .ZN(n5413) );
  NAND2_X1 U6928 ( .A1(n6722), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5412) );
  NAND4_X1 U6929 ( .A1(n5415), .A2(n5414), .A3(n5413), .A4(n5412), .ZN(n9046)
         );
  AND2_X1 U6930 ( .A1(n9532), .A2(n9046), .ZN(n5431) );
  INV_X1 U6931 ( .A(n5431), .ZN(n8849) );
  INV_X1 U6932 ( .A(n9532), .ZN(n5681) );
  NAND2_X1 U6933 ( .A1(n5681), .A2(n9790), .ZN(n8852) );
  NAND2_X1 U6934 ( .A1(n8849), .A2(n8852), .ZN(n9002) );
  INV_X1 U6935 ( .A(n5417), .ZN(n5418) );
  MUX2_X1 U6936 ( .A(n7102), .B(n7104), .S(n7856), .Z(n5433) );
  XNOR2_X1 U6937 ( .A(n5433), .B(SI_16_), .ZN(n5419) );
  XNOR2_X1 U6938 ( .A(n5437), .B(n5419), .ZN(n7101) );
  NAND2_X1 U6939 ( .A1(n7101), .A2(n8888), .ZN(n5424) );
  NAND2_X1 U6940 ( .A1(n5420), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5421) );
  MUX2_X1 U6941 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5421), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n5422) );
  AND2_X1 U6942 ( .A1(n5422), .A2(n5443), .ZN(n7776) );
  AOI22_X1 U6943 ( .A1(n5485), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5484), .B2(
        n7776), .ZN(n5423) );
  INV_X1 U6944 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U6945 ( .A1(n5425), .A2(n7723), .ZN(n5426) );
  AND2_X1 U6946 ( .A1(n5447), .A2(n5426), .ZN(n8709) );
  NAND2_X1 U6947 ( .A1(n5537), .A2(n8709), .ZN(n5430) );
  NAND2_X1 U6948 ( .A1(n5665), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U6949 ( .A1(n6722), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6950 ( .A1(n5647), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5427) );
  OR2_X1 U6951 ( .A1(n9431), .A2(n9329), .ZN(n8855) );
  NAND2_X1 U6952 ( .A1(n9431), .A2(n9329), .ZN(n8853) );
  NAND2_X1 U6953 ( .A1(n8855), .A2(n8853), .ZN(n9004) );
  NAND2_X1 U6954 ( .A1(n8853), .A2(n5431), .ZN(n5432) );
  AND2_X1 U6955 ( .A1(n5432), .A2(n8855), .ZN(n8929) );
  NOR2_X1 U6956 ( .A1(n5434), .A2(SI_16_), .ZN(n5436) );
  NAND2_X1 U6957 ( .A1(n5434), .A2(SI_16_), .ZN(n5435) );
  INV_X1 U6958 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7260) );
  INV_X1 U6959 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7258) );
  MUX2_X1 U6960 ( .A(n7260), .B(n7258), .S(n8014), .Z(n5439) );
  INV_X1 U6961 ( .A(SI_17_), .ZN(n5438) );
  NAND2_X1 U6962 ( .A1(n5439), .A2(n5438), .ZN(n5472) );
  INV_X1 U6963 ( .A(n5439), .ZN(n5440) );
  NAND2_X1 U6964 ( .A1(n5440), .A2(SI_17_), .ZN(n5441) );
  NAND2_X1 U6965 ( .A1(n5472), .A2(n5441), .ZN(n5471) );
  XNOR2_X1 U6966 ( .A(n5500), .B(n5471), .ZN(n7257) );
  NAND2_X1 U6967 ( .A1(n7257), .A2(n8888), .ZN(n5446) );
  NAND2_X1 U6968 ( .A1(n5443), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5442) );
  MUX2_X1 U6969 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5442), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n5444) );
  NAND2_X1 U6970 ( .A1(n5444), .A2(n5456), .ZN(n7783) );
  INV_X1 U6971 ( .A(n7783), .ZN(n7877) );
  AOI22_X1 U6972 ( .A1(n5485), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5484), .B2(
        n7877), .ZN(n5445) );
  INV_X1 U6973 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7780) );
  AND2_X1 U6974 ( .A1(n5447), .A2(n7780), .ZN(n5448) );
  OR2_X1 U6975 ( .A1(n5448), .A2(n5462), .ZN(n8717) );
  NAND2_X1 U6976 ( .A1(n5665), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6977 ( .A1(n6722), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5449) );
  AND2_X1 U6978 ( .A1(n5450), .A2(n5449), .ZN(n5452) );
  NAND2_X1 U6979 ( .A1(n5647), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5451) );
  OAI211_X1 U6980 ( .C1(n8717), .C2(n5199), .A(n5452), .B(n5451), .ZN(n9044)
         );
  NAND2_X1 U6981 ( .A1(n9426), .A2(n9418), .ZN(n8857) );
  INV_X1 U6982 ( .A(n9317), .ZN(n9327) );
  INV_X1 U6983 ( .A(n9298), .ZN(n5467) );
  OR2_X1 U6984 ( .A1(n5500), .A2(n5471), .ZN(n5453) );
  NAND2_X1 U6985 ( .A1(n5453), .A2(n5472), .ZN(n5455) );
  INV_X1 U6986 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7300) );
  INV_X1 U6987 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5454) );
  MUX2_X1 U6988 ( .A(n7300), .B(n5454), .S(n8014), .Z(n5469) );
  XNOR2_X1 U6989 ( .A(n5469), .B(SI_18_), .ZN(n5473) );
  NAND2_X1 U6990 ( .A1(n7285), .A2(n8888), .ZN(n5461) );
  INV_X1 U6991 ( .A(n5458), .ZN(n5457) );
  NAND2_X1 U6992 ( .A1(n5457), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U6993 ( .A1(n5458), .A2(n5656), .ZN(n5482) );
  AND2_X1 U6994 ( .A1(n5459), .A2(n5482), .ZN(n9121) );
  AOI22_X1 U6995 ( .A1(n5485), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5484), .B2(
        n9121), .ZN(n5460) );
  OR2_X1 U6996 ( .A1(n5462), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5463) );
  AND2_X1 U6997 ( .A1(n5463), .A2(n5488), .ZN(n9305) );
  NAND2_X1 U6998 ( .A1(n9305), .A2(n5537), .ZN(n5466) );
  AOI22_X1 U6999 ( .A1(n5647), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n5665), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U7000 ( .A1(n6722), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5464) );
  OR2_X1 U7001 ( .A1(n9421), .A2(n9330), .ZN(n8843) );
  NAND2_X1 U7002 ( .A1(n9421), .A2(n9330), .ZN(n8858) );
  NAND2_X1 U7003 ( .A1(n8843), .A2(n8858), .ZN(n9302) );
  INV_X1 U7004 ( .A(n8858), .ZN(n5468) );
  INV_X1 U7005 ( .A(n5469), .ZN(n5470) );
  OR2_X1 U7006 ( .A1(n5500), .A2(n5493), .ZN(n5476) );
  MUX2_X1 U7007 ( .A(n7305), .B(n7307), .S(n7856), .Z(n5478) );
  INV_X1 U7008 ( .A(SI_19_), .ZN(n5477) );
  NAND2_X1 U7009 ( .A1(n5478), .A2(n5477), .ZN(n5496) );
  INV_X1 U7010 ( .A(n5478), .ZN(n5479) );
  NAND2_X1 U7011 ( .A1(n5479), .A2(SI_19_), .ZN(n5480) );
  NAND2_X1 U7012 ( .A1(n7304), .A2(n8888), .ZN(n5487) );
  AOI22_X1 U7013 ( .A1(n5485), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9021), .B2(
        n5484), .ZN(n5486) );
  NAND2_X1 U7014 ( .A1(n5665), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7015 ( .A1(n5647), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5491) );
  INV_X1 U7016 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7885) );
  AOI21_X1 U7017 ( .B1(n7885), .B2(n5488), .A(n5504), .ZN(n9292) );
  NAND2_X1 U7018 ( .A1(n5537), .A2(n9292), .ZN(n5490) );
  NAND2_X1 U7019 ( .A1(n6722), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U7020 ( .A1(n9413), .A2(n9417), .ZN(n8902) );
  NAND2_X1 U7021 ( .A1(n9287), .A2(n9286), .ZN(n9285) );
  INV_X1 U7022 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10317) );
  INV_X1 U7023 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7299) );
  MUX2_X1 U7024 ( .A(n10317), .B(n7299), .S(n7856), .Z(n5509) );
  XNOR2_X1 U7025 ( .A(n5509), .B(SI_20_), .ZN(n5501) );
  XNOR2_X1 U7026 ( .A(n5511), .B(n5501), .ZN(n7302) );
  NAND2_X1 U7027 ( .A1(n7302), .A2(n8888), .ZN(n5503) );
  OR2_X1 U7028 ( .A1(n8890), .A2(n7299), .ZN(n5502) );
  NAND2_X1 U7029 ( .A1(n5647), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U7030 ( .A1(n5665), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7031 ( .A1(n5504), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5518) );
  OAI21_X1 U7032 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n5504), .A(n5518), .ZN(
        n8738) );
  INV_X1 U7033 ( .A(n8738), .ZN(n9271) );
  NAND2_X1 U7034 ( .A1(n5537), .A2(n9271), .ZN(n5506) );
  NAND2_X1 U7035 ( .A1(n6722), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7036 ( .A1(n9406), .A2(n9288), .ZN(n8839) );
  NAND2_X1 U7037 ( .A1(n8863), .A2(n8839), .ZN(n9275) );
  INV_X1 U7038 ( .A(SI_20_), .ZN(n5510) );
  NAND2_X1 U7039 ( .A1(n5511), .A2(n5510), .ZN(n5512) );
  MUX2_X1 U7040 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7856), .Z(n5525) );
  INV_X1 U7041 ( .A(SI_21_), .ZN(n5514) );
  XNOR2_X1 U7042 ( .A(n5525), .B(n5514), .ZN(n5515) );
  XNOR2_X1 U7043 ( .A(n5528), .B(n5515), .ZN(n7394) );
  NAND2_X1 U7044 ( .A1(n7394), .A2(n8888), .ZN(n5517) );
  INV_X1 U7045 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7422) );
  OR2_X1 U7046 ( .A1(n8890), .A2(n7422), .ZN(n5516) );
  NAND2_X1 U7047 ( .A1(n5665), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7048 ( .A1(n5647), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5523) );
  NOR2_X1 U7049 ( .A1(P1_REG3_REG_21__SCAN_IN), .A2(n5519), .ZN(n5520) );
  NOR2_X1 U7050 ( .A1(n5535), .A2(n5520), .ZN(n9258) );
  NAND2_X1 U7051 ( .A1(n5537), .A2(n9258), .ZN(n5522) );
  NAND2_X1 U7052 ( .A1(n6722), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5521) );
  INV_X1 U7053 ( .A(n9277), .ZN(n9389) );
  XNOR2_X1 U7054 ( .A(n9262), .B(n9389), .ZN(n9254) );
  NAND2_X1 U7055 ( .A1(n9262), .A2(n9277), .ZN(n8865) );
  NOR2_X1 U7056 ( .A1(n5525), .A2(SI_21_), .ZN(n5527) );
  NAND2_X1 U7057 ( .A1(n5525), .A2(SI_21_), .ZN(n5526) );
  INV_X1 U7058 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7541) );
  MUX2_X1 U7059 ( .A(n7541), .B(n10379), .S(n7856), .Z(n5530) );
  INV_X1 U7060 ( .A(SI_22_), .ZN(n5529) );
  NAND2_X1 U7061 ( .A1(n5530), .A2(n5529), .ZN(n5543) );
  INV_X1 U7062 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U7063 ( .A1(n5531), .A2(SI_22_), .ZN(n5532) );
  NAND2_X1 U7064 ( .A1(n5543), .A2(n5532), .ZN(n5544) );
  XNOR2_X1 U7065 ( .A(n5545), .B(n5544), .ZN(n7539) );
  NAND2_X1 U7066 ( .A1(n7539), .A2(n8888), .ZN(n5534) );
  OR2_X1 U7067 ( .A1(n8890), .A2(n10379), .ZN(n5533) );
  NAND2_X1 U7068 ( .A1(n5665), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7069 ( .A1(n5647), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5540) );
  NOR2_X1 U7070 ( .A1(n5535), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5536) );
  NOR2_X1 U7071 ( .A1(n5553), .A2(n5536), .ZN(n8748) );
  NAND2_X1 U7072 ( .A1(n5537), .A2(n8748), .ZN(n5539) );
  NAND2_X1 U7073 ( .A1(n6722), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5538) );
  OR2_X1 U7074 ( .A1(n9248), .A2(n9381), .ZN(n8794) );
  NAND2_X1 U7075 ( .A1(n9248), .A2(n9381), .ZN(n8793) );
  NAND2_X1 U7076 ( .A1(n8794), .A2(n8793), .ZN(n9236) );
  INV_X1 U7077 ( .A(n9236), .ZN(n9238) );
  INV_X1 U7078 ( .A(n8793), .ZN(n5542) );
  INV_X1 U7079 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5546) );
  INV_X1 U7080 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7573) );
  MUX2_X1 U7081 ( .A(n5546), .B(n7573), .S(n7856), .Z(n5548) );
  INV_X1 U7082 ( .A(SI_23_), .ZN(n5547) );
  NAND2_X1 U7083 ( .A1(n5548), .A2(n5547), .ZN(n5561) );
  INV_X1 U7084 ( .A(n5548), .ZN(n5549) );
  NAND2_X1 U7085 ( .A1(n5549), .A2(SI_23_), .ZN(n5550) );
  XNOR2_X1 U7086 ( .A(n5560), .B(n5559), .ZN(n7571) );
  NAND2_X1 U7087 ( .A1(n7571), .A2(n8888), .ZN(n5552) );
  OR2_X1 U7088 ( .A1(n8890), .A2(n7573), .ZN(n5551) );
  NAND2_X1 U7089 ( .A1(n5665), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7090 ( .A1(n6722), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5557) );
  NOR2_X1 U7091 ( .A1(n5553), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5554) );
  NOR2_X1 U7092 ( .A1(n5569), .A2(n5554), .ZN(n9229) );
  NAND2_X1 U7093 ( .A1(n5537), .A2(n9229), .ZN(n5556) );
  NAND2_X1 U7094 ( .A1(n5647), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5555) );
  OR2_X1 U7095 ( .A1(n9384), .A2(n9216), .ZN(n8866) );
  NAND2_X1 U7096 ( .A1(n9384), .A2(n9216), .ZN(n8936) );
  NOR2_X1 U7097 ( .A1(n9223), .A2(n9224), .ZN(n9213) );
  INV_X1 U7098 ( .A(n8936), .ZN(n9215) );
  INV_X1 U7099 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7662) );
  INV_X1 U7100 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7675) );
  MUX2_X1 U7101 ( .A(n7662), .B(n7675), .S(n7856), .Z(n5564) );
  INV_X1 U7102 ( .A(SI_24_), .ZN(n5563) );
  NAND2_X1 U7103 ( .A1(n5564), .A2(n5563), .ZN(n5576) );
  INV_X1 U7104 ( .A(n5564), .ZN(n5565) );
  NAND2_X1 U7105 ( .A1(n5565), .A2(SI_24_), .ZN(n5566) );
  XNOR2_X1 U7106 ( .A(n5575), .B(n5574), .ZN(n7661) );
  NAND2_X1 U7107 ( .A1(n7661), .A2(n8888), .ZN(n5568) );
  OR2_X1 U7108 ( .A1(n8890), .A2(n7675), .ZN(n5567) );
  NAND2_X1 U7109 ( .A1(n5665), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7110 ( .A1(n6722), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5572) );
  OAI21_X1 U7111 ( .B1(n5569), .B2(P1_REG3_REG_24__SCAN_IN), .A(n5583), .ZN(
        n8725) );
  INV_X1 U7112 ( .A(n8725), .ZN(n9209) );
  NAND2_X1 U7113 ( .A1(n5537), .A2(n9209), .ZN(n5571) );
  NAND2_X1 U7114 ( .A1(n5647), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7115 ( .A1(n9375), .A2(n9380), .ZN(n8939) );
  INV_X1 U7116 ( .A(n9191), .ZN(n5589) );
  INV_X1 U7117 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7731) );
  INV_X1 U7118 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7752) );
  MUX2_X1 U7119 ( .A(n7731), .B(n7752), .S(n7856), .Z(n5578) );
  INV_X1 U7120 ( .A(SI_25_), .ZN(n5577) );
  NAND2_X1 U7121 ( .A1(n5578), .A2(n5577), .ZN(n5593) );
  INV_X1 U7122 ( .A(n5578), .ZN(n5579) );
  NAND2_X1 U7123 ( .A1(n5579), .A2(SI_25_), .ZN(n5580) );
  NAND2_X1 U7124 ( .A1(n7730), .A2(n8888), .ZN(n5582) );
  OR2_X1 U7125 ( .A1(n8890), .A2(n7752), .ZN(n5581) );
  NAND2_X1 U7126 ( .A1(n5665), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7127 ( .A1(n6722), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5587) );
  INV_X1 U7128 ( .A(n5600), .ZN(n5602) );
  OAI21_X1 U7129 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n5584), .A(n5602), .ZN(
        n8698) );
  INV_X1 U7130 ( .A(n8698), .ZN(n9196) );
  NAND2_X1 U7131 ( .A1(n5537), .A2(n9196), .ZN(n5586) );
  NAND2_X1 U7132 ( .A1(n5647), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5585) );
  OR2_X1 U7133 ( .A1(n9370), .A2(n9358), .ZN(n8872) );
  NAND2_X1 U7134 ( .A1(n9370), .A2(n9358), .ZN(n8949) );
  NAND2_X1 U7135 ( .A1(n8872), .A2(n8949), .ZN(n9193) );
  INV_X1 U7136 ( .A(n8949), .ZN(n5590) );
  INV_X1 U7137 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10369) );
  INV_X1 U7138 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7768) );
  MUX2_X1 U7139 ( .A(n10369), .B(n7768), .S(n7856), .Z(n5595) );
  INV_X1 U7140 ( .A(SI_26_), .ZN(n5594) );
  NAND2_X1 U7141 ( .A1(n5595), .A2(n5594), .ZN(n5628) );
  INV_X1 U7142 ( .A(n5595), .ZN(n5596) );
  NAND2_X1 U7143 ( .A1(n5596), .A2(SI_26_), .ZN(n5597) );
  NAND2_X1 U7144 ( .A1(n7766), .A2(n8888), .ZN(n5599) );
  OR2_X1 U7145 ( .A1(n8890), .A2(n7768), .ZN(n5598) );
  NAND2_X1 U7146 ( .A1(n5665), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U7147 ( .A1(n6722), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5606) );
  INV_X1 U7148 ( .A(n5618), .ZN(n5620) );
  INV_X1 U7149 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U7150 ( .A1(n5602), .A2(n5601), .ZN(n5603) );
  NAND2_X1 U7151 ( .A1(n5537), .A2(n9184), .ZN(n5605) );
  NAND2_X1 U7152 ( .A1(n5647), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5604) );
  XNOR2_X1 U7153 ( .A(n9362), .B(n9367), .ZN(n9179) );
  NAND2_X1 U7154 ( .A1(n9362), .A2(n9367), .ZN(n9163) );
  INV_X1 U7155 ( .A(n9163), .ZN(n5626) );
  NAND2_X1 U7156 ( .A1(n5630), .A2(n5628), .ZN(n5615) );
  INV_X1 U7157 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5610) );
  INV_X1 U7158 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7869) );
  MUX2_X1 U7159 ( .A(n5610), .B(n7869), .S(n7856), .Z(n5612) );
  INV_X1 U7160 ( .A(SI_27_), .ZN(n5611) );
  NAND2_X1 U7161 ( .A1(n5612), .A2(n5611), .ZN(n5627) );
  INV_X1 U7162 ( .A(n5612), .ZN(n5613) );
  NAND2_X1 U7163 ( .A1(n5613), .A2(SI_27_), .ZN(n5631) );
  AND2_X1 U7164 ( .A1(n5627), .A2(n5631), .ZN(n5614) );
  NAND2_X1 U7165 ( .A1(n7787), .A2(n8888), .ZN(n5617) );
  OR2_X1 U7166 ( .A1(n8890), .A2(n7869), .ZN(n5616) );
  NAND2_X1 U7167 ( .A1(n5665), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7168 ( .A1(n5647), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U7169 ( .A1(n5618), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5649) );
  INV_X1 U7170 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7171 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  NAND2_X1 U7172 ( .A1(n5537), .A2(n9168), .ZN(n5623) );
  NAND2_X1 U7173 ( .A1(n6722), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5622) );
  NAND4_X1 U7174 ( .A1(n5625), .A2(n5624), .A3(n5623), .A4(n5622), .ZN(n9183)
         );
  NAND2_X1 U7175 ( .A1(n9352), .A2(n9359), .ZN(n9145) );
  AND2_X1 U7176 ( .A1(n5628), .A2(n5627), .ZN(n5629) );
  INV_X1 U7177 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5632) );
  INV_X1 U7178 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10378) );
  MUX2_X1 U7179 ( .A(n5632), .B(n10378), .S(n7856), .Z(n5643) );
  XNOR2_X1 U7180 ( .A(n5643), .B(SI_28_), .ZN(n5640) );
  NAND2_X1 U7181 ( .A1(n7808), .A2(n8888), .ZN(n5634) );
  OR2_X1 U7182 ( .A1(n8890), .A2(n10378), .ZN(n5633) );
  NAND2_X1 U7183 ( .A1(n5665), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7184 ( .A1(n5647), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5637) );
  XNOR2_X1 U7185 ( .A(n5649), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9151) );
  NAND2_X1 U7186 ( .A1(n5537), .A2(n9151), .ZN(n5636) );
  NAND2_X1 U7187 ( .A1(n6722), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5635) );
  NAND4_X1 U7188 ( .A1(n5638), .A2(n5637), .A3(n5636), .A4(n5635), .ZN(n9171)
         );
  NAND2_X1 U7189 ( .A1(n9152), .A2(n9349), .ZN(n8876) );
  AND2_X1 U7190 ( .A1(n8876), .A2(n9145), .ZN(n8960) );
  INV_X1 U7191 ( .A(n8961), .ZN(n5639) );
  AOI21_X1 U7192 ( .B1(n9165), .B2(n8960), .A(n5639), .ZN(n5654) );
  INV_X1 U7193 ( .A(SI_28_), .ZN(n5642) );
  NAND2_X1 U7194 ( .A1(n5643), .A2(n5642), .ZN(n5644) );
  INV_X1 U7195 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10301) );
  INV_X1 U7196 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10361) );
  MUX2_X1 U7197 ( .A(n10301), .B(n10361), .S(n7856), .Z(n7852) );
  XNOR2_X2 U7198 ( .A(n7851), .B(SI_29_), .ZN(n7848) );
  NOR2_X1 U7199 ( .A1(n8890), .A2(n10361), .ZN(n5646) );
  AOI21_X2 U7200 ( .B1(n7848), .B2(n8888), .A(n5646), .ZN(n9142) );
  NAND2_X1 U7201 ( .A1(n5665), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7202 ( .A1(n5647), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5652) );
  INV_X1 U7203 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5648) );
  NOR2_X1 U7204 ( .A1(n5649), .A2(n5648), .ZN(n9139) );
  NAND2_X1 U7205 ( .A1(n5537), .A2(n9139), .ZN(n5651) );
  NAND2_X1 U7206 ( .A1(n6722), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5650) );
  NAND4_X1 U7207 ( .A1(n5653), .A2(n5652), .A3(n5651), .A4(n5650), .ZN(n9041)
         );
  AND2_X1 U7208 ( .A1(n9142), .A2(n9041), .ZN(n8882) );
  INV_X1 U7209 ( .A(n9041), .ZN(n9148) );
  XNOR2_X1 U7210 ( .A(n5654), .B(n8984), .ZN(n5672) );
  INV_X1 U7211 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7212 ( .A1(n5082), .A2(n4759), .ZN(n5661) );
  INV_X1 U7213 ( .A(n5661), .ZN(n5659) );
  INV_X1 U7214 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7215 ( .A1(n5659), .A2(n5658), .ZN(n5660) );
  OR2_X1 U7216 ( .A1(n7542), .A2(n5702), .ZN(n5663) );
  NAND2_X1 U7217 ( .A1(n5661), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7218 ( .A1(n8988), .A2(n5701), .ZN(n9032) );
  NAND2_X1 U7219 ( .A1(n5663), .A2(n9032), .ZN(n9777) );
  INV_X1 U7220 ( .A(n7542), .ZN(n9033) );
  AND2_X1 U7221 ( .A1(n9033), .A2(n8988), .ZN(n9017) );
  INV_X1 U7222 ( .A(n9017), .ZN(n5997) );
  NAND2_X1 U7223 ( .A1(n5647), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7224 ( .A1(n5665), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U7225 ( .A1(n6722), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5666) );
  AND3_X1 U7226 ( .A1(n5668), .A2(n5667), .A3(n5666), .ZN(n8965) );
  NAND2_X1 U7227 ( .A1(n4502), .A2(n9017), .ZN(n9789) );
  INV_X1 U7228 ( .A(P1_B_REG_SCAN_IN), .ZN(n5725) );
  NOR2_X1 U7229 ( .A1(n7867), .A2(n5725), .ZN(n5670) );
  OR2_X1 U7230 ( .A1(n9789), .A2(n5670), .ZN(n9127) );
  OAI22_X1 U7231 ( .A1(n9349), .A2(n9787), .B1(n8965), .B2(n9127), .ZN(n5671)
         );
  AOI21_X1 U7232 ( .B1(n5672), .B2(n9777), .A(n5671), .ZN(n9136) );
  INV_X1 U7233 ( .A(n9793), .ZN(n8665) );
  INV_X1 U7234 ( .A(n9612), .ZN(n9047) );
  INV_X1 U7235 ( .A(n6889), .ZN(n9683) );
  AND2_X1 U7236 ( .A1(n6712), .A2(n9683), .ZN(n6873) );
  INV_X1 U7237 ( .A(n5761), .ZN(n8905) );
  NAND2_X1 U7238 ( .A1(n6795), .A2(n8905), .ZN(n5673) );
  NAND2_X1 U7239 ( .A1(n6888), .A2(n8987), .ZN(n5676) );
  NAND2_X1 U7240 ( .A1(n5239), .A2(n9691), .ZN(n5675) );
  NOR2_X1 U7241 ( .A1(n9050), .A2(n6958), .ZN(n5679) );
  INV_X1 U7242 ( .A(n7293), .ZN(n9646) );
  INV_X1 U7243 ( .A(n9653), .ZN(n9723) );
  INV_X1 U7244 ( .A(n7582), .ZN(n9739) );
  NAND2_X1 U7245 ( .A1(n8824), .A2(n8819), .ZN(n7390) );
  INV_X1 U7246 ( .A(n8993), .ZN(n7361) );
  INV_X1 U7247 ( .A(n7704), .ZN(n9629) );
  INV_X1 U7248 ( .A(n9636), .ZN(n9759) );
  INV_X1 U7249 ( .A(n9611), .ZN(n9630) );
  NAND2_X1 U7250 ( .A1(n9609), .A2(n8847), .ZN(n9617) );
  INV_X1 U7251 ( .A(n9616), .ZN(n9782) );
  OAI21_X1 U7252 ( .B1(n9046), .B2(n5681), .A(n7802), .ZN(n5683) );
  NAND2_X1 U7253 ( .A1(n5681), .A2(n9046), .ZN(n5682) );
  INV_X1 U7254 ( .A(n9329), .ZN(n9045) );
  INV_X1 U7255 ( .A(n9426), .ZN(n9325) );
  NAND2_X1 U7256 ( .A1(n9325), .A2(n9418), .ZN(n5685) );
  INV_X1 U7257 ( .A(n9330), .ZN(n9043) );
  INV_X1 U7258 ( .A(n9421), .ZN(n9312) );
  NAND2_X1 U7259 ( .A1(n4657), .A2(n9417), .ZN(n5686) );
  NAND2_X1 U7260 ( .A1(n9284), .A2(n5686), .ZN(n5688) );
  INV_X1 U7261 ( .A(n9417), .ZN(n9309) );
  NAND2_X1 U7262 ( .A1(n9413), .A2(n9309), .ZN(n5687) );
  NAND2_X1 U7263 ( .A1(n5688), .A2(n5687), .ZN(n9268) );
  INV_X1 U7264 ( .A(n9406), .ZN(n9273) );
  INV_X1 U7265 ( .A(n9288), .ZN(n9398) );
  NOR2_X1 U7266 ( .A1(n9262), .A2(n9389), .ZN(n5691) );
  INV_X1 U7267 ( .A(n9262), .ZN(n9401) );
  INV_X1 U7268 ( .A(n9248), .ZN(n9392) );
  NOR2_X1 U7269 ( .A1(n9392), .A2(n9381), .ZN(n5692) );
  INV_X1 U7270 ( .A(n9381), .ZN(n9397) );
  INV_X1 U7271 ( .A(n9216), .ZN(n9388) );
  INV_X1 U7272 ( .A(n9384), .ZN(n9227) );
  INV_X1 U7273 ( .A(n9375), .ZN(n9211) );
  NOR2_X1 U7274 ( .A1(n9211), .A2(n9380), .ZN(n5693) );
  INV_X1 U7275 ( .A(n9358), .ZN(n9042) );
  NAND2_X1 U7276 ( .A1(n9370), .A2(n9042), .ZN(n5694) );
  NOR2_X1 U7277 ( .A1(n5696), .A2(n9367), .ZN(n5698) );
  INV_X1 U7278 ( .A(n9367), .ZN(n9199) );
  INV_X1 U7279 ( .A(n9352), .ZN(n9174) );
  NAND2_X1 U7280 ( .A1(n8961), .A2(n8876), .ZN(n9156) );
  NAND2_X1 U7281 ( .A1(n9157), .A2(n9156), .ZN(n9158) );
  NAND2_X1 U7282 ( .A1(n9158), .A2(n5699), .ZN(n5700) );
  AND2_X1 U7283 ( .A1(n9017), .A2(n5750), .ZN(n9025) );
  INV_X1 U7284 ( .A(n8988), .ZN(n7420) );
  NAND2_X1 U7285 ( .A1(n7542), .A2(n7420), .ZN(n6002) );
  INV_X1 U7286 ( .A(n6002), .ZN(n9682) );
  NOR2_X1 U7287 ( .A1(n9025), .A2(n9682), .ZN(n6788) );
  INV_X1 U7288 ( .A(n5750), .ZN(n5710) );
  NAND2_X1 U7289 ( .A1(n5755), .A2(n5710), .ZN(n5705) );
  NAND2_X1 U7290 ( .A1(n6788), .A2(n5705), .ZN(n9626) );
  NAND2_X1 U7291 ( .A1(n7542), .A2(n9021), .ZN(n9031) );
  OR2_X1 U7292 ( .A1(n9031), .A2(n5701), .ZN(n9796) );
  NAND2_X1 U7293 ( .A1(n9137), .A2(n9784), .ZN(n5708) );
  NAND2_X1 U7294 ( .A1(n7143), .A2(n9713), .ZN(n7265) );
  NAND2_X1 U7295 ( .A1(n9211), .A2(n9226), .ZN(n9206) );
  AOI211_X1 U7296 ( .C1(n5706), .C2(n9150), .A(n9321), .B(n9132), .ZN(n9138)
         );
  AOI21_X1 U7297 ( .B1(n9344), .B2(n5706), .A(n9138), .ZN(n5707) );
  NAND2_X1 U7298 ( .A1(n9136), .A2(n5709), .ZN(n6541) );
  AND2_X1 U7299 ( .A1(n9017), .A2(n5710), .ZN(n6008) );
  INV_X1 U7300 ( .A(n6008), .ZN(n5724) );
  NAND2_X1 U7301 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  NAND2_X1 U7302 ( .A1(n5713), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5714) );
  XNOR2_X1 U7303 ( .A(n5714), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6678) );
  INV_X1 U7304 ( .A(n6678), .ZN(n6706) );
  NAND2_X1 U7305 ( .A1(n4532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5715) );
  MUX2_X1 U7306 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5716), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5717) );
  INV_X1 U7307 ( .A(n5717), .ZN(n5720) );
  INV_X1 U7308 ( .A(n5718), .ZN(n5719) );
  NAND2_X1 U7309 ( .A1(n5718), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5721) );
  MUX2_X1 U7310 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5721), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5722) );
  AND2_X1 U7311 ( .A1(n6007), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5723) );
  INV_X1 U7312 ( .A(n6003), .ZN(n5743) );
  NOR2_X1 U7313 ( .A1(n7751), .A2(n5725), .ZN(n5726) );
  MUX2_X1 U7314 ( .A(n5726), .B(n5725), .S(n5745), .Z(n5727) );
  INV_X1 U7315 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U7316 ( .A1(n6698), .A2(n6702), .ZN(n5729) );
  OR2_X1 U7317 ( .A1(n7751), .A2(n5728), .ZN(n6700) );
  NAND2_X1 U7318 ( .A1(n5729), .A2(n6700), .ZN(n5742) );
  NOR4_X1 U7319 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5733) );
  NOR4_X1 U7320 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5732) );
  NOR4_X1 U7321 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5731) );
  NOR4_X1 U7322 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5730) );
  NAND4_X1 U7323 ( .A1(n5733), .A2(n5732), .A3(n5731), .A4(n5730), .ZN(n5739)
         );
  NOR2_X1 U7324 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .ZN(
        n5737) );
  NOR4_X1 U7325 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5736) );
  NOR4_X1 U7326 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5735) );
  NOR4_X1 U7327 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5734) );
  NAND4_X1 U7328 ( .A1(n5737), .A2(n5736), .A3(n5735), .A4(n5734), .ZN(n5738)
         );
  NOR2_X1 U7329 ( .A1(n5739), .A2(n5738), .ZN(n5994) );
  INV_X1 U7330 ( .A(n5994), .ZN(n5740) );
  NAND2_X1 U7331 ( .A1(n6698), .A2(n5740), .ZN(n5741) );
  NAND4_X1 U7332 ( .A1(n6784), .A2(n5743), .A3(n5742), .A4(n5741), .ZN(n6540)
         );
  INV_X1 U7333 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7334 ( .A1(n6698), .A2(n5744), .ZN(n5746) );
  INV_X1 U7335 ( .A(n5745), .ZN(n7677) );
  NAND2_X1 U7336 ( .A1(n7770), .A2(n7677), .ZN(n9450) );
  NAND2_X1 U7337 ( .A1(n5746), .A2(n9450), .ZN(n6783) );
  NAND2_X1 U7338 ( .A1(n6541), .A2(n9825), .ZN(n5748) );
  INV_X1 U7339 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U7340 ( .A1(n5748), .A2(n5079), .ZN(P1_U3551) );
  INV_X2 U7341 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U7342 ( .A1(n6001), .A2(n8988), .ZN(n5752) );
  INV_X2 U7343 ( .A(n5754), .ZN(n5967) );
  NAND2_X1 U7344 ( .A1(n5704), .A2(n5750), .ZN(n5751) );
  OR2_X2 U7345 ( .A1(n5752), .A2(n5702), .ZN(n6886) );
  NAND2_X4 U7346 ( .A1(n5753), .A2(n6886), .ZN(n5971) );
  OAI22_X1 U7347 ( .A1(n9392), .A2(n5967), .B1(n9381), .B2(n5971), .ZN(n8746)
         );
  NAND2_X1 U7348 ( .A1(n5755), .A2(n7420), .ZN(n5756) );
  NAND2_X2 U7349 ( .A1(n5971), .A2(n5988), .ZN(n5792) );
  NAND2_X1 U7350 ( .A1(n5792), .A2(n5761), .ZN(n5758) );
  NAND2_X1 U7351 ( .A1(n5759), .A2(n5758), .ZN(n5760) );
  INV_X4 U7352 ( .A(n5988), .ZN(n5981) );
  INV_X1 U7353 ( .A(n5766), .ZN(n5764) );
  AND2_X1 U7354 ( .A1(n5761), .A2(n5754), .ZN(n5762) );
  INV_X1 U7355 ( .A(n5765), .ZN(n5763) );
  NAND2_X1 U7356 ( .A1(n5764), .A2(n5763), .ZN(n5767) );
  NAND2_X1 U7357 ( .A1(n5766), .A2(n5765), .ZN(n6895) );
  NAND2_X1 U7358 ( .A1(n5767), .A2(n6895), .ZN(n7842) );
  INV_X1 U7359 ( .A(n7842), .ZN(n5778) );
  NAND2_X1 U7360 ( .A1(n6712), .A2(n5754), .ZN(n5769) );
  AND2_X1 U7361 ( .A1(n5769), .A2(n5768), .ZN(n5774) );
  INV_X1 U7362 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U7363 ( .A1(n6712), .A2(n5990), .ZN(n5773) );
  OAI22_X1 U7364 ( .A1(n6889), .A2(n5967), .B1(n9072), .B2(n6007), .ZN(n5771)
         );
  INV_X1 U7365 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7366 ( .A1(n5773), .A2(n5772), .ZN(n6761) );
  NAND2_X1 U7367 ( .A1(n6760), .A2(n6761), .ZN(n5776) );
  NAND2_X1 U7368 ( .A1(n5774), .A2(n5981), .ZN(n5775) );
  INV_X1 U7369 ( .A(n7841), .ZN(n5777) );
  NAND2_X1 U7370 ( .A1(n5778), .A2(n5777), .ZN(n6898) );
  NAND2_X1 U7371 ( .A1(n6898), .A2(n6895), .ZN(n5790) );
  NAND2_X1 U7372 ( .A1(n5779), .A2(n5754), .ZN(n5781) );
  INV_X1 U7373 ( .A(n5792), .ZN(n5798) );
  NAND2_X1 U7374 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  XNOR2_X1 U7375 ( .A(n5782), .B(n5981), .ZN(n5788) );
  INV_X1 U7376 ( .A(n5788), .ZN(n5786) );
  NAND2_X1 U7377 ( .A1(n5779), .A2(n5990), .ZN(n5784) );
  OR2_X1 U7378 ( .A1(n9691), .A2(n5967), .ZN(n5783) );
  INV_X1 U7379 ( .A(n5787), .ZN(n5785) );
  NAND2_X1 U7380 ( .A1(n5786), .A2(n5785), .ZN(n5789) );
  NAND2_X1 U7381 ( .A1(n5788), .A2(n5787), .ZN(n5791) );
  NAND2_X1 U7382 ( .A1(n5790), .A2(n6897), .ZN(n6899) );
  NAND2_X1 U7383 ( .A1(n6899), .A2(n5791), .ZN(n6953) );
  NAND2_X1 U7384 ( .A1(n9050), .A2(n5754), .ZN(n5794) );
  NAND2_X1 U7385 ( .A1(n6958), .A2(n5948), .ZN(n5793) );
  NAND2_X1 U7386 ( .A1(n5794), .A2(n5793), .ZN(n5795) );
  XNOR2_X1 U7387 ( .A(n5795), .B(n5981), .ZN(n5804) );
  NAND2_X1 U7388 ( .A1(n9050), .A2(n5990), .ZN(n5797) );
  NAND2_X1 U7389 ( .A1(n6958), .A2(n5991), .ZN(n5796) );
  NAND2_X1 U7390 ( .A1(n5797), .A2(n5796), .ZN(n5802) );
  XNOR2_X1 U7391 ( .A(n5804), .B(n5802), .ZN(n6955) );
  NAND2_X1 U7392 ( .A1(n9662), .A2(n5754), .ZN(n5799) );
  NAND2_X1 U7393 ( .A1(n9662), .A2(n5990), .ZN(n5801) );
  OR2_X1 U7394 ( .A1(n9705), .A2(n5967), .ZN(n5800) );
  NAND2_X1 U7395 ( .A1(n5801), .A2(n5800), .ZN(n5807) );
  INV_X1 U7396 ( .A(n5802), .ZN(n5803) );
  NAND2_X1 U7397 ( .A1(n5804), .A2(n5803), .ZN(n6966) );
  AND2_X1 U7398 ( .A1(n6965), .A2(n6966), .ZN(n5805) );
  INV_X1 U7399 ( .A(n5806), .ZN(n5808) );
  NAND2_X1 U7400 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  NAND2_X1 U7401 ( .A1(n9049), .A2(n5991), .ZN(n5810) );
  OAI21_X1 U7402 ( .B1(n9713), .B2(n5798), .A(n5810), .ZN(n5811) );
  XNOR2_X1 U7403 ( .A(n5811), .B(n5988), .ZN(n5814) );
  NAND2_X1 U7404 ( .A1(n7163), .A2(n5991), .ZN(n5813) );
  NAND2_X1 U7405 ( .A1(n9049), .A2(n5990), .ZN(n5812) );
  AND2_X1 U7406 ( .A1(n5813), .A2(n5812), .ZN(n7161) );
  OR2_X1 U7407 ( .A1(n7293), .A2(n5971), .ZN(n5818) );
  NAND2_X1 U7408 ( .A1(n7268), .A2(n5991), .ZN(n5817) );
  AND2_X1 U7409 ( .A1(n5818), .A2(n5817), .ZN(n5820) );
  INV_X1 U7410 ( .A(n5819), .ZN(n5822) );
  INV_X1 U7411 ( .A(n5820), .ZN(n5821) );
  NAND2_X1 U7412 ( .A1(n5822), .A2(n5821), .ZN(n7170) );
  NAND2_X1 U7413 ( .A1(n9653), .A2(n5991), .ZN(n5824) );
  OR2_X1 U7414 ( .A1(n9729), .A2(n5971), .ZN(n5823) );
  NAND2_X1 U7415 ( .A1(n5824), .A2(n5823), .ZN(n7288) );
  NAND2_X1 U7416 ( .A1(n9653), .A2(n5948), .ZN(n5826) );
  OR2_X1 U7417 ( .A1(n9729), .A2(n5967), .ZN(n5825) );
  NAND2_X1 U7418 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  XNOR2_X1 U7419 ( .A(n5827), .B(n5988), .ZN(n7289) );
  NAND2_X1 U7420 ( .A1(n9732), .A2(n5948), .ZN(n5829) );
  OR2_X1 U7421 ( .A1(n7582), .A2(n5967), .ZN(n5828) );
  NAND2_X1 U7422 ( .A1(n5829), .A2(n5828), .ZN(n5830) );
  XNOR2_X1 U7423 ( .A(n5830), .B(n5981), .ZN(n7559) );
  NOR2_X1 U7424 ( .A1(n7582), .A2(n5971), .ZN(n5831) );
  AOI21_X1 U7425 ( .B1(n9732), .B2(n5991), .A(n5831), .ZN(n5837) );
  NAND2_X1 U7426 ( .A1(n7559), .A2(n5837), .ZN(n5832) );
  NAND2_X1 U7427 ( .A1(n7558), .A2(n5832), .ZN(n5841) );
  NAND2_X1 U7428 ( .A1(n9740), .A2(n5948), .ZN(n5834) );
  OR2_X1 U7429 ( .A1(n9747), .A2(n5967), .ZN(n5833) );
  NAND2_X1 U7430 ( .A1(n5834), .A2(n5833), .ZN(n5835) );
  XNOR2_X1 U7431 ( .A(n5835), .B(n5988), .ZN(n5842) );
  NOR2_X1 U7432 ( .A1(n9747), .A2(n5971), .ZN(n5836) );
  AOI21_X1 U7433 ( .B1(n9740), .B2(n5991), .A(n5836), .ZN(n5843) );
  XNOR2_X1 U7434 ( .A(n5842), .B(n5843), .ZN(n7576) );
  INV_X1 U7435 ( .A(n7559), .ZN(n5838) );
  INV_X1 U7436 ( .A(n5837), .ZN(n7562) );
  NAND2_X1 U7437 ( .A1(n5838), .A2(n7562), .ZN(n5839) );
  AND2_X1 U7438 ( .A1(n7576), .A2(n5839), .ZN(n5840) );
  INV_X1 U7439 ( .A(n5842), .ZN(n5844) );
  NAND2_X1 U7440 ( .A1(n5844), .A2(n5843), .ZN(n5845) );
  NAND2_X1 U7441 ( .A1(n9751), .A2(n5948), .ZN(n5847) );
  OR2_X1 U7442 ( .A1(n7704), .A2(n5967), .ZN(n5846) );
  NAND2_X1 U7443 ( .A1(n5847), .A2(n5846), .ZN(n5848) );
  XNOR2_X1 U7444 ( .A(n5848), .B(n5981), .ZN(n5849) );
  NAND2_X1 U7445 ( .A1(n9751), .A2(n5991), .ZN(n5852) );
  OR2_X1 U7446 ( .A1(n7704), .A2(n5971), .ZN(n5851) );
  NAND2_X1 U7447 ( .A1(n5852), .A2(n5851), .ZN(n7640) );
  NAND2_X1 U7448 ( .A1(n7638), .A2(n7698), .ZN(n5861) );
  NAND2_X1 U7449 ( .A1(n9636), .A2(n5948), .ZN(n5855) );
  OR2_X1 U7450 ( .A1(n9748), .A2(n5967), .ZN(n5854) );
  NAND2_X1 U7451 ( .A1(n5855), .A2(n5854), .ZN(n5856) );
  XNOR2_X1 U7452 ( .A(n5856), .B(n5981), .ZN(n5859) );
  NOR2_X1 U7453 ( .A1(n9748), .A2(n5971), .ZN(n5857) );
  AOI21_X1 U7454 ( .B1(n9636), .B2(n5991), .A(n5857), .ZN(n5858) );
  NAND2_X1 U7455 ( .A1(n5859), .A2(n5858), .ZN(n7755) );
  OR2_X1 U7456 ( .A1(n5859), .A2(n5858), .ZN(n5860) );
  AND2_X1 U7457 ( .A1(n7755), .A2(n5860), .ZN(n7699) );
  NAND2_X1 U7458 ( .A1(n5861), .A2(n7699), .ZN(n7702) );
  NAND2_X1 U7459 ( .A1(n7469), .A2(n5948), .ZN(n5863) );
  OR2_X1 U7460 ( .A1(n9611), .A2(n5967), .ZN(n5862) );
  NAND2_X1 U7461 ( .A1(n5863), .A2(n5862), .ZN(n5864) );
  XNOR2_X1 U7462 ( .A(n5864), .B(n5981), .ZN(n5867) );
  NOR2_X1 U7463 ( .A1(n9611), .A2(n5971), .ZN(n5865) );
  AOI21_X1 U7464 ( .B1(n7469), .B2(n5991), .A(n5865), .ZN(n5866) );
  NAND2_X1 U7465 ( .A1(n5867), .A2(n5866), .ZN(n5869) );
  OR2_X1 U7466 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  AND2_X1 U7467 ( .A1(n5869), .A2(n5868), .ZN(n7756) );
  NAND2_X1 U7468 ( .A1(n9616), .A2(n5948), .ZN(n5871) );
  OR2_X1 U7469 ( .A1(n9788), .A2(n5967), .ZN(n5870) );
  NAND2_X1 U7470 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  XNOR2_X1 U7471 ( .A(n5872), .B(n5988), .ZN(n5874) );
  NOR2_X1 U7472 ( .A1(n9788), .A2(n5971), .ZN(n5873) );
  AOI21_X1 U7473 ( .B1(n9616), .B2(n5991), .A(n5873), .ZN(n5875) );
  XNOR2_X1 U7474 ( .A(n5874), .B(n5875), .ZN(n7792) );
  INV_X1 U7475 ( .A(n5874), .ZN(n5876) );
  NAND2_X1 U7476 ( .A1(n5876), .A2(n5875), .ZN(n5883) );
  NAND2_X1 U7477 ( .A1(n9793), .A2(n5948), .ZN(n5878) );
  OR2_X1 U7478 ( .A1(n9612), .A2(n5967), .ZN(n5877) );
  NAND2_X1 U7479 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  XNOR2_X1 U7480 ( .A(n5879), .B(n5981), .ZN(n5889) );
  INV_X1 U7481 ( .A(n5889), .ZN(n5880) );
  NAND2_X1 U7482 ( .A1(n5881), .A2(n5880), .ZN(n8655) );
  NOR2_X1 U7483 ( .A1(n9612), .A2(n5971), .ZN(n5882) );
  AOI21_X1 U7484 ( .B1(n9793), .B2(n5991), .A(n5882), .ZN(n8658) );
  AND2_X1 U7485 ( .A1(n5883), .A2(n8658), .ZN(n5884) );
  INV_X1 U7486 ( .A(n8658), .ZN(n5885) );
  OR2_X1 U7487 ( .A1(n5885), .A2(n5889), .ZN(n5886) );
  NAND2_X1 U7488 ( .A1(n5888), .A2(n5889), .ZN(n8654) );
  OAI22_X1 U7489 ( .A1(n9532), .A2(n5798), .B1(n9790), .B2(n5967), .ZN(n5890)
         );
  XNOR2_X1 U7490 ( .A(n5890), .B(n5981), .ZN(n5891) );
  OR2_X1 U7491 ( .A1(n9532), .A2(n5967), .ZN(n5894) );
  NAND2_X1 U7492 ( .A1(n9046), .A2(n5990), .ZN(n5893) );
  AND2_X1 U7493 ( .A1(n5894), .A2(n5893), .ZN(n8775) );
  NAND2_X1 U7494 ( .A1(n8774), .A2(n5895), .ZN(n8704) );
  NAND2_X1 U7495 ( .A1(n9431), .A2(n5948), .ZN(n5897) );
  OR2_X1 U7496 ( .A1(n9329), .A2(n5967), .ZN(n5896) );
  NAND2_X1 U7497 ( .A1(n5897), .A2(n5896), .ZN(n5898) );
  XNOR2_X1 U7498 ( .A(n5898), .B(n5981), .ZN(n5901) );
  NOR2_X1 U7499 ( .A1(n9329), .A2(n5971), .ZN(n5899) );
  AOI21_X1 U7500 ( .B1(n9431), .B2(n5991), .A(n5899), .ZN(n5900) );
  NAND2_X1 U7501 ( .A1(n5901), .A2(n5900), .ZN(n5903) );
  OR2_X1 U7502 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  AND2_X1 U7503 ( .A1(n5903), .A2(n5902), .ZN(n8705) );
  NAND2_X1 U7504 ( .A1(n8704), .A2(n8705), .ZN(n8703) );
  NAND2_X1 U7505 ( .A1(n9426), .A2(n5948), .ZN(n5905) );
  NAND2_X1 U7506 ( .A1(n9044), .A2(n5991), .ZN(n5904) );
  NAND2_X1 U7507 ( .A1(n5905), .A2(n5904), .ZN(n5906) );
  XNOR2_X1 U7508 ( .A(n5906), .B(n5988), .ZN(n5908) );
  AND2_X1 U7509 ( .A1(n9044), .A2(n5990), .ZN(n5907) );
  AOI21_X1 U7510 ( .B1(n9426), .B2(n5991), .A(n5907), .ZN(n5909) );
  XNOR2_X1 U7511 ( .A(n5908), .B(n5909), .ZN(n8715) );
  INV_X1 U7512 ( .A(n5908), .ZN(n5910) );
  NAND2_X1 U7513 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  NAND2_X1 U7514 ( .A1(n9413), .A2(n5948), .ZN(n5913) );
  OR2_X1 U7515 ( .A1(n9417), .A2(n5967), .ZN(n5912) );
  NAND2_X1 U7516 ( .A1(n5913), .A2(n5912), .ZN(n5914) );
  XNOR2_X1 U7517 ( .A(n5914), .B(n5981), .ZN(n8679) );
  INV_X1 U7518 ( .A(n8679), .ZN(n5917) );
  NAND2_X1 U7519 ( .A1(n9413), .A2(n5991), .ZN(n5916) );
  OR2_X1 U7520 ( .A1(n9417), .A2(n5971), .ZN(n5915) );
  NAND2_X1 U7521 ( .A1(n5916), .A2(n5915), .ZN(n8678) );
  NAND2_X1 U7522 ( .A1(n5917), .A2(n8678), .ZN(n8730) );
  NAND2_X1 U7523 ( .A1(n9421), .A2(n5948), .ZN(n5919) );
  OR2_X1 U7524 ( .A1(n9330), .A2(n5967), .ZN(n5918) );
  NAND2_X1 U7525 ( .A1(n5919), .A2(n5918), .ZN(n5920) );
  XNOR2_X1 U7526 ( .A(n5920), .B(n5981), .ZN(n8676) );
  INV_X1 U7527 ( .A(n8676), .ZN(n8675) );
  NOR2_X1 U7528 ( .A1(n9330), .A2(n5971), .ZN(n5921) );
  AOI21_X1 U7529 ( .B1(n9421), .B2(n5991), .A(n5921), .ZN(n8758) );
  INV_X1 U7530 ( .A(n8758), .ZN(n5929) );
  NAND2_X1 U7531 ( .A1(n8675), .A2(n5929), .ZN(n5922) );
  AND2_X1 U7532 ( .A1(n8730), .A2(n5922), .ZN(n5923) );
  NAND2_X1 U7533 ( .A1(n9406), .A2(n5948), .ZN(n5925) );
  OR2_X1 U7534 ( .A1(n9288), .A2(n5967), .ZN(n5924) );
  NAND2_X1 U7535 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  XNOR2_X1 U7536 ( .A(n5926), .B(n5981), .ZN(n5934) );
  NOR2_X1 U7537 ( .A1(n9288), .A2(n5971), .ZN(n5927) );
  AOI21_X1 U7538 ( .B1(n9406), .B2(n5991), .A(n5927), .ZN(n5935) );
  NAND2_X1 U7539 ( .A1(n5934), .A2(n5935), .ZN(n8732) );
  NAND2_X1 U7540 ( .A1(n8676), .A2(n8758), .ZN(n5928) );
  NAND2_X1 U7541 ( .A1(n5928), .A2(n8678), .ZN(n5931) );
  NOR2_X1 U7542 ( .A1(n8678), .A2(n5929), .ZN(n5930) );
  AOI22_X1 U7543 ( .A1(n8679), .A2(n5931), .B1(n5930), .B2(n8676), .ZN(n5932)
         );
  INV_X1 U7544 ( .A(n5934), .ZN(n5937) );
  INV_X1 U7545 ( .A(n5935), .ZN(n5936) );
  AND2_X1 U7546 ( .A1(n5937), .A2(n5936), .ZN(n8733) );
  NAND2_X1 U7547 ( .A1(n9262), .A2(n5948), .ZN(n5941) );
  OR2_X1 U7548 ( .A1(n9277), .A2(n5967), .ZN(n5940) );
  NAND2_X1 U7549 ( .A1(n5941), .A2(n5940), .ZN(n5942) );
  XNOR2_X1 U7550 ( .A(n5942), .B(n5981), .ZN(n5946) );
  NOR2_X1 U7551 ( .A1(n9277), .A2(n5971), .ZN(n5943) );
  AOI21_X1 U7552 ( .B1(n9262), .B2(n5991), .A(n5943), .ZN(n5945) );
  XNOR2_X1 U7553 ( .A(n5946), .B(n5945), .ZN(n8690) );
  INV_X1 U7554 ( .A(n8690), .ZN(n5944) );
  NAND2_X1 U7555 ( .A1(n5946), .A2(n5945), .ZN(n5947) );
  NAND2_X1 U7556 ( .A1(n9248), .A2(n5948), .ZN(n5950) );
  OR2_X1 U7557 ( .A1(n9381), .A2(n5967), .ZN(n5949) );
  NAND2_X1 U7558 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  XNOR2_X1 U7559 ( .A(n5951), .B(n5981), .ZN(n5952) );
  NAND2_X1 U7560 ( .A1(n9384), .A2(n5948), .ZN(n5955) );
  OR2_X1 U7561 ( .A1(n9216), .A2(n5967), .ZN(n5954) );
  NAND2_X1 U7562 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  XNOR2_X1 U7563 ( .A(n5956), .B(n5981), .ZN(n5959) );
  NOR2_X1 U7564 ( .A1(n9216), .A2(n5971), .ZN(n5957) );
  AOI21_X1 U7565 ( .B1(n9384), .B2(n5991), .A(n5957), .ZN(n5958) );
  OR2_X1 U7566 ( .A1(n5959), .A2(n5958), .ZN(n8666) );
  AOI22_X1 U7567 ( .A1(n9375), .A2(n5948), .B1(n5991), .B2(n9228), .ZN(n5960)
         );
  XNOR2_X1 U7568 ( .A(n5960), .B(n5988), .ZN(n5962) );
  AOI22_X1 U7569 ( .A1(n9375), .A2(n5991), .B1(n5990), .B2(n9228), .ZN(n5961)
         );
  NAND2_X1 U7570 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  OAI21_X1 U7571 ( .B1(n5962), .B2(n5961), .A(n5963), .ZN(n8723) );
  NAND2_X1 U7572 ( .A1(n9370), .A2(n5948), .ZN(n5965) );
  OR2_X1 U7573 ( .A1(n9358), .A2(n5967), .ZN(n5964) );
  NAND2_X1 U7574 ( .A1(n5965), .A2(n5964), .ZN(n5966) );
  XNOR2_X1 U7575 ( .A(n5966), .B(n5988), .ZN(n5974) );
  INV_X1 U7576 ( .A(n9370), .ZN(n9201) );
  OAI22_X1 U7577 ( .A1(n9201), .A2(n5967), .B1(n9358), .B2(n5971), .ZN(n5973)
         );
  XNOR2_X1 U7578 ( .A(n5974), .B(n5973), .ZN(n8696) );
  NAND2_X1 U7579 ( .A1(n9362), .A2(n5948), .ZN(n5969) );
  OR2_X1 U7580 ( .A1(n9367), .A2(n5967), .ZN(n5968) );
  NAND2_X1 U7581 ( .A1(n5969), .A2(n5968), .ZN(n5970) );
  XNOR2_X1 U7582 ( .A(n5970), .B(n5981), .ZN(n5975) );
  NOR2_X1 U7583 ( .A1(n9367), .A2(n5971), .ZN(n5972) );
  AOI21_X1 U7584 ( .B1(n9362), .B2(n5991), .A(n5972), .ZN(n5976) );
  XNOR2_X1 U7585 ( .A(n5975), .B(n5976), .ZN(n8764) );
  NOR2_X1 U7586 ( .A1(n5974), .A2(n5973), .ZN(n8765) );
  INV_X1 U7587 ( .A(n5975), .ZN(n5978) );
  INV_X1 U7588 ( .A(n5976), .ZN(n5977) );
  NAND2_X1 U7589 ( .A1(n9352), .A2(n5948), .ZN(n5980) );
  NAND2_X1 U7590 ( .A1(n9183), .A2(n5991), .ZN(n5979) );
  NAND2_X1 U7591 ( .A1(n5980), .A2(n5979), .ZN(n5982) );
  XNOR2_X1 U7592 ( .A(n5982), .B(n5981), .ZN(n5985) );
  AND2_X1 U7593 ( .A1(n9183), .A2(n5990), .ZN(n5983) );
  AOI21_X1 U7594 ( .B1(n9352), .B2(n5991), .A(n5983), .ZN(n5984) );
  NAND2_X1 U7595 ( .A1(n5985), .A2(n5984), .ZN(n6016) );
  OAI21_X1 U7596 ( .B1(n5985), .B2(n5984), .A(n6016), .ZN(n6532) );
  NAND2_X1 U7597 ( .A1(n9152), .A2(n5948), .ZN(n5987) );
  NAND2_X1 U7598 ( .A1(n9171), .A2(n5991), .ZN(n5986) );
  NAND2_X1 U7599 ( .A1(n5987), .A2(n5986), .ZN(n5989) );
  XNOR2_X1 U7600 ( .A(n5989), .B(n5988), .ZN(n5993) );
  AOI22_X1 U7601 ( .A1(n9152), .A2(n5991), .B1(n5990), .B2(n9171), .ZN(n5992)
         );
  XNOR2_X1 U7602 ( .A(n5993), .B(n5992), .ZN(n6000) );
  INV_X1 U7603 ( .A(n6000), .ZN(n6017) );
  NAND2_X1 U7604 ( .A1(n5994), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7605 ( .A1(n6698), .A2(n5995), .ZN(n5996) );
  NAND2_X1 U7606 ( .A1(n5996), .A2(n6700), .ZN(n6782) );
  OR2_X1 U7607 ( .A1(n6783), .A2(n6782), .ZN(n6005) );
  INV_X1 U7608 ( .A(n9026), .ZN(n6705) );
  NOR2_X1 U7609 ( .A1(n6005), .A2(n6705), .ZN(n6011) );
  AND2_X1 U7610 ( .A1(n5997), .A2(n9781), .ZN(n5998) );
  NAND3_X1 U7611 ( .A1(n6017), .A2(n8777), .A3(n6016), .ZN(n5999) );
  INV_X1 U7612 ( .A(n6011), .ZN(n6004) );
  OR2_X1 U7613 ( .A1(n6002), .A2(n6001), .ZN(n6791) );
  OAI21_X2 U7614 ( .B1(n6004), .B2(n6791), .A(n9664), .ZN(n8769) );
  NAND2_X1 U7615 ( .A1(n5701), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7297) );
  INV_X1 U7616 ( .A(n6005), .ZN(n6006) );
  AOI21_X1 U7617 ( .B1(n9344), .B2(n7297), .A(n6006), .ZN(n6762) );
  AND2_X1 U7618 ( .A1(n6678), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9024) );
  INV_X1 U7619 ( .A(n6007), .ZN(n6677) );
  NOR4_X1 U7620 ( .A1(n6762), .A2(n9024), .A3(n6677), .A4(n6008), .ZN(n6009)
         );
  AOI22_X1 U7621 ( .A1(n6010), .A2(n9151), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6015) );
  NAND2_X1 U7622 ( .A1(n6011), .A2(n9025), .ZN(n6012) );
  NOR2_X1 U7623 ( .A1(n6012), .A2(n7068), .ZN(n8768) );
  INV_X1 U7624 ( .A(n6012), .ZN(n6013) );
  AOI22_X1 U7625 ( .A1(n8768), .A2(n9041), .B1(n8767), .B2(n9183), .ZN(n6014)
         );
  NAND2_X1 U7626 ( .A1(n6015), .A2(n6014), .ZN(n6019) );
  NOR3_X1 U7627 ( .A1(n6017), .A2(n8754), .A3(n6016), .ZN(n6018) );
  AOI211_X1 U7628 ( .C1(n9152), .C2(n8769), .A(n6019), .B(n6018), .ZN(n6020)
         );
  NOR2_X4 U7629 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6070) );
  NAND4_X1 U7630 ( .A1(n6026), .A2(n6025), .A3(n6024), .A4(n10333), .ZN(n6029)
         );
  NAND4_X1 U7631 ( .A1(n6280), .A2(n6238), .A3(n6233), .A4(n6027), .ZN(n6028)
         );
  NOR2_X1 U7632 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6030) );
  NAND2_X1 U7633 ( .A1(n6490), .A2(n6038), .ZN(n6032) );
  NOR2_X1 U7634 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6036) );
  NAND4_X1 U7635 ( .A1(n6036), .A2(n10184), .A3(n6475), .A4(n6035), .ZN(n6040)
         );
  INV_X1 U7636 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6037) );
  NAND4_X1 U7637 ( .A1(n6464), .A2(n6038), .A3(n6338), .A4(n6037), .ZN(n6039)
         );
  NOR2_X1 U7638 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  NAND2_X1 U7639 ( .A1(n6063), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7640 ( .A1(n6044), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6045) );
  MUX2_X1 U7641 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6045), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6047) );
  NAND2_X1 U7642 ( .A1(n6047), .A2(n6046), .ZN(n8026) );
  NAND2_X1 U7643 ( .A1(n4560), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6048) );
  XNOR2_X1 U7644 ( .A(n8026), .B(n6661), .ZN(n6057) );
  INV_X1 U7645 ( .A(n6054), .ZN(n6052) );
  NOR2_X1 U7646 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6049) );
  INV_X1 U7647 ( .A(P2_B_REG_SCAN_IN), .ZN(n6638) );
  AOI22_X1 U7648 ( .A1(n6049), .A2(P2_B_REG_SCAN_IN), .B1(n6638), .B2(
        P2_IR_REG_24__SCAN_IN), .ZN(n6050) );
  INV_X1 U7649 ( .A(n6050), .ZN(n6051) );
  XNOR2_X1 U7650 ( .A(P2_IR_REG_24__SCAN_IN), .B(P2_B_REG_SCAN_IN), .ZN(n6053)
         );
  NAND3_X1 U7651 ( .A1(n6054), .A2(P2_IR_REG_25__SCAN_IN), .A3(n6053), .ZN(
        n6055) );
  INV_X1 U7652 ( .A(n7767), .ZN(n6466) );
  INV_X1 U7653 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10318) );
  NAND3_X1 U7654 ( .A1(n6735), .A2(n6057), .A3(n6471), .ZN(n6062) );
  INV_X1 U7655 ( .A(n6058), .ZN(n6059) );
  NAND2_X1 U7656 ( .A1(n6059), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U7657 ( .A1(n6339), .A2(n6338), .ZN(n6341) );
  NAND2_X1 U7658 ( .A1(n6341), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6061) );
  INV_X1 U7659 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7660 ( .A1(n8251), .A2(n8203), .ZN(n6518) );
  NAND2_X2 U7661 ( .A1(n6062), .A2(n6518), .ZN(n6157) );
  NOR2_X1 U7662 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n6066) );
  INV_X1 U7663 ( .A(n6066), .ZN(n6067) );
  INV_X1 U7664 ( .A(n6074), .ZN(n6675) );
  NAND2_X1 U7665 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6069) );
  INV_X1 U7666 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6068) );
  MUX2_X1 U7667 ( .A(n6069), .B(P2_IR_REG_31__SCAN_IN), .S(n6068), .Z(n6072)
         );
  INV_X1 U7668 ( .A(n6070), .ZN(n6071) );
  NOR2_X1 U7669 ( .A1(n6074), .A2(n8014), .ZN(n6099) );
  NAND2_X1 U7670 ( .A1(n6099), .A2(n6073), .ZN(n6076) );
  NAND2_X1 U7671 ( .A1(n6297), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6075) );
  OAI211_X1 U7672 ( .C1(n6675), .C2(n6805), .A(n6076), .B(n6075), .ZN(n6549)
         );
  XNOR2_X1 U7673 ( .A(n6157), .B(n6549), .ZN(n6096) );
  INV_X1 U7674 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6079) );
  INV_X1 U7675 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6081) );
  INV_X1 U7676 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7183) );
  OR2_X1 U7677 ( .A1(n6147), .A2(n7183), .ZN(n6545) );
  NAND2_X2 U7678 ( .A1(n4498), .A2(n6083), .ZN(n6429) );
  NAND2_X1 U7679 ( .A1(n6117), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6547) );
  INV_X1 U7680 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6085) );
  OR2_X1 U7681 ( .A1(n6118), .A2(n6085), .ZN(n6546) );
  INV_X1 U7682 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7189) );
  OR2_X1 U7683 ( .A1(n6120), .A2(n7189), .ZN(n6544) );
  INV_X1 U7684 ( .A(n9996), .ZN(n8234) );
  XNOR2_X1 U7685 ( .A(n6096), .B(n8234), .ZN(n6939) );
  NAND2_X1 U7686 ( .A1(n6680), .A2(SI_0_), .ZN(n6087) );
  XNOR2_X1 U7687 ( .A(n6087), .B(n6086), .ZN(n8652) );
  INV_X1 U7688 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6806) );
  INV_X2 U7689 ( .A(n6675), .ZN(n6639) );
  MUX2_X1 U7690 ( .A(n8652), .B(n6806), .S(n6639), .Z(n6932) );
  NAND2_X1 U7691 ( .A1(n6157), .A2(n6932), .ZN(n6095) );
  INV_X1 U7692 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6088) );
  INV_X1 U7693 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6935) );
  OR2_X1 U7694 ( .A1(n6147), .A2(n6935), .ZN(n6093) );
  INV_X1 U7695 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6089) );
  OR2_X1 U7696 ( .A1(n6120), .A2(n6089), .ZN(n6092) );
  INV_X1 U7697 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6090) );
  OR2_X1 U7698 ( .A1(n6429), .A2(n6090), .ZN(n6091) );
  INV_X1 U7699 ( .A(n6932), .ZN(n7215) );
  NAND2_X1 U7700 ( .A1(n6939), .A2(n6940), .ZN(n6938) );
  NAND2_X1 U7701 ( .A1(n6096), .A2(n9996), .ZN(n6097) );
  NAND2_X1 U7702 ( .A1(n6938), .A2(n6097), .ZN(n6974) );
  INV_X1 U7703 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7704 ( .A1(n6070), .A2(n6098), .ZN(n6110) );
  INV_X1 U7705 ( .A(n6099), .ZN(n6279) );
  NAND2_X1 U7706 ( .A1(n6099), .A2(n6100), .ZN(n6101) );
  XNOR2_X1 U7707 ( .A(n6157), .B(n6553), .ZN(n6107) );
  INV_X1 U7708 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6804) );
  OR2_X1 U7709 ( .A1(n6429), .A2(n6804), .ZN(n6105) );
  INV_X1 U7710 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9988) );
  OR2_X1 U7711 ( .A1(n6147), .A2(n9988), .ZN(n6104) );
  INV_X1 U7712 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6102) );
  OR2_X1 U7713 ( .A1(n6118), .A2(n6102), .ZN(n6103) );
  XNOR2_X1 U7714 ( .A(n6107), .B(n8232), .ZN(n6973) );
  NAND2_X1 U7715 ( .A1(n6974), .A2(n6973), .ZN(n6109) );
  NAND2_X1 U7716 ( .A1(n6107), .A2(n4755), .ZN(n6108) );
  NAND2_X1 U7717 ( .A1(n6110), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6111) );
  MUX2_X1 U7718 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6111), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n6113) );
  NAND2_X1 U7719 ( .A1(n6113), .A2(n6112), .ZN(n6849) );
  NAND2_X1 U7720 ( .A1(n4499), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7721 ( .A1(n6099), .A2(n6114), .ZN(n6115) );
  OAI211_X1 U7722 ( .C1(n6675), .C2(n6849), .A(n6116), .B(n6115), .ZN(n7194)
         );
  XNOR2_X1 U7723 ( .A(n6157), .B(n7194), .ZN(n6126) );
  NAND2_X1 U7724 ( .A1(n7347), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6125) );
  OR2_X1 U7725 ( .A1(n6344), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6124) );
  INV_X1 U7726 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6119) );
  OR2_X1 U7727 ( .A1(n7349), .A2(n6119), .ZN(n6123) );
  INV_X1 U7728 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6121) );
  XNOR2_X1 U7729 ( .A(n6126), .B(n9994), .ZN(n6996) );
  INV_X1 U7730 ( .A(n6126), .ZN(n6127) );
  NAND2_X1 U7731 ( .A1(n6127), .A2(n4841), .ZN(n6128) );
  NAND2_X1 U7732 ( .A1(n6112), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6130) );
  INV_X1 U7733 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6129) );
  XNOR2_X1 U7734 ( .A(n6130), .B(n6129), .ZN(n9863) );
  NAND2_X1 U7735 ( .A1(n4499), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7736 ( .A1(n6099), .A2(n6688), .ZN(n6131) );
  OAI211_X1 U7737 ( .C1(n6675), .C2(n9863), .A(n6132), .B(n6131), .ZN(n8095)
         );
  XNOR2_X1 U7738 ( .A(n6157), .B(n8095), .ZN(n6142) );
  NAND2_X1 U7739 ( .A1(n6133), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6141) );
  INV_X1 U7740 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6839) );
  OR2_X1 U7741 ( .A1(n6429), .A2(n6839), .ZN(n6140) );
  NAND2_X1 U7742 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6136) );
  AND2_X1 U7743 ( .A1(n6150), .A2(n6136), .ZN(n7004) );
  OR2_X1 U7744 ( .A1(n6344), .A2(n7004), .ZN(n6139) );
  INV_X1 U7745 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6137) );
  OR2_X1 U7746 ( .A1(n7349), .A2(n6137), .ZN(n6138) );
  XNOR2_X1 U7747 ( .A(n6142), .B(n8096), .ZN(n7003) );
  NAND2_X1 U7748 ( .A1(n6142), .A2(n8096), .ZN(n7042) );
  OR2_X1 U7749 ( .A1(n6694), .A2(n6279), .ZN(n6146) );
  OR2_X1 U7750 ( .A1(n6143), .A2(n8644), .ZN(n6144) );
  XNOR2_X1 U7751 ( .A(n6144), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9888) );
  AOI22_X1 U7752 ( .A1(n4499), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9888), .B2(
        n6639), .ZN(n6145) );
  NAND2_X1 U7753 ( .A1(n6146), .A2(n6145), .ZN(n6607) );
  XNOR2_X1 U7754 ( .A(n6157), .B(n6607), .ZN(n6174) );
  NAND2_X1 U7755 ( .A1(n7347), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6156) );
  INV_X1 U7756 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U7757 ( .A1(n6150), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6151) );
  AND2_X1 U7758 ( .A1(n6163), .A2(n6151), .ZN(n7122) );
  OR2_X1 U7759 ( .A1(n6344), .A2(n7122), .ZN(n6154) );
  INV_X1 U7760 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6152) );
  OR2_X1 U7761 ( .A1(n7349), .A2(n6152), .ZN(n6153) );
  INV_X1 U7762 ( .A(n8230), .ZN(n7200) );
  NAND2_X1 U7763 ( .A1(n6174), .A2(n7200), .ZN(n6173) );
  AND2_X1 U7764 ( .A1(n7042), .A2(n6173), .ZN(n7126) );
  OR2_X1 U7765 ( .A1(n6697), .A2(n6279), .ZN(n6162) );
  AND2_X1 U7766 ( .A1(n6143), .A2(n6158), .ZN(n6159) );
  AOI22_X1 U7767 ( .A1(n6451), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6917), .B2(
        n6639), .ZN(n6161) );
  XNOR2_X1 U7768 ( .A(n6410), .B(n10032), .ZN(n6172) );
  NAND2_X1 U7769 ( .A1(n6133), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6169) );
  INV_X1 U7770 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6916) );
  OR2_X1 U7771 ( .A1(n6429), .A2(n6916), .ZN(n6168) );
  NAND2_X1 U7772 ( .A1(n6163), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6164) );
  AND2_X1 U7773 ( .A1(n6185), .A2(n6164), .ZN(n7225) );
  OR2_X1 U7774 ( .A1(n6344), .A2(n7225), .ZN(n6167) );
  INV_X1 U7775 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6165) );
  OR2_X1 U7776 ( .A1(n7349), .A2(n6165), .ZN(n6166) );
  NAND4_X1 U7777 ( .A1(n6169), .A2(n6168), .A3(n6167), .A4(n6166), .ZN(n8229)
         );
  XNOR2_X1 U7778 ( .A(n6172), .B(n8229), .ZN(n7134) );
  INV_X1 U7779 ( .A(n7134), .ZN(n6170) );
  AND2_X1 U7780 ( .A1(n7126), .A2(n6170), .ZN(n6171) );
  NAND2_X1 U7781 ( .A1(n6172), .A2(n8229), .ZN(n6176) );
  INV_X1 U7782 ( .A(n6173), .ZN(n6175) );
  XNOR2_X1 U7783 ( .A(n6174), .B(n8230), .ZN(n7044) );
  OR2_X1 U7784 ( .A1(n6175), .A2(n7044), .ZN(n7128) );
  OR2_X1 U7785 ( .A1(n7134), .A2(n7128), .ZN(n7130) );
  AND2_X1 U7786 ( .A1(n6176), .A2(n7130), .ZN(n6177) );
  OR2_X1 U7787 ( .A1(n6703), .A2(n6279), .ZN(n6181) );
  NAND2_X1 U7788 ( .A1(n6178), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6179) );
  XNOR2_X1 U7789 ( .A(n6179), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7016) );
  AOI22_X1 U7790 ( .A1(n6451), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7016), .B2(
        n6639), .ZN(n6180) );
  NAND2_X1 U7791 ( .A1(n6181), .A2(n6180), .ZN(n7153) );
  XNOR2_X1 U7792 ( .A(n6410), .B(n7153), .ZN(n6192) );
  NAND2_X1 U7793 ( .A1(n7347), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6191) );
  INV_X1 U7794 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6182) );
  OR2_X1 U7795 ( .A1(n7352), .A2(n6182), .ZN(n6190) );
  NAND2_X1 U7796 ( .A1(n6185), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6186) );
  AND2_X1 U7797 ( .A1(n6198), .A2(n6186), .ZN(n7281) );
  OR2_X1 U7798 ( .A1(n6344), .A2(n7281), .ZN(n6189) );
  INV_X1 U7799 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6187) );
  OR2_X1 U7800 ( .A1(n7349), .A2(n6187), .ZN(n6188) );
  NAND4_X1 U7801 ( .A1(n6191), .A2(n6190), .A3(n6189), .A4(n6188), .ZN(n8228)
         );
  XNOR2_X1 U7802 ( .A(n6192), .B(n8228), .ZN(n7150) );
  NAND2_X1 U7803 ( .A1(n6192), .A2(n6609), .ZN(n6193) );
  NAND2_X1 U7804 ( .A1(n6709), .A2(n8048), .ZN(n6196) );
  NAND2_X1 U7805 ( .A1(n6206), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6194) );
  XNOR2_X1 U7806 ( .A(n6194), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7035) );
  AOI22_X1 U7807 ( .A1(n6451), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7035), .B2(
        n6639), .ZN(n6195) );
  NAND2_X1 U7808 ( .A1(n6196), .A2(n6195), .ZN(n10044) );
  XNOR2_X1 U7809 ( .A(n10044), .B(n6410), .ZN(n6204) );
  NAND2_X1 U7810 ( .A1(n6133), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6203) );
  INV_X1 U7811 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7017) );
  OR2_X1 U7812 ( .A1(n6429), .A2(n7017), .ZN(n6202) );
  INV_X1 U7813 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6197) );
  OR2_X1 U7814 ( .A1(n7349), .A2(n6197), .ZN(n6201) );
  NAND2_X1 U7815 ( .A1(n6198), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6199) );
  AND2_X1 U7816 ( .A1(n6212), .A2(n6199), .ZN(n7373) );
  OR2_X1 U7817 ( .A1(n6344), .A2(n7373), .ZN(n6200) );
  NAND4_X1 U7818 ( .A1(n6203), .A2(n6202), .A3(n6201), .A4(n6200), .ZN(n8227)
         );
  XNOR2_X1 U7819 ( .A(n6204), .B(n8227), .ZN(n7230) );
  NAND2_X1 U7820 ( .A1(n6204), .A2(n7549), .ZN(n6205) );
  NAND2_X1 U7821 ( .A1(n6721), .A2(n8048), .ZN(n6208) );
  NAND2_X1 U7822 ( .A1(n6236), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6225) );
  XNOR2_X1 U7823 ( .A(n6225), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7339) );
  AOI22_X1 U7824 ( .A1(n6451), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7339), .B2(
        n6639), .ZN(n6207) );
  NAND2_X1 U7825 ( .A1(n6208), .A2(n6207), .ZN(n7552) );
  XNOR2_X1 U7826 ( .A(n7552), .B(n7829), .ZN(n6218) );
  NAND2_X1 U7827 ( .A1(n7347), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6217) );
  INV_X1 U7828 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6209) );
  OR2_X1 U7829 ( .A1(n7349), .A2(n6209), .ZN(n6216) );
  NAND2_X1 U7830 ( .A1(n6212), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6213) );
  AND2_X1 U7831 ( .A1(n6219), .A2(n6213), .ZN(n7550) );
  OR2_X1 U7832 ( .A1(n6344), .A2(n7550), .ZN(n6215) );
  INV_X1 U7833 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7551) );
  OR2_X1 U7834 ( .A1(n7352), .A2(n7551), .ZN(n6214) );
  NAND4_X1 U7835 ( .A1(n6217), .A2(n6216), .A3(n6215), .A4(n6214), .ZN(n8226)
         );
  XNOR2_X1 U7836 ( .A(n6218), .B(n8226), .ZN(n7411) );
  NAND2_X1 U7837 ( .A1(n6593), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6224) );
  INV_X1 U7838 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7434) );
  OR2_X1 U7839 ( .A1(n6429), .A2(n7434), .ZN(n6223) );
  NAND2_X1 U7840 ( .A1(n6219), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6220) );
  AND2_X1 U7841 ( .A1(n6245), .A2(n6220), .ZN(n7594) );
  OR2_X1 U7842 ( .A1(n6344), .A2(n7594), .ZN(n6222) );
  INV_X1 U7843 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7595) );
  OR2_X1 U7844 ( .A1(n7352), .A2(n7595), .ZN(n6221) );
  OR2_X1 U7845 ( .A1(n6717), .A2(n6279), .ZN(n6229) );
  INV_X1 U7846 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7847 ( .A1(n6225), .A2(n6234), .ZN(n6226) );
  NAND2_X1 U7848 ( .A1(n6226), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6227) );
  XNOR2_X1 U7849 ( .A(n6227), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7445) );
  AOI22_X1 U7850 ( .A1(n6451), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7445), .B2(
        n6639), .ZN(n6228) );
  NAND2_X1 U7851 ( .A1(n6229), .A2(n6228), .ZN(n7597) );
  XNOR2_X1 U7852 ( .A(n7597), .B(n6410), .ZN(n7454) );
  INV_X1 U7853 ( .A(n6230), .ZN(n6231) );
  NAND2_X1 U7854 ( .A1(n6231), .A2(n7682), .ZN(n6232) );
  NAND2_X1 U7855 ( .A1(n6738), .A2(n8048), .ZN(n6243) );
  NAND2_X1 U7856 ( .A1(n6234), .A2(n6233), .ZN(n6235) );
  NOR2_X1 U7857 ( .A1(n6239), .A2(n8644), .ZN(n6237) );
  MUX2_X1 U7858 ( .A(n8644), .B(n6237), .S(P2_IR_REG_11__SCAN_IN), .Z(n6241)
         );
  NAND2_X1 U7859 ( .A1(n6239), .A2(n6238), .ZN(n6262) );
  INV_X1 U7860 ( .A(n6262), .ZN(n6240) );
  AOI22_X1 U7861 ( .A1(n6451), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7613), .B2(
        n6639), .ZN(n6242) );
  NAND2_X1 U7862 ( .A1(n6593), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6250) );
  INV_X1 U7863 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6244) );
  OR2_X1 U7864 ( .A1(n7352), .A2(n6244), .ZN(n6249) );
  OR2_X1 U7865 ( .A1(n6429), .A2(n10077), .ZN(n6248) );
  NAND2_X1 U7866 ( .A1(n6245), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6246) );
  AND2_X1 U7867 ( .A1(n6253), .A2(n6246), .ZN(n7683) );
  OR2_X1 U7868 ( .A1(n6344), .A2(n7683), .ZN(n6247) );
  OR2_X1 U7869 ( .A1(n10054), .A2(n8116), .ZN(n8113) );
  NAND2_X1 U7870 ( .A1(n10054), .A2(n8116), .ZN(n8091) );
  NAND2_X1 U7871 ( .A1(n8113), .A2(n8091), .ZN(n7679) );
  XNOR2_X1 U7872 ( .A(n7679), .B(n6410), .ZN(n7666) );
  INV_X1 U7873 ( .A(n7666), .ZN(n6251) );
  INV_X1 U7874 ( .A(n8116), .ZN(n8224) );
  NAND2_X1 U7875 ( .A1(n7666), .A2(n8224), .ZN(n6252) );
  NAND2_X1 U7876 ( .A1(n7663), .A2(n6252), .ZN(n7654) );
  NAND2_X1 U7877 ( .A1(n6593), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6258) );
  INV_X1 U7878 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7615) );
  OR2_X1 U7879 ( .A1(n7352), .A2(n7615), .ZN(n6257) );
  INV_X1 U7880 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7614) );
  OR2_X1 U7881 ( .A1(n6429), .A2(n7614), .ZN(n6256) );
  NAND2_X1 U7882 ( .A1(n6253), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6254) );
  AND2_X1 U7883 ( .A1(n6270), .A2(n6254), .ZN(n7746) );
  OR2_X1 U7884 ( .A1(n6344), .A2(n7746), .ZN(n6255) );
  NAND4_X1 U7885 ( .A1(n6258), .A2(n6257), .A3(n6256), .A4(n6255), .ZN(n8223)
         );
  NAND2_X1 U7886 ( .A1(n6262), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6259) );
  XNOR2_X1 U7887 ( .A(n6259), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8244) );
  AOI22_X1 U7888 ( .A1(n6451), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8244), .B2(
        n6639), .ZN(n6260) );
  XNOR2_X1 U7889 ( .A(n7748), .B(n7829), .ZN(n7652) );
  NAND2_X1 U7890 ( .A1(n6263), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6281) );
  XNOR2_X1 U7891 ( .A(n6281), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U7892 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n6451), .B1(n9899), .B2(
        n6639), .ZN(n6264) );
  XNOR2_X1 U7893 ( .A(n8129), .B(n7829), .ZN(n7733) );
  NAND2_X1 U7894 ( .A1(n6593), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6275) );
  INV_X1 U7895 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6266) );
  OR2_X1 U7896 ( .A1(n7352), .A2(n6266), .ZN(n6274) );
  INV_X1 U7897 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6267) );
  OR2_X1 U7898 ( .A1(n6429), .A2(n6267), .ZN(n6273) );
  INV_X1 U7899 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7900 ( .A1(n6270), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6271) );
  AND2_X1 U7901 ( .A1(n6287), .A2(n6271), .ZN(n8498) );
  OR2_X1 U7902 ( .A1(n6344), .A2(n8498), .ZN(n6272) );
  NAND4_X1 U7903 ( .A1(n6275), .A2(n6274), .A3(n6273), .A4(n6272), .ZN(n8482)
         );
  INV_X1 U7904 ( .A(n7733), .ZN(n6276) );
  NAND2_X1 U7905 ( .A1(n6276), .A2(n8127), .ZN(n6277) );
  NAND2_X1 U7906 ( .A1(n6927), .A2(n8048), .ZN(n6286) );
  NAND2_X1 U7907 ( .A1(n6281), .A2(n6280), .ZN(n6282) );
  NAND2_X1 U7908 ( .A1(n6282), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6283) );
  OR2_X1 U7909 ( .A1(n6283), .A2(n10333), .ZN(n6284) );
  NAND2_X1 U7910 ( .A1(n6283), .A2(n10333), .ZN(n6295) );
  AOI22_X1 U7911 ( .A1(n9914), .A2(n6639), .B1(P1_DATAO_REG_14__SCAN_IN), .B2(
        n6451), .ZN(n6285) );
  XNOR2_X1 U7912 ( .A(n8637), .B(n6410), .ZN(n6293) );
  NAND2_X1 U7913 ( .A1(n6593), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6292) );
  INV_X1 U7914 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8548) );
  OR2_X1 U7915 ( .A1(n6429), .A2(n8548), .ZN(n6291) );
  NAND2_X1 U7916 ( .A1(n6287), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6288) );
  AND2_X1 U7917 ( .A1(n6301), .A2(n6288), .ZN(n8489) );
  OR2_X1 U7918 ( .A1(n6344), .A2(n8489), .ZN(n6290) );
  INV_X1 U7919 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8490) );
  OR2_X1 U7920 ( .A1(n7352), .A2(n8490), .ZN(n6289) );
  NAND4_X1 U7921 ( .A1(n6292), .A2(n6291), .A3(n6290), .A4(n6289), .ZN(n8467)
         );
  XNOR2_X1 U7922 ( .A(n6293), .B(n8467), .ZN(n7891) );
  AND2_X1 U7923 ( .A1(n6293), .A2(n8497), .ZN(n6294) );
  NAND2_X1 U7924 ( .A1(n7009), .A2(n8048), .ZN(n6299) );
  NAND2_X1 U7925 ( .A1(n6295), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6296) );
  XNOR2_X1 U7926 ( .A(n6296), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9931) );
  AOI22_X1 U7927 ( .A1(n9931), .A2(n6639), .B1(P1_DATAO_REG_15__SCAN_IN), .B2(
        n6451), .ZN(n6298) );
  XNOR2_X1 U7928 ( .A(n8631), .B(n6410), .ZN(n6307) );
  NAND2_X1 U7929 ( .A1(n6593), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6306) );
  INV_X1 U7930 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9940) );
  OR2_X1 U7931 ( .A1(n7352), .A2(n9940), .ZN(n6305) );
  INV_X1 U7932 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8545) );
  OR2_X1 U7933 ( .A1(n6429), .A2(n8545), .ZN(n6304) );
  INV_X1 U7934 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7935 ( .A1(n6301), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6302) );
  AND2_X1 U7936 ( .A1(n6314), .A2(n6302), .ZN(n8470) );
  OR2_X1 U7937 ( .A1(n6344), .A2(n8470), .ZN(n6303) );
  NAND4_X1 U7938 ( .A1(n6306), .A2(n6305), .A3(n6304), .A4(n6303), .ZN(n8480)
         );
  XNOR2_X1 U7939 ( .A(n6307), .B(n8480), .ZN(n7999) );
  NAND2_X1 U7940 ( .A1(n8000), .A2(n7999), .ZN(n7998) );
  INV_X1 U7941 ( .A(n6307), .ZN(n6308) );
  NAND2_X1 U7942 ( .A1(n6308), .A2(n8480), .ZN(n6309) );
  NAND2_X1 U7943 ( .A1(n7998), .A2(n6309), .ZN(n7931) );
  NAND2_X1 U7944 ( .A1(n7101), .A2(n8048), .ZN(n6313) );
  NAND2_X1 U7945 ( .A1(n6310), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6311) );
  XNOR2_X1 U7946 ( .A(n6311), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U7947 ( .A1(n6451), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9947), .B2(
        n6639), .ZN(n6312) );
  XNOR2_X1 U7948 ( .A(n8625), .B(n6410), .ZN(n6320) );
  NAND2_X1 U7949 ( .A1(n6593), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6319) );
  INV_X1 U7950 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8457) );
  OR2_X1 U7951 ( .A1(n7352), .A2(n8457), .ZN(n6318) );
  INV_X1 U7952 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8542) );
  OR2_X1 U7953 ( .A1(n6429), .A2(n8542), .ZN(n6317) );
  NAND2_X1 U7954 ( .A1(n6314), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6315) );
  AND2_X1 U7955 ( .A1(n6330), .A2(n6315), .ZN(n8458) );
  OR2_X1 U7956 ( .A1(n6344), .A2(n8458), .ZN(n6316) );
  NAND4_X1 U7957 ( .A1(n6319), .A2(n6318), .A3(n6317), .A4(n6316), .ZN(n8468)
         );
  XNOR2_X1 U7958 ( .A(n6320), .B(n8468), .ZN(n7930) );
  INV_X1 U7959 ( .A(n6320), .ZN(n6321) );
  NAND2_X1 U7960 ( .A1(n6321), .A2(n8468), .ZN(n6322) );
  NAND2_X1 U7961 ( .A1(n7257), .A2(n8048), .ZN(n6326) );
  INV_X1 U7962 ( .A(n6042), .ZN(n6323) );
  NAND2_X1 U7963 ( .A1(n6323), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6324) );
  XNOR2_X1 U7964 ( .A(n6324), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9965) );
  AOI22_X1 U7965 ( .A1(n6451), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9965), .B2(
        n6639), .ZN(n6325) );
  XNOR2_X1 U7966 ( .A(n8538), .B(n7829), .ZN(n6336) );
  NAND2_X1 U7967 ( .A1(n6593), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6335) );
  INV_X1 U7968 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9977) );
  OR2_X1 U7969 ( .A1(n7352), .A2(n9977), .ZN(n6334) );
  INV_X1 U7970 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6327) );
  OR2_X1 U7971 ( .A1(n6429), .A2(n6327), .ZN(n6333) );
  INV_X1 U7972 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U7973 ( .A1(n6330), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6331) );
  AND2_X1 U7974 ( .A1(n6345), .A2(n6331), .ZN(n8444) );
  OR2_X1 U7975 ( .A1(n6344), .A2(n8444), .ZN(n6332) );
  NAND4_X1 U7976 ( .A1(n6335), .A2(n6334), .A3(n6333), .A4(n6332), .ZN(n8454)
         );
  XNOR2_X1 U7977 ( .A(n6336), .B(n8454), .ZN(n7939) );
  INV_X1 U7978 ( .A(n6336), .ZN(n6337) );
  NAND2_X1 U7979 ( .A1(n6337), .A2(n8423), .ZN(n7972) );
  NAND2_X1 U7980 ( .A1(n7937), .A2(n7972), .ZN(n6351) );
  NAND2_X1 U7981 ( .A1(n7285), .A2(n8048), .ZN(n6343) );
  OR2_X1 U7982 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  AND2_X1 U7983 ( .A1(n6341), .A2(n6340), .ZN(n9467) );
  AOI22_X1 U7984 ( .A1(n4499), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9467), .B2(
        n6639), .ZN(n6342) );
  XNOR2_X1 U7985 ( .A(n6618), .B(n6410), .ZN(n6352) );
  NAND2_X1 U7986 ( .A1(n6345), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U7987 ( .A1(n6358), .A2(n6346), .ZN(n8429) );
  NAND2_X1 U7988 ( .A1(n6591), .A2(n8429), .ZN(n6350) );
  INV_X1 U7989 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8267) );
  OR2_X1 U7990 ( .A1(n7352), .A2(n8267), .ZN(n6349) );
  INV_X1 U7991 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8535) );
  OR2_X1 U7992 ( .A1(n6429), .A2(n8535), .ZN(n6348) );
  INV_X1 U7993 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8618) );
  OR2_X1 U7994 ( .A1(n7349), .A2(n8618), .ZN(n6347) );
  NAND4_X1 U7995 ( .A1(n6350), .A2(n6349), .A3(n6348), .A4(n6347), .ZN(n8437)
         );
  XNOR2_X1 U7996 ( .A(n6352), .B(n8437), .ZN(n7973) );
  NAND2_X1 U7997 ( .A1(n6352), .A2(n7907), .ZN(n6353) );
  NAND2_X1 U7998 ( .A1(n7304), .A2(n8048), .ZN(n6355) );
  AOI22_X1 U7999 ( .A1(n6451), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8279), .B2(
        n6639), .ZN(n6354) );
  XNOR2_X1 U8000 ( .A(n8612), .B(n6410), .ZN(n6364) );
  INV_X1 U8001 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8002 ( .A1(n6358), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U8003 ( .A1(n6367), .A2(n6359), .ZN(n8418) );
  NAND2_X1 U8004 ( .A1(n8418), .A2(n6591), .ZN(n6363) );
  INV_X1 U8005 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8417) );
  OR2_X1 U8006 ( .A1(n7352), .A2(n8417), .ZN(n6362) );
  INV_X1 U8007 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10295) );
  OR2_X1 U8008 ( .A1(n6429), .A2(n10295), .ZN(n6361) );
  NAND2_X1 U8009 ( .A1(n6593), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6360) );
  NAND4_X1 U8010 ( .A1(n6363), .A2(n6362), .A3(n6361), .A4(n6360), .ZN(n8405)
         );
  XNOR2_X1 U8011 ( .A(n6364), .B(n8405), .ZN(n7904) );
  NAND2_X1 U8012 ( .A1(n7302), .A2(n8048), .ZN(n6366) );
  NAND2_X1 U8013 ( .A1(n6451), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6365) );
  XNOR2_X1 U8014 ( .A(n8606), .B(n6410), .ZN(n6371) );
  INV_X1 U8015 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U8016 ( .A1(n6367), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U8017 ( .A1(n6377), .A2(n6368), .ZN(n8409) );
  NAND2_X1 U8018 ( .A1(n8409), .A2(n6591), .ZN(n6370) );
  AOI22_X1 U8019 ( .A1(n7347), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6593), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6369) );
  OAI211_X1 U8020 ( .C1(n7352), .C2(n8408), .A(n6370), .B(n6369), .ZN(n8415)
         );
  XNOR2_X1 U8021 ( .A(n6371), .B(n8415), .ZN(n7953) );
  NAND2_X1 U8022 ( .A1(n7954), .A2(n7953), .ZN(n6373) );
  INV_X1 U8023 ( .A(n8415), .ZN(n7915) );
  NAND2_X1 U8024 ( .A1(n6371), .A2(n7915), .ZN(n6372) );
  NAND2_X1 U8025 ( .A1(n6373), .A2(n6372), .ZN(n7912) );
  NAND2_X1 U8026 ( .A1(n7394), .A2(n8048), .ZN(n6375) );
  NAND2_X1 U8027 ( .A1(n4499), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6374) );
  XNOR2_X1 U8028 ( .A(n8600), .B(n6410), .ZN(n6381) );
  INV_X1 U8029 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8599) );
  INV_X1 U8030 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U8031 ( .A1(n6377), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U8032 ( .A1(n6386), .A2(n6378), .ZN(n8398) );
  NAND2_X1 U8033 ( .A1(n8398), .A2(n6591), .ZN(n6380) );
  AOI22_X1 U8034 ( .A1(n6133), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n7347), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n6379) );
  OAI211_X1 U8035 ( .C1(n7349), .C2(n8599), .A(n6380), .B(n6379), .ZN(n8406)
         );
  XNOR2_X1 U8036 ( .A(n6381), .B(n8406), .ZN(n7911) );
  NAND2_X1 U8037 ( .A1(n7912), .A2(n7911), .ZN(n6383) );
  INV_X1 U8038 ( .A(n8406), .ZN(n6574) );
  NAND2_X1 U8039 ( .A1(n6381), .A2(n6574), .ZN(n6382) );
  NAND2_X1 U8040 ( .A1(n6383), .A2(n6382), .ZN(n7963) );
  NAND2_X1 U8041 ( .A1(n7539), .A2(n8048), .ZN(n6385) );
  NAND2_X1 U8042 ( .A1(n6451), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6384) );
  XNOR2_X1 U8043 ( .A(n8594), .B(n6410), .ZN(n7961) );
  NAND2_X1 U8044 ( .A1(n6386), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U8045 ( .A1(n6401), .A2(n6387), .ZN(n8383) );
  NAND2_X1 U8046 ( .A1(n8383), .A2(n6591), .ZN(n6392) );
  INV_X1 U8047 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U8048 ( .A1(n7347), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U8049 ( .A1(n6593), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6388) );
  OAI211_X1 U8050 ( .C1(n8382), .C2(n7352), .A(n6389), .B(n6388), .ZN(n6390)
         );
  INV_X1 U8051 ( .A(n6390), .ZN(n6391) );
  AND2_X1 U8052 ( .A1(n7961), .A2(n7960), .ZN(n6395) );
  INV_X1 U8053 ( .A(n7961), .ZN(n6393) );
  NAND2_X1 U8054 ( .A1(n6393), .A2(n8395), .ZN(n6394) );
  OAI21_X2 U8055 ( .B1(n7963), .B2(n6395), .A(n6394), .ZN(n6399) );
  NAND2_X1 U8056 ( .A1(n7571), .A2(n8048), .ZN(n6397) );
  NAND2_X1 U8057 ( .A1(n4499), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6396) );
  XNOR2_X1 U8058 ( .A(n8588), .B(n7829), .ZN(n6398) );
  NAND2_X1 U8059 ( .A1(n6399), .A2(n6398), .ZN(n6400) );
  NAND2_X1 U8060 ( .A1(n6401), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U8061 ( .A1(n6412), .A2(n6402), .ZN(n8372) );
  NAND2_X1 U8062 ( .A1(n8372), .A2(n6591), .ZN(n6407) );
  INV_X1 U8063 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U8064 ( .A1(n6133), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U8065 ( .A1(n6593), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6403) );
  OAI211_X1 U8066 ( .C1(n6429), .C2(n10211), .A(n6404), .B(n6403), .ZN(n6405)
         );
  INV_X1 U8067 ( .A(n6405), .ZN(n6406) );
  NAND2_X1 U8068 ( .A1(n7661), .A2(n8048), .ZN(n6409) );
  NAND2_X1 U8069 ( .A1(n6451), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6408) );
  XNOR2_X1 U8070 ( .A(n6623), .B(n6410), .ZN(n6420) );
  INV_X1 U8071 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U8072 ( .A1(n6412), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U8073 ( .A1(n6427), .A2(n6413), .ZN(n8363) );
  NAND2_X1 U8074 ( .A1(n8363), .A2(n6591), .ZN(n6419) );
  INV_X1 U8075 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8076 ( .A1(n6593), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8077 ( .A1(n7347), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6414) );
  OAI211_X1 U8078 ( .C1(n7352), .C2(n6416), .A(n6415), .B(n6414), .ZN(n6417)
         );
  INV_X1 U8079 ( .A(n6417), .ZN(n6418) );
  NAND2_X1 U8080 ( .A1(n6420), .A2(n8347), .ZN(n7920) );
  INV_X1 U8081 ( .A(n6420), .ZN(n6421) );
  NAND2_X1 U8082 ( .A1(n6421), .A2(n8369), .ZN(n6422) );
  NAND2_X1 U8083 ( .A1(n7919), .A2(n7920), .ZN(n6438) );
  NAND2_X1 U8084 ( .A1(n7730), .A2(n8048), .ZN(n6424) );
  NAND2_X1 U8085 ( .A1(n4499), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6423) );
  XNOR2_X1 U8086 ( .A(n8172), .B(n6410), .ZN(n6435) );
  INV_X1 U8087 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U8088 ( .A1(n6427), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U8089 ( .A1(n6441), .A2(n6428), .ZN(n8349) );
  NAND2_X1 U8090 ( .A1(n8349), .A2(n6591), .ZN(n6434) );
  INV_X1 U8091 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8356) );
  NAND2_X1 U8092 ( .A1(n6593), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6431) );
  INV_X1 U8093 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10304) );
  OR2_X1 U8094 ( .A1(n6429), .A2(n10304), .ZN(n6430) );
  OAI211_X1 U8095 ( .C1(n7352), .C2(n8356), .A(n6431), .B(n6430), .ZN(n6432)
         );
  INV_X1 U8096 ( .A(n6432), .ZN(n6433) );
  NAND2_X1 U8097 ( .A1(n6435), .A2(n8332), .ZN(n7985) );
  INV_X1 U8098 ( .A(n6435), .ZN(n6436) );
  NAND2_X1 U8099 ( .A1(n6436), .A2(n8360), .ZN(n6437) );
  NAND2_X1 U8100 ( .A1(n6438), .A2(n7921), .ZN(n7923) );
  NAND2_X1 U8101 ( .A1(n7923), .A2(n7985), .ZN(n6448) );
  NAND2_X1 U8102 ( .A1(n7766), .A2(n8048), .ZN(n6440) );
  NAND2_X1 U8103 ( .A1(n6451), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6439) );
  XNOR2_X1 U8104 ( .A(n8340), .B(n6410), .ZN(n6449) );
  NAND2_X1 U8105 ( .A1(n6441), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8106 ( .A1(n8339), .A2(n6591), .ZN(n6447) );
  INV_X1 U8107 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U8108 ( .A1(n7347), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8109 ( .A1(n6593), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6443) );
  OAI211_X1 U8110 ( .C1(n8338), .C2(n7352), .A(n6444), .B(n6443), .ZN(n6445)
         );
  INV_X1 U8111 ( .A(n6445), .ZN(n6446) );
  XNOR2_X1 U8112 ( .A(n6449), .B(n8319), .ZN(n7986) );
  NAND2_X1 U8113 ( .A1(n6448), .A2(n7986), .ZN(n7989) );
  NAND2_X1 U8114 ( .A1(n6449), .A2(n8348), .ZN(n6450) );
  NAND2_X1 U8115 ( .A1(n7787), .A2(n8048), .ZN(n6453) );
  NAND2_X1 U8116 ( .A1(n6451), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6452) );
  XNOR2_X1 U8117 ( .A(n8511), .B(n7829), .ZN(n7828) );
  INV_X1 U8118 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U8119 ( .A1(n6456), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U8120 ( .A1(n6501), .A2(n6457), .ZN(n8325) );
  NAND2_X1 U8121 ( .A1(n8325), .A2(n6591), .ZN(n6462) );
  INV_X1 U8122 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8324) );
  NAND2_X1 U8123 ( .A1(n6593), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U8124 ( .A1(n7347), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6458) );
  OAI211_X1 U8125 ( .C1(n7352), .C2(n8324), .A(n6459), .B(n6458), .ZN(n6460)
         );
  INV_X1 U8126 ( .A(n6460), .ZN(n6461) );
  XNOR2_X1 U8127 ( .A(n7828), .B(n8297), .ZN(n6498) );
  NAND2_X1 U8128 ( .A1(n6463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U8129 ( .A1(n7732), .A2(n7767), .ZN(n6470) );
  INV_X1 U8130 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U8131 ( .A1(n6477), .A2(n6468), .ZN(n6469) );
  NAND2_X1 U8132 ( .A1(n6471), .A2(n6735), .ZN(n7111) );
  NOR2_X1 U8133 ( .A1(n6472), .A2(n7767), .ZN(n6473) );
  XNOR2_X1 U8134 ( .A(n6476), .B(n6475), .ZN(n6673) );
  NOR2_X1 U8135 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .ZN(
        n6481) );
  NOR4_X1 U8136 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6480) );
  NOR4_X1 U8137 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6479) );
  NOR4_X1 U8138 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6478) );
  NAND4_X1 U8139 ( .A1(n6481), .A2(n6480), .A3(n6479), .A4(n6478), .ZN(n6487)
         );
  NOR4_X1 U8140 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6485) );
  NOR4_X1 U8141 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6484) );
  NOR4_X1 U8142 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n6483) );
  NOR4_X1 U8143 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6482) );
  NAND4_X1 U8144 ( .A1(n6485), .A2(n6484), .A3(n6483), .A4(n6482), .ZN(n6486)
         );
  NOR2_X1 U8145 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  NOR2_X1 U8146 ( .A1(n6718), .A2(n6658), .ZN(n6489) );
  NAND2_X1 U8147 ( .A1(n6659), .A2(n6489), .ZN(n6649) );
  NAND2_X1 U8148 ( .A1(n7540), .A2(n8026), .ZN(n10057) );
  AND2_X1 U8149 ( .A1(n8182), .A2(n10057), .ZN(n6492) );
  NAND2_X1 U8150 ( .A1(n8218), .A2(n8279), .ZN(n6601) );
  NAND2_X1 U8151 ( .A1(n8026), .A2(n6661), .ZN(n6491) );
  OR2_X1 U8152 ( .A1(n6601), .A2(n6491), .ZN(n6647) );
  NAND2_X1 U8153 ( .A1(n6492), .A2(n6647), .ZN(n6515) );
  OR2_X1 U8154 ( .A1(n6649), .A2(n6515), .ZN(n6496) );
  INV_X1 U8155 ( .A(n6658), .ZN(n6493) );
  AND2_X1 U8156 ( .A1(n7111), .A2(n6493), .ZN(n6494) );
  NAND2_X1 U8157 ( .A1(n6494), .A2(n7109), .ZN(n6522) );
  NOR2_X1 U8158 ( .A1(n6522), .A2(n6718), .ZN(n6646) );
  INV_X1 U8159 ( .A(n6647), .ZN(n6517) );
  NAND2_X1 U8160 ( .A1(n6646), .A2(n6517), .ZN(n6495) );
  OR2_X1 U8161 ( .A1(n6649), .A2(n10057), .ZN(n6500) );
  AND2_X1 U8162 ( .A1(n8279), .A2(n8203), .ZN(n7116) );
  NAND2_X1 U8163 ( .A1(n7540), .A2(n7116), .ZN(n10046) );
  OR2_X1 U8164 ( .A1(n10046), .A2(n8064), .ZN(n6663) );
  NAND2_X1 U8165 ( .A1(n8511), .A2(n7968), .ZN(n6529) );
  NAND2_X1 U8166 ( .A1(n6501), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U8167 ( .A1(n7822), .A2(n6502), .ZN(n8303) );
  NAND2_X1 U8168 ( .A1(n8303), .A2(n6591), .ZN(n6507) );
  INV_X1 U8169 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U8170 ( .A1(n6593), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U8171 ( .A1(n7347), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6503) );
  OAI211_X1 U8172 ( .C1(n7352), .C2(n8302), .A(n6504), .B(n6503), .ZN(n6505)
         );
  INV_X1 U8173 ( .A(n6505), .ZN(n6506) );
  INV_X1 U8174 ( .A(n8320), .ZN(n6627) );
  INV_X1 U8175 ( .A(n6646), .ZN(n6509) );
  INV_X1 U8176 ( .A(n6518), .ZN(n6508) );
  NAND2_X1 U8177 ( .A1(n8199), .A2(n6508), .ZN(n7209) );
  NOR2_X1 U8178 ( .A1(n6509), .A2(n7209), .ZN(n6514) );
  NAND2_X1 U8179 ( .A1(n4529), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6510) );
  XNOR2_X1 U8180 ( .A(n6510), .B(P2_IR_REG_28__SCAN_IN), .ZN(n8215) );
  MUX2_X1 U8181 ( .A(n6511), .B(P2_IR_REG_31__SCAN_IN), .S(n5028), .Z(n6512)
         );
  INV_X1 U8182 ( .A(n8273), .ZN(n6766) );
  NAND2_X1 U8183 ( .A1(n8215), .A2(n6766), .ZN(n6513) );
  NAND2_X1 U8184 ( .A1(n6513), .A2(n6675), .ZN(n6632) );
  AND2_X2 U8185 ( .A1(n6514), .A2(n6632), .ZN(n7979) );
  INV_X1 U8186 ( .A(n7979), .ZN(n8002) );
  INV_X1 U8187 ( .A(n6632), .ZN(n6637) );
  NAND2_X1 U8188 ( .A1(n6514), .A2(n6637), .ZN(n7981) );
  AOI22_X1 U8189 ( .A1(n8319), .A2(n8006), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6526) );
  INV_X1 U8190 ( .A(n6659), .ZN(n6516) );
  NAND2_X1 U8191 ( .A1(n6515), .A2(n9987), .ZN(n6645) );
  OAI21_X1 U8192 ( .B1(n6516), .B2(n6658), .A(n6645), .ZN(n6520) );
  NAND2_X1 U8193 ( .A1(n6522), .A2(n6517), .ZN(n6519) );
  NAND2_X1 U8194 ( .A1(n8199), .A2(n6518), .ZN(n6656) );
  NAND4_X1 U8195 ( .A1(n6520), .A2(n6776), .A3(n6519), .A4(n6656), .ZN(n6521)
         );
  NAND2_X1 U8196 ( .A1(n6521), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6524) );
  NOR2_X1 U8197 ( .A1(n6718), .A2(n7209), .ZN(n8216) );
  NAND2_X1 U8198 ( .A1(n8216), .A2(n6522), .ZN(n6523) );
  NAND2_X1 U8199 ( .A1(n6524), .A2(n6523), .ZN(n6931) );
  INV_X1 U8200 ( .A(n6673), .ZN(n6775) );
  AND2_X1 U8201 ( .A1(n6775), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8214) );
  NAND2_X1 U8202 ( .A1(n8325), .A2(n7994), .ZN(n6525) );
  OAI211_X1 U8203 ( .C1(n6627), .C2(n8002), .A(n6526), .B(n6525), .ZN(n6527)
         );
  INV_X1 U8204 ( .A(n6527), .ZN(n6528) );
  OAI21_X1 U8205 ( .B1(n6533), .B2(n5059), .A(n8777), .ZN(n6538) );
  NAND2_X1 U8206 ( .A1(n9352), .A2(n8769), .ZN(n6537) );
  AOI22_X1 U8207 ( .A1(n8768), .A2(n9171), .B1(n8767), .B2(n9199), .ZN(n6535)
         );
  AOI22_X1 U8208 ( .A1(n6010), .A2(n9168), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6534) );
  AND2_X1 U8209 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  NAND3_X1 U8210 ( .A1(n6538), .A2(n6537), .A3(n6536), .ZN(P1_U3214) );
  INV_X1 U8211 ( .A(n6783), .ZN(n6539) );
  NAND2_X1 U8212 ( .A1(n6541), .A2(n9802), .ZN(n6543) );
  NAND2_X1 U8213 ( .A1(n6543), .A2(n6542), .ZN(P1_U3519) );
  INV_X1 U8214 ( .A(n7748), .ZN(n10058) );
  INV_X1 U8215 ( .A(n10032), .ZN(n7217) );
  INV_X1 U8216 ( .A(n6549), .ZN(n10007) );
  NAND2_X1 U8217 ( .A1(n7186), .A2(n7185), .ZN(n6552) );
  OR2_X1 U8218 ( .A1(n6550), .A2(n6549), .ZN(n6551) );
  NAND2_X1 U8219 ( .A1(n6552), .A2(n6551), .ZN(n9991) );
  NAND2_X1 U8220 ( .A1(n8232), .A2(n10013), .ZN(n8069) );
  OR2_X1 U8221 ( .A1(n8232), .A2(n6553), .ZN(n6554) );
  INV_X1 U8222 ( .A(n7194), .ZN(n10019) );
  AND2_X1 U8223 ( .A1(n9994), .A2(n10019), .ZN(n6555) );
  INV_X1 U8224 ( .A(n8095), .ZN(n10022) );
  NAND2_X1 U8225 ( .A1(n8096), .A2(n10022), .ZN(n6605) );
  OR2_X1 U8226 ( .A1(n8096), .A2(n10022), .ZN(n6606) );
  NAND2_X1 U8227 ( .A1(n6556), .A2(n6606), .ZN(n7117) );
  OR2_X1 U8228 ( .A1(n8230), .A2(n6607), .ZN(n6558) );
  AND2_X1 U8229 ( .A1(n8230), .A2(n6607), .ZN(n6557) );
  INV_X1 U8230 ( .A(n7153), .ZN(n10036) );
  INV_X1 U8231 ( .A(n7371), .ZN(n6563) );
  AOI21_X1 U8232 ( .B1(n7371), .B2(n8227), .A(n10044), .ZN(n6562) );
  INV_X1 U8233 ( .A(n8226), .ZN(n6564) );
  OR2_X1 U8234 ( .A1(n7552), .A2(n6564), .ZN(n8086) );
  NAND2_X1 U8235 ( .A1(n7552), .A2(n6564), .ZN(n8110) );
  INV_X1 U8236 ( .A(n7682), .ZN(n8225) );
  NOR2_X1 U8237 ( .A1(n7597), .A2(n8225), .ZN(n6565) );
  INV_X1 U8238 ( .A(n7597), .ZN(n10045) );
  AOI21_X1 U8239 ( .B1(n7680), .B2(n7679), .A(n6566), .ZN(n7744) );
  XNOR2_X1 U8240 ( .A(n8129), .B(n8127), .ZN(n8500) );
  INV_X1 U8241 ( .A(n8637), .ZN(n6569) );
  NOR2_X1 U8242 ( .A1(n6569), .A2(n8497), .ZN(n6570) );
  INV_X1 U8243 ( .A(n8480), .ZN(n6615) );
  INV_X1 U8244 ( .A(n8631), .ZN(n8010) );
  NAND2_X1 U8245 ( .A1(n8625), .A2(n8001), .ZN(n8136) );
  NAND2_X1 U8246 ( .A1(n8146), .A2(n8136), .ZN(n8452) );
  INV_X1 U8247 ( .A(n8625), .ZN(n7936) );
  OR2_X1 U8248 ( .A1(n8538), .A2(n8423), .ZN(n8150) );
  NAND2_X1 U8249 ( .A1(n8538), .A2(n8423), .ZN(n8139) );
  NAND2_X1 U8250 ( .A1(n8150), .A2(n8139), .ZN(n8435) );
  INV_X1 U8251 ( .A(n8538), .ZN(n8443) );
  NAND2_X1 U8252 ( .A1(n8434), .A2(n5072), .ZN(n8421) );
  OAI21_X1 U8253 ( .B1(n6618), .B2(n8437), .A(n8421), .ZN(n6571) );
  NAND2_X1 U8254 ( .A1(n8612), .A2(n8424), .ZN(n8156) );
  NAND2_X1 U8255 ( .A1(n8154), .A2(n8156), .ZN(n6620) );
  NAND2_X1 U8256 ( .A1(n8606), .A2(n7915), .ZN(n8387) );
  NAND2_X1 U8257 ( .A1(n8058), .A2(n8387), .ZN(n8403) );
  INV_X1 U8258 ( .A(n8606), .ZN(n6573) );
  NAND2_X1 U8259 ( .A1(n6573), .A2(n7915), .ZN(n8391) );
  NAND2_X1 U8260 ( .A1(n8600), .A2(n6574), .ZN(n8164) );
  NOR2_X1 U8261 ( .A1(n8600), .A2(n8406), .ZN(n8377) );
  NAND2_X1 U8262 ( .A1(n8594), .A2(n7960), .ZN(n8056) );
  NAND2_X1 U8263 ( .A1(n8168), .A2(n8056), .ZN(n8376) );
  OAI21_X1 U8264 ( .B1(n8594), .B2(n8395), .A(n8379), .ZN(n8368) );
  INV_X1 U8265 ( .A(n8588), .ZN(n6575) );
  NAND2_X1 U8266 ( .A1(n8368), .A2(n5071), .ZN(n6577) );
  NAND2_X1 U8267 ( .A1(n8172), .A2(n8332), .ZN(n8179) );
  NOR2_X1 U8268 ( .A1(n8511), .A2(n8297), .ZN(n6580) );
  NAND2_X1 U8269 ( .A1(n8340), .A2(n8319), .ZN(n8313) );
  NOR2_X1 U8270 ( .A1(n6580), .A2(n8313), .ZN(n6583) );
  OR2_X1 U8271 ( .A1(n8352), .A2(n6583), .ZN(n8309) );
  OR2_X1 U8272 ( .A1(n8309), .A2(n5086), .ZN(n6578) );
  NAND2_X1 U8273 ( .A1(n8576), .A2(n8332), .ZN(n8329) );
  NAND2_X1 U8274 ( .A1(n8571), .A2(n8348), .ZN(n6579) );
  AND2_X1 U8275 ( .A1(n8329), .A2(n6579), .ZN(n8312) );
  INV_X1 U8276 ( .A(n6580), .ZN(n6581) );
  AND2_X1 U8277 ( .A1(n8312), .A2(n6581), .ZN(n6582) );
  OR2_X1 U8278 ( .A1(n6583), .A2(n6582), .ZN(n8310) );
  NOR2_X1 U8279 ( .A1(n5086), .A2(n8310), .ZN(n6584) );
  NAND2_X1 U8280 ( .A1(n7808), .A2(n8048), .ZN(n6586) );
  NAND2_X1 U8281 ( .A1(n6451), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6585) );
  INV_X1 U8282 ( .A(n8304), .ZN(n8561) );
  NAND2_X1 U8283 ( .A1(n8561), .A2(n6627), .ZN(n6588) );
  AOI21_X1 U8284 ( .B1(n8295), .B2(n6588), .A(n6587), .ZN(n6600) );
  NAND2_X1 U8285 ( .A1(n7848), .A2(n8048), .ZN(n6590) );
  NAND2_X1 U8286 ( .A1(n4499), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6589) );
  INV_X1 U8287 ( .A(n7822), .ZN(n6592) );
  NAND2_X1 U8288 ( .A1(n6592), .A2(n6591), .ZN(n7355) );
  INV_X1 U8289 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U8290 ( .A1(n7347), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U8291 ( .A1(n6593), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6594) );
  OAI211_X1 U8292 ( .C1(n6596), .C2(n7352), .A(n6595), .B(n6594), .ZN(n6597)
         );
  INV_X1 U8293 ( .A(n6597), .ZN(n6598) );
  NAND2_X1 U8294 ( .A1(n7355), .A2(n6598), .ZN(n8298) );
  INV_X1 U8295 ( .A(n8298), .ZN(n6599) );
  NAND2_X1 U8296 ( .A1(n6654), .A2(n6599), .ZN(n8193) );
  NAND2_X1 U8297 ( .A1(n8064), .A2(n6661), .ZN(n8209) );
  NAND2_X1 U8298 ( .A1(n8024), .A2(n7179), .ZN(n7181) );
  NAND2_X1 U8299 ( .A1(n7181), .A2(n8067), .ZN(n9986) );
  NAND2_X1 U8300 ( .A1(n9994), .A2(n7194), .ZN(n8098) );
  AND2_X1 U8301 ( .A1(n8074), .A2(n8098), .ZN(n8023) );
  INV_X1 U8302 ( .A(n6604), .ZN(n7202) );
  NAND2_X1 U8303 ( .A1(n6606), .A2(n6605), .ZN(n8073) );
  NAND2_X1 U8304 ( .A1(n7202), .A2(n8073), .ZN(n7201) );
  NAND2_X1 U8305 ( .A1(n8096), .A2(n8095), .ZN(n8076) );
  INV_X1 U8306 ( .A(n6607), .ZN(n10026) );
  NAND2_X1 U8307 ( .A1(n8230), .A2(n10026), .ZN(n8094) );
  NAND2_X1 U8308 ( .A1(n7106), .A2(n8094), .ZN(n7223) );
  OR2_X1 U8309 ( .A1(n8230), .A2(n10026), .ZN(n8075) );
  OR2_X1 U8310 ( .A1(n8229), .A2(n10032), .ZN(n8079) );
  NAND2_X1 U8311 ( .A1(n8075), .A2(n8079), .ZN(n8102) );
  INV_X1 U8312 ( .A(n8102), .ZN(n6608) );
  NAND2_X1 U8313 ( .A1(n7223), .A2(n6608), .ZN(n7275) );
  NAND2_X1 U8314 ( .A1(n8229), .A2(n10032), .ZN(n8100) );
  NAND2_X1 U8315 ( .A1(n7275), .A2(n8100), .ZN(n6610) );
  OR2_X1 U8316 ( .A1(n6609), .A2(n7153), .ZN(n7374) );
  NAND2_X1 U8317 ( .A1(n6609), .A2(n7153), .ZN(n8105) );
  OR2_X1 U8318 ( .A1(n10044), .A2(n7549), .ZN(n8085) );
  AND2_X1 U8319 ( .A1(n8085), .A2(n7374), .ZN(n8082) );
  NAND2_X1 U8320 ( .A1(n10044), .A2(n7549), .ZN(n8104) );
  OR2_X1 U8321 ( .A1(n7597), .A2(n7682), .ZN(n8114) );
  AND2_X1 U8322 ( .A1(n8114), .A2(n8086), .ZN(n8089) );
  NAND2_X1 U8323 ( .A1(n7587), .A2(n8089), .ZN(n6611) );
  NAND2_X1 U8324 ( .A1(n7597), .A2(n7682), .ZN(n8111) );
  NAND2_X1 U8325 ( .A1(n6611), .A2(n8111), .ZN(n7678) );
  INV_X1 U8326 ( .A(n7679), .ZN(n8037) );
  NAND2_X1 U8327 ( .A1(n7678), .A2(n8037), .ZN(n6612) );
  NAND2_X1 U8328 ( .A1(n6612), .A2(n8091), .ZN(n7742) );
  OR2_X1 U8329 ( .A1(n7748), .A2(n8496), .ZN(n8123) );
  NAND2_X1 U8330 ( .A1(n7748), .A2(n8496), .ZN(n8124) );
  NAND2_X1 U8331 ( .A1(n8123), .A2(n8124), .ZN(n7743) );
  OAI21_X2 U8332 ( .B1(n7742), .B2(n7743), .A(n8123), .ZN(n8501) );
  NOR2_X1 U8333 ( .A1(n8129), .A2(n8127), .ZN(n6613) );
  NAND2_X1 U8334 ( .A1(n8129), .A2(n8127), .ZN(n6614) );
  OR2_X1 U8335 ( .A1(n8637), .A2(n8497), .ZN(n8130) );
  NAND2_X1 U8336 ( .A1(n8637), .A2(n8497), .ZN(n8131) );
  OR2_X1 U8337 ( .A1(n8631), .A2(n6615), .ZN(n8135) );
  NAND2_X1 U8338 ( .A1(n8631), .A2(n6615), .ZN(n8448) );
  AND2_X1 U8339 ( .A1(n8136), .A2(n8448), .ZN(n8144) );
  INV_X1 U8340 ( .A(n8146), .ZN(n6616) );
  NAND2_X1 U8341 ( .A1(n6618), .A2(n7907), .ZN(n8140) );
  NAND2_X1 U8342 ( .A1(n8151), .A2(n8140), .ZN(n8428) );
  AND2_X1 U8343 ( .A1(n8164), .A2(n8387), .ZN(n8059) );
  NAND2_X1 U8344 ( .A1(n8588), .A2(n7966), .ZN(n8169) );
  AND2_X1 U8345 ( .A1(n6623), .A2(n8347), .ZN(n8022) );
  NOR2_X1 U8346 ( .A1(n8340), .A2(n8348), .ZN(n8053) );
  NAND2_X1 U8347 ( .A1(n8294), .A2(n8296), .ZN(n6629) );
  OR2_X1 U8348 ( .A1(n8304), .A2(n6627), .ZN(n6628) );
  NAND2_X1 U8349 ( .A1(n6629), .A2(n6628), .ZN(n8204) );
  XNOR2_X2 U8350 ( .A(n8204), .B(n8188), .ZN(n6644) );
  OAI211_X1 U8351 ( .C1(n8218), .C2(n8203), .A(n10057), .B(n8251), .ZN(n6630)
         );
  INV_X1 U8352 ( .A(n6630), .ZN(n6631) );
  NAND2_X1 U8353 ( .A1(n6631), .A2(n7209), .ZN(n9992) );
  INV_X1 U8354 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U8355 ( .A1(n7347), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6634) );
  INV_X1 U8356 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10335) );
  OR2_X1 U8357 ( .A1(n7349), .A2(n10335), .ZN(n6633) );
  OAI211_X1 U8358 ( .C1(n7352), .C2(n8293), .A(n6634), .B(n6633), .ZN(n6635)
         );
  INV_X1 U8359 ( .A(n6635), .ZN(n6636) );
  NAND2_X1 U8360 ( .A1(n7355), .A2(n6636), .ZN(n8222) );
  NOR2_X1 U8361 ( .A1(n6639), .A2(n6638), .ZN(n6640) );
  NOR2_X1 U8362 ( .A1(n9993), .A2(n6640), .ZN(n8285) );
  AOI22_X1 U8363 ( .A1(n8481), .A2(n8320), .B1(n8222), .B2(n8285), .ZN(n6641)
         );
  OAI21_X1 U8364 ( .B1(n6644), .B2(n9992), .A(n6641), .ZN(n6642) );
  NAND2_X1 U8365 ( .A1(n6646), .A2(n6645), .ZN(n6651) );
  AND2_X1 U8366 ( .A1(n7209), .A2(n6647), .ZN(n6648) );
  INV_X1 U8367 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6652) );
  NAND2_X1 U8368 ( .A1(n10065), .A2(n6652), .ZN(n6653) );
  NAND2_X1 U8369 ( .A1(n6655), .A2(n5078), .ZN(P2_U3456) );
  INV_X1 U8370 ( .A(n6656), .ZN(n6657) );
  OR2_X1 U8371 ( .A1(n6658), .A2(n6657), .ZN(n6660) );
  NAND3_X1 U8372 ( .A1(n8218), .A2(n6661), .A3(n8251), .ZN(n6662) );
  NAND2_X1 U8373 ( .A1(n8182), .A2(n6662), .ZN(n7110) );
  NAND2_X1 U8374 ( .A1(n7109), .A2(n7110), .ZN(n6666) );
  INV_X1 U8375 ( .A(n6663), .ZN(n6664) );
  INV_X1 U8376 ( .A(n7110), .ZN(n7108) );
  OAI21_X1 U8377 ( .B1(n7111), .B2(n6664), .A(n7108), .ZN(n6665) );
  NAND2_X1 U8378 ( .A1(n6666), .A2(n6665), .ZN(n6667) );
  NOR2_X4 U8379 ( .A1(n7107), .A2(n6667), .ZN(n10081) );
  INV_X1 U8380 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U8381 ( .A1(n10079), .A2(n6669), .ZN(n6670) );
  NAND2_X1 U8382 ( .A1(n6671), .A2(n6670), .ZN(n6672) );
  INV_X1 U8383 ( .A(n10057), .ZN(n10055) );
  NAND2_X1 U8384 ( .A1(n6672), .A2(n5070), .ZN(P2_U3488) );
  INV_X1 U8385 ( .A(n6737), .ZN(n6930) );
  OR2_X2 U8386 ( .A1(n6776), .A2(n6930), .ZN(n8233) );
  NAND2_X1 U8387 ( .A1(n6776), .A2(n8182), .ZN(n6674) );
  NAND2_X1 U8388 ( .A1(n6674), .A2(n6673), .ZN(n6771) );
  NAND2_X1 U8389 ( .A1(n6771), .A2(n6675), .ZN(n6676) );
  NAND2_X1 U8390 ( .A1(n6676), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U8391 ( .A1(n6677), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6679) );
  INV_X2 U8392 ( .A(n9051), .ZN(P1_U3973) );
  INV_X1 U8393 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6681) );
  AND2_X1 U8394 ( .A1(n7856), .A2(P2_U3151), .ZN(n8647) );
  INV_X1 U8395 ( .A(n8647), .ZN(n7863) );
  OAI222_X1 U8396 ( .A1(n8650), .A2(n6682), .B1(n6846), .B2(P2_U3151), .C1(
        n6681), .C2(n7863), .ZN(P2_U3293) );
  OAI222_X1 U8397 ( .A1(n7863), .A2(n5088), .B1(n6805), .B2(P2_U3151), .C1(
        n8650), .C2(n6684), .ZN(P2_U3294) );
  NOR2_X1 U8398 ( .A1(n7856), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9455) );
  INV_X2 U8399 ( .A(n9455), .ZN(n7889) );
  AND2_X1 U8400 ( .A1(n7856), .A2(P1_U3086), .ZN(n7570) );
  INV_X2 U8401 ( .A(n7570), .ZN(n9457) );
  OAI222_X1 U8402 ( .A1(n7889), .A2(n6683), .B1(n9457), .B2(n6682), .C1(n7072), 
        .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U8403 ( .A1(n7889), .A2(n5002), .B1(n9457), .B2(n6684), .C1(n7073), 
        .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U8404 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6685) );
  OAI222_X1 U8405 ( .A1(n8650), .A2(n6686), .B1(n6849), .B2(P2_U3151), .C1(
        n6685), .C2(n7863), .ZN(P2_U3292) );
  OAI222_X1 U8406 ( .A1(n7889), .A2(n6687), .B1(n9457), .B2(n6686), .C1(n7076), 
        .C2(P1_U3086), .ZN(P1_U3352) );
  INV_X1 U8407 ( .A(n6688), .ZN(n6691) );
  INV_X1 U8408 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6689) );
  OAI222_X1 U8409 ( .A1(n8650), .A2(n6691), .B1(n9863), .B2(P2_U3151), .C1(
        n6689), .C2(n7863), .ZN(P2_U3291) );
  OAI222_X1 U8410 ( .A1(n7889), .A2(n6692), .B1(n9457), .B2(n6691), .C1(n6690), 
        .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U8411 ( .A(n9888), .ZN(n6853) );
  INV_X1 U8412 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6693) );
  OAI222_X1 U8413 ( .A1(n8650), .A2(n6694), .B1(n6853), .B2(P2_U3151), .C1(
        n6693), .C2(n7863), .ZN(P2_U3290) );
  INV_X1 U8414 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6695) );
  INV_X1 U8415 ( .A(n7082), .ZN(n9566) );
  OAI222_X1 U8416 ( .A1(n7889), .A2(n6695), .B1(n9457), .B2(n6694), .C1(n9566), 
        .C2(P1_U3086), .ZN(P1_U3350) );
  AOI22_X1 U8417 ( .A1(n6917), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n8647), .ZN(n6696) );
  OAI21_X1 U8418 ( .B1(n6697), .B2(n8650), .A(n6696), .ZN(P2_U3289) );
  INV_X1 U8419 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10390) );
  INV_X1 U8420 ( .A(n7084), .ZN(n9580) );
  OAI222_X1 U8421 ( .A1(n7889), .A2(n10390), .B1(n9457), .B2(n6697), .C1(n9580), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U8422 ( .A(n6698), .ZN(n6699) );
  NAND2_X1 U8423 ( .A1(n9681), .A2(n6700), .ZN(n6701) );
  OAI21_X1 U8424 ( .B1(n9681), .B2(n6702), .A(n6701), .ZN(P1_U3440) );
  INV_X1 U8425 ( .A(n7016), .ZN(n7027) );
  INV_X1 U8426 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10186) );
  OAI222_X1 U8427 ( .A1(n8650), .A2(n6703), .B1(n7027), .B2(P2_U3151), .C1(
        n10186), .C2(n7863), .ZN(P2_U3288) );
  INV_X1 U8428 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6704) );
  INV_X1 U8429 ( .A(n7087), .ZN(n9503) );
  OAI222_X1 U8430 ( .A1(n7889), .A2(n6704), .B1(n9457), .B2(n6703), .C1(n9503), 
        .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U8431 ( .A(n9024), .ZN(n9034) );
  NAND2_X1 U8432 ( .A1(n9034), .A2(n6705), .ZN(n6751) );
  NAND2_X1 U8433 ( .A1(n6706), .A2(n9017), .ZN(n6708) );
  NAND2_X1 U8434 ( .A1(n6708), .A2(n6707), .ZN(n6749) );
  NAND2_X1 U8435 ( .A1(n6751), .A2(n6749), .ZN(n9604) );
  INV_X1 U8436 ( .A(n9604), .ZN(n9553) );
  NOR2_X1 U8437 ( .A1(n9553), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8438 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10350) );
  INV_X1 U8439 ( .A(n6709), .ZN(n6710) );
  INV_X1 U8440 ( .A(n7090), .ZN(n9519) );
  OAI222_X1 U8441 ( .A1(n7889), .A2(n10350), .B1(n9457), .B2(n6710), .C1(
        P1_U3086), .C2(n9519), .ZN(P1_U3347) );
  INV_X1 U8442 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6711) );
  INV_X1 U8443 ( .A(n7035), .ZN(n7322) );
  OAI222_X1 U8444 ( .A1(n7863), .A2(n6711), .B1(n8650), .B2(n6710), .C1(
        P2_U3151), .C2(n7322), .ZN(P2_U3287) );
  NAND2_X1 U8445 ( .A1(n6712), .A2(P1_U3973), .ZN(n6713) );
  OAI21_X1 U8446 ( .B1(P1_U3973), .B2(n6086), .A(n6713), .ZN(P1_U3554) );
  NAND2_X1 U8447 ( .A1(n9051), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6714) );
  OAI21_X1 U8448 ( .B1(n8965), .B2(n9051), .A(n6714), .ZN(P1_U3584) );
  AOI22_X1 U8449 ( .A1(n9489), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9455), .ZN(n6715) );
  OAI21_X1 U8450 ( .B1(n6717), .B2(n9457), .A(n6715), .ZN(P1_U3345) );
  INV_X1 U8451 ( .A(n7445), .ZN(n7473) );
  INV_X1 U8452 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6716) );
  OAI222_X1 U8453 ( .A1(n8650), .A2(n6717), .B1(n7473), .B2(P2_U3151), .C1(
        n6716), .C2(n7863), .ZN(P2_U3285) );
  INV_X1 U8454 ( .A(n6718), .ZN(n6734) );
  INV_X1 U8455 ( .A(n7109), .ZN(n6719) );
  NAND2_X1 U8456 ( .A1(n6734), .A2(n6719), .ZN(n6720) );
  OAI21_X1 U8457 ( .B1(n6734), .B2(n6468), .A(n6720), .ZN(P2_U3377) );
  INV_X1 U8458 ( .A(n6721), .ZN(n6729) );
  INV_X1 U8459 ( .A(n7339), .ZN(n7429) );
  OAI222_X1 U8460 ( .A1(n8650), .A2(n6729), .B1(n7429), .B2(P2_U3151), .C1(
        n6731), .C2(n7863), .ZN(P2_U3286) );
  INV_X1 U8461 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6728) );
  INV_X1 U8462 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U8463 ( .A1(n5647), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U8464 ( .A1(n6722), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6723) );
  OAI211_X1 U8465 ( .C1(n6726), .C2(n6725), .A(n6724), .B(n6723), .ZN(n8983)
         );
  NAND2_X1 U8466 ( .A1(n8983), .A2(P1_U3973), .ZN(n6727) );
  OAI21_X1 U8467 ( .B1(P1_U3973), .B2(n6728), .A(n6727), .ZN(P1_U3585) );
  INV_X1 U8468 ( .A(n9108), .ZN(n6730) );
  OAI222_X1 U8469 ( .A1(n7889), .A2(n10251), .B1(P1_U3086), .B2(n6730), .C1(
        n6729), .C2(n9457), .ZN(P1_U3346) );
  MUX2_X1 U8470 ( .A(n6731), .B(n9747), .S(P1_U3973), .Z(n6732) );
  INV_X1 U8471 ( .A(n6732), .ZN(P1_U3563) );
  INV_X1 U8472 ( .A(n6735), .ZN(n6736) );
  AOI22_X1 U8473 ( .A1(n10105), .A2(n10318), .B1(n6737), .B2(n6736), .ZN(
        P2_U3376) );
  INV_X1 U8474 ( .A(n6738), .ZN(n6741) );
  AOI22_X1 U8475 ( .A1(n9585), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9455), .ZN(n6739) );
  OAI21_X1 U8476 ( .B1(n6741), .B2(n9457), .A(n6739), .ZN(P1_U3344) );
  NAND2_X1 U8477 ( .A1(P2_U3893), .A2(n7187), .ZN(n6740) );
  OAI21_X1 U8478 ( .B1(P2_U3893), .B2(n5219), .A(n6740), .ZN(P2_U3491) );
  AND2_X1 U8479 ( .A1(n10105), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8480 ( .A1(n10105), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8481 ( .A1(n10105), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8482 ( .A1(n10105), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8483 ( .A1(n10105), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8484 ( .A1(n10105), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8485 ( .A1(n10105), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8486 ( .A1(n10105), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8487 ( .A1(n10105), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8488 ( .A1(n10105), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8489 ( .A1(n10105), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8490 ( .A1(n10105), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8491 ( .A1(n10105), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8492 ( .A1(n10105), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8493 ( .A1(n10105), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8494 ( .A1(n10105), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8495 ( .A1(n10105), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8496 ( .A1(n10105), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8497 ( .A1(n10105), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8498 ( .A1(n10105), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  INV_X1 U8499 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10363) );
  INV_X1 U8500 ( .A(n7613), .ZN(n7604) );
  OAI222_X1 U8501 ( .A1(n7863), .A2(n10363), .B1(n8650), .B2(n6741), .C1(
        P2_U3151), .C2(n7604), .ZN(P2_U3284) );
  INV_X1 U8502 ( .A(n8244), .ZN(n8236) );
  INV_X1 U8503 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6742) );
  OAI222_X1 U8504 ( .A1(n8650), .A2(n6743), .B1(n8236), .B2(P2_U3151), .C1(
        n6742), .C2(n7863), .ZN(P2_U3283) );
  INV_X1 U8505 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6744) );
  OAI222_X1 U8506 ( .A1(n7889), .A2(n6744), .B1(n9457), .B2(n6743), .C1(n7097), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8507 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10196) );
  NOR2_X1 U8508 ( .A1(n6748), .A2(n10196), .ZN(P2_U3256) );
  INV_X1 U8509 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10315) );
  NOR2_X1 U8510 ( .A1(n6748), .A2(n10315), .ZN(P2_U3248) );
  INV_X1 U8511 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6745) );
  NOR2_X1 U8512 ( .A1(n6748), .A2(n6745), .ZN(P2_U3262) );
  INV_X1 U8513 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10242) );
  NOR2_X1 U8514 ( .A1(n6748), .A2(n10242), .ZN(P2_U3259) );
  INV_X1 U8515 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6746) );
  NOR2_X1 U8516 ( .A1(n6748), .A2(n6746), .ZN(P2_U3257) );
  INV_X1 U8517 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10237) );
  NOR2_X1 U8518 ( .A1(n6748), .A2(n10237), .ZN(P2_U3242) );
  INV_X1 U8519 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6747) );
  NOR2_X1 U8520 ( .A1(n6748), .A2(n6747), .ZN(P2_U3263) );
  INV_X1 U8521 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10392) );
  NOR2_X1 U8522 ( .A1(n6748), .A2(n10392), .ZN(P2_U3236) );
  INV_X1 U8523 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10275) );
  NOR2_X1 U8524 ( .A1(n6748), .A2(n10275), .ZN(P2_U3235) );
  INV_X1 U8525 ( .A(n6749), .ZN(n6750) );
  NOR2_X1 U8526 ( .A1(n7867), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6752) );
  OR2_X1 U8527 ( .A1(n4502), .A2(n6752), .ZN(n9071) );
  AOI21_X1 U8528 ( .B1(n5770), .B2(n7867), .A(n9071), .ZN(n6753) );
  MUX2_X1 U8529 ( .A(n9071), .B(n6753), .S(n9072), .Z(n6758) );
  INV_X1 U8530 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6755) );
  INV_X1 U8531 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6754) );
  OAI22_X1 U8532 ( .A1(n9604), .A2(n6755), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6754), .ZN(n6757) );
  AND2_X1 U8533 ( .A1(n7067), .A2(n7867), .ZN(n9595) );
  AND3_X1 U8534 ( .A1(n9595), .A2(P1_IR_REG_0__SCAN_IN), .A3(n5770), .ZN(n6756) );
  AOI211_X1 U8535 ( .C1(n7067), .C2(n6758), .A(n6757), .B(n6756), .ZN(n6759)
         );
  INV_X1 U8536 ( .A(n6759), .ZN(P1_U3243) );
  XOR2_X1 U8537 ( .A(n6760), .B(n6761), .Z(n9068) );
  NAND2_X1 U8538 ( .A1(n9068), .A2(n8777), .ZN(n6765) );
  INV_X1 U8539 ( .A(n6762), .ZN(n6763) );
  NAND2_X1 U8540 ( .A1(n6763), .A2(n6784), .ZN(n7844) );
  AOI22_X1 U8541 ( .A1(n7844), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9683), .B2(
        n8769), .ZN(n6764) );
  OAI211_X1 U8542 ( .C1(n6795), .C2(n8780), .A(n6765), .B(n6764), .ZN(P1_U3232) );
  NAND2_X1 U8543 ( .A1(n6766), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7789) );
  NOR2_X1 U8544 ( .A1(n7789), .A2(n8215), .ZN(n6767) );
  NAND2_X1 U8545 ( .A1(n6771), .A2(n6767), .ZN(n6770) );
  INV_X1 U8546 ( .A(n8215), .ZN(n6768) );
  OR2_X1 U8547 ( .A1(n8233), .A2(n6768), .ZN(n6769) );
  INV_X1 U8548 ( .A(n9964), .ZN(n9864) );
  AND2_X1 U8549 ( .A1(n8215), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7809) );
  INV_X1 U8550 ( .A(n6803), .ZN(n6798) );
  AOI21_X1 U8551 ( .B1(n6806), .B2(n6772), .A(n9837), .ZN(n6773) );
  AOI21_X1 U8552 ( .B1(n6798), .B2(n9875), .A(n6773), .ZN(n6774) );
  AOI21_X1 U8553 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6774), .ZN(
        n6779) );
  NOR2_X1 U8554 ( .A1(n6776), .A2(n6775), .ZN(n6777) );
  INV_X1 U8555 ( .A(n9897), .ZN(n9966) );
  NAND2_X1 U8556 ( .A1(n9966), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n6778) );
  OAI211_X1 U8557 ( .C1(n9864), .C2(n6806), .A(n6779), .B(n6778), .ZN(P2_U3182) );
  INV_X1 U8558 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6780) );
  OAI222_X1 U8559 ( .A1(n8650), .A2(n6781), .B1(n4923), .B2(P2_U3151), .C1(
        n6780), .C2(n7863), .ZN(P2_U3282) );
  INV_X1 U8560 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10199) );
  INV_X1 U8561 ( .A(n7312), .ZN(n7253) );
  OAI222_X1 U8562 ( .A1(n7889), .A2(n10199), .B1(n9457), .B2(n6781), .C1(n7253), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U8563 ( .A(n6782), .ZN(n6785) );
  NAND3_X1 U8564 ( .A1(n6785), .A2(n6784), .A3(n6783), .ZN(n6792) );
  OR2_X1 U8565 ( .A1(n9666), .A2(n9789), .ZN(n7364) );
  INV_X1 U8566 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6786) );
  NOR2_X1 U8567 ( .A1(n9296), .A2(n6786), .ZN(n6790) );
  INV_X1 U8568 ( .A(n6876), .ZN(n6787) );
  NAND2_X1 U8569 ( .A1(n6712), .A2(n6889), .ZN(n8907) );
  NAND2_X1 U8570 ( .A1(n6787), .A2(n8907), .ZN(n9684) );
  AND3_X1 U8571 ( .A1(n9684), .A2(n6788), .A3(n9296), .ZN(n6789) );
  AOI211_X1 U8572 ( .C1(n9651), .C2(P1_REG3_REG_0__SCAN_IN), .A(n6790), .B(
        n6789), .ZN(n6794) );
  NOR2_X1 U8573 ( .A1(n9264), .A2(n9321), .ZN(n9282) );
  OAI21_X1 U8574 ( .B1(n9652), .B2(n9282), .A(n9683), .ZN(n6793) );
  OAI211_X1 U8575 ( .C1(n6795), .C2(n7364), .A(n6794), .B(n6793), .ZN(P1_U3293) );
  INV_X1 U8576 ( .A(n6805), .ZN(n9832) );
  INV_X1 U8577 ( .A(n6796), .ZN(n6797) );
  MUX2_X1 U8578 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8273), .Z(n6823) );
  INV_X1 U8579 ( .A(n6846), .ZN(n6819) );
  XNOR2_X1 U8580 ( .A(n6823), .B(n6819), .ZN(n6824) );
  XNOR2_X1 U8581 ( .A(n6825), .B(n6824), .ZN(n6822) );
  INV_X1 U8582 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7498) );
  INV_X1 U8583 ( .A(n9980), .ZN(n6924) );
  INV_X1 U8584 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10004) );
  MUX2_X1 U8585 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10004), .S(n6846), .Z(n6802)
         );
  AND2_X1 U8586 ( .A1(n6806), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6799) );
  NAND2_X1 U8587 ( .A1(n6070), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6800) );
  OAI21_X1 U8588 ( .B1(n6805), .B2(n6799), .A(n6800), .ZN(n9828) );
  OR2_X1 U8589 ( .A1(n9828), .A2(n7189), .ZN(n9830) );
  NAND2_X1 U8590 ( .A1(n9830), .A2(n6800), .ZN(n6801) );
  OAI21_X1 U8591 ( .B1(n6802), .B2(n6801), .A(n6848), .ZN(n6815) );
  MUX2_X1 U8592 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6804), .S(n6846), .Z(n6813)
         );
  NAND2_X1 U8593 ( .A1(n6070), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U8594 ( .A1(n6805), .A2(n6810), .ZN(n6809) );
  NAND2_X1 U8595 ( .A1(n6806), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6807) );
  OR2_X1 U8596 ( .A1(n6807), .A2(n6070), .ZN(n6808) );
  NAND2_X1 U8597 ( .A1(n6809), .A2(n6808), .ZN(n9826) );
  NAND2_X1 U8598 ( .A1(n9826), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6811) );
  NAND2_X1 U8599 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  NAND2_X1 U8600 ( .A1(n6813), .A2(n6812), .ZN(n6835) );
  OAI21_X1 U8601 ( .B1(n6813), .B2(n6812), .A(n6835), .ZN(n6814) );
  AOI22_X1 U8602 ( .A1(n6924), .A2(n6815), .B1(n9974), .B2(n6814), .ZN(n6816)
         );
  OAI21_X1 U8603 ( .B1(n7498), .B2(n9897), .A(n6816), .ZN(n6817) );
  INV_X1 U8604 ( .A(n6817), .ZN(n6821) );
  NOR2_X1 U8605 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9988), .ZN(n6818) );
  AOI21_X1 U8606 ( .B1(n9964), .B2(n6819), .A(n6818), .ZN(n6820) );
  OAI211_X1 U8607 ( .C1(n9875), .C2(n6822), .A(n6821), .B(n6820), .ZN(P2_U3184) );
  MUX2_X1 U8608 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8273), .Z(n6827) );
  MUX2_X1 U8609 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8273), .Z(n6826) );
  AOI22_X1 U8610 ( .A1(n6825), .A2(n6824), .B1(n6823), .B2(n6846), .ZN(n9854)
         );
  XOR2_X1 U8611 ( .A(n6826), .B(n6849), .Z(n9853) );
  NAND2_X1 U8612 ( .A1(n9854), .A2(n9853), .ZN(n9852) );
  OAI21_X1 U8613 ( .B1(n6826), .B2(n6849), .A(n9852), .ZN(n9876) );
  XNOR2_X1 U8614 ( .A(n6827), .B(n9863), .ZN(n9877) );
  INV_X1 U8615 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6828) );
  MUX2_X1 U8616 ( .A(n6829), .B(n6828), .S(n8273), .Z(n6830) );
  XNOR2_X1 U8617 ( .A(n6830), .B(n9888), .ZN(n9893) );
  INV_X1 U8618 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6911) );
  MUX2_X1 U8619 ( .A(n6911), .B(n6916), .S(n8273), .Z(n6831) );
  NAND2_X1 U8620 ( .A1(n6831), .A2(n6917), .ZN(n6906) );
  OAI21_X1 U8621 ( .B1(n6917), .B2(n6831), .A(n6906), .ZN(n6832) );
  AOI21_X1 U8622 ( .B1(n6833), .B2(n6832), .A(n6908), .ZN(n6867) );
  INV_X1 U8623 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7507) );
  MUX2_X1 U8624 ( .A(n6916), .B(P2_REG1_REG_6__SCAN_IN), .S(n6917), .Z(n6845)
         );
  NAND2_X1 U8625 ( .A1(n6846), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6834) );
  NAND2_X1 U8626 ( .A1(n6835), .A2(n6834), .ZN(n6836) );
  INV_X1 U8627 ( .A(n6849), .ZN(n9847) );
  XNOR2_X1 U8628 ( .A(n6836), .B(n9847), .ZN(n9844) );
  NAND2_X1 U8629 ( .A1(n9844), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U8630 ( .A1(n6836), .A2(n6849), .ZN(n6837) );
  NAND2_X1 U8631 ( .A1(n6838), .A2(n6837), .ZN(n9860) );
  MUX2_X1 U8632 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6839), .S(n9863), .Z(n9861)
         );
  NAND2_X1 U8633 ( .A1(n9860), .A2(n9861), .ZN(n9859) );
  NAND2_X1 U8634 ( .A1(n9863), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U8635 ( .A1(n9859), .A2(n6840), .ZN(n6841) );
  XNOR2_X1 U8636 ( .A(n6841), .B(n9888), .ZN(n9885) );
  NAND2_X1 U8637 ( .A1(n9885), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U8638 ( .A1(n6841), .A2(n6853), .ZN(n6842) );
  NAND2_X1 U8639 ( .A1(n6843), .A2(n6842), .ZN(n6844) );
  NAND2_X1 U8640 ( .A1(n6844), .A2(n6845), .ZN(n6919) );
  OAI21_X1 U8641 ( .B1(n6845), .B2(n6844), .A(n6919), .ZN(n6862) );
  NAND2_X1 U8642 ( .A1(n6846), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6847) );
  NAND2_X1 U8643 ( .A1(n6850), .A2(n6849), .ZN(n9866) );
  NAND2_X1 U8644 ( .A1(n9868), .A2(n9866), .ZN(n6851) );
  INV_X1 U8645 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7205) );
  MUX2_X1 U8646 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7205), .S(n9863), .Z(n9865)
         );
  NAND2_X1 U8647 ( .A1(n6851), .A2(n9865), .ZN(n9870) );
  NAND2_X1 U8648 ( .A1(n9863), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U8649 ( .A1(n9870), .A2(n6852), .ZN(n6854) );
  NAND2_X1 U8650 ( .A1(n6854), .A2(n6853), .ZN(n6858) );
  NAND2_X1 U8651 ( .A1(n9882), .A2(n6858), .ZN(n6856) );
  XNOR2_X1 U8652 ( .A(n6917), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6857) );
  NAND2_X1 U8653 ( .A1(n6856), .A2(n6857), .ZN(n6913) );
  INV_X1 U8654 ( .A(n6857), .ZN(n6859) );
  NAND3_X1 U8655 ( .A1(n9882), .A2(n6859), .A3(n6858), .ZN(n6860) );
  AOI21_X1 U8656 ( .B1(n6913), .B2(n6860), .A(n9980), .ZN(n6861) );
  AOI21_X1 U8657 ( .B1(n9974), .B2(n6862), .A(n6861), .ZN(n6864) );
  AND2_X1 U8658 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7135) );
  AOI21_X1 U8659 ( .B1(n9964), .B2(n6917), .A(n7135), .ZN(n6863) );
  OAI211_X1 U8660 ( .C1(n7507), .C2(n9897), .A(n6864), .B(n6863), .ZN(n6865)
         );
  INV_X1 U8661 ( .A(n6865), .ZN(n6866) );
  OAI21_X1 U8662 ( .B1(n6867), .B2(n9875), .A(n6866), .ZN(P2_U3188) );
  NAND2_X1 U8663 ( .A1(n7187), .A2(n6932), .ZN(n8062) );
  INV_X1 U8664 ( .A(n8062), .ZN(n6868) );
  OR2_X1 U8665 ( .A1(n6868), .A2(n7179), .ZN(n7210) );
  NAND2_X1 U8666 ( .A1(n9992), .A2(n10046), .ZN(n10030) );
  OR2_X1 U8667 ( .A1(n10030), .A2(n8484), .ZN(n6869) );
  NAND2_X1 U8668 ( .A1(n7210), .A2(n6869), .ZN(n6870) );
  NAND2_X1 U8669 ( .A1(n8234), .A2(n8479), .ZN(n7211) );
  OAI211_X1 U8670 ( .C1(n10057), .C2(n6932), .A(n6870), .B(n7211), .ZN(n8553)
         );
  NAND2_X1 U8671 ( .A1(n10063), .A2(n8553), .ZN(n6871) );
  OAI21_X1 U8672 ( .B1(n10063), .B2(n6088), .A(n6871), .ZN(P2_U3390) );
  INV_X1 U8673 ( .A(n9796), .ZN(n9764) );
  INV_X1 U8674 ( .A(n6872), .ZN(n8985) );
  XNOR2_X1 U8675 ( .A(n6873), .B(n8985), .ZN(n6880) );
  INV_X1 U8676 ( .A(n6880), .ZN(n6950) );
  XNOR2_X1 U8677 ( .A(n5761), .B(n6889), .ZN(n6874) );
  NAND2_X1 U8678 ( .A1(n6874), .A2(n9673), .ZN(n6948) );
  OAI21_X1 U8679 ( .B1(n8905), .B2(n9781), .A(n6948), .ZN(n6881) );
  INV_X1 U8680 ( .A(n9787), .ZN(n9766) );
  INV_X1 U8681 ( .A(n9789), .ZN(n9769) );
  AOI22_X1 U8682 ( .A1(n9766), .A2(n6712), .B1(n5779), .B2(n9769), .ZN(n6879)
         );
  OAI21_X1 U8683 ( .B1(n6876), .B2(n6872), .A(n6875), .ZN(n6877) );
  NAND2_X1 U8684 ( .A1(n6877), .A2(n9777), .ZN(n6878) );
  OAI211_X1 U8685 ( .C1(n6880), .C2(n9626), .A(n6879), .B(n6878), .ZN(n6944)
         );
  AOI211_X1 U8686 ( .C1(n9764), .C2(n6950), .A(n6881), .B(n6944), .ZN(n9688)
         );
  NAND2_X1 U8687 ( .A1(n9823), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6882) );
  OAI21_X1 U8688 ( .B1(n9688), .B2(n9823), .A(n6882), .ZN(P1_U3523) );
  XOR2_X1 U8689 ( .A(n8987), .B(n6883), .Z(n6885) );
  AOI222_X1 U8690 ( .A1(n9777), .A2(n6885), .B1(n9050), .B2(n9769), .C1(n6884), 
        .C2(n9766), .ZN(n9692) );
  OR2_X1 U8691 ( .A1(n9634), .A2(n6886), .ZN(n6945) );
  OR2_X1 U8692 ( .A1(n9666), .A2(n9626), .ZN(n6887) );
  XNOR2_X1 U8693 ( .A(n8987), .B(n6888), .ZN(n9695) );
  AOI21_X1 U8694 ( .B1(n8905), .B2(n6889), .A(n9691), .ZN(n6890) );
  NOR3_X1 U8695 ( .A1(n9674), .A2(n6890), .A3(n9321), .ZN(n9689) );
  INV_X1 U8696 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7054) );
  INV_X1 U8697 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9073) );
  OAI22_X1 U8698 ( .A1(n9296), .A2(n7054), .B1(n9073), .B2(n9664), .ZN(n6891)
         );
  AOI21_X1 U8699 ( .B1(n9689), .B2(n9676), .A(n6891), .ZN(n6892) );
  OAI21_X1 U8700 ( .B1(n9691), .B2(n9668), .A(n6892), .ZN(n6893) );
  AOI21_X1 U8701 ( .B1(n9677), .B2(n9695), .A(n6893), .ZN(n6894) );
  OAI21_X1 U8702 ( .B1(n9692), .B2(n9634), .A(n6894), .ZN(P1_U3291) );
  INV_X1 U8703 ( .A(n6895), .ZN(n6896) );
  NOR2_X1 U8704 ( .A1(n6897), .A2(n6896), .ZN(n6901) );
  INV_X1 U8705 ( .A(n6899), .ZN(n6900) );
  AOI21_X1 U8706 ( .B1(n6901), .B2(n6898), .A(n6900), .ZN(n6905) );
  INV_X1 U8707 ( .A(n9691), .ZN(n6902) );
  AOI22_X1 U8708 ( .A1(n7844), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n6902), .B2(
        n8769), .ZN(n6904) );
  AOI22_X1 U8709 ( .A1(n8768), .A2(n9050), .B1(n8767), .B2(n6884), .ZN(n6903)
         );
  OAI211_X1 U8710 ( .C1(n6905), .C2(n8754), .A(n6904), .B(n6903), .ZN(P1_U3237) );
  INV_X1 U8711 ( .A(n6906), .ZN(n6907) );
  NOR2_X1 U8712 ( .A1(n6908), .A2(n6907), .ZN(n6910) );
  MUX2_X1 U8713 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8273), .Z(n7013) );
  XOR2_X1 U8714 ( .A(n7016), .B(n7013), .Z(n6909) );
  AOI21_X1 U8715 ( .B1(n6910), .B2(n6909), .A(n7014), .ZN(n6926) );
  OR2_X1 U8716 ( .A1(n6917), .A2(n6911), .ZN(n6912) );
  NAND2_X1 U8717 ( .A1(n6913), .A2(n6912), .ZN(n7028) );
  XNOR2_X1 U8718 ( .A(n7028), .B(n7016), .ZN(n6914) );
  OAI21_X1 U8719 ( .B1(n6914), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7030), .ZN(
        n6923) );
  INV_X1 U8720 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7510) );
  AND2_X1 U8721 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7152) );
  AOI21_X1 U8722 ( .B1(n9964), .B2(n7016), .A(n7152), .ZN(n6915) );
  OAI21_X1 U8723 ( .B1(n9897), .B2(n7510), .A(n6915), .ZN(n6922) );
  INV_X1 U8724 ( .A(n9974), .ZN(n7345) );
  OR2_X1 U8725 ( .A1(n6917), .A2(n6916), .ZN(n6918) );
  NAND2_X1 U8726 ( .A1(n6919), .A2(n6918), .ZN(n7022) );
  XNOR2_X1 U8727 ( .A(n7022), .B(n7016), .ZN(n7021) );
  XOR2_X1 U8728 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7021), .Z(n6920) );
  NOR2_X1 U8729 ( .A1(n7345), .A2(n6920), .ZN(n6921) );
  AOI211_X1 U8730 ( .C1(n6924), .C2(n6923), .A(n6922), .B(n6921), .ZN(n6925)
         );
  OAI21_X1 U8731 ( .B1(n6926), .B2(n9875), .A(n6925), .ZN(P2_U3189) );
  INV_X1 U8732 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6928) );
  INV_X1 U8733 ( .A(n6927), .ZN(n6929) );
  INV_X1 U8734 ( .A(n9914), .ZN(n8257) );
  OAI222_X1 U8735 ( .A1(n7863), .A2(n6928), .B1(n8650), .B2(n6929), .C1(
        P2_U3151), .C2(n8257), .ZN(P2_U3281) );
  INV_X1 U8736 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10262) );
  INV_X1 U8737 ( .A(n7630), .ZN(n7318) );
  OAI222_X1 U8738 ( .A1(n7889), .A2(n10262), .B1(n9457), .B2(n6929), .C1(
        P1_U3086), .C2(n7318), .ZN(P1_U3341) );
  NOR2_X1 U8739 ( .A1(n6931), .A2(n6930), .ZN(n6975) );
  INV_X1 U8740 ( .A(n7210), .ZN(n8025) );
  INV_X1 U8741 ( .A(n7968), .ZN(n8009) );
  OAI22_X1 U8742 ( .A1(n8025), .A2(n7970), .B1(n8009), .B2(n6932), .ZN(n6933)
         );
  AOI21_X1 U8743 ( .B1(n7979), .B2(n8234), .A(n6933), .ZN(n6934) );
  OAI21_X1 U8744 ( .B1(n6975), .B2(n6935), .A(n6934), .ZN(P2_U3172) );
  INV_X1 U8745 ( .A(n7187), .ZN(n6936) );
  OAI22_X1 U8746 ( .A1(n10007), .A2(n8009), .B1(n7981), .B2(n6936), .ZN(n6937)
         );
  AOI21_X1 U8747 ( .B1(n7979), .B2(n8232), .A(n6937), .ZN(n6943) );
  OAI21_X1 U8748 ( .B1(n6940), .B2(n6939), .A(n6938), .ZN(n6941) );
  NAND2_X1 U8749 ( .A1(n6941), .A2(n7997), .ZN(n6942) );
  OAI211_X1 U8750 ( .C1(n6975), .C2(n7183), .A(n6943), .B(n6942), .ZN(P2_U3162) );
  INV_X1 U8751 ( .A(n6944), .ZN(n6952) );
  INV_X2 U8752 ( .A(n9296), .ZN(n9634) );
  INV_X1 U8753 ( .A(n6945), .ZN(n9658) );
  NAND2_X1 U8754 ( .A1(n9652), .A2(n5761), .ZN(n6947) );
  AOI22_X1 U8755 ( .A1(n9666), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9651), .ZN(n6946) );
  OAI211_X1 U8756 ( .C1(n6948), .C2(n9264), .A(n6947), .B(n6946), .ZN(n6949)
         );
  AOI21_X1 U8757 ( .B1(n6950), .B2(n9658), .A(n6949), .ZN(n6951) );
  OAI21_X1 U8758 ( .B1(n6952), .B2(n9634), .A(n6951), .ZN(P1_U3292) );
  OAI21_X1 U8759 ( .B1(n6955), .B2(n6953), .A(n6954), .ZN(n6962) );
  NAND2_X1 U8760 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9087) );
  INV_X1 U8761 ( .A(n9087), .ZN(n6956) );
  AOI21_X1 U8762 ( .B1(n6010), .B2(n6957), .A(n6956), .ZN(n6960) );
  AOI22_X1 U8763 ( .A1(n8768), .A2(n9662), .B1(n6958), .B2(n8769), .ZN(n6959)
         );
  OAI211_X1 U8764 ( .C1(n5239), .C2(n8779), .A(n6960), .B(n6959), .ZN(n6961)
         );
  AOI21_X1 U8765 ( .B1(n6962), .B2(n8777), .A(n6961), .ZN(n6963) );
  INV_X1 U8766 ( .A(n6963), .ZN(P1_U3218) );
  NAND2_X1 U8767 ( .A1(n6964), .A2(n8777), .ZN(n6972) );
  AOI21_X1 U8768 ( .B1(n6954), .B2(n6966), .A(n6965), .ZN(n6971) );
  AOI22_X1 U8769 ( .A1(n8768), .A2(n9049), .B1(n6988), .B2(n8769), .ZN(n6970)
         );
  AND2_X1 U8770 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9552) );
  INV_X1 U8771 ( .A(n9050), .ZN(n6967) );
  NOR2_X1 U8772 ( .A1(n8779), .A2(n6967), .ZN(n6968) );
  AOI211_X1 U8773 ( .C1(n6010), .C2(n6987), .A(n9552), .B(n6968), .ZN(n6969)
         );
  OAI211_X1 U8774 ( .C1(n6972), .C2(n6971), .A(n6970), .B(n6969), .ZN(P1_U3230) );
  XOR2_X1 U8775 ( .A(n6974), .B(n6973), .Z(n6979) );
  OAI22_X1 U8776 ( .A1(n10013), .A2(n8009), .B1(n7981), .B2(n9996), .ZN(n6977)
         );
  NOR2_X1 U8777 ( .A1(n6975), .A2(n9988), .ZN(n6976) );
  AOI211_X1 U8778 ( .C1(n7979), .C2(n4841), .A(n6977), .B(n6976), .ZN(n6978)
         );
  OAI21_X1 U8779 ( .B1(n7970), .B2(n6979), .A(n6978), .ZN(P2_U3177) );
  XNOR2_X1 U8780 ( .A(n6980), .B(n4528), .ZN(n6981) );
  NAND2_X1 U8781 ( .A1(n6981), .A2(n9777), .ZN(n6983) );
  AOI22_X1 U8782 ( .A1(n9766), .A2(n9050), .B1(n9049), .B2(n9769), .ZN(n6982)
         );
  AND2_X1 U8783 ( .A1(n6983), .A2(n6982), .ZN(n9709) );
  XNOR2_X1 U8784 ( .A(n6984), .B(n4528), .ZN(n9707) );
  NAND2_X1 U8785 ( .A1(n9672), .A2(n6988), .ZN(n6985) );
  NAND2_X1 U8786 ( .A1(n6985), .A2(n9673), .ZN(n6986) );
  OR2_X1 U8787 ( .A1(n6986), .A2(n7143), .ZN(n9704) );
  AOI22_X1 U8788 ( .A1(n9666), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n6987), .B2(
        n9651), .ZN(n6990) );
  NAND2_X1 U8789 ( .A1(n9652), .A2(n6988), .ZN(n6989) );
  OAI211_X1 U8790 ( .C1(n9704), .C2(n9264), .A(n6990), .B(n6989), .ZN(n6991)
         );
  AOI21_X1 U8791 ( .B1(n9707), .B2(n9677), .A(n6991), .ZN(n6992) );
  OAI21_X1 U8792 ( .B1(n9709), .B2(n9666), .A(n6992), .ZN(P1_U3289) );
  INV_X1 U8793 ( .A(n6993), .ZN(n6994) );
  AOI211_X1 U8794 ( .C1(n6996), .C2(n6995), .A(n7970), .B(n6994), .ZN(n7000)
         );
  INV_X1 U8795 ( .A(n8096), .ZN(n8231) );
  AOI22_X1 U8796 ( .A1(n8006), .A2(n8232), .B1(n7979), .B2(n8231), .ZN(n6998)
         );
  NOR2_X1 U8797 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6135), .ZN(n9846) );
  AOI21_X1 U8798 ( .B1(n7968), .B2(n7194), .A(n9846), .ZN(n6997) );
  OAI211_X1 U8799 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8003), .A(n6998), .B(
        n6997), .ZN(n6999) );
  OR2_X1 U8800 ( .A1(n7000), .A2(n6999), .ZN(P2_U3158) );
  INV_X1 U8801 ( .A(n7127), .ZN(n7001) );
  AOI21_X1 U8802 ( .B1(n7003), .B2(n7002), .A(n7001), .ZN(n7008) );
  INV_X1 U8803 ( .A(n7004), .ZN(n7203) );
  AOI22_X1 U8804 ( .A1(n8006), .A2(n4841), .B1(n7979), .B2(n8230), .ZN(n7005)
         );
  NAND2_X1 U8805 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9862) );
  OAI211_X1 U8806 ( .C1(n10022), .C2(n8009), .A(n7005), .B(n9862), .ZN(n7006)
         );
  AOI21_X1 U8807 ( .B1(n7203), .B2(n7994), .A(n7006), .ZN(n7007) );
  OAI21_X1 U8808 ( .B1(n7008), .B2(n7970), .A(n7007), .ZN(P2_U3170) );
  INV_X1 U8809 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7010) );
  INV_X1 U8810 ( .A(n7009), .ZN(n7011) );
  OAI222_X1 U8811 ( .A1(n7889), .A2(n7010), .B1(n9457), .B2(n7011), .C1(
        P1_U3086), .C2(n7716), .ZN(P1_U3340) );
  INV_X1 U8812 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7012) );
  INV_X1 U8813 ( .A(n9931), .ZN(n8255) );
  OAI222_X1 U8814 ( .A1(n7863), .A2(n7012), .B1(n8650), .B2(n7011), .C1(
        P2_U3151), .C2(n8255), .ZN(P2_U3280) );
  INV_X1 U8815 ( .A(n7013), .ZN(n7015) );
  INV_X1 U8816 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7031) );
  MUX2_X1 U8817 ( .A(n7031), .B(n7017), .S(n8273), .Z(n7018) );
  NAND2_X1 U8818 ( .A1(n7018), .A2(n7035), .ZN(n7335) );
  OAI21_X1 U8819 ( .B1(n7018), .B2(n7035), .A(n7335), .ZN(n7019) );
  AOI21_X1 U8820 ( .B1(n7020), .B2(n7019), .A(n7333), .ZN(n7041) );
  NAND2_X1 U8821 ( .A1(n7021), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7024) );
  NAND2_X1 U8822 ( .A1(n7022), .A2(n7027), .ZN(n7023) );
  NAND2_X1 U8823 ( .A1(n7024), .A2(n7023), .ZN(n7026) );
  AOI22_X1 U8824 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7322), .B1(n7035), .B2(
        n7017), .ZN(n7025) );
  NAND2_X1 U8825 ( .A1(n7025), .A2(n7026), .ZN(n7323) );
  OAI21_X1 U8826 ( .B1(n7026), .B2(n7025), .A(n7323), .ZN(n7039) );
  NAND2_X1 U8827 ( .A1(n7028), .A2(n7027), .ZN(n7029) );
  OR2_X1 U8828 ( .A1(n7035), .A2(n7031), .ZN(n7326) );
  OAI21_X1 U8829 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7322), .A(n7326), .ZN(
        n7032) );
  AOI21_X1 U8830 ( .B1(n7033), .B2(n7032), .A(n7325), .ZN(n7034) );
  NOR2_X1 U8831 ( .A1(n7034), .A2(n9980), .ZN(n7038) );
  INV_X1 U8832 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10353) );
  AND2_X1 U8833 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7232) );
  AOI21_X1 U8834 ( .B1(n9964), .B2(n7035), .A(n7232), .ZN(n7036) );
  OAI21_X1 U8835 ( .B1(n9897), .B2(n10353), .A(n7036), .ZN(n7037) );
  AOI211_X1 U8836 ( .C1(n9974), .C2(n7039), .A(n7038), .B(n7037), .ZN(n7040)
         );
  OAI21_X1 U8837 ( .B1(n7041), .B2(n9875), .A(n7040), .ZN(P2_U3190) );
  NAND2_X1 U8838 ( .A1(n7127), .A2(n7042), .ZN(n7043) );
  XOR2_X1 U8839 ( .A(n7044), .B(n7043), .Z(n7050) );
  INV_X1 U8840 ( .A(n7122), .ZN(n7048) );
  AOI22_X1 U8841 ( .A1(n8006), .A2(n8231), .B1(n7979), .B2(n8229), .ZN(n7046)
         );
  AND2_X1 U8842 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9887) );
  INV_X1 U8843 ( .A(n9887), .ZN(n7045) );
  OAI211_X1 U8844 ( .C1(n10026), .C2(n8009), .A(n7046), .B(n7045), .ZN(n7047)
         );
  AOI21_X1 U8845 ( .B1(n7048), .B2(n7994), .A(n7047), .ZN(n7049) );
  OAI21_X1 U8846 ( .B1(n7050), .B2(n7970), .A(n7049), .ZN(P2_U3167) );
  NOR2_X1 U8847 ( .A1(n7246), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7051) );
  AOI21_X1 U8848 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7246), .A(n7051), .ZN(
        n7066) );
  NAND2_X1 U8849 ( .A1(n9489), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7052) );
  OAI21_X1 U8850 ( .B1(n9489), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7052), .ZN(
        n9485) );
  NOR2_X1 U8851 ( .A1(n9108), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7053) );
  AOI21_X1 U8852 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9108), .A(n7053), .ZN(
        n9101) );
  MUX2_X1 U8853 ( .A(n7054), .B(P1_REG2_REG_2__SCAN_IN), .S(n7072), .Z(n9082)
         );
  XNOR2_X1 U8854 ( .A(n7073), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9060) );
  NAND2_X1 U8855 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9065) );
  INV_X1 U8856 ( .A(n9065), .ZN(n9059) );
  NAND2_X1 U8857 ( .A1(n9060), .A2(n9059), .ZN(n9058) );
  INV_X1 U8858 ( .A(n7073), .ZN(n9054) );
  NAND2_X1 U8859 ( .A1(n9054), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U8860 ( .A1(n9058), .A2(n7055), .ZN(n9081) );
  NAND2_X1 U8861 ( .A1(n9082), .A2(n9081), .ZN(n9080) );
  INV_X1 U8862 ( .A(n7072), .ZN(n9076) );
  NAND2_X1 U8863 ( .A1(n9076), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7056) );
  NAND2_X1 U8864 ( .A1(n9080), .A2(n7056), .ZN(n9091) );
  XNOR2_X1 U8865 ( .A(n7076), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U8866 ( .A1(n9091), .A2(n9092), .ZN(n9090) );
  INV_X1 U8867 ( .A(n7076), .ZN(n9089) );
  NAND2_X1 U8868 ( .A1(n9089), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7057) );
  NAND2_X1 U8869 ( .A1(n9090), .A2(n7057), .ZN(n9537) );
  NAND2_X1 U8870 ( .A1(n9549), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7058) );
  OAI21_X1 U8871 ( .B1(n9549), .B2(P1_REG2_REG_4__SCAN_IN), .A(n7058), .ZN(
        n9540) );
  INV_X1 U8872 ( .A(n9540), .ZN(n7059) );
  AND2_X1 U8873 ( .A1(n9537), .A2(n7059), .ZN(n9539) );
  INV_X1 U8874 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7060) );
  AOI22_X1 U8875 ( .A1(n7082), .A2(n7060), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n9566), .ZN(n9558) );
  NOR2_X1 U8876 ( .A1(n9557), .A2(n9558), .ZN(n9556) );
  AOI21_X1 U8877 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n7082), .A(n9556), .ZN(
        n9571) );
  INV_X1 U8878 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7061) );
  AOI22_X1 U8879 ( .A1(n7084), .A2(n7061), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n9580), .ZN(n9572) );
  NOR2_X1 U8880 ( .A1(n9571), .A2(n9572), .ZN(n9570) );
  NAND2_X1 U8881 ( .A1(n7087), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7062) );
  OAI21_X1 U8882 ( .B1(n7087), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7062), .ZN(
        n9495) );
  NOR2_X1 U8883 ( .A1(n9494), .A2(n9495), .ZN(n9493) );
  NAND2_X1 U8884 ( .A1(n7090), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7063) );
  OAI21_X1 U8885 ( .B1(n7090), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7063), .ZN(
        n9511) );
  NOR2_X1 U8886 ( .A1(n9510), .A2(n9511), .ZN(n9509) );
  AOI21_X1 U8887 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7090), .A(n9509), .ZN(
        n9100) );
  NAND2_X1 U8888 ( .A1(n9101), .A2(n9100), .ZN(n9099) );
  OAI21_X1 U8889 ( .B1(n9108), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9099), .ZN(
        n9486) );
  NOR2_X1 U8890 ( .A1(n9485), .A2(n9486), .ZN(n9484) );
  NAND2_X1 U8891 ( .A1(n9585), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7064) );
  OAI21_X1 U8892 ( .B1(n9585), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7064), .ZN(
        n9588) );
  NOR2_X1 U8893 ( .A1(n9587), .A2(n9588), .ZN(n9586) );
  AOI21_X1 U8894 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9585), .A(n9586), .ZN(
        n7065) );
  NAND2_X1 U8895 ( .A1(n7066), .A2(n7065), .ZN(n7242) );
  OAI21_X1 U8896 ( .B1(n7066), .B2(n7065), .A(n7242), .ZN(n7099) );
  INV_X1 U8897 ( .A(n7867), .ZN(n9067) );
  AND2_X1 U8898 ( .A1(n7068), .A2(n9067), .ZN(n9064) );
  INV_X1 U8899 ( .A(n7067), .ZN(n7069) );
  NAND2_X1 U8900 ( .A1(n9489), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7070) );
  OAI21_X1 U8901 ( .B1(n9489), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7070), .ZN(
        n9482) );
  NOR2_X1 U8902 ( .A1(n9108), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7071) );
  AOI21_X1 U8903 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9108), .A(n7071), .ZN(
        n9106) );
  INV_X1 U8904 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9804) );
  MUX2_X1 U8905 ( .A(n9804), .B(P1_REG1_REG_2__SCAN_IN), .S(n7072), .Z(n9079)
         );
  XNOR2_X1 U8906 ( .A(n7073), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9057) );
  AND2_X1 U8907 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9056) );
  NAND2_X1 U8908 ( .A1(n9057), .A2(n9056), .ZN(n9055) );
  NAND2_X1 U8909 ( .A1(n9054), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7074) );
  NAND2_X1 U8910 ( .A1(n9055), .A2(n7074), .ZN(n9078) );
  NAND2_X1 U8911 ( .A1(n9079), .A2(n9078), .ZN(n9077) );
  NAND2_X1 U8912 ( .A1(n9076), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7075) );
  NAND2_X1 U8913 ( .A1(n9077), .A2(n7075), .ZN(n9094) );
  XNOR2_X1 U8914 ( .A(n7076), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U8915 ( .A1(n9094), .A2(n9095), .ZN(n9093) );
  NAND2_X1 U8916 ( .A1(n9089), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7077) );
  NAND2_X1 U8917 ( .A1(n9093), .A2(n7077), .ZN(n9542) );
  NAND2_X1 U8918 ( .A1(n9549), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7078) );
  OAI21_X1 U8919 ( .B1(n9549), .B2(P1_REG1_REG_4__SCAN_IN), .A(n7078), .ZN(
        n9545) );
  INV_X1 U8920 ( .A(n9545), .ZN(n7079) );
  AND2_X1 U8921 ( .A1(n9542), .A2(n7079), .ZN(n9544) );
  AND2_X1 U8922 ( .A1(n9549), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7080) );
  INV_X1 U8923 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7081) );
  MUX2_X1 U8924 ( .A(n7081), .B(P1_REG1_REG_5__SCAN_IN), .S(n7082), .Z(n9561)
         );
  NOR2_X1 U8925 ( .A1(n9562), .A2(n9561), .ZN(n9560) );
  AOI21_X1 U8926 ( .B1(n7082), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9560), .ZN(
        n9576) );
  INV_X1 U8927 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7083) );
  MUX2_X1 U8928 ( .A(n7083), .B(P1_REG1_REG_6__SCAN_IN), .S(n7084), .Z(n9575)
         );
  NOR2_X1 U8929 ( .A1(n9576), .A2(n9575), .ZN(n9574) );
  OR2_X1 U8930 ( .A1(n7087), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7086) );
  NAND2_X1 U8931 ( .A1(n7087), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7085) );
  NAND2_X1 U8932 ( .A1(n7086), .A2(n7085), .ZN(n9499) );
  NOR2_X1 U8933 ( .A1(n9498), .A2(n9499), .ZN(n9497) );
  AOI21_X1 U8934 ( .B1(n7087), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9497), .ZN(
        n9514) );
  OR2_X1 U8935 ( .A1(n7090), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7089) );
  NAND2_X1 U8936 ( .A1(n7090), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7088) );
  NAND2_X1 U8937 ( .A1(n7089), .A2(n7088), .ZN(n9515) );
  NOR2_X1 U8938 ( .A1(n9514), .A2(n9515), .ZN(n9513) );
  NAND2_X1 U8939 ( .A1(n9106), .A2(n9105), .ZN(n9104) );
  OAI21_X1 U8940 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9108), .A(n9104), .ZN(
        n9483) );
  NOR2_X1 U8941 ( .A1(n9482), .A2(n9483), .ZN(n9481) );
  INV_X1 U8942 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7091) );
  MUX2_X1 U8943 ( .A(n7091), .B(P1_REG1_REG_11__SCAN_IN), .S(n9585), .Z(n9593)
         );
  NOR2_X1 U8944 ( .A1(n9592), .A2(n9593), .ZN(n9591) );
  AOI21_X1 U8945 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9585), .A(n9591), .ZN(
        n7093) );
  INV_X1 U8946 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9819) );
  AOI22_X1 U8947 ( .A1(n7246), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n9819), .B2(
        n7097), .ZN(n7092) );
  NAND2_X1 U8948 ( .A1(n7093), .A2(n7092), .ZN(n7245) );
  OAI21_X1 U8949 ( .B1(n7093), .B2(n7092), .A(n7245), .ZN(n7094) );
  NAND2_X1 U8950 ( .A1(n7094), .A2(n9595), .ZN(n7096) );
  AND2_X1 U8951 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7762) );
  AOI21_X1 U8952 ( .B1(n9553), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7762), .ZN(
        n7095) );
  OAI211_X1 U8953 ( .C1(n9599), .C2(n7097), .A(n7096), .B(n7095), .ZN(n7098)
         );
  AOI21_X1 U8954 ( .B1(n7099), .B2(n9590), .A(n7098), .ZN(n7100) );
  INV_X1 U8955 ( .A(n7100), .ZN(P1_U3255) );
  INV_X1 U8956 ( .A(n7101), .ZN(n7103) );
  INV_X1 U8957 ( .A(n9947), .ZN(n8253) );
  OAI222_X1 U8958 ( .A1(n8650), .A2(n7103), .B1(n8253), .B2(P2_U3151), .C1(
        n7102), .C2(n7863), .ZN(P2_U3279) );
  INV_X1 U8959 ( .A(n7776), .ZN(n7726) );
  OAI222_X1 U8960 ( .A1(n7889), .A2(n7104), .B1(n9457), .B2(n7103), .C1(n7726), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  AND2_X1 U8961 ( .A1(n8075), .A2(n8094), .ZN(n8027) );
  INV_X1 U8962 ( .A(n8027), .ZN(n7105) );
  XNOR2_X1 U8963 ( .A(n7106), .B(n7105), .ZN(n10027) );
  INV_X1 U8964 ( .A(n7107), .ZN(n7115) );
  NAND2_X1 U8965 ( .A1(n7109), .A2(n7108), .ZN(n7113) );
  NAND2_X1 U8966 ( .A1(n7111), .A2(n7110), .ZN(n7112) );
  AND2_X1 U8967 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  NAND2_X1 U8968 ( .A1(n7115), .A2(n7114), .ZN(n7121) );
  AND2_X1 U8969 ( .A1(n8064), .A2(n7116), .ZN(n10002) );
  NAND2_X1 U8970 ( .A1(n4500), .A2(n10002), .ZN(n7827) );
  XNOR2_X1 U8971 ( .A(n7117), .B(n8027), .ZN(n7119) );
  OAI22_X1 U8972 ( .A1(n4891), .A2(n9993), .B1(n8096), .B2(n9995), .ZN(n7118)
         );
  AOI21_X1 U8973 ( .B1(n7119), .B2(n8484), .A(n7118), .ZN(n7120) );
  OAI21_X1 U8974 ( .B1(n10027), .B2(n9992), .A(n7120), .ZN(n10029) );
  NAND2_X1 U8975 ( .A1(n10029), .A2(n4500), .ZN(n7125) );
  OAI22_X1 U8976 ( .A1(n8442), .A2(n10026), .B1(n7122), .B2(n9989), .ZN(n7123)
         );
  AOI21_X1 U8977 ( .B1(n10005), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7123), .ZN(
        n7124) );
  OAI211_X1 U8978 ( .C1(n10027), .C2(n7827), .A(n7125), .B(n7124), .ZN(
        P2_U3228) );
  NAND2_X1 U8979 ( .A1(n7127), .A2(n7126), .ZN(n7129) );
  AND2_X1 U8980 ( .A1(n7129), .A2(n7128), .ZN(n7133) );
  NAND2_X1 U8981 ( .A1(n7131), .A2(n7130), .ZN(n7132) );
  AOI211_X1 U8982 ( .C1(n7134), .C2(n7133), .A(n7970), .B(n7132), .ZN(n7139)
         );
  AOI22_X1 U8983 ( .A1(n8006), .A2(n8230), .B1(n7979), .B2(n8228), .ZN(n7137)
         );
  AOI21_X1 U8984 ( .B1(n7968), .B2(n7217), .A(n7135), .ZN(n7136) );
  OAI211_X1 U8985 ( .C1(n7225), .C2(n8003), .A(n7137), .B(n7136), .ZN(n7138)
         );
  OR2_X1 U8986 ( .A1(n7139), .A2(n7138), .ZN(P2_U3179) );
  NAND3_X1 U8987 ( .A1(n8797), .A2(n8802), .A3(n8986), .ZN(n7141) );
  NAND2_X1 U8988 ( .A1(n7141), .A2(n7140), .ZN(n7142) );
  AOI222_X1 U8989 ( .A1(n9777), .A2(n7142), .B1(n9662), .B2(n9766), .C1(n9646), 
        .C2(n9769), .ZN(n9712) );
  OAI22_X1 U8990 ( .A1(n9296), .A2(n7060), .B1(n7164), .B2(n9664), .ZN(n7145)
         );
  OAI211_X1 U8991 ( .C1(n7143), .C2(n9713), .A(n9673), .B(n7265), .ZN(n9711)
         );
  NOR2_X1 U8992 ( .A1(n9711), .A2(n9264), .ZN(n7144) );
  AOI211_X1 U8993 ( .C1(n9652), .C2(n7163), .A(n7145), .B(n7144), .ZN(n7148)
         );
  XNOR2_X1 U8994 ( .A(n8986), .B(n7146), .ZN(n9715) );
  NAND2_X1 U8995 ( .A1(n9715), .A2(n9677), .ZN(n7147) );
  OAI211_X1 U8996 ( .C1(n9712), .C2(n9666), .A(n7148), .B(n7147), .ZN(P1_U3288) );
  OAI21_X1 U8997 ( .B1(n7151), .B2(n7150), .A(n7149), .ZN(n7157) );
  AOI22_X1 U8998 ( .A1(n8006), .A2(n8229), .B1(n7979), .B2(n8227), .ZN(n7155)
         );
  AOI21_X1 U8999 ( .B1(n7968), .B2(n7153), .A(n7152), .ZN(n7154) );
  OAI211_X1 U9000 ( .C1(n7281), .C2(n8003), .A(n7155), .B(n7154), .ZN(n7156)
         );
  AOI21_X1 U9001 ( .B1(n7157), .B2(n7997), .A(n7156), .ZN(n7158) );
  INV_X1 U9002 ( .A(n7158), .ZN(P2_U3153) );
  NAND2_X1 U9003 ( .A1(n7160), .A2(n7159), .ZN(n7162) );
  XNOR2_X1 U9004 ( .A(n7162), .B(n7161), .ZN(n7168) );
  AOI22_X1 U9005 ( .A1(n8767), .A2(n9662), .B1(n8769), .B2(n7163), .ZN(n7167)
         );
  NAND2_X1 U9006 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9568) );
  OAI21_X1 U9007 ( .B1(n8750), .B2(n7164), .A(n9568), .ZN(n7165) );
  AOI21_X1 U9008 ( .B1(n8768), .B2(n9646), .A(n7165), .ZN(n7166) );
  OAI211_X1 U9009 ( .C1(n7168), .C2(n8754), .A(n7167), .B(n7166), .ZN(P1_U3227) );
  NAND2_X1 U9010 ( .A1(n5046), .A2(n7170), .ZN(n7171) );
  XNOR2_X1 U9011 ( .A(n7169), .B(n7171), .ZN(n7176) );
  INV_X1 U9012 ( .A(n9729), .ZN(n9048) );
  AOI22_X1 U9013 ( .A1(n8768), .A2(n9048), .B1(n8767), .B2(n9049), .ZN(n7175)
         );
  NOR2_X1 U9014 ( .A1(n8786), .A2(n4789), .ZN(n7173) );
  NAND2_X1 U9015 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9582) );
  INV_X1 U9016 ( .A(n9582), .ZN(n7172) );
  AOI211_X1 U9017 ( .C1(n6010), .C2(n7267), .A(n7173), .B(n7172), .ZN(n7174)
         );
  OAI211_X1 U9018 ( .C1(n7176), .C2(n8754), .A(n7175), .B(n7174), .ZN(P1_U3239) );
  INV_X1 U9019 ( .A(n10002), .ZN(n7177) );
  NAND2_X1 U9020 ( .A1(n9992), .A2(n7177), .ZN(n7178) );
  INV_X1 U9021 ( .A(n7179), .ZN(n7180) );
  NAND2_X1 U9022 ( .A1(n7180), .A2(n7186), .ZN(n7182) );
  NAND2_X1 U9023 ( .A1(n7182), .A2(n7181), .ZN(n10011) );
  OAI22_X1 U9024 ( .A1(n8442), .A2(n10007), .B1(n7183), .B2(n9989), .ZN(n7184)
         );
  AOI21_X1 U9025 ( .B1(n8502), .B2(n10011), .A(n7184), .ZN(n7191) );
  XNOR2_X1 U9026 ( .A(n7186), .B(n7185), .ZN(n7188) );
  AOI222_X1 U9027 ( .A1(n8484), .A2(n7188), .B1(n8232), .B2(n8479), .C1(n7187), 
        .C2(n8481), .ZN(n10008) );
  MUX2_X1 U9028 ( .A(n7189), .B(n10008), .S(n4500), .Z(n7190) );
  NAND2_X1 U9029 ( .A1(n7191), .A2(n7190), .ZN(P2_U3232) );
  XOR2_X1 U9030 ( .A(n8023), .B(n7192), .Z(n7193) );
  AOI222_X1 U9031 ( .A1(n8484), .A2(n7193), .B1(n8231), .B2(n8479), .C1(n8232), 
        .C2(n8481), .ZN(n10018) );
  XNOR2_X1 U9032 ( .A(n8061), .B(n8023), .ZN(n10021) );
  AOI22_X1 U9033 ( .A1(n8473), .A2(n7194), .B1(n6135), .B2(n8472), .ZN(n7195)
         );
  OAI21_X1 U9034 ( .B1(n6121), .B2(n4500), .A(n7195), .ZN(n7196) );
  AOI21_X1 U9035 ( .B1(n8502), .B2(n10021), .A(n7196), .ZN(n7197) );
  OAI21_X1 U9036 ( .B1(n10018), .B2(n10005), .A(n7197), .ZN(P2_U3230) );
  XOR2_X1 U9037 ( .A(n8073), .B(n7198), .Z(n7199) );
  OAI222_X1 U9038 ( .A1(n9995), .A2(n9994), .B1(n9993), .B2(n7200), .C1(n10000), .C2(n7199), .ZN(n10023) );
  INV_X1 U9039 ( .A(n10023), .ZN(n7208) );
  OAI21_X1 U9040 ( .B1(n7202), .B2(n8073), .A(n7201), .ZN(n10025) );
  AOI22_X1 U9041 ( .A1(n8473), .A2(n8095), .B1(n8472), .B2(n7203), .ZN(n7204)
         );
  OAI21_X1 U9042 ( .B1(n7205), .B2(n4500), .A(n7204), .ZN(n7206) );
  AOI21_X1 U9043 ( .B1(n8502), .B2(n10025), .A(n7206), .ZN(n7207) );
  OAI21_X1 U9044 ( .B1(n7208), .B2(n10005), .A(n7207), .ZN(P2_U3229) );
  NAND3_X1 U9045 ( .A1(n7210), .A2(n7209), .A3(n10057), .ZN(n7212) );
  OAI211_X1 U9046 ( .C1(n9989), .C2(n6935), .A(n7212), .B(n7211), .ZN(n7213)
         );
  MUX2_X1 U9047 ( .A(P2_REG2_REG_0__SCAN_IN), .B(n7213), .S(n4500), .Z(n7214)
         );
  AOI21_X1 U9048 ( .B1(n8473), .B2(n7215), .A(n7214), .ZN(n7216) );
  INV_X1 U9049 ( .A(n7216), .ZN(P2_U3233) );
  XNOR2_X1 U9050 ( .A(n8229), .B(n7217), .ZN(n8030) );
  INV_X1 U9051 ( .A(n8030), .ZN(n7218) );
  XNOR2_X1 U9052 ( .A(n7219), .B(n7218), .ZN(n7220) );
  NAND2_X1 U9053 ( .A1(n7220), .A2(n8484), .ZN(n7222) );
  AOI22_X1 U9054 ( .A1(n8479), .A2(n8228), .B1(n8230), .B2(n8481), .ZN(n7221)
         );
  NAND2_X1 U9055 ( .A1(n7222), .A2(n7221), .ZN(n10034) );
  INV_X1 U9056 ( .A(n10034), .ZN(n7229) );
  NAND2_X1 U9057 ( .A1(n7223), .A2(n8075), .ZN(n7224) );
  XNOR2_X1 U9058 ( .A(n7224), .B(n8030), .ZN(n10031) );
  NOR2_X1 U9059 ( .A1(n4500), .A2(n6911), .ZN(n7227) );
  OAI22_X1 U9060 ( .A1(n8442), .A2(n10032), .B1(n7225), .B2(n9989), .ZN(n7226)
         );
  AOI211_X1 U9061 ( .C1(n10031), .C2(n8502), .A(n7227), .B(n7226), .ZN(n7228)
         );
  OAI21_X1 U9062 ( .B1(n7229), .B2(n10005), .A(n7228), .ZN(P2_U3227) );
  XNOR2_X1 U9063 ( .A(n7231), .B(n7230), .ZN(n7239) );
  AOI21_X1 U9064 ( .B1(n8006), .B2(n8228), .A(n7232), .ZN(n7237) );
  INV_X1 U9065 ( .A(n7373), .ZN(n7233) );
  NAND2_X1 U9066 ( .A1(n7994), .A2(n7233), .ZN(n7236) );
  NAND2_X1 U9067 ( .A1(n7968), .A2(n10044), .ZN(n7235) );
  NAND2_X1 U9068 ( .A1(n7979), .A2(n8226), .ZN(n7234) );
  NAND4_X1 U9069 ( .A1(n7237), .A2(n7236), .A3(n7235), .A4(n7234), .ZN(n7238)
         );
  AOI21_X1 U9070 ( .B1(n7239), .B2(n7997), .A(n7238), .ZN(n7240) );
  INV_X1 U9071 ( .A(n7240), .ZN(P2_U3161) );
  NAND2_X1 U9072 ( .A1(n7312), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7241) );
  OAI21_X1 U9073 ( .B1(n7312), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7241), .ZN(
        n7244) );
  OAI21_X1 U9074 ( .B1(n7246), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7242), .ZN(
        n7243) );
  NOR2_X1 U9075 ( .A1(n7244), .A2(n7243), .ZN(n7308) );
  AOI21_X1 U9076 ( .B1(n7244), .B2(n7243), .A(n7308), .ZN(n7255) );
  INV_X1 U9077 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9821) );
  AOI22_X1 U9078 ( .A1(n7312), .A2(n9821), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n7253), .ZN(n7248) );
  OAI21_X1 U9079 ( .B1(n7246), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7245), .ZN(
        n7247) );
  NOR2_X1 U9080 ( .A1(n7248), .A2(n7247), .ZN(n7311) );
  AOI21_X1 U9081 ( .B1(n7248), .B2(n7247), .A(n7311), .ZN(n7249) );
  NAND2_X1 U9082 ( .A1(n7249), .A2(n9595), .ZN(n7252) );
  NOR2_X1 U9083 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7250), .ZN(n7795) );
  AOI21_X1 U9084 ( .B1(n9553), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7795), .ZN(
        n7251) );
  OAI211_X1 U9085 ( .C1(n9599), .C2(n7253), .A(n7252), .B(n7251), .ZN(n7254)
         );
  AOI21_X1 U9086 ( .B1(n7255), .B2(n9590), .A(n7254), .ZN(n7256) );
  INV_X1 U9087 ( .A(n7256), .ZN(P1_U3256) );
  INV_X1 U9088 ( .A(n7257), .ZN(n7259) );
  OAI222_X1 U9089 ( .A1(n7889), .A2(n7258), .B1(n9457), .B2(n7259), .C1(
        P1_U3086), .C2(n7783), .ZN(P1_U3338) );
  INV_X1 U9090 ( .A(n9965), .ZN(n8265) );
  OAI222_X1 U9091 ( .A1(n7863), .A2(n7260), .B1(n8650), .B2(n7259), .C1(
        P2_U3151), .C2(n8265), .ZN(P2_U3278) );
  XOR2_X1 U9092 ( .A(n7264), .B(n7387), .Z(n7261) );
  OAI222_X1 U9093 ( .A1(n9787), .A2(n7262), .B1(n9789), .B2(n9729), .C1(n7261), 
        .C2(n9754), .ZN(n9718) );
  INV_X1 U9094 ( .A(n9718), .ZN(n7273) );
  XNOR2_X1 U9095 ( .A(n7263), .B(n7264), .ZN(n9720) );
  INV_X1 U9096 ( .A(n7265), .ZN(n7266) );
  OAI211_X1 U9097 ( .C1(n7266), .C2(n4789), .A(n9673), .B(n9654), .ZN(n9717)
         );
  AOI22_X1 U9098 ( .A1(n9634), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7267), .B2(
        n9651), .ZN(n7270) );
  NAND2_X1 U9099 ( .A1(n9652), .A2(n7268), .ZN(n7269) );
  OAI211_X1 U9100 ( .C1(n9717), .C2(n9264), .A(n7270), .B(n7269), .ZN(n7271)
         );
  AOI21_X1 U9101 ( .B1(n9720), .B2(n9677), .A(n7271), .ZN(n7272) );
  OAI21_X1 U9102 ( .B1(n7273), .B2(n9634), .A(n7272), .ZN(P1_U3287) );
  INV_X1 U9103 ( .A(n8101), .ZN(n7274) );
  NAND3_X1 U9104 ( .A1(n7275), .A2(n8100), .A3(n7274), .ZN(n7276) );
  NAND2_X1 U9105 ( .A1(n7375), .A2(n7276), .ZN(n10037) );
  XOR2_X1 U9106 ( .A(n7277), .B(n8101), .Z(n7278) );
  NAND2_X1 U9107 ( .A1(n7278), .A2(n8484), .ZN(n7280) );
  AOI22_X1 U9108 ( .A1(n8479), .A2(n8227), .B1(n8229), .B2(n8481), .ZN(n7279)
         );
  OAI211_X1 U9109 ( .C1(n9992), .C2(n10037), .A(n7280), .B(n7279), .ZN(n10039)
         );
  NAND2_X1 U9110 ( .A1(n10039), .A2(n4500), .ZN(n7284) );
  OAI22_X1 U9111 ( .A1(n8442), .A2(n10036), .B1(n7281), .B2(n9989), .ZN(n7282)
         );
  AOI21_X1 U9112 ( .B1(n10005), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7282), .ZN(
        n7283) );
  OAI211_X1 U9113 ( .C1(n10037), .C2(n7827), .A(n7284), .B(n7283), .ZN(
        P2_U3226) );
  INV_X1 U9114 ( .A(n7285), .ZN(n7301) );
  AOI22_X1 U9115 ( .A1(n9121), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9455), .ZN(n7286) );
  OAI21_X1 U9116 ( .B1(n7301), .B2(n9457), .A(n7286), .ZN(P1_U3337) );
  XNOR2_X1 U9117 ( .A(n7289), .B(n7288), .ZN(n7290) );
  XNOR2_X1 U9118 ( .A(n7287), .B(n7290), .ZN(n7291) );
  NAND2_X1 U9119 ( .A1(n7291), .A2(n8777), .ZN(n7296) );
  INV_X1 U9120 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7292) );
  NOR2_X1 U9121 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7292), .ZN(n9505) );
  OAI22_X1 U9122 ( .A1(n7582), .A2(n8780), .B1(n8779), .B2(n7293), .ZN(n7294)
         );
  AOI211_X1 U9123 ( .C1(n6010), .C2(n9650), .A(n9505), .B(n7294), .ZN(n7295)
         );
  OAI211_X1 U9124 ( .C1(n9723), .C2(n8786), .A(n7296), .B(n7295), .ZN(P1_U3213) );
  NAND2_X1 U9125 ( .A1(n7302), .A2(n7570), .ZN(n7298) );
  OAI211_X1 U9126 ( .C1(n7299), .C2(n7889), .A(n7298), .B(n7297), .ZN(P1_U3335) );
  INV_X1 U9127 ( .A(n9467), .ZN(n9468) );
  OAI222_X1 U9128 ( .A1(n8650), .A2(n7301), .B1(n9468), .B2(P2_U3151), .C1(
        n7300), .C2(n7863), .ZN(P2_U3277) );
  INV_X1 U9129 ( .A(n7302), .ZN(n7303) );
  OAI222_X1 U9130 ( .A1(n8650), .A2(n7303), .B1(n8203), .B2(P2_U3151), .C1(
        n10317), .C2(n7863), .ZN(P2_U3275) );
  INV_X1 U9131 ( .A(n7304), .ZN(n7306) );
  OAI222_X1 U9132 ( .A1(n7863), .A2(n7305), .B1(n8650), .B2(n7306), .C1(
        P2_U3151), .C2(n8251), .ZN(P2_U3276) );
  OAI222_X1 U9133 ( .A1(n7889), .A2(n7307), .B1(n9457), .B2(n7306), .C1(
        P1_U3086), .C2(n5702), .ZN(P1_U3336) );
  XNOR2_X1 U9134 ( .A(n7630), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n7309) );
  INV_X1 U9135 ( .A(n9590), .ZN(n9538) );
  NOR2_X1 U9136 ( .A1(n7310), .A2(n7309), .ZN(n7627) );
  AOI211_X1 U9137 ( .C1(n7310), .C2(n7309), .A(n9538), .B(n7627), .ZN(n7321)
         );
  INV_X1 U9138 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10397) );
  NOR2_X1 U9139 ( .A1(n7630), .A2(n10397), .ZN(n7313) );
  AOI21_X1 U9140 ( .B1(n7630), .B2(n10397), .A(n7313), .ZN(n7314) );
  INV_X1 U9141 ( .A(n9595), .ZN(n9543) );
  NOR2_X1 U9142 ( .A1(n7315), .A2(n7314), .ZN(n7629) );
  AOI211_X1 U9143 ( .C1(n7315), .C2(n7314), .A(n9543), .B(n7629), .ZN(n7320)
         );
  NOR2_X1 U9144 ( .A1(n7316), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8661) );
  AOI21_X1 U9145 ( .B1(n9553), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n8661), .ZN(
        n7317) );
  OAI21_X1 U9146 ( .B1(n7318), .B2(n9599), .A(n7317), .ZN(n7319) );
  OR3_X1 U9147 ( .A1(n7321), .A2(n7320), .A3(n7319), .ZN(P1_U3257) );
  NAND2_X1 U9148 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7322), .ZN(n7324) );
  NAND2_X1 U9149 ( .A1(n7324), .A2(n7323), .ZN(n7423) );
  XNOR2_X1 U9150 ( .A(n7423), .B(n7339), .ZN(n7424) );
  INV_X1 U9151 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7329) );
  XNOR2_X1 U9152 ( .A(n7424), .B(n7329), .ZN(n7346) );
  XNOR2_X1 U9153 ( .A(n7428), .B(n7339), .ZN(n7327) );
  OAI21_X1 U9154 ( .B1(n7327), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7431), .ZN(
        n7328) );
  INV_X1 U9155 ( .A(n7328), .ZN(n7342) );
  MUX2_X1 U9156 ( .A(n7551), .B(n7329), .S(n8273), .Z(n7330) );
  NAND2_X1 U9157 ( .A1(n7330), .A2(n7339), .ZN(n7441) );
  INV_X1 U9158 ( .A(n7330), .ZN(n7331) );
  NAND2_X1 U9159 ( .A1(n7331), .A2(n7429), .ZN(n7332) );
  AND2_X1 U9160 ( .A1(n7441), .A2(n7332), .ZN(n7337) );
  NAND2_X1 U9161 ( .A1(n7335), .A2(n7334), .ZN(n7336) );
  NAND2_X1 U9162 ( .A1(n7337), .A2(n7336), .ZN(n7442) );
  OAI21_X1 U9163 ( .B1(n7337), .B2(n7336), .A(n7442), .ZN(n7338) );
  AND2_X1 U9164 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7412) );
  AOI21_X1 U9165 ( .B1(n9973), .B2(n7338), .A(n7412), .ZN(n7341) );
  NAND2_X1 U9166 ( .A1(n9964), .A2(n7339), .ZN(n7340) );
  OAI211_X1 U9167 ( .C1(n7342), .C2(n9980), .A(n7341), .B(n7340), .ZN(n7343)
         );
  AOI21_X1 U9168 ( .B1(n9966), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7343), .ZN(
        n7344) );
  OAI21_X1 U9169 ( .B1(n7346), .B2(n7345), .A(n7344), .ZN(P2_U3191) );
  INV_X1 U9170 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10332) );
  INV_X1 U9171 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U9172 ( .A1(n7347), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7351) );
  INV_X1 U9173 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7348) );
  OR2_X1 U9174 ( .A1(n7349), .A2(n7348), .ZN(n7350) );
  OAI211_X1 U9175 ( .C1(n7352), .C2(n8290), .A(n7351), .B(n7350), .ZN(n7353)
         );
  INV_X1 U9176 ( .A(n7353), .ZN(n7354) );
  INV_X1 U9177 ( .A(n8287), .ZN(n7356) );
  NAND2_X1 U9178 ( .A1(n7356), .A2(P2_U3893), .ZN(n7357) );
  OAI21_X1 U9179 ( .B1(P2_U3893), .B2(n10332), .A(n7357), .ZN(P2_U3522) );
  INV_X1 U9180 ( .A(n7358), .ZN(n7359) );
  AOI21_X1 U9181 ( .B1(n8993), .B2(n7360), .A(n7359), .ZN(n9753) );
  NOR2_X1 U9182 ( .A1(n9634), .A2(n9754), .ZN(n9266) );
  INV_X1 U9183 ( .A(n9266), .ZN(n9316) );
  XNOR2_X1 U9184 ( .A(n7362), .B(n7361), .ZN(n9756) );
  NAND2_X1 U9185 ( .A1(n9756), .A2(n9677), .ZN(n7370) );
  INV_X1 U9186 ( .A(n7363), .ZN(n9639) );
  AOI211_X1 U9187 ( .C1(n9751), .C2(n7383), .A(n9321), .B(n9639), .ZN(n9749)
         );
  NOR2_X1 U9188 ( .A1(n4664), .A2(n9668), .ZN(n7368) );
  OR2_X1 U9189 ( .A1(n9666), .A2(n9787), .ZN(n9307) );
  INV_X1 U9190 ( .A(n7364), .ZN(n9310) );
  INV_X1 U9191 ( .A(n9748), .ZN(n9767) );
  NAND2_X1 U9192 ( .A1(n9310), .A2(n9767), .ZN(n7366) );
  AOI22_X1 U9193 ( .A1(n9634), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n5080), .B2(
        n9651), .ZN(n7365) );
  OAI211_X1 U9194 ( .C1(n9747), .C2(n9307), .A(n7366), .B(n7365), .ZN(n7367)
         );
  AOI211_X1 U9195 ( .C1(n9749), .C2(n9676), .A(n7368), .B(n7367), .ZN(n7369)
         );
  OAI211_X1 U9196 ( .C1(n9753), .C2(n9316), .A(n7370), .B(n7369), .ZN(P1_U3283) );
  AND2_X1 U9197 ( .A1(n8085), .A2(n8104), .ZN(n8031) );
  XNOR2_X1 U9198 ( .A(n7371), .B(n8031), .ZN(n7372) );
  AOI222_X1 U9199 ( .A1(n8484), .A2(n7372), .B1(n8228), .B2(n8481), .C1(n8226), 
        .C2(n8479), .ZN(n10041) );
  OAI22_X1 U9200 ( .A1(n4500), .A2(n7031), .B1(n7373), .B2(n9989), .ZN(n7378)
         );
  NAND2_X1 U9201 ( .A1(n7375), .A2(n7374), .ZN(n7376) );
  XNOR2_X1 U9202 ( .A(n7376), .B(n8031), .ZN(n10040) );
  NOR2_X1 U9203 ( .A1(n10040), .A2(n8476), .ZN(n7377) );
  AOI211_X1 U9204 ( .C1(n8473), .C2(n10044), .A(n7378), .B(n7377), .ZN(n7379)
         );
  OAI21_X1 U9205 ( .B1(n10041), .B2(n10005), .A(n7379), .ZN(P2_U3225) );
  XOR2_X1 U9206 ( .A(n7390), .B(n7380), .Z(n9743) );
  AOI22_X1 U9207 ( .A1(n9634), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7584), .B2(
        n9651), .ZN(n7381) );
  OAI21_X1 U9208 ( .B1(n9307), .B2(n7582), .A(n7381), .ZN(n7386) );
  INV_X1 U9209 ( .A(n7404), .ZN(n7382) );
  AOI21_X1 U9210 ( .B1(n7382), .B2(n9740), .A(n9321), .ZN(n7384) );
  AOI22_X1 U9211 ( .A1(n7384), .A2(n7383), .B1(n9769), .B2(n9629), .ZN(n9742)
         );
  NOR2_X1 U9212 ( .A1(n9742), .A2(n9264), .ZN(n7385) );
  AOI211_X1 U9213 ( .C1(n9652), .C2(n9740), .A(n7386), .B(n7385), .ZN(n7393)
         );
  OAI21_X1 U9214 ( .B1(n7387), .B2(n8800), .A(n8799), .ZN(n9645) );
  NOR2_X1 U9215 ( .A1(n9645), .A2(n4561), .ZN(n9644) );
  INV_X1 U9216 ( .A(n7388), .ZN(n7389) );
  NOR2_X1 U9217 ( .A1(n9644), .A2(n7389), .ZN(n7398) );
  NAND2_X1 U9218 ( .A1(n7398), .A2(n7397), .ZN(n7396) );
  NAND2_X1 U9219 ( .A1(n7396), .A2(n8809), .ZN(n7391) );
  XNOR2_X1 U9220 ( .A(n7391), .B(n7390), .ZN(n9745) );
  NAND2_X1 U9221 ( .A1(n9745), .A2(n9266), .ZN(n7392) );
  OAI211_X1 U9222 ( .C1(n9743), .C2(n9336), .A(n7393), .B(n7392), .ZN(P1_U3284) );
  INV_X1 U9223 ( .A(n7394), .ZN(n7421) );
  INV_X1 U9224 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10198) );
  OAI222_X1 U9225 ( .A1(n8650), .A2(n7421), .B1(n8026), .B2(P2_U3151), .C1(
        n10198), .C2(n7863), .ZN(P2_U3274) );
  XOR2_X1 U9226 ( .A(n7395), .B(n7397), .Z(n9735) );
  INV_X1 U9227 ( .A(n9735), .ZN(n9737) );
  OAI211_X1 U9228 ( .C1(n7398), .C2(n7397), .A(n9777), .B(n7396), .ZN(n9733)
         );
  NAND2_X1 U9229 ( .A1(n9310), .A2(n4892), .ZN(n7402) );
  INV_X1 U9230 ( .A(n7399), .ZN(n7563) );
  NOR2_X1 U9231 ( .A1(n9664), .A2(n7563), .ZN(n7400) );
  AOI21_X1 U9232 ( .B1(n9666), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7400), .ZN(
        n7401) );
  OAI211_X1 U9233 ( .C1(n9729), .C2(n9307), .A(n7402), .B(n7401), .ZN(n7403)
         );
  AOI21_X1 U9234 ( .B1(n9652), .B2(n9732), .A(n7403), .ZN(n7407) );
  OAI21_X1 U9235 ( .B1(n9655), .B2(n4794), .A(n9673), .ZN(n7405) );
  NOR2_X1 U9236 ( .A1(n7405), .A2(n7404), .ZN(n9730) );
  NAND2_X1 U9237 ( .A1(n9730), .A2(n9676), .ZN(n7406) );
  OAI211_X1 U9238 ( .C1(n9733), .C2(n9634), .A(n7407), .B(n7406), .ZN(n7408)
         );
  AOI21_X1 U9239 ( .B1(n9677), .B2(n9737), .A(n7408), .ZN(n7409) );
  INV_X1 U9240 ( .A(n7409), .ZN(P1_U3285) );
  AOI211_X1 U9241 ( .C1(n7411), .C2(n7410), .A(n7970), .B(n4590), .ZN(n7419)
         );
  AOI21_X1 U9242 ( .B1(n8006), .B2(n8227), .A(n7412), .ZN(n7417) );
  NAND2_X1 U9243 ( .A1(n7968), .A2(n7552), .ZN(n7416) );
  INV_X1 U9244 ( .A(n7550), .ZN(n7413) );
  NAND2_X1 U9245 ( .A1(n7994), .A2(n7413), .ZN(n7415) );
  NAND2_X1 U9246 ( .A1(n7979), .A2(n8225), .ZN(n7414) );
  NAND4_X1 U9247 ( .A1(n7417), .A2(n7416), .A3(n7415), .A4(n7414), .ZN(n7418)
         );
  OR2_X1 U9248 ( .A1(n7419), .A2(n7418), .ZN(P2_U3171) );
  OAI222_X1 U9249 ( .A1(n7889), .A2(n7422), .B1(n9457), .B2(n7421), .C1(n7420), 
        .C2(P1_U3086), .ZN(P1_U3334) );
  AOI22_X1 U9250 ( .A1(n7424), .A2(P2_REG1_REG_9__SCAN_IN), .B1(n7423), .B2(
        n7429), .ZN(n7425) );
  INV_X1 U9251 ( .A(n7425), .ZN(n7427) );
  AOI22_X1 U9252 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7473), .B1(n7445), .B2(
        n7434), .ZN(n7426) );
  NAND2_X1 U9253 ( .A1(n7426), .A2(n7427), .ZN(n7474) );
  OAI21_X1 U9254 ( .B1(n7427), .B2(n7426), .A(n7474), .ZN(n7451) );
  INV_X1 U9255 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7518) );
  NOR2_X1 U9256 ( .A1(n9897), .A2(n7518), .ZN(n7450) );
  OR2_X1 U9257 ( .A1(n7445), .A2(n7595), .ZN(n7479) );
  OAI21_X1 U9258 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7473), .A(n7479), .ZN(
        n7433) );
  NAND2_X1 U9259 ( .A1(n7429), .A2(n7428), .ZN(n7430) );
  AOI21_X1 U9260 ( .B1(n7433), .B2(n7432), .A(n7477), .ZN(n7448) );
  NAND2_X1 U9261 ( .A1(n7442), .A2(n7441), .ZN(n7439) );
  MUX2_X1 U9262 ( .A(n7595), .B(n7434), .S(n8273), .Z(n7435) );
  NAND2_X1 U9263 ( .A1(n7435), .A2(n7445), .ZN(n7483) );
  INV_X1 U9264 ( .A(n7435), .ZN(n7436) );
  NAND2_X1 U9265 ( .A1(n7436), .A2(n7473), .ZN(n7437) );
  NAND2_X1 U9266 ( .A1(n7483), .A2(n7437), .ZN(n7440) );
  INV_X1 U9267 ( .A(n7440), .ZN(n7438) );
  NAND2_X1 U9268 ( .A1(n7439), .A2(n7438), .ZN(n7484) );
  NAND3_X1 U9269 ( .A1(n7442), .A2(n7441), .A3(n7440), .ZN(n7443) );
  NAND2_X1 U9270 ( .A1(n7484), .A2(n7443), .ZN(n7444) );
  AND2_X1 U9271 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7455) );
  AOI21_X1 U9272 ( .B1(n9973), .B2(n7444), .A(n7455), .ZN(n7447) );
  NAND2_X1 U9273 ( .A1(n9964), .A2(n7445), .ZN(n7446) );
  OAI211_X1 U9274 ( .C1(n7448), .C2(n9980), .A(n7447), .B(n7446), .ZN(n7449)
         );
  AOI211_X1 U9275 ( .C1(n7451), .C2(n9974), .A(n7450), .B(n7449), .ZN(n7452)
         );
  INV_X1 U9276 ( .A(n7452), .ZN(P2_U3192) );
  XNOR2_X1 U9277 ( .A(n7453), .B(n7454), .ZN(n7462) );
  AOI21_X1 U9278 ( .B1(n8006), .B2(n8226), .A(n7455), .ZN(n7460) );
  NAND2_X1 U9279 ( .A1(n7968), .A2(n7597), .ZN(n7459) );
  INV_X1 U9280 ( .A(n7594), .ZN(n7456) );
  NAND2_X1 U9281 ( .A1(n7994), .A2(n7456), .ZN(n7458) );
  NAND2_X1 U9282 ( .A1(n7979), .A2(n8224), .ZN(n7457) );
  NAND4_X1 U9283 ( .A1(n7460), .A2(n7459), .A3(n7458), .A4(n7457), .ZN(n7461)
         );
  AOI21_X1 U9284 ( .B1(n7462), .B2(n7997), .A(n7461), .ZN(n7463) );
  INV_X1 U9285 ( .A(n7463), .ZN(P2_U3157) );
  XOR2_X1 U9286 ( .A(n8999), .B(n7464), .Z(n9773) );
  OAI21_X1 U9287 ( .B1(n7465), .B2(n8999), .A(n9607), .ZN(n9776) );
  OAI211_X1 U9288 ( .C1(n4820), .C2(n9637), .A(n9673), .B(n9619), .ZN(n9771)
         );
  INV_X1 U9289 ( .A(n9788), .ZN(n9768) );
  NAND2_X1 U9290 ( .A1(n9310), .A2(n9768), .ZN(n7467) );
  AOI22_X1 U9291 ( .A1(n9634), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7763), .B2(
        n9651), .ZN(n7466) );
  OAI211_X1 U9292 ( .C1(n9748), .C2(n9307), .A(n7467), .B(n7466), .ZN(n7468)
         );
  AOI21_X1 U9293 ( .B1(n7469), .B2(n9652), .A(n7468), .ZN(n7470) );
  OAI21_X1 U9294 ( .B1(n9771), .B2(n9264), .A(n7470), .ZN(n7471) );
  AOI21_X1 U9295 ( .B1(n9776), .B2(n9266), .A(n7471), .ZN(n7472) );
  OAI21_X1 U9296 ( .B1(n9773), .B2(n9336), .A(n7472), .ZN(P1_U3281) );
  NAND2_X1 U9297 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7473), .ZN(n7475) );
  NAND2_X1 U9298 ( .A1(n7475), .A2(n7474), .ZN(n7605) );
  XNOR2_X1 U9299 ( .A(n7605), .B(n7613), .ZN(n7476) );
  NAND2_X1 U9300 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7476), .ZN(n7606) );
  OAI21_X1 U9301 ( .B1(n7476), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7606), .ZN(
        n7494) );
  INV_X1 U9302 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7519) );
  NOR2_X1 U9303 ( .A1(n9897), .A2(n7519), .ZN(n7493) );
  NAND2_X1 U9304 ( .A1(n7479), .A2(n7478), .ZN(n7480) );
  AOI21_X1 U9305 ( .B1(n7481), .B2(n6244), .A(n7600), .ZN(n7482) );
  OR2_X1 U9306 ( .A1(n9980), .A2(n7482), .ZN(n7491) );
  AND2_X1 U9307 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7667) );
  INV_X1 U9308 ( .A(n7667), .ZN(n7490) );
  NAND2_X1 U9309 ( .A1(n9964), .A2(n7613), .ZN(n7489) );
  NAND2_X1 U9310 ( .A1(n7484), .A2(n7483), .ZN(n7486) );
  MUX2_X1 U9311 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8273), .Z(n7610) );
  XNOR2_X1 U9312 ( .A(n7610), .B(n7613), .ZN(n7485) );
  NOR2_X1 U9313 ( .A1(n7486), .A2(n7485), .ZN(n7487) );
  OAI21_X1 U9314 ( .B1(n7611), .B2(n7487), .A(n9973), .ZN(n7488) );
  NAND4_X1 U9315 ( .A1(n7491), .A2(n7490), .A3(n7489), .A4(n7488), .ZN(n7492)
         );
  AOI211_X1 U9316 ( .C1(n7494), .C2(n9974), .A(n7493), .B(n7492), .ZN(n7495)
         );
  INV_X1 U9317 ( .A(n7495), .ZN(P2_U3193) );
  NOR2_X1 U9318 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7534) );
  NOR2_X1 U9319 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7532) );
  NOR2_X1 U9320 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7530) );
  NOR2_X1 U9321 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7528) );
  NOR2_X1 U9322 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7526) );
  NOR2_X1 U9323 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7524) );
  NOR2_X1 U9324 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7521) );
  INV_X1 U9325 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9492) );
  INV_X1 U9326 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7516) );
  INV_X1 U9327 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10168) );
  NOR2_X1 U9328 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7514) );
  NOR2_X1 U9329 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7512) );
  NOR2_X1 U9330 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7509) );
  NOR2_X1 U9331 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7506) );
  NOR2_X1 U9332 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7504) );
  NAND2_X1 U9333 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7502) );
  XNOR2_X1 U9334 ( .A(n10367), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10500) );
  NAND2_X1 U9335 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7500) );
  AOI21_X1 U9336 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10082) );
  INV_X1 U9337 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10322) );
  NAND2_X1 U9338 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7496) );
  NOR2_X1 U9339 ( .A1(n10322), .A2(n7496), .ZN(n10083) );
  NOR2_X1 U9340 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10083), .ZN(n7497) );
  NOR2_X1 U9341 ( .A1(n10082), .A2(n7497), .ZN(n10498) );
  XNOR2_X1 U9342 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n7498), .ZN(n10497) );
  NAND2_X1 U9343 ( .A1(n10498), .A2(n10497), .ZN(n7499) );
  NAND2_X1 U9344 ( .A1(n7500), .A2(n7499), .ZN(n10499) );
  NAND2_X1 U9345 ( .A1(n10500), .A2(n10499), .ZN(n7501) );
  NAND2_X1 U9346 ( .A1(n7502), .A2(n7501), .ZN(n10502) );
  INV_X1 U9347 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9881) );
  XOR2_X1 U9348 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n9881), .Z(n10501) );
  NOR2_X1 U9349 ( .A1(n10502), .A2(n10501), .ZN(n7503) );
  NOR2_X1 U9350 ( .A1(n7504), .A2(n7503), .ZN(n10490) );
  INV_X1 U9351 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9898) );
  XOR2_X1 U9352 ( .A(n9898), .B(P1_ADDR_REG_5__SCAN_IN), .Z(n10489) );
  NOR2_X1 U9353 ( .A1(n10490), .A2(n10489), .ZN(n7505) );
  NOR2_X1 U9354 ( .A1(n7506), .A2(n7505), .ZN(n10488) );
  XOR2_X1 U9355 ( .A(n7507), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10487) );
  NOR2_X1 U9356 ( .A1(n10488), .A2(n10487), .ZN(n7508) );
  NOR2_X1 U9357 ( .A1(n7509), .A2(n7508), .ZN(n10494) );
  XOR2_X1 U9358 ( .A(n7510), .B(P1_ADDR_REG_7__SCAN_IN), .Z(n10493) );
  NOR2_X1 U9359 ( .A1(n10494), .A2(n10493), .ZN(n7511) );
  NOR2_X1 U9360 ( .A1(n7512), .A2(n7511), .ZN(n10496) );
  INV_X1 U9361 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9523) );
  AOI22_X1 U9362 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9523), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n10353), .ZN(n10495) );
  NOR2_X1 U9363 ( .A1(n10496), .A2(n10495), .ZN(n7513) );
  NOR2_X1 U9364 ( .A1(n7514), .A2(n7513), .ZN(n10492) );
  AOI22_X1 U9365 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10168), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7516), .ZN(n10491) );
  NOR2_X1 U9366 ( .A1(n10492), .A2(n10491), .ZN(n7515) );
  AOI21_X1 U9367 ( .B1(n7516), .B2(n10168), .A(n7515), .ZN(n10104) );
  AOI22_X1 U9368 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n9492), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n7518), .ZN(n10103) );
  NOR2_X1 U9369 ( .A1(n10104), .A2(n10103), .ZN(n7517) );
  AOI21_X1 U9370 ( .B1(n7518), .B2(n9492), .A(n7517), .ZN(n10102) );
  INV_X1 U9371 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9603) );
  AOI22_X1 U9372 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n9603), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7519), .ZN(n10101) );
  NOR2_X1 U9373 ( .A1(n10102), .A2(n10101), .ZN(n7520) );
  NOR2_X1 U9374 ( .A1(n7521), .A2(n7520), .ZN(n10100) );
  INV_X1 U9375 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7522) );
  INV_X1 U9376 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7622) );
  AOI22_X1 U9377 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7522), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n7622), .ZN(n10099) );
  NOR2_X1 U9378 ( .A1(n10100), .A2(n10099), .ZN(n7523) );
  NOR2_X1 U9379 ( .A1(n7524), .A2(n7523), .ZN(n10098) );
  XNOR2_X1 U9380 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10097) );
  NOR2_X1 U9381 ( .A1(n10098), .A2(n10097), .ZN(n7525) );
  NOR2_X1 U9382 ( .A1(n7526), .A2(n7525), .ZN(n10096) );
  XNOR2_X1 U9383 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10095) );
  NOR2_X1 U9384 ( .A1(n10096), .A2(n10095), .ZN(n7527) );
  NOR2_X1 U9385 ( .A1(n7528), .A2(n7527), .ZN(n10094) );
  INV_X1 U9386 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10239) );
  XOR2_X1 U9387 ( .A(n10239), .B(P1_ADDR_REG_15__SCAN_IN), .Z(n10093) );
  NOR2_X1 U9388 ( .A1(n10094), .A2(n10093), .ZN(n7529) );
  NOR2_X1 U9389 ( .A1(n7530), .A2(n7529), .ZN(n10092) );
  XNOR2_X1 U9390 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10091) );
  NOR2_X1 U9391 ( .A1(n10092), .A2(n10091), .ZN(n7531) );
  NOR2_X1 U9392 ( .A1(n7532), .A2(n7531), .ZN(n10090) );
  XNOR2_X1 U9393 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10089) );
  NOR2_X1 U9394 ( .A1(n10090), .A2(n10089), .ZN(n7533) );
  NOR2_X1 U9395 ( .A1(n7534), .A2(n7533), .ZN(n7535) );
  AND2_X1 U9396 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7535), .ZN(n10086) );
  NOR2_X1 U9397 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10086), .ZN(n7536) );
  NOR2_X1 U9398 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7535), .ZN(n10087) );
  NOR2_X1 U9399 ( .A1(n7536), .A2(n10087), .ZN(n7538) );
  XNOR2_X1 U9400 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7537) );
  XNOR2_X1 U9401 ( .A(n7538), .B(n7537), .ZN(ADD_1068_U4) );
  INV_X1 U9402 ( .A(n7539), .ZN(n7543) );
  OAI222_X1 U9403 ( .A1(n7863), .A2(n7541), .B1(n8650), .B2(n7543), .C1(
        P2_U3151), .C2(n7540), .ZN(P2_U3273) );
  OAI222_X1 U9404 ( .A1(n7889), .A2(n10379), .B1(n9457), .B2(n7543), .C1(
        P1_U3086), .C2(n7542), .ZN(P1_U3333) );
  NAND2_X1 U9405 ( .A1(n7544), .A2(n7546), .ZN(n7545) );
  AND2_X1 U9406 ( .A1(n7587), .A2(n7545), .ZN(n7647) );
  INV_X1 U9407 ( .A(n7647), .ZN(n7557) );
  XNOR2_X1 U9408 ( .A(n7547), .B(n7546), .ZN(n7548) );
  OAI222_X1 U9409 ( .A1(n9993), .A2(n7682), .B1(n9995), .B2(n7549), .C1(n10000), .C2(n7548), .ZN(n7646) );
  NAND2_X1 U9410 ( .A1(n7646), .A2(n4500), .ZN(n7556) );
  OAI22_X1 U9411 ( .A1(n4500), .A2(n7551), .B1(n7550), .B2(n9989), .ZN(n7554)
         );
  INV_X1 U9412 ( .A(n7552), .ZN(n7651) );
  NOR2_X1 U9413 ( .A1(n8442), .A2(n7651), .ZN(n7553) );
  NOR2_X1 U9414 ( .A1(n7554), .A2(n7553), .ZN(n7555) );
  OAI211_X1 U9415 ( .C1(n7557), .C2(n8476), .A(n7556), .B(n7555), .ZN(P2_U3224) );
  INV_X1 U9416 ( .A(n7558), .ZN(n7560) );
  NAND2_X1 U9417 ( .A1(n7560), .A2(n7559), .ZN(n7574) );
  OAI21_X1 U9418 ( .B1(n7560), .B2(n7559), .A(n7574), .ZN(n7561) );
  NOR2_X1 U9419 ( .A1(n7561), .A2(n7562), .ZN(n7577) );
  AOI21_X1 U9420 ( .B1(n7562), .B2(n7561), .A(n7577), .ZN(n7567) );
  OAI22_X1 U9421 ( .A1(n9747), .A2(n8780), .B1(n8779), .B2(n9729), .ZN(n7565)
         );
  OAI22_X1 U9422 ( .A1(n8750), .A2(n7563), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5161), .ZN(n7564) );
  AOI211_X1 U9423 ( .C1(n9732), .C2(n8769), .A(n7565), .B(n7564), .ZN(n7566)
         );
  OAI21_X1 U9424 ( .B1(n7567), .B2(n8754), .A(n7566), .ZN(P1_U3221) );
  INV_X1 U9425 ( .A(n7571), .ZN(n7569) );
  AOI21_X1 U9426 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8647), .A(n8214), .ZN(
        n7568) );
  OAI21_X1 U9427 ( .B1(n7569), .B2(n8650), .A(n7568), .ZN(P2_U3272) );
  NAND2_X1 U9428 ( .A1(n7571), .A2(n7570), .ZN(n7572) );
  OAI211_X1 U9429 ( .C1(n7573), .C2(n7889), .A(n7572), .B(n9034), .ZN(P1_U3332) );
  INV_X1 U9430 ( .A(n7574), .ZN(n7575) );
  NOR3_X1 U9431 ( .A1(n7577), .A2(n7576), .A3(n7575), .ZN(n7580) );
  INV_X1 U9432 ( .A(n7578), .ZN(n7579) );
  OAI21_X1 U9433 ( .B1(n7580), .B2(n7579), .A(n8777), .ZN(n7586) );
  NOR2_X1 U9434 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7581), .ZN(n9103) );
  OAI22_X1 U9435 ( .A1(n7704), .A2(n8780), .B1(n8779), .B2(n7582), .ZN(n7583)
         );
  AOI211_X1 U9436 ( .C1(n6010), .C2(n7584), .A(n9103), .B(n7583), .ZN(n7585)
         );
  OAI211_X1 U9437 ( .C1(n4893), .C2(n8786), .A(n7586), .B(n7585), .ZN(P1_U3231) );
  NAND2_X1 U9438 ( .A1(n7587), .A2(n8086), .ZN(n7589) );
  NAND2_X1 U9439 ( .A1(n8114), .A2(n8111), .ZN(n8034) );
  INV_X1 U9440 ( .A(n8034), .ZN(n7588) );
  XNOR2_X1 U9441 ( .A(n7589), .B(n7588), .ZN(n10047) );
  XNOR2_X1 U9442 ( .A(n7590), .B(n8034), .ZN(n7591) );
  NAND2_X1 U9443 ( .A1(n7591), .A2(n8484), .ZN(n7593) );
  AOI22_X1 U9444 ( .A1(n8224), .A2(n8479), .B1(n8481), .B2(n8226), .ZN(n7592)
         );
  OAI211_X1 U9445 ( .C1(n10047), .C2(n9992), .A(n7593), .B(n7592), .ZN(n10049)
         );
  NAND2_X1 U9446 ( .A1(n10049), .A2(n4500), .ZN(n7599) );
  OAI22_X1 U9447 ( .A1(n4500), .A2(n7595), .B1(n7594), .B2(n9989), .ZN(n7596)
         );
  AOI21_X1 U9448 ( .B1(n8473), .B2(n7597), .A(n7596), .ZN(n7598) );
  OAI211_X1 U9449 ( .C1(n10047), .C2(n7827), .A(n7599), .B(n7598), .ZN(
        P2_U3223) );
  NOR2_X1 U9450 ( .A1(n7601), .A2(n7600), .ZN(n7603) );
  AOI22_X1 U9451 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8244), .B1(n8236), .B2(
        n7615), .ZN(n7602) );
  AOI21_X1 U9452 ( .B1(n7603), .B2(n7602), .A(n8235), .ZN(n7626) );
  AOI22_X1 U9453 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8236), .B1(n8244), .B2(
        n7614), .ZN(n7609) );
  NAND2_X1 U9454 ( .A1(n7605), .A2(n7604), .ZN(n7607) );
  NAND2_X1 U9455 ( .A1(n7607), .A2(n7606), .ZN(n7608) );
  NAND2_X1 U9456 ( .A1(n7609), .A2(n7608), .ZN(n8243) );
  OAI21_X1 U9457 ( .B1(n7609), .B2(n7608), .A(n8243), .ZN(n7624) );
  INV_X1 U9458 ( .A(n7610), .ZN(n7612) );
  MUX2_X1 U9459 ( .A(n7615), .B(n7614), .S(n8273), .Z(n7616) );
  NOR2_X1 U9460 ( .A1(n7616), .A2(n8244), .ZN(n8259) );
  NOR2_X1 U9461 ( .A1(n8259), .A2(n4594), .ZN(n7618) );
  NAND2_X1 U9462 ( .A1(n8260), .A2(n7618), .ZN(n7617) );
  OAI211_X1 U9463 ( .C1(n8260), .C2(n7618), .A(n9973), .B(n7617), .ZN(n7621)
         );
  NOR2_X1 U9464 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7619), .ZN(n7656) );
  AOI21_X1 U9465 ( .B1(n9964), .B2(n8244), .A(n7656), .ZN(n7620) );
  OAI211_X1 U9466 ( .C1(n7622), .C2(n9897), .A(n7621), .B(n7620), .ZN(n7623)
         );
  AOI21_X1 U9467 ( .B1(n7624), .B2(n9974), .A(n7623), .ZN(n7625) );
  OAI21_X1 U9468 ( .B1(n7626), .B2(n9980), .A(n7625), .ZN(P2_U3194) );
  INV_X1 U9469 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10272) );
  XNOR2_X1 U9470 ( .A(n7716), .B(n7709), .ZN(n7628) );
  NOR2_X1 U9471 ( .A1(n10272), .A2(n7628), .ZN(n7710) );
  AOI21_X1 U9472 ( .B1(n10272), .B2(n7628), .A(n7710), .ZN(n7636) );
  INV_X1 U9473 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9535) );
  XNOR2_X1 U9474 ( .A(n7716), .B(n7717), .ZN(n7631) );
  NOR2_X1 U9475 ( .A1(n9535), .A2(n7631), .ZN(n7718) );
  AOI21_X1 U9476 ( .B1(n9535), .B2(n7631), .A(n7718), .ZN(n7632) );
  NAND2_X1 U9477 ( .A1(n7632), .A2(n9595), .ZN(n7634) );
  AND2_X1 U9478 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8782) );
  AOI21_X1 U9479 ( .B1(n9553), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n8782), .ZN(
        n7633) );
  OAI211_X1 U9480 ( .C1(n9599), .C2(n7716), .A(n7634), .B(n7633), .ZN(n7635)
         );
  AOI21_X1 U9481 ( .B1(n7636), .B2(n9590), .A(n7635), .ZN(n7637) );
  INV_X1 U9482 ( .A(n7637), .ZN(P1_U3258) );
  INV_X1 U9483 ( .A(n7638), .ZN(n7701) );
  AOI21_X1 U9484 ( .B1(n7640), .B2(n7639), .A(n7701), .ZN(n7645) );
  NAND2_X1 U9485 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9490) );
  INV_X1 U9486 ( .A(n9490), .ZN(n7642) );
  OAI22_X1 U9487 ( .A1(n9748), .A2(n8780), .B1(n8779), .B2(n9747), .ZN(n7641)
         );
  AOI211_X1 U9488 ( .C1(n6010), .C2(n5080), .A(n7642), .B(n7641), .ZN(n7644)
         );
  NAND2_X1 U9489 ( .A1(n9751), .A2(n8769), .ZN(n7643) );
  OAI211_X1 U9490 ( .C1(n7645), .C2(n8754), .A(n7644), .B(n7643), .ZN(P1_U3217) );
  AOI21_X1 U9491 ( .B1(n7647), .B2(n10030), .A(n7646), .ZN(n7649) );
  MUX2_X1 U9492 ( .A(n6209), .B(n7649), .S(n10063), .Z(n7648) );
  OAI21_X1 U9493 ( .B1(n7651), .B2(n8620), .A(n7648), .ZN(P2_U3417) );
  MUX2_X1 U9494 ( .A(n7329), .B(n7649), .S(n10081), .Z(n7650) );
  OAI21_X1 U9495 ( .B1(n7651), .B2(n8537), .A(n7650), .ZN(P2_U3468) );
  XNOR2_X1 U9496 ( .A(n7652), .B(n8496), .ZN(n7653) );
  XNOR2_X1 U9497 ( .A(n7654), .B(n7653), .ZN(n7660) );
  NOR2_X1 U9498 ( .A1(n7981), .A2(n8116), .ZN(n7655) );
  AOI211_X1 U9499 ( .C1(n7979), .C2(n8482), .A(n7656), .B(n7655), .ZN(n7657)
         );
  OAI21_X1 U9500 ( .B1(n7746), .B2(n8003), .A(n7657), .ZN(n7658) );
  AOI21_X1 U9501 ( .B1(n7748), .B2(n7968), .A(n7658), .ZN(n7659) );
  OAI21_X1 U9502 ( .B1(n7660), .B2(n7970), .A(n7659), .ZN(P2_U3164) );
  INV_X1 U9503 ( .A(n7661), .ZN(n7676) );
  OAI222_X1 U9504 ( .A1(n8650), .A2(n7676), .B1(P2_U3151), .B2(n6472), .C1(
        n7662), .C2(n7863), .ZN(P2_U3271) );
  INV_X1 U9505 ( .A(n7663), .ZN(n7664) );
  AOI211_X1 U9506 ( .C1(n7666), .C2(n7665), .A(n7970), .B(n7664), .ZN(n7674)
         );
  AOI21_X1 U9507 ( .B1(n8006), .B2(n8225), .A(n7667), .ZN(n7672) );
  NAND2_X1 U9508 ( .A1(n10054), .A2(n7968), .ZN(n7671) );
  INV_X1 U9509 ( .A(n7683), .ZN(n7668) );
  NAND2_X1 U9510 ( .A1(n7994), .A2(n7668), .ZN(n7670) );
  NAND2_X1 U9511 ( .A1(n7979), .A2(n8223), .ZN(n7669) );
  NAND4_X1 U9512 ( .A1(n7672), .A2(n7671), .A3(n7670), .A4(n7669), .ZN(n7673)
         );
  OR2_X1 U9513 ( .A1(n7674), .A2(n7673), .ZN(P2_U3176) );
  OAI222_X1 U9514 ( .A1(n7677), .A2(P1_U3086), .B1(n9457), .B2(n7676), .C1(
        n7675), .C2(n7889), .ZN(P1_U3331) );
  XNOR2_X1 U9515 ( .A(n7678), .B(n7679), .ZN(n10051) );
  XNOR2_X1 U9516 ( .A(n7680), .B(n7679), .ZN(n7681) );
  OAI222_X1 U9517 ( .A1(n9993), .A2(n8496), .B1(n9995), .B2(n7682), .C1(n7681), 
        .C2(n10000), .ZN(n10052) );
  NAND2_X1 U9518 ( .A1(n10052), .A2(n4500), .ZN(n7686) );
  OAI22_X1 U9519 ( .A1(n4500), .A2(n6244), .B1(n7683), .B2(n9989), .ZN(n7684)
         );
  AOI21_X1 U9520 ( .B1(n8473), .B2(n10054), .A(n7684), .ZN(n7685) );
  OAI211_X1 U9521 ( .C1(n8476), .C2(n10051), .A(n7686), .B(n7685), .ZN(
        P2_U3222) );
  XNOR2_X1 U9522 ( .A(n7687), .B(n9001), .ZN(n9797) );
  AOI211_X1 U9523 ( .C1(n9793), .C2(n9620), .A(n9321), .B(n4589), .ZN(n9791)
         );
  AOI22_X1 U9524 ( .A1(n9634), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8662), .B2(
        n9651), .ZN(n7688) );
  OAI21_X1 U9525 ( .B1(n9307), .B2(n9788), .A(n7688), .ZN(n7689) );
  AOI21_X1 U9526 ( .B1(n9310), .B2(n9046), .A(n7689), .ZN(n7690) );
  OAI21_X1 U9527 ( .B1(n8665), .B2(n9668), .A(n7690), .ZN(n7696) );
  NAND2_X1 U9528 ( .A1(n7691), .A2(n9001), .ZN(n7692) );
  NAND2_X1 U9529 ( .A1(n7693), .A2(n7692), .ZN(n7694) );
  NAND2_X1 U9530 ( .A1(n7694), .A2(n9777), .ZN(n9794) );
  NOR2_X1 U9531 ( .A1(n9794), .A2(n9634), .ZN(n7695) );
  AOI211_X1 U9532 ( .C1(n9791), .C2(n9676), .A(n7696), .B(n7695), .ZN(n7697)
         );
  OAI21_X1 U9533 ( .B1(n9797), .B2(n9336), .A(n7697), .ZN(P1_U3279) );
  INV_X1 U9534 ( .A(n7698), .ZN(n7700) );
  NOR3_X1 U9535 ( .A1(n7701), .A2(n7700), .A3(n7699), .ZN(n7703) );
  INV_X1 U9536 ( .A(n7702), .ZN(n7757) );
  OAI21_X1 U9537 ( .B1(n7703), .B2(n7757), .A(n8777), .ZN(n7708) );
  NAND2_X1 U9538 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9601) );
  INV_X1 U9539 ( .A(n9601), .ZN(n7706) );
  OAI22_X1 U9540 ( .A1(n9611), .A2(n8780), .B1(n8779), .B2(n7704), .ZN(n7705)
         );
  AOI211_X1 U9541 ( .C1(n6010), .C2(n9635), .A(n7706), .B(n7705), .ZN(n7707)
         );
  OAI211_X1 U9542 ( .C1(n9759), .C2(n8786), .A(n7708), .B(n7707), .ZN(P1_U3236) );
  NOR2_X1 U9543 ( .A1(n7709), .A2(n7716), .ZN(n7711) );
  NAND2_X1 U9544 ( .A1(n7776), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7712) );
  OAI21_X1 U9545 ( .B1(n7776), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7712), .ZN(
        n7713) );
  NOR2_X1 U9546 ( .A1(n7714), .A2(n7713), .ZN(n7771) );
  AOI21_X1 U9547 ( .B1(n7714), .B2(n7713), .A(n7771), .ZN(n7728) );
  INV_X1 U9548 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7715) );
  AOI22_X1 U9549 ( .A1(n7776), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n7715), .B2(
        n7726), .ZN(n7721) );
  NOR2_X1 U9550 ( .A1(n7717), .A2(n7716), .ZN(n7719) );
  OAI21_X1 U9551 ( .B1(n7721), .B2(n7720), .A(n7775), .ZN(n7722) );
  NAND2_X1 U9552 ( .A1(n7722), .A2(n9595), .ZN(n7725) );
  NOR2_X1 U9553 ( .A1(n7723), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8708) );
  AOI21_X1 U9554 ( .B1(n9553), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n8708), .ZN(
        n7724) );
  OAI211_X1 U9555 ( .C1(n9599), .C2(n7726), .A(n7725), .B(n7724), .ZN(n7727)
         );
  AOI21_X1 U9556 ( .B1(n7728), .B2(n9590), .A(n7727), .ZN(n7729) );
  INV_X1 U9557 ( .A(n7729), .ZN(P1_U3259) );
  INV_X1 U9558 ( .A(n7730), .ZN(n7753) );
  OAI222_X1 U9559 ( .A1(n8650), .A2(n7753), .B1(P2_U3151), .B2(n7732), .C1(
        n7731), .C2(n7863), .ZN(P2_U3270) );
  XNOR2_X1 U9560 ( .A(n7733), .B(n8127), .ZN(n7734) );
  XNOR2_X1 U9561 ( .A(n7735), .B(n7734), .ZN(n7741) );
  NAND2_X1 U9562 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9911) );
  INV_X1 U9563 ( .A(n9911), .ZN(n7737) );
  NOR2_X1 U9564 ( .A1(n7981), .A2(n8496), .ZN(n7736) );
  AOI211_X1 U9565 ( .C1(n7979), .C2(n8467), .A(n7737), .B(n7736), .ZN(n7738)
         );
  OAI21_X1 U9566 ( .B1(n8498), .B2(n8003), .A(n7738), .ZN(n7739) );
  AOI21_X1 U9567 ( .B1(n8129), .B2(n7968), .A(n7739), .ZN(n7740) );
  OAI21_X1 U9568 ( .B1(n7741), .B2(n7970), .A(n7740), .ZN(P2_U3174) );
  XNOR2_X1 U9569 ( .A(n7742), .B(n7743), .ZN(n10060) );
  INV_X1 U9570 ( .A(n7743), .ZN(n8121) );
  XNOR2_X1 U9571 ( .A(n7744), .B(n8121), .ZN(n7745) );
  OAI222_X1 U9572 ( .A1(n9993), .A2(n8127), .B1(n9995), .B2(n8116), .C1(n7745), 
        .C2(n10000), .ZN(n10062) );
  NAND2_X1 U9573 ( .A1(n10062), .A2(n4500), .ZN(n7750) );
  OAI22_X1 U9574 ( .A1(n4500), .A2(n7615), .B1(n7746), .B2(n9989), .ZN(n7747)
         );
  AOI21_X1 U9575 ( .B1(n7748), .B2(n8473), .A(n7747), .ZN(n7749) );
  OAI211_X1 U9576 ( .C1(n8476), .C2(n10060), .A(n7750), .B(n7749), .ZN(
        P2_U3221) );
  INV_X1 U9577 ( .A(n7751), .ZN(n7754) );
  OAI222_X1 U9578 ( .A1(n7754), .A2(P1_U3086), .B1(n9457), .B2(n7753), .C1(
        n7752), .C2(n7889), .ZN(P1_U3330) );
  NOR3_X1 U9579 ( .A1(n7757), .A2(n4615), .A3(n7756), .ZN(n7760) );
  INV_X1 U9580 ( .A(n7758), .ZN(n7759) );
  OAI21_X1 U9581 ( .B1(n7760), .B2(n7759), .A(n8777), .ZN(n7765) );
  OAI22_X1 U9582 ( .A1(n9788), .A2(n8780), .B1(n8779), .B2(n9748), .ZN(n7761)
         );
  AOI211_X1 U9583 ( .C1(n6010), .C2(n7763), .A(n7762), .B(n7761), .ZN(n7764)
         );
  OAI211_X1 U9584 ( .C1(n4820), .C2(n8786), .A(n7765), .B(n7764), .ZN(P1_U3224) );
  INV_X1 U9585 ( .A(n7766), .ZN(n7769) );
  OAI222_X1 U9586 ( .A1(n8650), .A2(n7769), .B1(P2_U3151), .B2(n7767), .C1(
        n10369), .C2(n7863), .ZN(P2_U3269) );
  OAI222_X1 U9587 ( .A1(n7770), .A2(P1_U3086), .B1(n9457), .B2(n7769), .C1(
        n7768), .C2(n7889), .ZN(P1_U3329) );
  INV_X1 U9588 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U9589 ( .A1(n7877), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10336), .B2(
        n7783), .ZN(n7773) );
  NAND2_X1 U9590 ( .A1(n7773), .A2(n7772), .ZN(n7870) );
  OAI21_X1 U9591 ( .B1(n7773), .B2(n7772), .A(n7870), .ZN(n7785) );
  INV_X1 U9592 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7774) );
  AOI22_X1 U9593 ( .A1(n7877), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n7774), .B2(
        n7783), .ZN(n7778) );
  OAI21_X1 U9594 ( .B1(n7776), .B2(P1_REG1_REG_16__SCAN_IN), .A(n7775), .ZN(
        n7777) );
  NAND2_X1 U9595 ( .A1(n7778), .A2(n7777), .ZN(n7876) );
  OAI21_X1 U9596 ( .B1(n7778), .B2(n7777), .A(n7876), .ZN(n7779) );
  NAND2_X1 U9597 ( .A1(n7779), .A2(n9595), .ZN(n7782) );
  NOR2_X1 U9598 ( .A1(n7780), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8719) );
  AOI21_X1 U9599 ( .B1(n9553), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n8719), .ZN(
        n7781) );
  OAI211_X1 U9600 ( .C1(n9599), .C2(n7783), .A(n7782), .B(n7781), .ZN(n7784)
         );
  AOI21_X1 U9601 ( .B1(n7785), .B2(n9590), .A(n7784), .ZN(n7786) );
  INV_X1 U9602 ( .A(n7786), .ZN(P1_U3260) );
  INV_X1 U9603 ( .A(n7787), .ZN(n7868) );
  NAND2_X1 U9604 ( .A1(n8647), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7788) );
  OAI211_X1 U9605 ( .C1(n7868), .C2(n8650), .A(n7789), .B(n7788), .ZN(P2_U3268) );
  OAI21_X1 U9606 ( .B1(n7792), .B2(n7791), .A(n7790), .ZN(n7793) );
  NAND2_X1 U9607 ( .A1(n7793), .A2(n8777), .ZN(n7797) );
  OAI22_X1 U9608 ( .A1(n9612), .A2(n8780), .B1(n8779), .B2(n9611), .ZN(n7794)
         );
  AOI211_X1 U9609 ( .C1(n6010), .C2(n9615), .A(n7795), .B(n7794), .ZN(n7796)
         );
  OAI211_X1 U9610 ( .C1(n9782), .C2(n8786), .A(n7797), .B(n7796), .ZN(P1_U3234) );
  AOI211_X1 U9611 ( .C1(n9002), .C2(n7799), .A(n9754), .B(n7798), .ZN(n7801)
         );
  OAI22_X1 U9612 ( .A1(n9329), .A2(n9789), .B1(n9612), .B2(n9787), .ZN(n7800)
         );
  NOR2_X1 U9613 ( .A1(n7801), .A2(n7800), .ZN(n9531) );
  XOR2_X1 U9614 ( .A(n7802), .B(n9002), .Z(n9534) );
  NAND2_X1 U9615 ( .A1(n9534), .A2(n9677), .ZN(n7807) );
  OAI211_X1 U9616 ( .C1(n9532), .C2(n4589), .A(n9673), .B(n7813), .ZN(n9530)
         );
  INV_X1 U9617 ( .A(n9530), .ZN(n7805) );
  AOI22_X1 U9618 ( .A1(n9634), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8783), .B2(
        n9651), .ZN(n7803) );
  OAI21_X1 U9619 ( .B1(n9532), .B2(n9668), .A(n7803), .ZN(n7804) );
  AOI21_X1 U9620 ( .B1(n7805), .B2(n9676), .A(n7804), .ZN(n7806) );
  OAI211_X1 U9621 ( .C1(n9666), .C2(n9531), .A(n7807), .B(n7806), .ZN(P1_U3278) );
  INV_X1 U9622 ( .A(n7808), .ZN(n7888) );
  AOI21_X1 U9623 ( .B1(n8647), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7809), .ZN(
        n7810) );
  OAI21_X1 U9624 ( .B1(n7888), .B2(n8650), .A(n7810), .ZN(P2_U3267) );
  XNOR2_X1 U9625 ( .A(n7811), .B(n9004), .ZN(n9434) );
  INV_X1 U9626 ( .A(n7812), .ZN(n9322) );
  AOI211_X1 U9627 ( .C1(n9431), .C2(n7813), .A(n9321), .B(n7812), .ZN(n9430)
         );
  INV_X1 U9628 ( .A(n9431), .ZN(n8712) );
  AOI22_X1 U9629 ( .A1(n9634), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8709), .B2(
        n9651), .ZN(n7814) );
  OAI21_X1 U9630 ( .B1(n8712), .B2(n9668), .A(n7814), .ZN(n7819) );
  AOI211_X1 U9631 ( .C1(n7815), .C2(n9004), .A(n9754), .B(n4584), .ZN(n7817)
         );
  OAI22_X1 U9632 ( .A1(n9418), .A2(n9789), .B1(n9790), .B2(n9787), .ZN(n7816)
         );
  NOR2_X1 U9633 ( .A1(n7817), .A2(n7816), .ZN(n9433) );
  NOR2_X1 U9634 ( .A1(n9433), .A2(n9634), .ZN(n7818) );
  AOI211_X1 U9635 ( .C1(n9430), .C2(n9676), .A(n7819), .B(n7818), .ZN(n7820)
         );
  OAI21_X1 U9636 ( .B1(n9434), .B2(n9336), .A(n7820), .ZN(P1_U3277) );
  NAND2_X1 U9637 ( .A1(n7821), .A2(n4500), .ZN(n7826) );
  NOR2_X1 U9638 ( .A1(n7822), .A2(n9989), .ZN(n8288) );
  NOR2_X1 U9639 ( .A1(n7823), .A2(n8442), .ZN(n7824) );
  AOI211_X1 U9640 ( .C1(n10005), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8288), .B(
        n7824), .ZN(n7825) );
  OAI211_X1 U9641 ( .C1(n6644), .C2(n7827), .A(n7826), .B(n7825), .ZN(P2_U3204) );
  INV_X1 U9642 ( .A(n7828), .ZN(n7834) );
  XNOR2_X1 U9643 ( .A(n8320), .B(n7829), .ZN(n7830) );
  XNOR2_X1 U9644 ( .A(n8304), .B(n7830), .ZN(n7831) );
  INV_X1 U9645 ( .A(n7831), .ZN(n7835) );
  OAI211_X1 U9646 ( .C1(n8333), .C2(n7834), .A(n7835), .B(n7997), .ZN(n7839)
         );
  AOI22_X1 U9647 ( .A1(n8298), .A2(n7979), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7833) );
  NAND2_X1 U9648 ( .A1(n8303), .A2(n7994), .ZN(n7832) );
  OAI211_X1 U9649 ( .C1(n8333), .C2(n7981), .A(n7833), .B(n7832), .ZN(n7837)
         );
  NOR4_X1 U9650 ( .A1(n7835), .A2(n7834), .A3(n8333), .A4(n7970), .ZN(n7836)
         );
  AOI211_X1 U9651 ( .C1(n8304), .C2(n7968), .A(n7837), .B(n7836), .ZN(n7838)
         );
  INV_X1 U9652 ( .A(n6898), .ZN(n7843) );
  AOI21_X1 U9653 ( .B1(n7841), .B2(n7842), .A(n7843), .ZN(n7847) );
  AOI22_X1 U9654 ( .A1(n7844), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n5761), .B2(
        n8769), .ZN(n7846) );
  AOI22_X1 U9655 ( .A1(n8768), .A2(n5779), .B1(n8767), .B2(n6712), .ZN(n7845)
         );
  OAI211_X1 U9656 ( .C1(n7847), .C2(n8754), .A(n7846), .B(n7845), .ZN(P1_U3222) );
  INV_X1 U9657 ( .A(n7848), .ZN(n7866) );
  OAI222_X1 U9658 ( .A1(n7889), .A2(n10361), .B1(n9457), .B2(n7866), .C1(n7849), .C2(P1_U3086), .ZN(P1_U3326) );
  INV_X1 U9659 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10398) );
  INV_X1 U9660 ( .A(SI_29_), .ZN(n7850) );
  INV_X1 U9661 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7857) );
  MUX2_X1 U9662 ( .A(n7857), .B(n10398), .S(n7856), .Z(n7859) );
  INV_X1 U9663 ( .A(SI_30_), .ZN(n7858) );
  NAND2_X1 U9664 ( .A1(n7859), .A2(n7858), .ZN(n8011) );
  INV_X1 U9665 ( .A(n7859), .ZN(n7860) );
  NAND2_X1 U9666 ( .A1(n7860), .A2(SI_30_), .ZN(n7861) );
  NAND2_X1 U9667 ( .A1(n8011), .A2(n7861), .ZN(n8012) );
  INV_X1 U9668 ( .A(n8885), .ZN(n8651) );
  OAI222_X1 U9669 ( .A1(n7889), .A2(n10398), .B1(n9457), .B2(n8651), .C1(
        P1_U3086), .C2(n7862), .ZN(P1_U3325) );
  OAI222_X1 U9670 ( .A1(n8650), .A2(n7866), .B1(n7865), .B2(P2_U3151), .C1(
        n10301), .C2(n7863), .ZN(P2_U3266) );
  OAI222_X1 U9671 ( .A1(n7889), .A2(n7869), .B1(n9457), .B2(n7868), .C1(n7867), 
        .C2(P1_U3086), .ZN(P1_U3328) );
  OAI21_X1 U9672 ( .B1(n7877), .B2(P1_REG2_REG_17__SCAN_IN), .A(n7870), .ZN(
        n7871) );
  INV_X1 U9673 ( .A(n7871), .ZN(n9115) );
  NAND2_X1 U9674 ( .A1(n9121), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7873) );
  OAI21_X1 U9675 ( .B1(n9121), .B2(P1_REG2_REG_18__SCAN_IN), .A(n7873), .ZN(
        n7872) );
  INV_X1 U9676 ( .A(n7872), .ZN(n9114) );
  NAND2_X1 U9677 ( .A1(n9115), .A2(n9114), .ZN(n9113) );
  NAND2_X1 U9678 ( .A1(n9113), .A2(n7873), .ZN(n7875) );
  INV_X1 U9679 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n7874) );
  INV_X1 U9680 ( .A(n7882), .ZN(n7880) );
  OAI21_X1 U9681 ( .B1(n7877), .B2(P1_REG1_REG_17__SCAN_IN), .A(n7876), .ZN(
        n9118) );
  NAND2_X1 U9682 ( .A1(n9121), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7878) );
  OAI21_X1 U9683 ( .B1(n9121), .B2(P1_REG1_REG_18__SCAN_IN), .A(n7878), .ZN(
        n9117) );
  OR2_X1 U9684 ( .A1(n9118), .A2(n9117), .ZN(n9119) );
  OAI21_X1 U9685 ( .B1(n7881), .B2(n9543), .A(n9599), .ZN(n7879) );
  AOI21_X1 U9686 ( .B1(n7880), .B2(n9590), .A(n7879), .ZN(n7884) );
  AOI22_X1 U9687 ( .A1(n7882), .A2(n9590), .B1(n9595), .B2(n7881), .ZN(n7883)
         );
  NOR2_X1 U9688 ( .A1(n7885), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8684) );
  INV_X1 U9689 ( .A(n8684), .ZN(n7886) );
  OAI222_X1 U9690 ( .A1(n7889), .A2(n10378), .B1(n9457), .B2(n7888), .C1(n4502), .C2(P1_U3086), .ZN(P1_U3327) );
  XOR2_X1 U9691 ( .A(n7891), .B(n7890), .Z(n7896) );
  AOI22_X1 U9692 ( .A1(n8006), .A2(n8482), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7893) );
  NAND2_X1 U9693 ( .A1(n7979), .A2(n8480), .ZN(n7892) );
  OAI211_X1 U9694 ( .C1(n8489), .C2(n8003), .A(n7893), .B(n7892), .ZN(n7894)
         );
  AOI21_X1 U9695 ( .B1(n8637), .B2(n7968), .A(n7894), .ZN(n7895) );
  OAI21_X1 U9696 ( .B1(n7896), .B2(n7970), .A(n7895), .ZN(P2_U3155) );
  AOI21_X1 U9697 ( .B1(n8380), .B2(n7897), .A(n4509), .ZN(n7902) );
  AOI22_X1 U9698 ( .A1(n8369), .A2(n7979), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7899) );
  NAND2_X1 U9699 ( .A1(n7994), .A2(n8372), .ZN(n7898) );
  OAI211_X1 U9700 ( .C1(n7960), .C2(n7981), .A(n7899), .B(n7898), .ZN(n7900)
         );
  AOI21_X1 U9701 ( .B1(n8588), .B2(n7968), .A(n7900), .ZN(n7901) );
  OAI21_X1 U9702 ( .B1(n7902), .B2(n7970), .A(n7901), .ZN(P2_U3156) );
  XOR2_X1 U9703 ( .A(n7904), .B(n7903), .Z(n7910) );
  AOI22_X1 U9704 ( .A1(n7979), .A2(n8415), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n7906) );
  NAND2_X1 U9705 ( .A1(n7994), .A2(n8418), .ZN(n7905) );
  OAI211_X1 U9706 ( .C1(n7907), .C2(n7981), .A(n7906), .B(n7905), .ZN(n7908)
         );
  AOI21_X1 U9707 ( .B1(n8612), .B2(n7968), .A(n7908), .ZN(n7909) );
  OAI21_X1 U9708 ( .B1(n7910), .B2(n7970), .A(n7909), .ZN(P2_U3159) );
  XOR2_X1 U9709 ( .A(n7912), .B(n7911), .Z(n7918) );
  AOI22_X1 U9710 ( .A1(n7979), .A2(n8395), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7914) );
  NAND2_X1 U9711 ( .A1(n7994), .A2(n8398), .ZN(n7913) );
  OAI211_X1 U9712 ( .C1(n7915), .C2(n7981), .A(n7914), .B(n7913), .ZN(n7916)
         );
  AOI21_X1 U9713 ( .B1(n8600), .B2(n7968), .A(n7916), .ZN(n7917) );
  OAI21_X1 U9714 ( .B1(n7918), .B2(n7970), .A(n7917), .ZN(P2_U3163) );
  INV_X1 U9715 ( .A(n7919), .ZN(n7947) );
  INV_X1 U9716 ( .A(n7920), .ZN(n7922) );
  NOR3_X1 U9717 ( .A1(n7947), .A2(n7922), .A3(n7921), .ZN(n7924) );
  INV_X1 U9718 ( .A(n7923), .ZN(n7988) );
  OAI21_X1 U9719 ( .B1(n7924), .B2(n7988), .A(n7997), .ZN(n7928) );
  AOI22_X1 U9720 ( .A1(n8319), .A2(n7979), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7925) );
  OAI21_X1 U9721 ( .B1(n8347), .B2(n7981), .A(n7925), .ZN(n7926) );
  AOI21_X1 U9722 ( .B1(n8349), .B2(n7994), .A(n7926), .ZN(n7927) );
  OAI211_X1 U9723 ( .C1(n8576), .C2(n8009), .A(n7928), .B(n7927), .ZN(P2_U3165) );
  OAI211_X1 U9724 ( .C1(n7931), .C2(n7930), .A(n7929), .B(n7997), .ZN(n7935)
         );
  NAND2_X1 U9725 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9961) );
  OAI21_X1 U9726 ( .B1(n8002), .B2(n8423), .A(n9961), .ZN(n7933) );
  NOR2_X1 U9727 ( .A1(n8003), .A2(n8458), .ZN(n7932) );
  AOI211_X1 U9728 ( .C1(n8006), .C2(n8480), .A(n7933), .B(n7932), .ZN(n7934)
         );
  OAI211_X1 U9729 ( .C1(n7936), .C2(n8009), .A(n7935), .B(n7934), .ZN(P2_U3166) );
  INV_X1 U9730 ( .A(n7937), .ZN(n7975) );
  AOI21_X1 U9731 ( .B1(n7939), .B2(n7938), .A(n7975), .ZN(n7944) );
  AOI22_X1 U9732 ( .A1(n7979), .A2(n8437), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n7941) );
  NAND2_X1 U9733 ( .A1(n8006), .A2(n8468), .ZN(n7940) );
  OAI211_X1 U9734 ( .C1(n8003), .C2(n8444), .A(n7941), .B(n7940), .ZN(n7942)
         );
  AOI21_X1 U9735 ( .B1(n8538), .B2(n7968), .A(n7942), .ZN(n7943) );
  OAI21_X1 U9736 ( .B1(n7944), .B2(n7970), .A(n7943), .ZN(P2_U3168) );
  NOR3_X1 U9737 ( .A1(n4509), .A2(n4942), .A3(n7946), .ZN(n7948) );
  OAI21_X1 U9738 ( .B1(n7948), .B2(n7947), .A(n7997), .ZN(n7952) );
  AOI22_X1 U9739 ( .A1(n8360), .A2(n7979), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7949) );
  OAI21_X1 U9740 ( .B1(n7966), .B2(n7981), .A(n7949), .ZN(n7950) );
  AOI21_X1 U9741 ( .B1(n8363), .B2(n7994), .A(n7950), .ZN(n7951) );
  OAI211_X1 U9742 ( .C1(n8585), .C2(n8009), .A(n7952), .B(n7951), .ZN(P2_U3169) );
  XOR2_X1 U9743 ( .A(n7954), .B(n7953), .Z(n7959) );
  AOI22_X1 U9744 ( .A1(n7979), .A2(n8406), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7956) );
  NAND2_X1 U9745 ( .A1(n7994), .A2(n8409), .ZN(n7955) );
  OAI211_X1 U9746 ( .C1(n8424), .C2(n7981), .A(n7956), .B(n7955), .ZN(n7957)
         );
  AOI21_X1 U9747 ( .B1(n8606), .B2(n7968), .A(n7957), .ZN(n7958) );
  OAI21_X1 U9748 ( .B1(n7959), .B2(n7970), .A(n7958), .ZN(P2_U3173) );
  XNOR2_X1 U9749 ( .A(n7961), .B(n7960), .ZN(n7962) );
  XNOR2_X1 U9750 ( .A(n4495), .B(n7962), .ZN(n7971) );
  AOI22_X1 U9751 ( .A1(n8006), .A2(n8406), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n7965) );
  NAND2_X1 U9752 ( .A1(n7994), .A2(n8383), .ZN(n7964) );
  OAI211_X1 U9753 ( .C1(n7966), .C2(n8002), .A(n7965), .B(n7964), .ZN(n7967)
         );
  AOI21_X1 U9754 ( .B1(n8594), .B2(n7968), .A(n7967), .ZN(n7969) );
  OAI21_X1 U9755 ( .B1(n7971), .B2(n7970), .A(n7969), .ZN(P2_U3175) );
  INV_X1 U9756 ( .A(n7972), .ZN(n7974) );
  NOR3_X1 U9757 ( .A1(n7975), .A2(n7974), .A3(n7973), .ZN(n7978) );
  INV_X1 U9758 ( .A(n7976), .ZN(n7977) );
  OAI21_X1 U9759 ( .B1(n7978), .B2(n7977), .A(n7997), .ZN(n7984) );
  AOI22_X1 U9760 ( .A1(n7979), .A2(n8405), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n7980) );
  OAI21_X1 U9761 ( .B1(n8423), .B2(n7981), .A(n7980), .ZN(n7982) );
  AOI21_X1 U9762 ( .B1(n8429), .B2(n7994), .A(n7982), .ZN(n7983) );
  OAI211_X1 U9763 ( .C1(n8621), .C2(n8009), .A(n7984), .B(n7983), .ZN(P2_U3178) );
  INV_X1 U9764 ( .A(n7985), .ZN(n7987) );
  NOR3_X1 U9765 ( .A1(n7988), .A2(n7987), .A3(n7986), .ZN(n7991) );
  INV_X1 U9766 ( .A(n7989), .ZN(n7990) );
  OAI21_X1 U9767 ( .B1(n7991), .B2(n7990), .A(n7997), .ZN(n7996) );
  AOI22_X1 U9768 ( .A1(n8360), .A2(n8006), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n7992) );
  OAI21_X1 U9769 ( .B1(n8333), .B2(n8002), .A(n7992), .ZN(n7993) );
  AOI21_X1 U9770 ( .B1(n8339), .B2(n7994), .A(n7993), .ZN(n7995) );
  OAI211_X1 U9771 ( .C1(n8571), .C2(n8009), .A(n7996), .B(n7995), .ZN(P2_U3180) );
  OAI211_X1 U9772 ( .C1(n8000), .C2(n7999), .A(n7998), .B(n7997), .ZN(n8008)
         );
  NAND2_X1 U9773 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9944) );
  OAI21_X1 U9774 ( .B1(n8002), .B2(n8001), .A(n9944), .ZN(n8005) );
  NOR2_X1 U9775 ( .A1(n8003), .A2(n8470), .ZN(n8004) );
  AOI211_X1 U9776 ( .C1(n8006), .C2(n8467), .A(n8005), .B(n8004), .ZN(n8007)
         );
  OAI211_X1 U9777 ( .C1(n8010), .C2(n8009), .A(n8008), .B(n8007), .ZN(P2_U3181) );
  MUX2_X1 U9778 ( .A(n6728), .B(n10332), .S(n7856), .Z(n8015) );
  XNOR2_X1 U9779 ( .A(n8015), .B(SI_31_), .ZN(n8016) );
  NAND2_X1 U9780 ( .A1(n8889), .A2(n8048), .ZN(n8019) );
  NAND2_X1 U9781 ( .A1(n4499), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8018) );
  INV_X1 U9782 ( .A(n8020), .ZN(n8183) );
  INV_X1 U9783 ( .A(n8307), .ZN(n8315) );
  INV_X1 U9784 ( .A(n8021), .ZN(n8054) );
  NAND2_X1 U9785 ( .A1(n8175), .A2(n8169), .ZN(n8367) );
  INV_X1 U9786 ( .A(n8376), .ZN(n8167) );
  INV_X1 U9787 ( .A(n8463), .ZN(n8465) );
  NAND4_X1 U9788 ( .A1(n8025), .A2(n8024), .A3(n9990), .A4(n8023), .ZN(n8029)
         );
  NAND3_X1 U9789 ( .A1(n8073), .A2(n8027), .A3(n8026), .ZN(n8028) );
  NOR2_X1 U9790 ( .A1(n8029), .A2(n8028), .ZN(n8032) );
  NAND4_X1 U9791 ( .A1(n8032), .A2(n8031), .A3(n8101), .A4(n8030), .ZN(n8033)
         );
  NOR2_X1 U9792 ( .A1(n8034), .A2(n8033), .ZN(n8035) );
  NAND4_X1 U9793 ( .A1(n8121), .A2(n8037), .A3(n8036), .A4(n8035), .ZN(n8038)
         );
  OR4_X1 U9794 ( .A1(n8465), .A2(n8500), .A3(n4744), .A4(n8038), .ZN(n8039) );
  NOR2_X1 U9795 ( .A1(n8452), .A2(n8039), .ZN(n8040) );
  NAND4_X1 U9796 ( .A1(n8413), .A2(n6619), .A3(n6617), .A4(n8040), .ZN(n8041)
         );
  NOR2_X1 U9797 ( .A1(n8041), .A2(n8403), .ZN(n8042) );
  NAND3_X1 U9798 ( .A1(n8167), .A2(n8392), .A3(n8042), .ZN(n8043) );
  NOR2_X1 U9799 ( .A1(n8367), .A2(n8043), .ZN(n8044) );
  NAND3_X1 U9800 ( .A1(n8352), .A2(n8359), .A3(n8044), .ZN(n8045) );
  NOR2_X1 U9801 ( .A1(n8330), .A2(n8045), .ZN(n8046) );
  NAND3_X1 U9802 ( .A1(n8315), .A2(n8296), .A3(n8046), .ZN(n8047) );
  NOR2_X1 U9803 ( .A1(n8185), .A2(n8047), .ZN(n8052) );
  NAND2_X1 U9804 ( .A1(n8885), .A2(n8048), .ZN(n8050) );
  NAND2_X1 U9805 ( .A1(n6451), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8049) );
  INV_X1 U9806 ( .A(n8222), .ZN(n8051) );
  NAND2_X1 U9807 ( .A1(n8557), .A2(n8051), .ZN(n8195) );
  MUX2_X1 U9808 ( .A(n8320), .B(n8304), .S(n8182), .Z(n8190) );
  MUX2_X1 U9809 ( .A(n8054), .B(n8053), .S(n8199), .Z(n8055) );
  NOR2_X1 U9810 ( .A1(n8307), .A2(n8055), .ZN(n8187) );
  NAND2_X1 U9811 ( .A1(n8169), .A2(n8056), .ZN(n8057) );
  AND2_X1 U9812 ( .A1(n8165), .A2(n8058), .ZN(n8060) );
  MUX2_X1 U9813 ( .A(n8060), .B(n8059), .S(n8182), .Z(n8163) );
  INV_X1 U9814 ( .A(n8140), .ZN(n8143) );
  AND2_X1 U9815 ( .A1(n8063), .A2(n8062), .ZN(n8066) );
  NAND3_X1 U9816 ( .A1(n9990), .A2(n8064), .A3(n8066), .ZN(n8065) );
  INV_X1 U9817 ( .A(n8066), .ZN(n8068) );
  NAND2_X1 U9818 ( .A1(n8068), .A2(n8067), .ZN(n8071) );
  OAI211_X1 U9819 ( .C1(n8071), .C2(n8070), .A(n8069), .B(n8074), .ZN(n8072)
         );
  INV_X1 U9820 ( .A(n8074), .ZN(n8077) );
  OAI211_X1 U9821 ( .C1(n8093), .C2(n8077), .A(n8076), .B(n8075), .ZN(n8078)
         );
  NAND2_X1 U9822 ( .A1(n8078), .A2(n8094), .ZN(n8080) );
  NAND2_X1 U9823 ( .A1(n8080), .A2(n8079), .ZN(n8081) );
  NAND2_X1 U9824 ( .A1(n8081), .A2(n8100), .ZN(n8084) );
  INV_X1 U9825 ( .A(n8082), .ZN(n8083) );
  AOI21_X1 U9826 ( .B1(n8084), .B2(n8101), .A(n8083), .ZN(n8090) );
  NAND2_X1 U9827 ( .A1(n8110), .A2(n8104), .ZN(n8088) );
  NAND2_X1 U9828 ( .A1(n8086), .A2(n8085), .ZN(n8087) );
  MUX2_X1 U9829 ( .A(n8088), .B(n8087), .S(n8199), .Z(n8107) );
  OAI21_X1 U9830 ( .B1(n8090), .B2(n8107), .A(n8089), .ZN(n8092) );
  NAND4_X1 U9831 ( .A1(n8092), .A2(n8182), .A3(n8091), .A4(n8111), .ZN(n8122)
         );
  INV_X1 U9832 ( .A(n8093), .ZN(n8099) );
  OAI21_X1 U9833 ( .B1(n8096), .B2(n8095), .A(n8094), .ZN(n8097) );
  AOI21_X1 U9834 ( .B1(n8099), .B2(n8098), .A(n8097), .ZN(n8103) );
  OAI211_X1 U9835 ( .C1(n8103), .C2(n8102), .A(n8101), .B(n8100), .ZN(n8106)
         );
  NAND3_X1 U9836 ( .A1(n8106), .A2(n8105), .A3(n8104), .ZN(n8109) );
  INV_X1 U9837 ( .A(n8107), .ZN(n8108) );
  NAND2_X1 U9838 ( .A1(n8109), .A2(n8108), .ZN(n8112) );
  NAND3_X1 U9839 ( .A1(n8112), .A2(n8111), .A3(n8110), .ZN(n8115) );
  NAND4_X1 U9840 ( .A1(n8115), .A2(n8199), .A3(n8114), .A4(n8113), .ZN(n8120)
         );
  NOR2_X1 U9841 ( .A1(n8116), .A2(n8199), .ZN(n8118) );
  OAI21_X1 U9842 ( .B1(n8182), .B2(n8224), .A(n10054), .ZN(n8117) );
  OAI21_X1 U9843 ( .B1(n8118), .B2(n10054), .A(n8117), .ZN(n8119) );
  NAND4_X1 U9844 ( .A1(n8122), .A2(n8121), .A3(n8120), .A4(n8119), .ZN(n8126)
         );
  MUX2_X1 U9845 ( .A(n8124), .B(n8123), .S(n8199), .Z(n8125) );
  INV_X1 U9846 ( .A(n8129), .ZN(n9524) );
  MUX2_X1 U9847 ( .A(n8127), .B(n9524), .S(n8199), .Z(n8128) );
  MUX2_X1 U9848 ( .A(n8131), .B(n8130), .S(n8199), .Z(n8132) );
  NAND2_X1 U9849 ( .A1(n8133), .A2(n8132), .ZN(n8134) );
  NAND2_X1 U9850 ( .A1(n8134), .A2(n8463), .ZN(n8145) );
  NAND3_X1 U9851 ( .A1(n8145), .A2(n8146), .A3(n8135), .ZN(n8137) );
  NAND3_X1 U9852 ( .A1(n8137), .A2(n8199), .A3(n8136), .ZN(n8138) );
  NAND2_X1 U9853 ( .A1(n8140), .A2(n8139), .ZN(n8141) );
  NAND2_X1 U9854 ( .A1(n8141), .A2(n8199), .ZN(n8142) );
  NAND2_X1 U9855 ( .A1(n8145), .A2(n8144), .ZN(n8147) );
  NAND3_X1 U9856 ( .A1(n8147), .A2(n8182), .A3(n8146), .ZN(n8148) );
  NAND2_X1 U9857 ( .A1(n8149), .A2(n8148), .ZN(n8152) );
  NAND3_X1 U9858 ( .A1(n8152), .A2(n8151), .A3(n8150), .ZN(n8153) );
  NAND2_X1 U9859 ( .A1(n8153), .A2(n8156), .ZN(n8160) );
  INV_X1 U9860 ( .A(n8154), .ZN(n8155) );
  NOR2_X1 U9861 ( .A1(n8403), .A2(n8155), .ZN(n8158) );
  AND2_X1 U9862 ( .A1(n8387), .A2(n8156), .ZN(n8157) );
  MUX2_X1 U9863 ( .A(n8158), .B(n8157), .S(n8199), .Z(n8159) );
  OAI21_X1 U9864 ( .B1(n8161), .B2(n8160), .A(n8159), .ZN(n8162) );
  MUX2_X1 U9865 ( .A(n8165), .B(n8164), .S(n8199), .Z(n8166) );
  NAND3_X1 U9866 ( .A1(n8170), .A2(n8199), .A3(n8176), .ZN(n8171) );
  NAND2_X1 U9867 ( .A1(n8171), .A2(n8352), .ZN(n8174) );
  OR3_X1 U9868 ( .A1(n8172), .A2(n8332), .A3(n8182), .ZN(n8173) );
  NAND2_X1 U9869 ( .A1(n8174), .A2(n8173), .ZN(n8181) );
  NAND3_X1 U9870 ( .A1(n8177), .A2(n8176), .A3(n8175), .ZN(n8178) );
  NAND3_X1 U9871 ( .A1(n8178), .A2(n5015), .A3(n8182), .ZN(n8180) );
  MUX2_X1 U9872 ( .A(n8184), .B(n8183), .S(n8182), .Z(n8186) );
  AOI21_X1 U9873 ( .B1(n8188), .B2(n8190), .A(n8189), .ZN(n8197) );
  INV_X1 U9874 ( .A(n8190), .ZN(n8191) );
  NAND2_X1 U9875 ( .A1(n8195), .A2(n8193), .ZN(n8205) );
  NOR2_X1 U9876 ( .A1(n8198), .A2(n8205), .ZN(n8194) );
  OAI211_X1 U9877 ( .C1(n8197), .C2(n8320), .A(n8194), .B(n8207), .ZN(n8202)
         );
  INV_X1 U9878 ( .A(n8212), .ZN(n8196) );
  OAI211_X1 U9879 ( .C1(n8196), .C2(n8199), .A(n8207), .B(n8195), .ZN(n8201)
         );
  INV_X1 U9880 ( .A(n8198), .ZN(n8200) );
  INV_X1 U9881 ( .A(n8557), .ZN(n8508) );
  AOI21_X1 U9882 ( .B1(n4496), .B2(n8206), .A(n8205), .ZN(n8208) );
  OAI211_X1 U9883 ( .C1(n8508), .C2(n8284), .A(n8208), .B(n8207), .ZN(n8211)
         );
  INV_X1 U9884 ( .A(n8209), .ZN(n8210) );
  XNOR2_X1 U9885 ( .A(n8213), .B(n8279), .ZN(n8221) );
  INV_X1 U9886 ( .A(n8214), .ZN(n8220) );
  NAND3_X1 U9887 ( .A1(n8216), .A2(n8215), .A3(n8273), .ZN(n8217) );
  OAI211_X1 U9888 ( .C1(n8218), .C2(n8220), .A(n8217), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8219) );
  OAI21_X1 U9889 ( .B1(n8221), .B2(n8220), .A(n8219), .ZN(P2_U3296) );
  MUX2_X1 U9890 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8222), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9891 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8298), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9892 ( .A(n8320), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8233), .Z(
        P2_U3519) );
  MUX2_X1 U9893 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8297), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9894 ( .A(n8319), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8233), .Z(
        P2_U3517) );
  MUX2_X1 U9895 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8360), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9896 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8369), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9897 ( .A(n8380), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8233), .Z(
        P2_U3514) );
  MUX2_X1 U9898 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8395), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9899 ( .A(n8406), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8233), .Z(
        P2_U3512) );
  MUX2_X1 U9900 ( .A(n8415), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8233), .Z(
        P2_U3511) );
  MUX2_X1 U9901 ( .A(n8405), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8233), .Z(
        P2_U3510) );
  MUX2_X1 U9902 ( .A(n8437), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8233), .Z(
        P2_U3509) );
  MUX2_X1 U9903 ( .A(n8454), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8233), .Z(
        P2_U3508) );
  MUX2_X1 U9904 ( .A(n8468), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8233), .Z(
        P2_U3507) );
  MUX2_X1 U9905 ( .A(n8480), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8233), .Z(
        P2_U3506) );
  MUX2_X1 U9906 ( .A(n8467), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8233), .Z(
        P2_U3505) );
  MUX2_X1 U9907 ( .A(n8482), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8233), .Z(
        P2_U3504) );
  MUX2_X1 U9908 ( .A(n8223), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8233), .Z(
        P2_U3503) );
  MUX2_X1 U9909 ( .A(n8224), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8233), .Z(
        P2_U3502) );
  MUX2_X1 U9910 ( .A(n8225), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8233), .Z(
        P2_U3501) );
  MUX2_X1 U9911 ( .A(n8226), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8233), .Z(
        P2_U3500) );
  MUX2_X1 U9912 ( .A(n8227), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8233), .Z(
        P2_U3499) );
  MUX2_X1 U9913 ( .A(n8228), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8233), .Z(
        P2_U3498) );
  MUX2_X1 U9914 ( .A(n8229), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8233), .Z(
        P2_U3497) );
  MUX2_X1 U9915 ( .A(n8230), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8233), .Z(
        P2_U3496) );
  MUX2_X1 U9916 ( .A(n8231), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8233), .Z(
        P2_U3495) );
  MUX2_X1 U9917 ( .A(n4841), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8233), .Z(
        P2_U3494) );
  MUX2_X1 U9918 ( .A(n8232), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8233), .Z(
        P2_U3493) );
  MUX2_X1 U9919 ( .A(n8234), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8233), .Z(
        P2_U3492) );
  NOR2_X1 U9920 ( .A1(n9899), .A2(n8237), .ZN(n8238) );
  XNOR2_X1 U9921 ( .A(n9914), .B(n8490), .ZN(n9924) );
  NOR2_X1 U9922 ( .A1(n9925), .A2(n9924), .ZN(n9923) );
  XNOR2_X1 U9923 ( .A(n9947), .B(n8457), .ZN(n9957) );
  NOR2_X1 U9924 ( .A1(n9958), .A2(n9957), .ZN(n9956) );
  AOI21_X1 U9925 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8253), .A(n9956), .ZN(
        n8240) );
  NOR2_X1 U9926 ( .A1(n9468), .A2(n8267), .ZN(n8241) );
  AOI21_X1 U9927 ( .B1(n8267), .B2(n9468), .A(n8241), .ZN(n9475) );
  MUX2_X1 U9928 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8417), .S(n8251), .Z(n8275)
         );
  XNOR2_X1 U9929 ( .A(n8242), .B(n8275), .ZN(n8283) );
  AOI22_X1 U9930 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8253), .B1(n9947), .B2(
        n8542), .ZN(n9950) );
  AOI22_X1 U9931 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8257), .B1(n9914), .B2(
        n8548), .ZN(n9917) );
  OAI21_X1 U9932 ( .B1(n8244), .B2(n7614), .A(n8243), .ZN(n8245) );
  NAND2_X1 U9933 ( .A1(n4923), .A2(n8245), .ZN(n8246) );
  XNOR2_X1 U9934 ( .A(n9899), .B(n8245), .ZN(n9901) );
  NAND2_X1 U9935 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9901), .ZN(n9900) );
  NAND2_X1 U9936 ( .A1(n8246), .A2(n9900), .ZN(n9916) );
  NAND2_X1 U9937 ( .A1(n9917), .A2(n9916), .ZN(n9915) );
  OAI21_X1 U9938 ( .B1(n9914), .B2(n8548), .A(n9915), .ZN(n8247) );
  NAND2_X1 U9939 ( .A1(n8255), .A2(n8247), .ZN(n8248) );
  XOR2_X1 U9940 ( .A(n8247), .B(n8255), .Z(n9933) );
  NAND2_X1 U9941 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9933), .ZN(n9932) );
  NAND2_X1 U9942 ( .A1(n8248), .A2(n9932), .ZN(n9949) );
  NAND2_X1 U9943 ( .A1(n9950), .A2(n9949), .ZN(n9948) );
  OAI21_X1 U9944 ( .B1(n9947), .B2(n8542), .A(n9948), .ZN(n8249) );
  NAND2_X1 U9945 ( .A1(n8265), .A2(n8249), .ZN(n8250) );
  XNOR2_X1 U9946 ( .A(n9965), .B(n8249), .ZN(n9968) );
  NAND2_X1 U9947 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n9968), .ZN(n9967) );
  NAND2_X1 U9948 ( .A1(n8250), .A2(n9967), .ZN(n9462) );
  XNOR2_X1 U9949 ( .A(n9467), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n9461) );
  AOI22_X1 U9950 ( .A1(n9462), .A2(n9461), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n9468), .ZN(n8252) );
  XNOR2_X1 U9951 ( .A(n8251), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8272) );
  XNOR2_X1 U9952 ( .A(n8252), .B(n8272), .ZN(n8281) );
  MUX2_X1 U9953 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8273), .Z(n8266) );
  XNOR2_X1 U9954 ( .A(n8266), .B(n9965), .ZN(n9971) );
  MUX2_X1 U9955 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8273), .Z(n8254) );
  OR2_X1 U9956 ( .A1(n8254), .A2(n8253), .ZN(n8264) );
  XNOR2_X1 U9957 ( .A(n8254), .B(n9947), .ZN(n9953) );
  MUX2_X1 U9958 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8273), .Z(n8256) );
  OR2_X1 U9959 ( .A1(n8256), .A2(n8255), .ZN(n8263) );
  XNOR2_X1 U9960 ( .A(n9931), .B(n8256), .ZN(n9936) );
  MUX2_X1 U9961 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8273), .Z(n8258) );
  OR2_X1 U9962 ( .A1(n8258), .A2(n8257), .ZN(n8262) );
  XNOR2_X1 U9963 ( .A(n8258), .B(n9914), .ZN(n9920) );
  MUX2_X1 U9964 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8273), .Z(n8261) );
  XNOR2_X1 U9965 ( .A(n8261), .B(n9899), .ZN(n9904) );
  NAND2_X1 U9966 ( .A1(n9920), .A2(n9919), .ZN(n9918) );
  NAND2_X1 U9967 ( .A1(n8262), .A2(n9918), .ZN(n9935) );
  NAND2_X1 U9968 ( .A1(n9936), .A2(n9935), .ZN(n9934) );
  NAND2_X1 U9969 ( .A1(n8263), .A2(n9934), .ZN(n9952) );
  NAND2_X1 U9970 ( .A1(n9953), .A2(n9952), .ZN(n9951) );
  NAND2_X1 U9971 ( .A1(n8264), .A2(n9951), .ZN(n9970) );
  NAND2_X1 U9972 ( .A1(n9971), .A2(n9970), .ZN(n9969) );
  OAI21_X1 U9973 ( .B1(n8266), .B2(n8265), .A(n9969), .ZN(n8268) );
  MUX2_X1 U9974 ( .A(n8267), .B(n8535), .S(n8273), .Z(n8269) );
  NAND2_X1 U9975 ( .A1(n8268), .A2(n8269), .ZN(n9465) );
  NAND2_X1 U9976 ( .A1(n9465), .A2(n9468), .ZN(n9471) );
  INV_X1 U9977 ( .A(n8268), .ZN(n8271) );
  INV_X1 U9978 ( .A(n8269), .ZN(n8270) );
  NAND2_X1 U9979 ( .A1(n8271), .A2(n8270), .ZN(n9464) );
  NAND2_X1 U9980 ( .A1(n9471), .A2(n9464), .ZN(n8277) );
  INV_X1 U9981 ( .A(n8272), .ZN(n8274) );
  MUX2_X1 U9982 ( .A(n8275), .B(n8274), .S(n8273), .Z(n8276) );
  NAND2_X1 U9983 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n8278) );
  AOI21_X1 U9984 ( .B1(n8281), .B2(n9974), .A(n8280), .ZN(n8282) );
  OAI21_X1 U9985 ( .B1(n8283), .B2(n9980), .A(n8282), .ZN(P2_U3201) );
  NAND2_X1 U9986 ( .A1(n8284), .A2(n8473), .ZN(n8289) );
  INV_X1 U9987 ( .A(n8285), .ZN(n8286) );
  NOR2_X1 U9988 ( .A1(n8287), .A2(n8286), .ZN(n8554) );
  OAI21_X1 U9989 ( .B1(n8554), .B2(n8288), .A(n4500), .ZN(n8291) );
  OAI211_X1 U9990 ( .C1(n4500), .C2(n8290), .A(n8289), .B(n8291), .ZN(P2_U3202) );
  NAND2_X1 U9991 ( .A1(n8557), .A2(n8473), .ZN(n8292) );
  OAI211_X1 U9992 ( .C1(n4500), .C2(n8293), .A(n8292), .B(n8291), .ZN(P2_U3203) );
  XNOR2_X1 U9993 ( .A(n4497), .B(n8296), .ZN(n8562) );
  XOR2_X1 U9994 ( .A(n8296), .B(n8295), .Z(n8300) );
  AOI22_X1 U9995 ( .A1(n8298), .A2(n8479), .B1(n8481), .B2(n8297), .ZN(n8299)
         );
  INV_X1 U9996 ( .A(n8560), .ZN(n8301) );
  MUX2_X1 U9997 ( .A(n8302), .B(n8301), .S(n4500), .Z(n8306) );
  AOI22_X1 U9998 ( .A1(n8304), .A2(n8473), .B1(n8472), .B2(n8303), .ZN(n8305)
         );
  OAI211_X1 U9999 ( .C1(n8562), .C2(n8476), .A(n8306), .B(n8305), .ZN(P2_U3205) );
  XNOR2_X1 U10000 ( .A(n8308), .B(n8307), .ZN(n8567) );
  OR2_X1 U10001 ( .A1(n8345), .A2(n8309), .ZN(n8311) );
  NAND2_X1 U10002 ( .A1(n8311), .A2(n8310), .ZN(n8318) );
  OR2_X2 U10003 ( .A1(n8345), .A2(n8352), .ZN(n8343) );
  NAND2_X1 U10004 ( .A1(n8343), .A2(n8312), .ZN(n8314) );
  AOI21_X1 U10005 ( .B1(n8316), .B2(n8315), .A(n10000), .ZN(n8317) );
  OAI21_X1 U10006 ( .B1(n8318), .B2(n5086), .A(n8317), .ZN(n8322) );
  AOI22_X1 U10007 ( .A1(n8320), .A2(n8479), .B1(n8481), .B2(n8319), .ZN(n8321)
         );
  NAND2_X1 U10008 ( .A1(n8322), .A2(n8321), .ZN(n8565) );
  INV_X1 U10009 ( .A(n8565), .ZN(n8323) );
  MUX2_X1 U10010 ( .A(n8324), .B(n8323), .S(n4500), .Z(n8327) );
  AOI22_X1 U10011 ( .A1(n8511), .A2(n8473), .B1(n8472), .B2(n8325), .ZN(n8326)
         );
  OAI211_X1 U10012 ( .C1(n8567), .C2(n8476), .A(n8327), .B(n8326), .ZN(
        P2_U3206) );
  XOR2_X1 U10013 ( .A(n8330), .B(n8328), .Z(n8572) );
  NAND2_X1 U10014 ( .A1(n8343), .A2(n8329), .ZN(n8331) );
  INV_X1 U10015 ( .A(n8570), .ZN(n8337) );
  MUX2_X1 U10016 ( .A(n8338), .B(n8337), .S(n4500), .Z(n8342) );
  AOI22_X1 U10017 ( .A1(n8340), .A2(n8473), .B1(n8472), .B2(n8339), .ZN(n8341)
         );
  OAI211_X1 U10018 ( .C1(n8572), .C2(n8476), .A(n8342), .B(n8341), .ZN(
        P2_U3207) );
  INV_X1 U10019 ( .A(n8343), .ZN(n8344) );
  AOI21_X1 U10020 ( .B1(n8352), .B2(n8345), .A(n8344), .ZN(n8346) );
  OAI222_X1 U10021 ( .A1(n9993), .A2(n8348), .B1(n9995), .B2(n8347), .C1(
        n10000), .C2(n8346), .ZN(n8575) );
  INV_X1 U10022 ( .A(n8349), .ZN(n8350) );
  OAI22_X1 U10023 ( .A1(n8576), .A2(n9987), .B1(n8350), .B2(n9989), .ZN(n8351)
         );
  OAI21_X1 U10024 ( .B1(n8575), .B2(n8351), .A(n4500), .ZN(n8355) );
  XNOR2_X1 U10025 ( .A(n8353), .B(n8352), .ZN(n8577) );
  OR2_X1 U10026 ( .A1(n8577), .A2(n8476), .ZN(n8354) );
  OAI211_X1 U10027 ( .C1(n4500), .C2(n8356), .A(n8355), .B(n8354), .ZN(
        P2_U3208) );
  XNOR2_X1 U10028 ( .A(n8357), .B(n8359), .ZN(n8582) );
  INV_X1 U10029 ( .A(n8582), .ZN(n8366) );
  XOR2_X1 U10030 ( .A(n8359), .B(n8358), .Z(n8361) );
  AOI222_X1 U10031 ( .A1(n8484), .A2(n8361), .B1(n8360), .B2(n8479), .C1(n8380), .C2(n8481), .ZN(n8580) );
  OAI21_X1 U10032 ( .B1(n8585), .B2(n9987), .A(n8580), .ZN(n8362) );
  NAND2_X1 U10033 ( .A1(n8362), .A2(n4500), .ZN(n8365) );
  AOI22_X1 U10034 ( .A1(n10005), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8472), 
        .B2(n8363), .ZN(n8364) );
  OAI211_X1 U10035 ( .C1(n8366), .C2(n8476), .A(n8365), .B(n8364), .ZN(
        P2_U3209) );
  XNOR2_X1 U10036 ( .A(n4571), .B(n8367), .ZN(n8591) );
  INV_X1 U10037 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8371) );
  XNOR2_X1 U10038 ( .A(n8368), .B(n8367), .ZN(n8370) );
  AOI222_X1 U10039 ( .A1(n8484), .A2(n8370), .B1(n8369), .B2(n8479), .C1(n8395), .C2(n8481), .ZN(n8586) );
  MUX2_X1 U10040 ( .A(n8371), .B(n8586), .S(n4500), .Z(n8374) );
  AOI22_X1 U10041 ( .A1(n8588), .A2(n8473), .B1(n8472), .B2(n8372), .ZN(n8373)
         );
  OAI211_X1 U10042 ( .C1(n8591), .C2(n8476), .A(n8374), .B(n8373), .ZN(
        P2_U3210) );
  XNOR2_X1 U10043 ( .A(n8375), .B(n8376), .ZN(n8595) );
  INV_X1 U10044 ( .A(n8595), .ZN(n8386) );
  OR3_X1 U10045 ( .A1(n8390), .A2(n8377), .A3(n8376), .ZN(n8378) );
  NAND2_X1 U10046 ( .A1(n8379), .A2(n8378), .ZN(n8381) );
  AOI222_X1 U10047 ( .A1(n8484), .A2(n8381), .B1(n8380), .B2(n8479), .C1(n8406), .C2(n8481), .ZN(n8592) );
  MUX2_X1 U10048 ( .A(n8382), .B(n8592), .S(n4500), .Z(n8385) );
  AOI22_X1 U10049 ( .A1(n8594), .A2(n8473), .B1(n8472), .B2(n8383), .ZN(n8384)
         );
  OAI211_X1 U10050 ( .C1(n8386), .C2(n8476), .A(n8385), .B(n8384), .ZN(
        P2_U3211) );
  NAND2_X1 U10051 ( .A1(n8388), .A2(n8387), .ZN(n8389) );
  XOR2_X1 U10052 ( .A(n8392), .B(n8389), .Z(n8603) );
  INV_X1 U10053 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8397) );
  INV_X1 U10054 ( .A(n8390), .ZN(n8394) );
  NAND3_X1 U10055 ( .A1(n8402), .A2(n8392), .A3(n8391), .ZN(n8393) );
  NAND2_X1 U10056 ( .A1(n8394), .A2(n8393), .ZN(n8396) );
  AOI222_X1 U10057 ( .A1(n8484), .A2(n8396), .B1(n8395), .B2(n8479), .C1(n8415), .C2(n8481), .ZN(n8598) );
  MUX2_X1 U10058 ( .A(n8397), .B(n8598), .S(n4500), .Z(n8400) );
  AOI22_X1 U10059 ( .A1(n8600), .A2(n8473), .B1(n8472), .B2(n8398), .ZN(n8399)
         );
  OAI211_X1 U10060 ( .C1(n8603), .C2(n8476), .A(n8400), .B(n8399), .ZN(
        P2_U3212) );
  XOR2_X1 U10061 ( .A(n8401), .B(n8403), .Z(n8609) );
  OAI21_X1 U10062 ( .B1(n8404), .B2(n8403), .A(n8402), .ZN(n8407) );
  AOI222_X1 U10063 ( .A1(n8484), .A2(n8407), .B1(n8406), .B2(n8479), .C1(n8405), .C2(n8481), .ZN(n8604) );
  MUX2_X1 U10064 ( .A(n8408), .B(n8604), .S(n4500), .Z(n8411) );
  AOI22_X1 U10065 ( .A1(n8606), .A2(n8473), .B1(n8472), .B2(n8409), .ZN(n8410)
         );
  OAI211_X1 U10066 ( .C1(n8609), .C2(n8476), .A(n8411), .B(n8410), .ZN(
        P2_U3213) );
  XNOR2_X1 U10067 ( .A(n8412), .B(n8413), .ZN(n8616) );
  XNOR2_X1 U10068 ( .A(n8414), .B(n8413), .ZN(n8416) );
  AOI222_X1 U10069 ( .A1(n8484), .A2(n8416), .B1(n8415), .B2(n8479), .C1(n8437), .C2(n8481), .ZN(n8610) );
  MUX2_X1 U10070 ( .A(n8417), .B(n8610), .S(n4500), .Z(n8420) );
  AOI22_X1 U10071 ( .A1(n8612), .A2(n8473), .B1(n8472), .B2(n8418), .ZN(n8419)
         );
  OAI211_X1 U10072 ( .C1(n8616), .C2(n8476), .A(n8420), .B(n8419), .ZN(
        P2_U3214) );
  XNOR2_X1 U10073 ( .A(n8421), .B(n8428), .ZN(n8422) );
  OAI222_X1 U10074 ( .A1(n9993), .A2(n8424), .B1(n9995), .B2(n8423), .C1(n8422), .C2(n10000), .ZN(n8533) );
  INV_X1 U10075 ( .A(n8533), .ZN(n8433) );
  INV_X1 U10076 ( .A(n8425), .ZN(n8426) );
  AOI21_X1 U10077 ( .B1(n8428), .B2(n8427), .A(n8426), .ZN(n8534) );
  AOI22_X1 U10078 ( .A1(n10005), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8472), 
        .B2(n8429), .ZN(n8430) );
  OAI21_X1 U10079 ( .B1(n8621), .B2(n8442), .A(n8430), .ZN(n8431) );
  AOI21_X1 U10080 ( .B1(n8534), .B2(n8502), .A(n8431), .ZN(n8432) );
  OAI21_X1 U10081 ( .B1(n8433), .B2(n10005), .A(n8432), .ZN(P2_U3215) );
  OAI211_X1 U10082 ( .C1(n8436), .C2(n8435), .A(n8434), .B(n8484), .ZN(n8439)
         );
  AOI22_X1 U10083 ( .A1(n8481), .A2(n8468), .B1(n8437), .B2(n8479), .ZN(n8438)
         );
  OAI21_X1 U10084 ( .B1(n6617), .B2(n8441), .A(n8440), .ZN(n8539) );
  NOR2_X1 U10085 ( .A1(n8443), .A2(n8442), .ZN(n8446) );
  OAI22_X1 U10086 ( .A1(n4500), .A2(n9977), .B1(n8444), .B2(n9989), .ZN(n8445)
         );
  AOI211_X1 U10087 ( .C1(n8539), .C2(n8502), .A(n8446), .B(n8445), .ZN(n8447)
         );
  OAI21_X1 U10088 ( .B1(n8541), .B2(n10005), .A(n8447), .ZN(P2_U3216) );
  NAND2_X1 U10089 ( .A1(n8449), .A2(n8448), .ZN(n8450) );
  XOR2_X1 U10090 ( .A(n8452), .B(n8450), .Z(n8626) );
  INV_X1 U10091 ( .A(n8626), .ZN(n8462) );
  OAI211_X1 U10092 ( .C1(n8453), .C2(n8452), .A(n8451), .B(n8484), .ZN(n8456)
         );
  AOI22_X1 U10093 ( .A1(n8481), .A2(n8480), .B1(n8454), .B2(n8479), .ZN(n8455)
         );
  MUX2_X1 U10094 ( .A(n8457), .B(n8623), .S(n4500), .Z(n8461) );
  INV_X1 U10095 ( .A(n8458), .ZN(n8459) );
  AOI22_X1 U10096 ( .A1(n8625), .A2(n8473), .B1(n8472), .B2(n8459), .ZN(n8460)
         );
  OAI211_X1 U10097 ( .C1(n8462), .C2(n8476), .A(n8461), .B(n8460), .ZN(
        P2_U3217) );
  XNOR2_X1 U10098 ( .A(n8464), .B(n8463), .ZN(n8632) );
  INV_X1 U10099 ( .A(n8632), .ZN(n8477) );
  XNOR2_X1 U10100 ( .A(n8466), .B(n8465), .ZN(n8469) );
  AOI222_X1 U10101 ( .A1(n8484), .A2(n8469), .B1(n8468), .B2(n8479), .C1(n8467), .C2(n8481), .ZN(n8629) );
  MUX2_X1 U10102 ( .A(n9940), .B(n8629), .S(n4500), .Z(n8475) );
  INV_X1 U10103 ( .A(n8470), .ZN(n8471) );
  AOI22_X1 U10104 ( .A1(n8631), .A2(n8473), .B1(n8472), .B2(n8471), .ZN(n8474)
         );
  OAI211_X1 U10105 ( .C1(n8477), .C2(n8476), .A(n8475), .B(n8474), .ZN(
        P2_U3218) );
  INV_X1 U10106 ( .A(n9987), .ZN(n8486) );
  XNOR2_X1 U10107 ( .A(n8478), .B(n8487), .ZN(n8483) );
  AOI222_X1 U10108 ( .A1(n8484), .A2(n8483), .B1(n8482), .B2(n8481), .C1(n8480), .C2(n8479), .ZN(n8635) );
  INV_X1 U10109 ( .A(n8635), .ZN(n8485) );
  AOI21_X1 U10110 ( .B1(n8486), .B2(n8637), .A(n8485), .ZN(n8493) );
  XNOR2_X1 U10111 ( .A(n8488), .B(n8487), .ZN(n8640) );
  OAI22_X1 U10112 ( .A1(n4500), .A2(n8490), .B1(n8489), .B2(n9989), .ZN(n8491)
         );
  AOI21_X1 U10113 ( .B1(n8640), .B2(n8502), .A(n8491), .ZN(n8492) );
  OAI21_X1 U10114 ( .B1(n8493), .B2(n10005), .A(n8492), .ZN(P2_U3219) );
  XOR2_X1 U10115 ( .A(n8500), .B(n8494), .Z(n8495) );
  OAI222_X1 U10116 ( .A1(n9993), .A2(n8497), .B1(n9995), .B2(n8496), .C1(n8495), .C2(n10000), .ZN(n9525) );
  OAI22_X1 U10117 ( .A1(n9524), .A2(n9987), .B1(n8498), .B2(n9989), .ZN(n8499)
         );
  OAI21_X1 U10118 ( .B1(n9525), .B2(n8499), .A(n4500), .ZN(n8504) );
  XNOR2_X1 U10119 ( .A(n8501), .B(n8500), .ZN(n9527) );
  NAND2_X1 U10120 ( .A1(n9527), .A2(n8502), .ZN(n8503) );
  OAI211_X1 U10121 ( .C1(n6266), .C2(n4500), .A(n8504), .B(n8503), .ZN(
        P2_U3220) );
  NAND2_X1 U10122 ( .A1(n8554), .A2(n10081), .ZN(n8506) );
  NAND2_X1 U10123 ( .A1(n10079), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8505) );
  OAI211_X1 U10124 ( .C1(n8556), .C2(n8537), .A(n8506), .B(n8505), .ZN(
        P2_U3490) );
  NAND2_X1 U10125 ( .A1(n10079), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8507) );
  OAI211_X1 U10126 ( .C1(n8508), .C2(n8537), .A(n8507), .B(n8506), .ZN(
        P2_U3489) );
  MUX2_X1 U10127 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8560), .S(n10081), .Z(
        n8510) );
  NAND2_X1 U10128 ( .A1(n10081), .A2(n10030), .ZN(n8532) );
  OAI22_X1 U10129 ( .A1(n8562), .A2(n8532), .B1(n8561), .B2(n8537), .ZN(n8509)
         );
  OR2_X1 U10130 ( .A1(n8510), .A2(n8509), .ZN(P2_U3487) );
  MUX2_X1 U10131 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8565), .S(n10081), .Z(
        n8513) );
  INV_X1 U10132 ( .A(n8511), .ZN(n8566) );
  OAI22_X1 U10133 ( .A1(n8567), .A2(n8532), .B1(n8566), .B2(n8537), .ZN(n8512)
         );
  OR2_X1 U10134 ( .A1(n8513), .A2(n8512), .ZN(P2_U3486) );
  MUX2_X1 U10135 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8570), .S(n10081), .Z(
        n8515) );
  OAI22_X1 U10136 ( .A1(n8572), .A2(n8532), .B1(n8571), .B2(n8537), .ZN(n8514)
         );
  OR2_X1 U10137 ( .A1(n8515), .A2(n8514), .ZN(P2_U3485) );
  MUX2_X1 U10138 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8575), .S(n10081), .Z(
        n8517) );
  OAI22_X1 U10139 ( .A1(n8577), .A2(n8532), .B1(n8576), .B2(n8537), .ZN(n8516)
         );
  OR2_X1 U10140 ( .A1(n8517), .A2(n8516), .ZN(P2_U3484) );
  INV_X1 U10141 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8518) );
  MUX2_X1 U10142 ( .A(n8518), .B(n8580), .S(n10081), .Z(n8520) );
  INV_X1 U10143 ( .A(n8532), .ZN(n8550) );
  NAND2_X1 U10144 ( .A1(n8582), .A2(n8550), .ZN(n8519) );
  OAI211_X1 U10145 ( .C1(n8585), .C2(n8537), .A(n8520), .B(n8519), .ZN(
        P2_U3483) );
  MUX2_X1 U10146 ( .A(n10211), .B(n8586), .S(n10081), .Z(n8522) );
  NAND2_X1 U10147 ( .A1(n8588), .A2(n8549), .ZN(n8521) );
  OAI211_X1 U10148 ( .C1(n8591), .C2(n8532), .A(n8522), .B(n8521), .ZN(
        P2_U3482) );
  INV_X1 U10149 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8523) );
  MUX2_X1 U10150 ( .A(n8523), .B(n8592), .S(n10081), .Z(n8525) );
  AOI22_X1 U10151 ( .A1(n8595), .A2(n8550), .B1(n8549), .B2(n8594), .ZN(n8524)
         );
  NAND2_X1 U10152 ( .A1(n8525), .A2(n8524), .ZN(P2_U3481) );
  INV_X1 U10153 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10187) );
  MUX2_X1 U10154 ( .A(n10187), .B(n8598), .S(n10081), .Z(n8527) );
  NAND2_X1 U10155 ( .A1(n8600), .A2(n8549), .ZN(n8526) );
  OAI211_X1 U10156 ( .C1(n8532), .C2(n8603), .A(n8527), .B(n8526), .ZN(
        P2_U3480) );
  INV_X1 U10157 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10352) );
  MUX2_X1 U10158 ( .A(n10352), .B(n8604), .S(n10081), .Z(n8529) );
  NAND2_X1 U10159 ( .A1(n8606), .A2(n8549), .ZN(n8528) );
  OAI211_X1 U10160 ( .C1(n8609), .C2(n8532), .A(n8529), .B(n8528), .ZN(
        P2_U3479) );
  MUX2_X1 U10161 ( .A(n10295), .B(n8610), .S(n10081), .Z(n8531) );
  NAND2_X1 U10162 ( .A1(n8612), .A2(n8549), .ZN(n8530) );
  OAI211_X1 U10163 ( .C1(n8616), .C2(n8532), .A(n8531), .B(n8530), .ZN(
        P2_U3478) );
  AOI21_X1 U10164 ( .B1(n8534), .B2(n10030), .A(n8533), .ZN(n8617) );
  MUX2_X1 U10165 ( .A(n8535), .B(n8617), .S(n10081), .Z(n8536) );
  OAI21_X1 U10166 ( .B1(n8621), .B2(n8537), .A(n8536), .ZN(P2_U3477) );
  AOI22_X1 U10167 ( .A1(n8539), .A2(n10030), .B1(n10055), .B2(n8538), .ZN(
        n8540) );
  NAND2_X1 U10168 ( .A1(n8541), .A2(n8540), .ZN(n8622) );
  MUX2_X1 U10169 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8622), .S(n10081), .Z(
        P2_U3476) );
  MUX2_X1 U10170 ( .A(n8542), .B(n8623), .S(n10081), .Z(n8544) );
  AOI22_X1 U10171 ( .A1(n8626), .A2(n8550), .B1(n8549), .B2(n8625), .ZN(n8543)
         );
  NAND2_X1 U10172 ( .A1(n8544), .A2(n8543), .ZN(P2_U3475) );
  MUX2_X1 U10173 ( .A(n8545), .B(n8629), .S(n10081), .Z(n8547) );
  AOI22_X1 U10174 ( .A1(n8632), .A2(n8550), .B1(n8549), .B2(n8631), .ZN(n8546)
         );
  NAND2_X1 U10175 ( .A1(n8547), .A2(n8546), .ZN(P2_U3474) );
  MUX2_X1 U10176 ( .A(n8548), .B(n8635), .S(n10081), .Z(n8552) );
  AOI22_X1 U10177 ( .A1(n8640), .A2(n8550), .B1(n8549), .B2(n8637), .ZN(n8551)
         );
  NAND2_X1 U10178 ( .A1(n8552), .A2(n8551), .ZN(P2_U3473) );
  MUX2_X1 U10179 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8553), .S(n10081), .Z(
        P2_U3459) );
  NAND2_X1 U10180 ( .A1(n8554), .A2(n10063), .ZN(n8558) );
  NAND2_X1 U10181 ( .A1(n10065), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8555) );
  OAI211_X1 U10182 ( .C1(n8556), .C2(n8620), .A(n8558), .B(n8555), .ZN(
        P2_U3458) );
  NAND2_X1 U10183 ( .A1(n8557), .A2(n8638), .ZN(n8559) );
  OAI211_X1 U10184 ( .C1(n10063), .C2(n10335), .A(n8559), .B(n8558), .ZN(
        P2_U3457) );
  MUX2_X1 U10185 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8560), .S(n10063), .Z(
        n8564) );
  INV_X1 U10186 ( .A(n10030), .ZN(n10059) );
  OAI22_X1 U10187 ( .A1(n8562), .A2(n8615), .B1(n8561), .B2(n8620), .ZN(n8563)
         );
  OR2_X1 U10188 ( .A1(n8564), .A2(n8563), .ZN(P2_U3455) );
  MUX2_X1 U10189 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8565), .S(n10063), .Z(
        n8569) );
  OAI22_X1 U10190 ( .A1(n8567), .A2(n8615), .B1(n8566), .B2(n8620), .ZN(n8568)
         );
  OR2_X1 U10191 ( .A1(n8569), .A2(n8568), .ZN(P2_U3454) );
  MUX2_X1 U10192 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8570), .S(n10063), .Z(
        n8574) );
  OAI22_X1 U10193 ( .A1(n8572), .A2(n8615), .B1(n8571), .B2(n8620), .ZN(n8573)
         );
  OR2_X1 U10194 ( .A1(n8574), .A2(n8573), .ZN(P2_U3453) );
  MUX2_X1 U10195 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8575), .S(n10063), .Z(
        n8579) );
  OAI22_X1 U10196 ( .A1(n8577), .A2(n8615), .B1(n8576), .B2(n8620), .ZN(n8578)
         );
  OR2_X1 U10197 ( .A1(n8579), .A2(n8578), .ZN(P2_U3452) );
  INV_X1 U10198 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8581) );
  MUX2_X1 U10199 ( .A(n8581), .B(n8580), .S(n10063), .Z(n8584) );
  INV_X1 U10200 ( .A(n8615), .ZN(n8639) );
  NAND2_X1 U10201 ( .A1(n8582), .A2(n8639), .ZN(n8583) );
  OAI211_X1 U10202 ( .C1(n8585), .C2(n8620), .A(n8584), .B(n8583), .ZN(
        P2_U3451) );
  INV_X1 U10203 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8587) );
  MUX2_X1 U10204 ( .A(n8587), .B(n8586), .S(n10063), .Z(n8590) );
  NAND2_X1 U10205 ( .A1(n8588), .A2(n8638), .ZN(n8589) );
  OAI211_X1 U10206 ( .C1(n8591), .C2(n8615), .A(n8590), .B(n8589), .ZN(
        P2_U3450) );
  INV_X1 U10207 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8593) );
  MUX2_X1 U10208 ( .A(n8593), .B(n8592), .S(n10063), .Z(n8597) );
  AOI22_X1 U10209 ( .A1(n8595), .A2(n8639), .B1(n8638), .B2(n8594), .ZN(n8596)
         );
  NAND2_X1 U10210 ( .A1(n8597), .A2(n8596), .ZN(P2_U3449) );
  MUX2_X1 U10211 ( .A(n8599), .B(n8598), .S(n10063), .Z(n8602) );
  NAND2_X1 U10212 ( .A1(n8600), .A2(n8638), .ZN(n8601) );
  OAI211_X1 U10213 ( .C1(n8603), .C2(n8615), .A(n8602), .B(n8601), .ZN(
        P2_U3448) );
  INV_X1 U10214 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8605) );
  MUX2_X1 U10215 ( .A(n8605), .B(n8604), .S(n10063), .Z(n8608) );
  NAND2_X1 U10216 ( .A1(n8606), .A2(n8638), .ZN(n8607) );
  OAI211_X1 U10217 ( .C1(n8609), .C2(n8615), .A(n8608), .B(n8607), .ZN(
        P2_U3447) );
  INV_X1 U10218 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8611) );
  MUX2_X1 U10219 ( .A(n8611), .B(n8610), .S(n10063), .Z(n8614) );
  NAND2_X1 U10220 ( .A1(n8612), .A2(n8638), .ZN(n8613) );
  OAI211_X1 U10221 ( .C1(n8616), .C2(n8615), .A(n8614), .B(n8613), .ZN(
        P2_U3446) );
  MUX2_X1 U10222 ( .A(n8618), .B(n8617), .S(n10063), .Z(n8619) );
  OAI21_X1 U10223 ( .B1(n8621), .B2(n8620), .A(n8619), .ZN(P2_U3444) );
  MUX2_X1 U10224 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8622), .S(n10063), .Z(
        P2_U3441) );
  INV_X1 U10225 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8624) );
  MUX2_X1 U10226 ( .A(n8624), .B(n8623), .S(n10063), .Z(n8628) );
  AOI22_X1 U10227 ( .A1(n8626), .A2(n8639), .B1(n8638), .B2(n8625), .ZN(n8627)
         );
  NAND2_X1 U10228 ( .A1(n8628), .A2(n8627), .ZN(P2_U3438) );
  INV_X1 U10229 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8630) );
  MUX2_X1 U10230 ( .A(n8630), .B(n8629), .S(n10063), .Z(n8634) );
  AOI22_X1 U10231 ( .A1(n8632), .A2(n8639), .B1(n8638), .B2(n8631), .ZN(n8633)
         );
  NAND2_X1 U10232 ( .A1(n8634), .A2(n8633), .ZN(P2_U3435) );
  INV_X1 U10233 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8636) );
  MUX2_X1 U10234 ( .A(n8636), .B(n8635), .S(n10063), .Z(n8642) );
  AOI22_X1 U10235 ( .A1(n8640), .A2(n8639), .B1(n8638), .B2(n8637), .ZN(n8641)
         );
  NAND2_X1 U10236 ( .A1(n8642), .A2(n8641), .ZN(P2_U3432) );
  INV_X1 U10237 ( .A(n8889), .ZN(n9458) );
  NOR4_X1 U10238 ( .A1(n8643), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8644), .ZN(n8645) );
  AOI21_X1 U10239 ( .B1(n8647), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8645), .ZN(
        n8646) );
  OAI21_X1 U10240 ( .B1(n9458), .B2(n8650), .A(n8646), .ZN(P2_U3264) );
  AOI22_X1 U10241 ( .A1(n8648), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8647), .ZN(n8649) );
  OAI21_X1 U10242 ( .B1(n8651), .B2(n8650), .A(n8649), .ZN(P2_U3265) );
  INV_X1 U10243 ( .A(n8652), .ZN(n8653) );
  MUX2_X1 U10244 ( .A(n8653), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AND2_X1 U10245 ( .A1(n8655), .A2(n8654), .ZN(n8657) );
  OAI21_X1 U10246 ( .B1(n8658), .B2(n8657), .A(n8656), .ZN(n8659) );
  NAND2_X1 U10247 ( .A1(n8659), .A2(n8777), .ZN(n8664) );
  OAI22_X1 U10248 ( .A1(n9790), .A2(n8780), .B1(n8779), .B2(n9788), .ZN(n8660)
         );
  AOI211_X1 U10249 ( .C1(n6010), .C2(n8662), .A(n8661), .B(n8660), .ZN(n8663)
         );
  OAI211_X1 U10250 ( .C1(n8665), .C2(n8786), .A(n8664), .B(n8663), .ZN(
        P1_U3215) );
  NAND2_X1 U10251 ( .A1(n4585), .A2(n8666), .ZN(n8667) );
  XNOR2_X1 U10252 ( .A(n8668), .B(n8667), .ZN(n8674) );
  INV_X1 U10253 ( .A(n9229), .ZN(n8670) );
  INV_X1 U10254 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8669) );
  OAI22_X1 U10255 ( .A1(n8750), .A2(n8670), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8669), .ZN(n8672) );
  OAI22_X1 U10256 ( .A1(n9380), .A2(n8780), .B1(n8779), .B2(n9381), .ZN(n8671)
         );
  AOI211_X1 U10257 ( .C1(n9384), .C2(n8769), .A(n8672), .B(n8671), .ZN(n8673)
         );
  OAI21_X1 U10258 ( .B1(n8674), .B2(n8754), .A(n8673), .ZN(P1_U3216) );
  XNOR2_X1 U10259 ( .A(n8677), .B(n8675), .ZN(n8757) );
  NAND2_X1 U10260 ( .A1(n8757), .A2(n8758), .ZN(n8756) );
  NAND2_X1 U10261 ( .A1(n8677), .A2(n8676), .ZN(n8680) );
  AND2_X1 U10262 ( .A1(n8756), .A2(n8680), .ZN(n8682) );
  XNOR2_X1 U10263 ( .A(n8679), .B(n8678), .ZN(n8681) );
  NAND3_X1 U10264 ( .A1(n8756), .A2(n8681), .A3(n8680), .ZN(n8731) );
  OAI211_X1 U10265 ( .C1(n8682), .C2(n8681), .A(n8777), .B(n8731), .ZN(n8686)
         );
  OAI22_X1 U10266 ( .A1(n9288), .A2(n8780), .B1(n8779), .B2(n9330), .ZN(n8683)
         );
  AOI211_X1 U10267 ( .C1(n6010), .C2(n9292), .A(n8684), .B(n8683), .ZN(n8685)
         );
  OAI211_X1 U10268 ( .C1(n4657), .C2(n8786), .A(n8686), .B(n8685), .ZN(
        P1_U3219) );
  INV_X1 U10269 ( .A(n8687), .ZN(n8688) );
  AOI21_X1 U10270 ( .B1(n8690), .B2(n8689), .A(n8688), .ZN(n8695) );
  INV_X1 U10271 ( .A(n9258), .ZN(n8691) );
  INV_X1 U10272 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n10314) );
  OAI22_X1 U10273 ( .A1(n8750), .A2(n8691), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10314), .ZN(n8693) );
  OAI22_X1 U10274 ( .A1(n9381), .A2(n8780), .B1(n8779), .B2(n9288), .ZN(n8692)
         );
  AOI211_X1 U10275 ( .C1(n9262), .C2(n8769), .A(n8693), .B(n8692), .ZN(n8694)
         );
  OAI21_X1 U10276 ( .B1(n8695), .B2(n8754), .A(n8694), .ZN(P1_U3223) );
  AOI21_X1 U10277 ( .B1(n8697), .B2(n8696), .A(n4542), .ZN(n8702) );
  INV_X1 U10278 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10321) );
  OAI22_X1 U10279 ( .A1(n8750), .A2(n8698), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10321), .ZN(n8700) );
  OAI22_X1 U10280 ( .A1(n9367), .A2(n8780), .B1(n8779), .B2(n9380), .ZN(n8699)
         );
  AOI211_X1 U10281 ( .C1(n9370), .C2(n8769), .A(n8700), .B(n8699), .ZN(n8701)
         );
  OAI21_X1 U10282 ( .B1(n8702), .B2(n8754), .A(n8701), .ZN(P1_U3225) );
  OAI21_X1 U10283 ( .B1(n8705), .B2(n8704), .A(n8703), .ZN(n8706) );
  NAND2_X1 U10284 ( .A1(n8706), .A2(n8777), .ZN(n8711) );
  OAI22_X1 U10285 ( .A1(n9418), .A2(n8780), .B1(n8779), .B2(n9790), .ZN(n8707)
         );
  AOI211_X1 U10286 ( .C1(n6010), .C2(n8709), .A(n8708), .B(n8707), .ZN(n8710)
         );
  OAI211_X1 U10287 ( .C1(n8712), .C2(n8786), .A(n8711), .B(n8710), .ZN(
        P1_U3226) );
  OAI21_X1 U10288 ( .B1(n8715), .B2(n8714), .A(n8713), .ZN(n8716) );
  NAND2_X1 U10289 ( .A1(n8716), .A2(n8777), .ZN(n8721) );
  INV_X1 U10290 ( .A(n8717), .ZN(n9323) );
  OAI22_X1 U10291 ( .A1(n9330), .A2(n8780), .B1(n8779), .B2(n9329), .ZN(n8718)
         );
  AOI211_X1 U10292 ( .C1(n6010), .C2(n9323), .A(n8719), .B(n8718), .ZN(n8720)
         );
  OAI211_X1 U10293 ( .C1(n9325), .C2(n8786), .A(n8721), .B(n8720), .ZN(
        P1_U3228) );
  AOI21_X1 U10294 ( .B1(n8724), .B2(n8723), .A(n8722), .ZN(n8729) );
  INV_X1 U10295 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n10171) );
  OAI22_X1 U10296 ( .A1(n8750), .A2(n8725), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10171), .ZN(n8727) );
  OAI22_X1 U10297 ( .A1(n9358), .A2(n8780), .B1(n8779), .B2(n9216), .ZN(n8726)
         );
  AOI211_X1 U10298 ( .C1(n9375), .C2(n8769), .A(n8727), .B(n8726), .ZN(n8728)
         );
  OAI21_X1 U10299 ( .B1(n8729), .B2(n8754), .A(n8728), .ZN(P1_U3229) );
  NAND2_X1 U10300 ( .A1(n8731), .A2(n8730), .ZN(n8736) );
  INV_X1 U10301 ( .A(n8732), .ZN(n8734) );
  NOR2_X1 U10302 ( .A1(n8734), .A2(n8733), .ZN(n8735) );
  XNOR2_X1 U10303 ( .A(n8736), .B(n8735), .ZN(n8742) );
  INV_X1 U10304 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8737) );
  OAI22_X1 U10305 ( .A1(n8750), .A2(n8738), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8737), .ZN(n8740) );
  OAI22_X1 U10306 ( .A1(n9277), .A2(n8780), .B1(n8779), .B2(n9417), .ZN(n8739)
         );
  AOI211_X1 U10307 ( .C1(n9406), .C2(n8769), .A(n8740), .B(n8739), .ZN(n8741)
         );
  OAI21_X1 U10308 ( .B1(n8742), .B2(n8754), .A(n8741), .ZN(P1_U3233) );
  INV_X1 U10309 ( .A(n8743), .ZN(n8744) );
  NOR2_X1 U10310 ( .A1(n8745), .A2(n8744), .ZN(n8747) );
  XNOR2_X1 U10311 ( .A(n8747), .B(n8746), .ZN(n8755) );
  INV_X1 U10312 ( .A(n8748), .ZN(n9243) );
  INV_X1 U10313 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8749) );
  OAI22_X1 U10314 ( .A1(n8750), .A2(n9243), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8749), .ZN(n8752) );
  OAI22_X1 U10315 ( .A1(n9216), .A2(n8780), .B1(n8779), .B2(n9277), .ZN(n8751)
         );
  AOI211_X1 U10316 ( .C1(n9248), .C2(n8769), .A(n8752), .B(n8751), .ZN(n8753)
         );
  OAI21_X1 U10317 ( .B1(n8755), .B2(n8754), .A(n8753), .ZN(P1_U3235) );
  OAI21_X1 U10318 ( .B1(n8758), .B2(n8757), .A(n8756), .ZN(n8759) );
  NAND2_X1 U10319 ( .A1(n8759), .A2(n8777), .ZN(n8763) );
  INV_X1 U10320 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8760) );
  NOR2_X1 U10321 ( .A1(n8760), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9116) );
  OAI22_X1 U10322 ( .A1(n9417), .A2(n8780), .B1(n8779), .B2(n9418), .ZN(n8761)
         );
  AOI211_X1 U10323 ( .C1(n6010), .C2(n9305), .A(n9116), .B(n8761), .ZN(n8762)
         );
  OAI211_X1 U10324 ( .C1(n9312), .C2(n8786), .A(n8763), .B(n8762), .ZN(
        P1_U3238) );
  OAI21_X1 U10325 ( .B1(n4542), .B2(n8765), .A(n8764), .ZN(n8766) );
  NAND3_X1 U10326 ( .A1(n5069), .A2(n8777), .A3(n8766), .ZN(n8773) );
  AOI22_X1 U10327 ( .A1(n6010), .A2(n9184), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8772) );
  AOI22_X1 U10328 ( .A1(n8768), .A2(n9183), .B1(n8767), .B2(n9042), .ZN(n8771)
         );
  NAND2_X1 U10329 ( .A1(n9362), .A2(n8769), .ZN(n8770) );
  NAND4_X1 U10330 ( .A1(n8773), .A2(n8772), .A3(n8771), .A4(n8770), .ZN(
        P1_U3240) );
  OAI21_X1 U10331 ( .B1(n8776), .B2(n8775), .A(n8774), .ZN(n8778) );
  NAND2_X1 U10332 ( .A1(n8778), .A2(n8777), .ZN(n8785) );
  OAI22_X1 U10333 ( .A1(n9329), .A2(n8780), .B1(n8779), .B2(n9612), .ZN(n8781)
         );
  AOI211_X1 U10334 ( .C1(n6010), .C2(n8783), .A(n8782), .B(n8781), .ZN(n8784)
         );
  OAI211_X1 U10335 ( .C1(n9532), .C2(n8786), .A(n8785), .B(n8784), .ZN(
        P1_U3241) );
  NOR2_X1 U10336 ( .A1(n9183), .A2(n9031), .ZN(n8787) );
  NAND2_X1 U10337 ( .A1(n9352), .A2(n8787), .ZN(n8791) );
  OAI21_X1 U10338 ( .B1(n9031), .B2(n9171), .A(n8791), .ZN(n8788) );
  NAND2_X1 U10339 ( .A1(n8788), .A2(n9152), .ZN(n8790) );
  INV_X1 U10340 ( .A(n9031), .ZN(n8899) );
  OR3_X1 U10341 ( .A1(n9152), .A2(n9349), .A3(n8899), .ZN(n8789) );
  OAI211_X1 U10342 ( .C1(n9171), .C2(n8791), .A(n8790), .B(n8789), .ZN(n8792)
         );
  AND2_X1 U10343 ( .A1(n9163), .A2(n9031), .ZN(n8875) );
  NAND2_X1 U10344 ( .A1(n8936), .A2(n8793), .ZN(n8953) );
  NAND2_X1 U10345 ( .A1(n8866), .A2(n8794), .ZN(n8937) );
  MUX2_X1 U10346 ( .A(n8953), .B(n8937), .S(n8899), .Z(n8869) );
  AOI21_X1 U10347 ( .B1(n8863), .B2(n8844), .A(n9031), .ZN(n8842) );
  NAND2_X1 U10348 ( .A1(n8839), .A2(n8902), .ZN(n8838) );
  AND2_X1 U10349 ( .A1(n8843), .A2(n9298), .ZN(n9007) );
  INV_X1 U10350 ( .A(n6980), .ZN(n8795) );
  NAND2_X1 U10351 ( .A1(n8795), .A2(n8802), .ZN(n8796) );
  NAND2_X1 U10352 ( .A1(n8796), .A2(n8904), .ZN(n8798) );
  MUX2_X1 U10353 ( .A(n8798), .B(n8915), .S(n9031), .Z(n8805) );
  NAND2_X1 U10354 ( .A1(n8805), .A2(n8803), .ZN(n8801) );
  AND2_X1 U10355 ( .A1(n8799), .A2(n8913), .ZN(n8804) );
  AOI21_X1 U10356 ( .B1(n8801), .B2(n8804), .A(n8800), .ZN(n8807) );
  NAND2_X1 U10357 ( .A1(n8803), .A2(n8802), .ZN(n8909) );
  AND2_X1 U10358 ( .A1(n8809), .A2(n8808), .ZN(n8811) );
  MUX2_X1 U10359 ( .A(n8811), .B(n8810), .S(n9031), .Z(n8812) );
  NAND2_X1 U10360 ( .A1(n8813), .A2(n8812), .ZN(n8818) );
  AND2_X1 U10361 ( .A1(n8819), .A2(n8814), .ZN(n8816) );
  MUX2_X1 U10362 ( .A(n8816), .B(n8815), .S(n9031), .Z(n8817) );
  NAND2_X1 U10363 ( .A1(n8818), .A2(n8817), .ZN(n8825) );
  NAND2_X1 U10364 ( .A1(n8825), .A2(n8819), .ZN(n8821) );
  NAND2_X1 U10365 ( .A1(n8827), .A2(n8820), .ZN(n8924) );
  AOI21_X1 U10366 ( .B1(n8821), .B2(n8916), .A(n8924), .ZN(n8822) );
  NAND2_X1 U10367 ( .A1(n8831), .A2(n8826), .ZN(n8922) );
  OAI21_X1 U10368 ( .B1(n8822), .B2(n8922), .A(n9606), .ZN(n8834) );
  AOI21_X1 U10369 ( .B1(n8825), .B2(n8824), .A(n8823), .ZN(n8829) );
  NAND2_X1 U10370 ( .A1(n8826), .A2(n8916), .ZN(n8828) );
  OAI21_X1 U10371 ( .B1(n8829), .B2(n8828), .A(n8827), .ZN(n8832) );
  AOI21_X1 U10372 ( .B1(n8832), .B2(n8831), .A(n8830), .ZN(n8833) );
  MUX2_X1 U10373 ( .A(n8834), .B(n8833), .S(n8899), .Z(n8845) );
  NAND2_X1 U10374 ( .A1(n8850), .A2(n9609), .ZN(n8926) );
  AND2_X1 U10375 ( .A1(n8852), .A2(n8846), .ZN(n8835) );
  NAND2_X1 U10376 ( .A1(n8853), .A2(n8835), .ZN(n8930) );
  NAND2_X1 U10377 ( .A1(n8902), .A2(n8858), .ZN(n8836) );
  MUX2_X1 U10378 ( .A(n8838), .B(n8837), .S(n8899), .Z(n8841) );
  NAND2_X1 U10379 ( .A1(n8865), .A2(n8839), .ZN(n8948) );
  NAND2_X1 U10380 ( .A1(n8948), .A2(n8899), .ZN(n8840) );
  OAI21_X1 U10381 ( .B1(n8842), .B2(n8841), .A(n8840), .ZN(n8862) );
  OR2_X1 U10382 ( .A1(n9277), .A2(n9262), .ZN(n8954) );
  AND2_X1 U10383 ( .A1(n8844), .A2(n8843), .ZN(n8932) );
  NAND2_X1 U10384 ( .A1(n8845), .A2(n9609), .ZN(n8848) );
  NAND3_X1 U10385 ( .A1(n8848), .A2(n8847), .A3(n8846), .ZN(n8851) );
  NAND3_X1 U10386 ( .A1(n8851), .A2(n8850), .A3(n8849), .ZN(n8854) );
  NAND3_X1 U10387 ( .A1(n8854), .A2(n8853), .A3(n8852), .ZN(n8856) );
  NAND3_X1 U10388 ( .A1(n8856), .A2(n9317), .A3(n8855), .ZN(n8859) );
  AND2_X1 U10389 ( .A1(n8858), .A2(n8857), .ZN(n9006) );
  NAND2_X1 U10390 ( .A1(n8859), .A2(n9006), .ZN(n8860) );
  NAND3_X1 U10391 ( .A1(n8932), .A2(n8860), .A3(n9031), .ZN(n8861) );
  NAND2_X1 U10392 ( .A1(n8954), .A2(n8863), .ZN(n8935) );
  NAND2_X1 U10393 ( .A1(n8935), .A2(n9031), .ZN(n8864) );
  MUX2_X1 U10394 ( .A(n8866), .B(n8936), .S(n8899), .Z(n8867) );
  OR2_X1 U10395 ( .A1(n9191), .A2(n9031), .ZN(n8870) );
  NAND2_X1 U10396 ( .A1(n8871), .A2(n8870), .ZN(n8877) );
  NAND2_X1 U10397 ( .A1(n8949), .A2(n8939), .ZN(n8955) );
  OR2_X1 U10398 ( .A1(n9362), .A2(n9367), .ZN(n8873) );
  AND2_X1 U10399 ( .A1(n8873), .A2(n8872), .ZN(n8957) );
  OAI21_X1 U10400 ( .B1(n8877), .B2(n8955), .A(n8957), .ZN(n8874) );
  NAND4_X1 U10401 ( .A1(n8876), .A2(n8875), .A3(n9145), .A4(n8874), .ZN(n8881)
         );
  NAND2_X1 U10402 ( .A1(n8877), .A2(n8949), .ZN(n8878) );
  NAND2_X1 U10403 ( .A1(n8957), .A2(n8878), .ZN(n8879) );
  NAND2_X1 U10404 ( .A1(n8879), .A2(n9163), .ZN(n8880) );
  MUX2_X1 U10405 ( .A(n8883), .B(n8882), .S(n9031), .Z(n8884) );
  NAND2_X1 U10406 ( .A1(n8885), .A2(n8888), .ZN(n8887) );
  OR2_X1 U10407 ( .A1(n8890), .A2(n10398), .ZN(n8886) );
  MUX2_X1 U10408 ( .A(n8894), .B(n9031), .S(n8979), .Z(n8893) );
  NAND2_X1 U10409 ( .A1(n8889), .A2(n8888), .ZN(n8892) );
  OR2_X1 U10410 ( .A1(n8890), .A2(n10332), .ZN(n8891) );
  INV_X1 U10411 ( .A(n8983), .ZN(n9128) );
  NOR2_X1 U10412 ( .A1(n9128), .A2(n8965), .ZN(n8977) );
  NOR3_X1 U10413 ( .A1(n8893), .A2(n9015), .A3(n8977), .ZN(n8898) );
  NOR3_X1 U10414 ( .A1(n8895), .A2(n9338), .A3(n8965), .ZN(n8897) );
  INV_X1 U10415 ( .A(n9338), .ZN(n8896) );
  NOR3_X1 U10416 ( .A1(n8898), .A2(n8897), .A3(n9018), .ZN(n9028) );
  AND2_X1 U10417 ( .A1(n8979), .A2(n8965), .ZN(n9013) );
  INV_X1 U10418 ( .A(n9013), .ZN(n8901) );
  NAND2_X1 U10419 ( .A1(n8901), .A2(n8900), .ZN(n8980) );
  INV_X1 U10420 ( .A(n8980), .ZN(n8967) );
  INV_X1 U10421 ( .A(n8902), .ZN(n8945) );
  INV_X1 U10422 ( .A(n8996), .ZN(n8921) );
  NAND2_X1 U10423 ( .A1(n8904), .A2(n8903), .ZN(n8912) );
  NAND2_X1 U10424 ( .A1(n6884), .A2(n8905), .ZN(n8906) );
  NAND4_X1 U10425 ( .A1(n8908), .A2(n8907), .A3(n8988), .A4(n8906), .ZN(n8911)
         );
  INV_X1 U10426 ( .A(n8909), .ZN(n8910) );
  OAI21_X1 U10427 ( .B1(n8912), .B2(n8911), .A(n8910), .ZN(n8914) );
  OAI21_X1 U10428 ( .B1(n8915), .B2(n8914), .A(n8913), .ZN(n8920) );
  INV_X1 U10429 ( .A(n8916), .ZN(n8919) );
  INV_X1 U10430 ( .A(n8917), .ZN(n8918) );
  AOI211_X1 U10431 ( .C1(n8921), .C2(n8920), .A(n8919), .B(n8918), .ZN(n8925)
         );
  INV_X1 U10432 ( .A(n8922), .ZN(n8923) );
  OAI21_X1 U10433 ( .B1(n8925), .B2(n8924), .A(n8923), .ZN(n8927) );
  AOI21_X1 U10434 ( .B1(n8928), .B2(n8927), .A(n8926), .ZN(n8931) );
  OAI211_X1 U10435 ( .C1(n8931), .C2(n8930), .A(n9007), .B(n8929), .ZN(n8934)
         );
  INV_X1 U10436 ( .A(n8932), .ZN(n8933) );
  AOI21_X1 U10437 ( .B1(n9006), .B2(n8934), .A(n8933), .ZN(n8944) );
  INV_X1 U10438 ( .A(n8935), .ZN(n8942) );
  NAND2_X1 U10439 ( .A1(n8937), .A2(n8936), .ZN(n8938) );
  NAND2_X1 U10440 ( .A1(n8938), .A2(n9191), .ZN(n8940) );
  AND2_X1 U10441 ( .A1(n8940), .A2(n8939), .ZN(n8950) );
  INV_X1 U10442 ( .A(n8950), .ZN(n8941) );
  NAND3_X1 U10443 ( .A1(n8957), .A2(n8942), .A3(n8941), .ZN(n8971) );
  INV_X1 U10444 ( .A(n8971), .ZN(n8943) );
  OAI21_X1 U10445 ( .B1(n8945), .B2(n8944), .A(n8943), .ZN(n8947) );
  INV_X1 U10446 ( .A(n8974), .ZN(n8946) );
  AOI21_X1 U10447 ( .B1(n8947), .B2(n9163), .A(n8946), .ZN(n8964) );
  INV_X1 U10448 ( .A(n8955), .ZN(n8952) );
  NOR2_X1 U10449 ( .A1(n8953), .A2(n8948), .ZN(n8951) );
  AOI22_X1 U10450 ( .A1(n8952), .A2(n8951), .B1(n8950), .B2(n8949), .ZN(n8958)
         );
  OR3_X1 U10451 ( .A1(n8955), .A2(n8954), .A3(n8953), .ZN(n8956) );
  NAND4_X1 U10452 ( .A1(n8974), .A2(n8958), .A3(n8957), .A4(n8956), .ZN(n8959)
         );
  NAND2_X1 U10453 ( .A1(n8960), .A2(n8959), .ZN(n8972) );
  NAND2_X1 U10454 ( .A1(n8962), .A2(n8961), .ZN(n8976) );
  INV_X1 U10455 ( .A(n8976), .ZN(n8963) );
  OAI21_X1 U10456 ( .B1(n8964), .B2(n8972), .A(n8963), .ZN(n8966) );
  NOR2_X1 U10457 ( .A1(n8979), .A2(n8965), .ZN(n9014) );
  AOI21_X1 U10458 ( .B1(n8967), .B2(n8966), .A(n9014), .ZN(n8968) );
  OAI21_X1 U10459 ( .B1(n8968), .B2(n9015), .A(n9030), .ZN(n8969) );
  XNOR2_X1 U10460 ( .A(n8969), .B(n9021), .ZN(n9023) );
  OAI21_X1 U10461 ( .B1(n8971), .B2(n8970), .A(n9163), .ZN(n8973) );
  AOI21_X1 U10462 ( .B1(n8974), .B2(n8973), .A(n8972), .ZN(n8975) );
  NOR2_X1 U10463 ( .A1(n8976), .A2(n8975), .ZN(n8981) );
  INV_X1 U10464 ( .A(n8977), .ZN(n8978) );
  OAI22_X1 U10465 ( .A1(n8981), .A2(n8980), .B1(n8979), .B2(n8978), .ZN(n8982)
         );
  INV_X1 U10466 ( .A(n9015), .ZN(n9037) );
  OAI211_X1 U10467 ( .C1(n9341), .C2(n8983), .A(n8982), .B(n9037), .ZN(n9016)
         );
  NOR2_X1 U10468 ( .A1(n8986), .A2(n8985), .ZN(n8991) );
  NOR2_X1 U10469 ( .A1(n8987), .A2(n9670), .ZN(n8990) );
  NOR2_X1 U10470 ( .A1(n9684), .A2(n8988), .ZN(n8989) );
  NAND4_X1 U10471 ( .A1(n8991), .A2(n8990), .A3(n4528), .A4(n8989), .ZN(n8992)
         );
  OR3_X1 U10472 ( .A1(n8994), .A2(n8993), .A3(n8992), .ZN(n8995) );
  NOR2_X1 U10473 ( .A1(n8996), .A2(n8995), .ZN(n8997) );
  NAND3_X1 U10474 ( .A1(n8999), .A2(n8998), .A3(n8997), .ZN(n9000) );
  OR4_X1 U10475 ( .A1(n9002), .A2(n9617), .A3(n9001), .A4(n9000), .ZN(n9003)
         );
  NOR2_X1 U10476 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  NAND4_X1 U10477 ( .A1(n9286), .A2(n9007), .A3(n9006), .A4(n9005), .ZN(n9008)
         );
  NOR2_X1 U10478 ( .A1(n9275), .A2(n9008), .ZN(n9009) );
  NAND4_X1 U10479 ( .A1(n9010), .A2(n9238), .A3(n9009), .A4(n9254), .ZN(n9011)
         );
  NOR4_X2 U10480 ( .A1(n9015), .A2(n9014), .A3(n9013), .A4(n9012), .ZN(n9020)
         );
  AOI21_X1 U10481 ( .B1(n9017), .B2(n9016), .A(n9020), .ZN(n9019) );
  NOR2_X1 U10482 ( .A1(n9019), .A2(n9018), .ZN(n9022) );
  NAND3_X1 U10483 ( .A1(n9026), .A2(n9064), .A3(n9025), .ZN(n9027) );
  OAI211_X1 U10484 ( .C1(n9033), .C2(n9034), .A(n9027), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9039) );
  INV_X1 U10485 ( .A(n9028), .ZN(n9029) );
  OAI21_X1 U10486 ( .B1(n9031), .B2(n9030), .A(n9029), .ZN(n9036) );
  NOR3_X1 U10487 ( .A1(n9034), .A2(n9033), .A3(n9032), .ZN(n9035) );
  OAI211_X1 U10488 ( .C1(n9037), .C2(n5702), .A(n9036), .B(n9035), .ZN(n9038)
         );
  NAND3_X1 U10489 ( .A1(n9040), .A2(n9039), .A3(n9038), .ZN(P1_U3242) );
  MUX2_X1 U10490 ( .A(n9041), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9051), .Z(
        P1_U3583) );
  MUX2_X1 U10491 ( .A(n9171), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9051), .Z(
        P1_U3582) );
  MUX2_X1 U10492 ( .A(n9183), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9051), .Z(
        P1_U3581) );
  MUX2_X1 U10493 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9199), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10494 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9042), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10495 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9228), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10496 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9388), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10497 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9397), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10498 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9389), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10499 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9398), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10500 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9309), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10501 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9043), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10502 ( .A(n9044), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9051), .Z(
        P1_U3571) );
  MUX2_X1 U10503 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9045), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10504 ( .A(n9046), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9051), .Z(
        P1_U3569) );
  MUX2_X1 U10505 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9047), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10506 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9768), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10507 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9630), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10508 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9767), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10509 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9629), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10510 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9739), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10511 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9048), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10512 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9646), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10513 ( .A(n9049), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9051), .Z(
        P1_U3559) );
  MUX2_X1 U10514 ( .A(n9662), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9051), .Z(
        P1_U3558) );
  MUX2_X1 U10515 ( .A(n9050), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9051), .Z(
        P1_U3557) );
  MUX2_X1 U10516 ( .A(n5779), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9051), .Z(
        P1_U3556) );
  MUX2_X1 U10517 ( .A(n6884), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9051), .Z(
        P1_U3555) );
  INV_X1 U10518 ( .A(n9599), .ZN(n9550) );
  INV_X1 U10519 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9052) );
  OAI22_X1 U10520 ( .A1(n9604), .A2(n10322), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9052), .ZN(n9053) );
  AOI21_X1 U10521 ( .B1(n9054), .B2(n9550), .A(n9053), .ZN(n9063) );
  OAI211_X1 U10522 ( .C1(n9057), .C2(n9056), .A(n9595), .B(n9055), .ZN(n9062)
         );
  OAI211_X1 U10523 ( .C1(n9060), .C2(n9059), .A(n9590), .B(n9058), .ZN(n9061)
         );
  NAND3_X1 U10524 ( .A1(n9063), .A2(n9062), .A3(n9061), .ZN(P1_U3244) );
  INV_X1 U10525 ( .A(n9064), .ZN(n9066) );
  OAI21_X1 U10526 ( .B1(n9066), .B2(n9065), .A(P1_U3973), .ZN(n9070) );
  NOR3_X1 U10527 ( .A1(n9068), .A2(n9067), .A3(n4502), .ZN(n9069) );
  AOI211_X1 U10528 ( .C1(n9072), .C2(n9071), .A(n9070), .B(n9069), .ZN(n9551)
         );
  INV_X1 U10529 ( .A(n9551), .ZN(n9086) );
  INV_X1 U10530 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9074) );
  OAI22_X1 U10531 ( .A1(n9604), .A2(n9074), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9073), .ZN(n9075) );
  AOI21_X1 U10532 ( .B1(n9076), .B2(n9550), .A(n9075), .ZN(n9085) );
  OAI211_X1 U10533 ( .C1(n9079), .C2(n9078), .A(n9595), .B(n9077), .ZN(n9084)
         );
  OAI211_X1 U10534 ( .C1(n9082), .C2(n9081), .A(n9590), .B(n9080), .ZN(n9083)
         );
  NAND4_X1 U10535 ( .A1(n9086), .A2(n9085), .A3(n9084), .A4(n9083), .ZN(
        P1_U3245) );
  OAI21_X1 U10536 ( .B1(n9604), .B2(n10367), .A(n9087), .ZN(n9088) );
  AOI21_X1 U10537 ( .B1(n9089), .B2(n9550), .A(n9088), .ZN(n9098) );
  OAI211_X1 U10538 ( .C1(n9092), .C2(n9091), .A(n9590), .B(n9090), .ZN(n9097)
         );
  OAI211_X1 U10539 ( .C1(n9095), .C2(n9094), .A(n9595), .B(n9093), .ZN(n9096)
         );
  NAND3_X1 U10540 ( .A1(n9098), .A2(n9097), .A3(n9096), .ZN(P1_U3246) );
  OAI21_X1 U10541 ( .B1(n9101), .B2(n9100), .A(n9099), .ZN(n9102) );
  NAND2_X1 U10542 ( .A1(n9102), .A2(n9590), .ZN(n9112) );
  AOI21_X1 U10543 ( .B1(n9553), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9103), .ZN(
        n9111) );
  OAI21_X1 U10544 ( .B1(n9106), .B2(n9105), .A(n9104), .ZN(n9107) );
  NAND2_X1 U10545 ( .A1(n9107), .A2(n9595), .ZN(n9110) );
  NAND2_X1 U10546 ( .A1(n9550), .A2(n9108), .ZN(n9109) );
  NAND4_X1 U10547 ( .A1(n9112), .A2(n9111), .A3(n9110), .A4(n9109), .ZN(
        P1_U3252) );
  OAI211_X1 U10548 ( .C1(n9115), .C2(n9114), .A(n9113), .B(n9590), .ZN(n9125)
         );
  AOI21_X1 U10549 ( .B1(n9553), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9116), .ZN(
        n9124) );
  AOI21_X1 U10550 ( .B1(n9118), .B2(n9117), .A(n9543), .ZN(n9120) );
  NAND2_X1 U10551 ( .A1(n9120), .A2(n9119), .ZN(n9123) );
  NAND2_X1 U10552 ( .A1(n9550), .A2(n9121), .ZN(n9122) );
  NAND4_X1 U10553 ( .A1(n9125), .A2(n9124), .A3(n9123), .A4(n9122), .ZN(
        P1_U3261) );
  NAND2_X1 U10554 ( .A1(n9132), .A2(n9341), .ZN(n9131) );
  XNOR2_X1 U10555 ( .A(n9131), .B(n9338), .ZN(n9126) );
  NAND2_X1 U10556 ( .A1(n9126), .A2(n9673), .ZN(n9337) );
  OR2_X1 U10557 ( .A1(n9128), .A2(n9127), .ZN(n9339) );
  NOR2_X1 U10558 ( .A1(n9339), .A2(n9634), .ZN(n9134) );
  NOR2_X1 U10559 ( .A1(n9338), .A2(n9668), .ZN(n9129) );
  AOI211_X1 U10560 ( .C1(n9666), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9134), .B(
        n9129), .ZN(n9130) );
  OAI21_X1 U10561 ( .B1(n9337), .B2(n9264), .A(n9130), .ZN(P1_U3263) );
  OAI211_X1 U10562 ( .C1(n9132), .C2(n9341), .A(n9673), .B(n9131), .ZN(n9340)
         );
  NOR2_X1 U10563 ( .A1(n9341), .A2(n9668), .ZN(n9133) );
  AOI211_X1 U10564 ( .C1(n9666), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9134), .B(
        n9133), .ZN(n9135) );
  OAI21_X1 U10565 ( .B1(n9264), .B2(n9340), .A(n9135), .ZN(P1_U3264) );
  NAND2_X1 U10566 ( .A1(n9138), .A2(n9676), .ZN(n9141) );
  AOI22_X1 U10567 ( .A1(n9634), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9139), .B2(
        n9651), .ZN(n9140) );
  OAI211_X1 U10568 ( .C1(n9142), .C2(n9668), .A(n9141), .B(n9140), .ZN(n9143)
         );
  AOI21_X1 U10569 ( .B1(n9137), .B2(n9677), .A(n9143), .ZN(n9144) );
  OAI21_X1 U10570 ( .B1(n9136), .B2(n9666), .A(n9144), .ZN(P1_U3356) );
  NAND2_X1 U10571 ( .A1(n9165), .A2(n9145), .ZN(n9147) );
  INV_X1 U10572 ( .A(n9156), .ZN(n9146) );
  OAI211_X1 U10573 ( .C1(n9343), .C2(n9167), .A(n9673), .B(n9150), .ZN(n9346)
         );
  AOI22_X1 U10574 ( .A1(n9634), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9151), .B2(
        n9651), .ZN(n9154) );
  NAND2_X1 U10575 ( .A1(n9152), .A2(n9652), .ZN(n9153) );
  OAI211_X1 U10576 ( .C1(n9346), .C2(n9264), .A(n9154), .B(n9153), .ZN(n9155)
         );
  INV_X1 U10577 ( .A(n9155), .ZN(n9160) );
  NAND3_X1 U10578 ( .A1(n9342), .A2(n9158), .A3(n9677), .ZN(n9159) );
  OAI211_X1 U10579 ( .C1(n9348), .C2(n9634), .A(n9160), .B(n9159), .ZN(
        P1_U3265) );
  XNOR2_X1 U10580 ( .A(n9161), .B(n4997), .ZN(n9356) );
  NAND2_X1 U10581 ( .A1(n9164), .A2(n9163), .ZN(n9166) );
  OAI21_X1 U10582 ( .B1(n9162), .B2(n9166), .A(n9165), .ZN(n9353) );
  AOI211_X1 U10583 ( .C1(n9352), .C2(n9181), .A(n9321), .B(n9167), .ZN(n9350)
         );
  NAND2_X1 U10584 ( .A1(n9350), .A2(n9676), .ZN(n9173) );
  AOI22_X1 U10585 ( .A1(n9634), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9168), .B2(
        n9651), .ZN(n9169) );
  OAI21_X1 U10586 ( .B1(n9307), .B2(n9367), .A(n9169), .ZN(n9170) );
  AOI21_X1 U10587 ( .B1(n9310), .B2(n9171), .A(n9170), .ZN(n9172) );
  OAI211_X1 U10588 ( .C1(n9174), .C2(n9668), .A(n9173), .B(n9172), .ZN(n9175)
         );
  AOI21_X1 U10589 ( .B1(n9353), .B2(n9266), .A(n9175), .ZN(n9176) );
  OAI21_X1 U10590 ( .B1(n9356), .B2(n9336), .A(n9176), .ZN(P1_U3266) );
  AOI21_X1 U10591 ( .B1(n9177), .B2(n9179), .A(n9162), .ZN(n9365) );
  XOR2_X1 U10592 ( .A(n9179), .B(n9178), .Z(n9357) );
  NAND2_X1 U10593 ( .A1(n9357), .A2(n9677), .ZN(n9190) );
  INV_X1 U10594 ( .A(n9181), .ZN(n9182) );
  AOI211_X1 U10595 ( .C1(n9362), .C2(n9195), .A(n9321), .B(n9182), .ZN(n9360)
         );
  NOR2_X1 U10596 ( .A1(n5696), .A2(n9668), .ZN(n9188) );
  NAND2_X1 U10597 ( .A1(n9310), .A2(n9183), .ZN(n9186) );
  AOI22_X1 U10598 ( .A1(n9666), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9184), .B2(
        n9651), .ZN(n9185) );
  OAI211_X1 U10599 ( .C1(n9358), .C2(n9307), .A(n9186), .B(n9185), .ZN(n9187)
         );
  AOI211_X1 U10600 ( .C1(n9360), .C2(n9676), .A(n9188), .B(n9187), .ZN(n9189)
         );
  OAI211_X1 U10601 ( .C1(n9365), .C2(n9316), .A(n9190), .B(n9189), .ZN(
        P1_U3267) );
  NAND2_X1 U10602 ( .A1(n4879), .A2(n9191), .ZN(n9192) );
  AOI21_X1 U10603 ( .B1(n9193), .B2(n9192), .A(n4576), .ZN(n9373) );
  XNOR2_X1 U10604 ( .A(n9194), .B(n9193), .ZN(n9366) );
  NAND2_X1 U10605 ( .A1(n9366), .A2(n9677), .ZN(n9204) );
  AOI211_X1 U10606 ( .C1(n9370), .C2(n9206), .A(n9321), .B(n9180), .ZN(n9368)
         );
  AOI22_X1 U10607 ( .A1(n9634), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9196), .B2(
        n9651), .ZN(n9197) );
  OAI21_X1 U10608 ( .B1(n9307), .B2(n9380), .A(n9197), .ZN(n9198) );
  AOI21_X1 U10609 ( .B1(n9310), .B2(n9199), .A(n9198), .ZN(n9200) );
  OAI21_X1 U10610 ( .B1(n9201), .B2(n9668), .A(n9200), .ZN(n9202) );
  AOI21_X1 U10611 ( .B1(n9368), .B2(n9676), .A(n9202), .ZN(n9203) );
  OAI211_X1 U10612 ( .C1(n9373), .C2(n9316), .A(n9204), .B(n9203), .ZN(
        P1_U3268) );
  XNOR2_X1 U10613 ( .A(n9205), .B(n9214), .ZN(n9378) );
  INV_X1 U10614 ( .A(n9226), .ZN(n9208) );
  INV_X1 U10615 ( .A(n9206), .ZN(n9207) );
  AOI211_X1 U10616 ( .C1(n9375), .C2(n9208), .A(n9321), .B(n9207), .ZN(n9374)
         );
  AOI22_X1 U10617 ( .A1(n9666), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9209), .B2(
        n9651), .ZN(n9210) );
  OAI21_X1 U10618 ( .B1(n9211), .B2(n9668), .A(n9210), .ZN(n9221) );
  NOR2_X1 U10619 ( .A1(n9212), .A2(n9754), .ZN(n9219) );
  OAI21_X1 U10620 ( .B1(n9213), .B2(n9215), .A(n9214), .ZN(n9218) );
  OAI22_X1 U10621 ( .A1(n9216), .A2(n9787), .B1(n9358), .B2(n9789), .ZN(n9217)
         );
  AOI21_X1 U10622 ( .B1(n9219), .B2(n9218), .A(n9217), .ZN(n9377) );
  NOR2_X1 U10623 ( .A1(n9377), .A2(n9634), .ZN(n9220) );
  AOI211_X1 U10624 ( .C1(n9374), .C2(n9676), .A(n9221), .B(n9220), .ZN(n9222)
         );
  OAI21_X1 U10625 ( .B1(n9336), .B2(n9378), .A(n9222), .ZN(P1_U3269) );
  AOI21_X1 U10626 ( .B1(n9223), .B2(n9224), .A(n9213), .ZN(n9387) );
  XNOR2_X1 U10627 ( .A(n9225), .B(n9224), .ZN(n9379) );
  NAND2_X1 U10628 ( .A1(n9379), .A2(n9677), .ZN(n9235) );
  AOI211_X1 U10629 ( .C1(n9384), .C2(n9241), .A(n9321), .B(n9226), .ZN(n9382)
         );
  NOR2_X1 U10630 ( .A1(n9227), .A2(n9668), .ZN(n9233) );
  NAND2_X1 U10631 ( .A1(n9310), .A2(n9228), .ZN(n9231) );
  AOI22_X1 U10632 ( .A1(n9634), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9229), .B2(
        n9651), .ZN(n9230) );
  OAI211_X1 U10633 ( .C1(n9381), .C2(n9307), .A(n9231), .B(n9230), .ZN(n9232)
         );
  AOI211_X1 U10634 ( .C1(n9382), .C2(n9676), .A(n9233), .B(n9232), .ZN(n9234)
         );
  OAI211_X1 U10635 ( .C1(n9387), .C2(n9316), .A(n9235), .B(n9234), .ZN(
        P1_U3270) );
  XNOR2_X1 U10636 ( .A(n9237), .B(n9236), .ZN(n9396) );
  XNOR2_X1 U10637 ( .A(n9239), .B(n9238), .ZN(n9394) );
  AOI21_X1 U10638 ( .B1(n9248), .B2(n9257), .A(n9321), .ZN(n9242) );
  NAND2_X1 U10639 ( .A1(n9242), .A2(n9241), .ZN(n9391) );
  NAND2_X1 U10640 ( .A1(n9310), .A2(n9388), .ZN(n9246) );
  NOR2_X1 U10641 ( .A1(n9664), .A2(n9243), .ZN(n9244) );
  AOI21_X1 U10642 ( .B1(n9666), .B2(P1_REG2_REG_22__SCAN_IN), .A(n9244), .ZN(
        n9245) );
  OAI211_X1 U10643 ( .C1(n9277), .C2(n9307), .A(n9246), .B(n9245), .ZN(n9247)
         );
  AOI21_X1 U10644 ( .B1(n9248), .B2(n9652), .A(n9247), .ZN(n9249) );
  OAI21_X1 U10645 ( .B1(n9391), .B2(n9264), .A(n9249), .ZN(n9250) );
  AOI21_X1 U10646 ( .B1(n9394), .B2(n9677), .A(n9250), .ZN(n9251) );
  OAI21_X1 U10647 ( .B1(n9316), .B2(n9396), .A(n9251), .ZN(P1_U3271) );
  XNOR2_X1 U10648 ( .A(n9252), .B(n9254), .ZN(n9405) );
  OAI21_X1 U10649 ( .B1(n9255), .B2(n9254), .A(n9253), .ZN(n9403) );
  INV_X1 U10650 ( .A(n9256), .ZN(n9270) );
  OAI211_X1 U10651 ( .C1(n9401), .C2(n9270), .A(n9673), .B(n9257), .ZN(n9400)
         );
  NAND2_X1 U10652 ( .A1(n9310), .A2(n9397), .ZN(n9260) );
  AOI22_X1 U10653 ( .A1(n9634), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9258), .B2(
        n9651), .ZN(n9259) );
  OAI211_X1 U10654 ( .C1(n9288), .C2(n9307), .A(n9260), .B(n9259), .ZN(n9261)
         );
  AOI21_X1 U10655 ( .B1(n9262), .B2(n9652), .A(n9261), .ZN(n9263) );
  OAI21_X1 U10656 ( .B1(n9400), .B2(n9264), .A(n9263), .ZN(n9265) );
  AOI21_X1 U10657 ( .B1(n9403), .B2(n9266), .A(n9265), .ZN(n9267) );
  OAI21_X1 U10658 ( .B1(n9405), .B2(n9336), .A(n9267), .ZN(P1_U3272) );
  XOR2_X1 U10659 ( .A(n9269), .B(n9275), .Z(n9410) );
  AOI21_X1 U10660 ( .B1(n9406), .B2(n4659), .A(n9270), .ZN(n9407) );
  AOI22_X1 U10661 ( .A1(n9634), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9271), .B2(
        n9651), .ZN(n9272) );
  OAI21_X1 U10662 ( .B1(n9273), .B2(n9668), .A(n9272), .ZN(n9281) );
  AOI211_X1 U10663 ( .C1(n9276), .C2(n9275), .A(n9754), .B(n9274), .ZN(n9279)
         );
  OAI22_X1 U10664 ( .A1(n9277), .A2(n9789), .B1(n9417), .B2(n9787), .ZN(n9278)
         );
  NOR2_X1 U10665 ( .A1(n9279), .A2(n9278), .ZN(n9409) );
  NOR2_X1 U10666 ( .A1(n9409), .A2(n9634), .ZN(n9280) );
  AOI211_X1 U10667 ( .C1(n9407), .C2(n9282), .A(n9281), .B(n9280), .ZN(n9283)
         );
  OAI21_X1 U10668 ( .B1(n9336), .B2(n9410), .A(n9283), .ZN(P1_U3273) );
  XOR2_X1 U10669 ( .A(n9284), .B(n9286), .Z(n9415) );
  OAI211_X1 U10670 ( .C1(n9287), .C2(n9286), .A(n9285), .B(n9777), .ZN(n9290)
         );
  OR2_X1 U10671 ( .A1(n9288), .A2(n9789), .ZN(n9289) );
  OAI211_X1 U10672 ( .C1(n9330), .C2(n9787), .A(n9290), .B(n9289), .ZN(n9411)
         );
  AOI211_X1 U10673 ( .C1(n9413), .C2(n9303), .A(n9321), .B(n9291), .ZN(n9412)
         );
  NAND2_X1 U10674 ( .A1(n9412), .A2(n9676), .ZN(n9294) );
  AOI22_X1 U10675 ( .A1(n9666), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9292), .B2(
        n9651), .ZN(n9293) );
  OAI211_X1 U10676 ( .C1(n4657), .C2(n9668), .A(n9294), .B(n9293), .ZN(n9295)
         );
  AOI21_X1 U10677 ( .B1(n9411), .B2(n9296), .A(n9295), .ZN(n9297) );
  OAI21_X1 U10678 ( .B1(n9415), .B2(n9336), .A(n9297), .ZN(P1_U3274) );
  INV_X1 U10679 ( .A(n9326), .ZN(n9299) );
  NAND2_X1 U10680 ( .A1(n9299), .A2(n9298), .ZN(n9301) );
  AOI21_X1 U10681 ( .B1(n9302), .B2(n9301), .A(n9300), .ZN(n9424) );
  XOR2_X1 U10682 ( .A(n9302), .B(n4582), .Z(n9416) );
  NAND2_X1 U10683 ( .A1(n9416), .A2(n9677), .ZN(n9315) );
  INV_X1 U10684 ( .A(n9303), .ZN(n9304) );
  AOI211_X1 U10685 ( .C1(n9421), .C2(n9319), .A(n9321), .B(n9304), .ZN(n9419)
         );
  AOI22_X1 U10686 ( .A1(n9634), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9305), .B2(
        n9651), .ZN(n9306) );
  OAI21_X1 U10687 ( .B1(n9307), .B2(n9418), .A(n9306), .ZN(n9308) );
  AOI21_X1 U10688 ( .B1(n9310), .B2(n9309), .A(n9308), .ZN(n9311) );
  OAI21_X1 U10689 ( .B1(n9312), .B2(n9668), .A(n9311), .ZN(n9313) );
  AOI21_X1 U10690 ( .B1(n9419), .B2(n9676), .A(n9313), .ZN(n9314) );
  OAI211_X1 U10691 ( .C1(n9424), .C2(n9316), .A(n9315), .B(n9314), .ZN(
        P1_U3275) );
  XNOR2_X1 U10692 ( .A(n9318), .B(n9317), .ZN(n9429) );
  INV_X1 U10693 ( .A(n9319), .ZN(n9320) );
  AOI211_X1 U10694 ( .C1(n9426), .C2(n9322), .A(n9321), .B(n9320), .ZN(n9425)
         );
  AOI22_X1 U10695 ( .A1(n9634), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9323), .B2(
        n9651), .ZN(n9324) );
  OAI21_X1 U10696 ( .B1(n9325), .B2(n9668), .A(n9324), .ZN(n9334) );
  AOI211_X1 U10697 ( .C1(n9328), .C2(n9327), .A(n9754), .B(n9326), .ZN(n9332)
         );
  OAI22_X1 U10698 ( .A1(n9330), .A2(n9789), .B1(n9329), .B2(n9787), .ZN(n9331)
         );
  NOR2_X1 U10699 ( .A1(n9332), .A2(n9331), .ZN(n9428) );
  NOR2_X1 U10700 ( .A1(n9428), .A2(n9666), .ZN(n9333) );
  AOI211_X1 U10701 ( .C1(n9425), .C2(n9676), .A(n9334), .B(n9333), .ZN(n9335)
         );
  OAI21_X1 U10702 ( .B1(n9429), .B2(n9336), .A(n9335), .ZN(P1_U3276) );
  OAI211_X1 U10703 ( .C1(n9338), .C2(n9781), .A(n9337), .B(n9339), .ZN(n9435)
         );
  MUX2_X1 U10704 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9435), .S(n9825), .Z(
        P1_U3553) );
  OAI211_X1 U10705 ( .C1(n9341), .C2(n9781), .A(n9340), .B(n9339), .ZN(n9436)
         );
  MUX2_X1 U10706 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9436), .S(n9825), .Z(
        P1_U3552) );
  NAND2_X1 U10707 ( .A1(n9152), .A2(n9344), .ZN(n9345) );
  OAI22_X1 U10708 ( .A1(n9349), .A2(n9789), .B1(n9367), .B2(n9787), .ZN(n9351)
         );
  AOI211_X1 U10709 ( .C1(n9344), .C2(n9352), .A(n9351), .B(n9350), .ZN(n9355)
         );
  NAND2_X1 U10710 ( .A1(n9353), .A2(n9777), .ZN(n9354) );
  OAI211_X1 U10711 ( .C1(n9356), .C2(n9772), .A(n9355), .B(n9354), .ZN(n9438)
         );
  MUX2_X1 U10712 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9438), .S(n9825), .Z(
        P1_U3549) );
  NAND2_X1 U10713 ( .A1(n9357), .A2(n9784), .ZN(n9364) );
  OAI22_X1 U10714 ( .A1(n9359), .A2(n9789), .B1(n9358), .B2(n9787), .ZN(n9361)
         );
  AOI211_X1 U10715 ( .C1(n9344), .C2(n9362), .A(n9361), .B(n9360), .ZN(n9363)
         );
  OAI211_X1 U10716 ( .C1(n9754), .C2(n9365), .A(n9364), .B(n9363), .ZN(n9439)
         );
  MUX2_X1 U10717 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9439), .S(n9825), .Z(
        P1_U3548) );
  NAND2_X1 U10718 ( .A1(n9366), .A2(n9784), .ZN(n9372) );
  OAI22_X1 U10719 ( .A1(n9380), .A2(n9787), .B1(n9367), .B2(n9789), .ZN(n9369)
         );
  AOI211_X1 U10720 ( .C1(n9344), .C2(n9370), .A(n9369), .B(n9368), .ZN(n9371)
         );
  OAI211_X1 U10721 ( .C1(n9754), .C2(n9373), .A(n9372), .B(n9371), .ZN(n9440)
         );
  MUX2_X1 U10722 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9440), .S(n9825), .Z(
        P1_U3547) );
  AOI21_X1 U10723 ( .B1(n9344), .B2(n9375), .A(n9374), .ZN(n9376) );
  OAI211_X1 U10724 ( .C1(n9378), .C2(n9772), .A(n9377), .B(n9376), .ZN(n9441)
         );
  MUX2_X1 U10725 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9441), .S(n9825), .Z(
        P1_U3546) );
  NAND2_X1 U10726 ( .A1(n9379), .A2(n9784), .ZN(n9386) );
  OAI22_X1 U10727 ( .A1(n9381), .A2(n9787), .B1(n9380), .B2(n9789), .ZN(n9383)
         );
  AOI211_X1 U10728 ( .C1(n9344), .C2(n9384), .A(n9383), .B(n9382), .ZN(n9385)
         );
  OAI211_X1 U10729 ( .C1(n9754), .C2(n9387), .A(n9386), .B(n9385), .ZN(n9442)
         );
  MUX2_X1 U10730 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9442), .S(n9825), .Z(
        P1_U3545) );
  AOI22_X1 U10731 ( .A1(n9766), .A2(n9389), .B1(n9388), .B2(n9769), .ZN(n9390)
         );
  OAI211_X1 U10732 ( .C1(n9392), .C2(n9781), .A(n9391), .B(n9390), .ZN(n9393)
         );
  AOI21_X1 U10733 ( .B1(n9394), .B2(n9784), .A(n9393), .ZN(n9395) );
  OAI21_X1 U10734 ( .B1(n9754), .B2(n9396), .A(n9395), .ZN(n9443) );
  MUX2_X1 U10735 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9443), .S(n9825), .Z(
        P1_U3544) );
  AOI22_X1 U10736 ( .A1(n9766), .A2(n9398), .B1(n9397), .B2(n9769), .ZN(n9399)
         );
  OAI211_X1 U10737 ( .C1(n9401), .C2(n9781), .A(n9400), .B(n9399), .ZN(n9402)
         );
  AOI21_X1 U10738 ( .B1(n9403), .B2(n9777), .A(n9402), .ZN(n9404) );
  OAI21_X1 U10739 ( .B1(n9405), .B2(n9772), .A(n9404), .ZN(n9444) );
  MUX2_X1 U10740 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9444), .S(n9825), .Z(
        P1_U3543) );
  AOI22_X1 U10741 ( .A1(n9407), .A2(n9673), .B1(n9344), .B2(n9406), .ZN(n9408)
         );
  OAI211_X1 U10742 ( .C1(n9410), .C2(n9772), .A(n9409), .B(n9408), .ZN(n9445)
         );
  MUX2_X1 U10743 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9445), .S(n9825), .Z(
        P1_U3542) );
  AOI211_X1 U10744 ( .C1(n9344), .C2(n9413), .A(n9412), .B(n9411), .ZN(n9414)
         );
  OAI21_X1 U10745 ( .B1(n9415), .B2(n9772), .A(n9414), .ZN(n9446) );
  MUX2_X1 U10746 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9446), .S(n9825), .Z(
        P1_U3541) );
  NAND2_X1 U10747 ( .A1(n9416), .A2(n9784), .ZN(n9423) );
  OAI22_X1 U10748 ( .A1(n9418), .A2(n9787), .B1(n9417), .B2(n9789), .ZN(n9420)
         );
  AOI211_X1 U10749 ( .C1(n9344), .C2(n9421), .A(n9420), .B(n9419), .ZN(n9422)
         );
  OAI211_X1 U10750 ( .C1(n9754), .C2(n9424), .A(n9423), .B(n9422), .ZN(n9447)
         );
  MUX2_X1 U10751 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9447), .S(n9825), .Z(
        P1_U3540) );
  AOI21_X1 U10752 ( .B1(n9344), .B2(n9426), .A(n9425), .ZN(n9427) );
  OAI211_X1 U10753 ( .C1(n9429), .C2(n9772), .A(n9428), .B(n9427), .ZN(n9448)
         );
  MUX2_X1 U10754 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9448), .S(n9825), .Z(
        P1_U3539) );
  AOI21_X1 U10755 ( .B1(n9344), .B2(n9431), .A(n9430), .ZN(n9432) );
  OAI211_X1 U10756 ( .C1(n9434), .C2(n9772), .A(n9433), .B(n9432), .ZN(n9449)
         );
  MUX2_X1 U10757 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9449), .S(n9825), .Z(
        P1_U3538) );
  MUX2_X1 U10758 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9435), .S(n9802), .Z(
        P1_U3521) );
  MUX2_X1 U10759 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9436), .S(n9802), .Z(
        P1_U3520) );
  MUX2_X1 U10760 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9438), .S(n9802), .Z(
        P1_U3517) );
  MUX2_X1 U10761 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9439), .S(n9802), .Z(
        P1_U3516) );
  MUX2_X1 U10762 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9440), .S(n9802), .Z(
        P1_U3515) );
  MUX2_X1 U10763 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9441), .S(n9802), .Z(
        P1_U3514) );
  MUX2_X1 U10764 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9442), .S(n9802), .Z(
        P1_U3513) );
  MUX2_X1 U10765 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9443), .S(n9802), .Z(
        P1_U3512) );
  MUX2_X1 U10766 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9444), .S(n9802), .Z(
        P1_U3511) );
  MUX2_X1 U10767 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9445), .S(n9802), .Z(
        P1_U3510) );
  MUX2_X1 U10768 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9446), .S(n9802), .Z(
        P1_U3509) );
  MUX2_X1 U10769 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9447), .S(n9802), .Z(
        P1_U3507) );
  MUX2_X1 U10770 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9448), .S(n9802), .Z(
        P1_U3504) );
  MUX2_X1 U10771 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9449), .S(n9802), .Z(
        P1_U3501) );
  MUX2_X1 U10772 ( .A(P1_D_REG_0__SCAN_IN), .B(n9450), .S(n9681), .Z(P1_U3439)
         );
  INV_X1 U10773 ( .A(n9451), .ZN(n9453) );
  NOR4_X1 U10774 ( .A1(n9453), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9452), .A4(
        P1_U3086), .ZN(n9454) );
  AOI21_X1 U10775 ( .B1(n9455), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9454), .ZN(
        n9456) );
  OAI21_X1 U10776 ( .B1(n9458), .B2(n9457), .A(n9456), .ZN(P1_U3324) );
  INV_X1 U10777 ( .A(n9459), .ZN(n9460) );
  MUX2_X1 U10778 ( .A(n9460), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U10779 ( .A(n9462), .B(n9461), .ZN(n9463) );
  AOI22_X1 U10780 ( .A1(n9463), .A2(n9974), .B1(n9966), .B2(
        P2_ADDR_REG_18__SCAN_IN), .ZN(n9480) );
  INV_X1 U10781 ( .A(n9464), .ZN(n9472) );
  NAND3_X1 U10782 ( .A1(P2_U3893), .A2(n9465), .A3(n9464), .ZN(n9466) );
  NAND3_X1 U10783 ( .A1(n9864), .A2(n9467), .A3(n9466), .ZN(n9470) );
  NAND2_X1 U10784 ( .A1(n9875), .A2(n9468), .ZN(n9469) );
  OAI211_X1 U10785 ( .C1(n9472), .C2(n9471), .A(n9470), .B(n9469), .ZN(n9479)
         );
  NAND2_X1 U10786 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n9478) );
  AOI21_X1 U10787 ( .B1(n9475), .B2(n9474), .A(n9473), .ZN(n9476) );
  OR2_X1 U10788 ( .A1(n9476), .A2(n9980), .ZN(n9477) );
  NAND4_X1 U10789 ( .A1(n9480), .A2(n9479), .A3(n9478), .A4(n9477), .ZN(
        P2_U3200) );
  AOI211_X1 U10790 ( .C1(n9483), .C2(n9482), .A(n9481), .B(n9543), .ZN(n9488)
         );
  AOI211_X1 U10791 ( .C1(n9486), .C2(n9485), .A(n9484), .B(n9538), .ZN(n9487)
         );
  AOI211_X1 U10792 ( .C1(n9550), .C2(n9489), .A(n9488), .B(n9487), .ZN(n9491)
         );
  OAI211_X1 U10793 ( .C1(n9604), .C2(n9492), .A(n9491), .B(n9490), .ZN(
        P1_U3253) );
  INV_X1 U10794 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9508) );
  AOI21_X1 U10795 ( .B1(n9495), .B2(n9494), .A(n9493), .ZN(n9496) );
  NAND2_X1 U10796 ( .A1(n9590), .A2(n9496), .ZN(n9502) );
  AOI21_X1 U10797 ( .B1(n9499), .B2(n9498), .A(n9497), .ZN(n9500) );
  NAND2_X1 U10798 ( .A1(n9595), .A2(n9500), .ZN(n9501) );
  OAI211_X1 U10799 ( .C1(n9599), .C2(n9503), .A(n9502), .B(n9501), .ZN(n9504)
         );
  INV_X1 U10800 ( .A(n9504), .ZN(n9507) );
  INV_X1 U10801 ( .A(n9505), .ZN(n9506) );
  OAI211_X1 U10802 ( .C1(n9604), .C2(n9508), .A(n9507), .B(n9506), .ZN(
        P1_U3250) );
  AOI21_X1 U10803 ( .B1(n9511), .B2(n9510), .A(n9509), .ZN(n9512) );
  NAND2_X1 U10804 ( .A1(n9590), .A2(n9512), .ZN(n9518) );
  AOI21_X1 U10805 ( .B1(n9515), .B2(n9514), .A(n9513), .ZN(n9516) );
  NAND2_X1 U10806 ( .A1(n9595), .A2(n9516), .ZN(n9517) );
  OAI211_X1 U10807 ( .C1(n9599), .C2(n9519), .A(n9518), .B(n9517), .ZN(n9520)
         );
  INV_X1 U10808 ( .A(n9520), .ZN(n9522) );
  NAND2_X1 U10809 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9521) );
  OAI211_X1 U10810 ( .C1(n9604), .C2(n9523), .A(n9522), .B(n9521), .ZN(
        P1_U3251) );
  NOR2_X1 U10811 ( .A1(n9524), .A2(n10057), .ZN(n9526) );
  AOI211_X1 U10812 ( .C1(n9527), .C2(n10030), .A(n9526), .B(n9525), .ZN(n9528)
         );
  AOI22_X1 U10813 ( .A1(n10081), .A2(n9528), .B1(n6267), .B2(n10079), .ZN(
        P2_U3472) );
  INV_X1 U10814 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9529) );
  AOI22_X1 U10815 ( .A1(n10065), .A2(n9529), .B1(n9528), .B2(n10063), .ZN(
        P2_U3429) );
  OAI211_X1 U10816 ( .C1(n9532), .C2(n9781), .A(n9531), .B(n9530), .ZN(n9533)
         );
  AOI21_X1 U10817 ( .B1(n9534), .B2(n9784), .A(n9533), .ZN(n9536) );
  AOI22_X1 U10818 ( .A1(n9825), .A2(n9536), .B1(n9535), .B2(n9823), .ZN(
        P1_U3537) );
  INV_X1 U10819 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U10820 ( .A1(n9802), .A2(n9536), .B1(n10188), .B2(n9801), .ZN(
        P1_U3498) );
  XNOR2_X1 U10821 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10822 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10823 ( .A(n9537), .ZN(n9541) );
  AOI211_X1 U10824 ( .C1(n9541), .C2(n9540), .A(n9539), .B(n9538), .ZN(n9548)
         );
  INV_X1 U10825 ( .A(n9542), .ZN(n9546) );
  AOI211_X1 U10826 ( .C1(n9546), .C2(n9545), .A(n9544), .B(n9543), .ZN(n9547)
         );
  AOI211_X1 U10827 ( .C1(n9550), .C2(n9549), .A(n9548), .B(n9547), .ZN(n9555)
         );
  AOI211_X1 U10828 ( .C1(n9553), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9552), .B(
        n9551), .ZN(n9554) );
  NAND2_X1 U10829 ( .A1(n9555), .A2(n9554), .ZN(P1_U3247) );
  INV_X1 U10830 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10209) );
  AOI21_X1 U10831 ( .B1(n9558), .B2(n9557), .A(n9556), .ZN(n9559) );
  NAND2_X1 U10832 ( .A1(n9590), .A2(n9559), .ZN(n9565) );
  AOI21_X1 U10833 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(n9563) );
  NAND2_X1 U10834 ( .A1(n9595), .A2(n9563), .ZN(n9564) );
  OAI211_X1 U10835 ( .C1(n9599), .C2(n9566), .A(n9565), .B(n9564), .ZN(n9567)
         );
  INV_X1 U10836 ( .A(n9567), .ZN(n9569) );
  OAI211_X1 U10837 ( .C1(n9604), .C2(n10209), .A(n9569), .B(n9568), .ZN(
        P1_U3248) );
  INV_X1 U10838 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9584) );
  AOI21_X1 U10839 ( .B1(n9572), .B2(n9571), .A(n9570), .ZN(n9573) );
  NAND2_X1 U10840 ( .A1(n9590), .A2(n9573), .ZN(n9579) );
  AOI21_X1 U10841 ( .B1(n9576), .B2(n9575), .A(n9574), .ZN(n9577) );
  NAND2_X1 U10842 ( .A1(n9595), .A2(n9577), .ZN(n9578) );
  OAI211_X1 U10843 ( .C1(n9599), .C2(n9580), .A(n9579), .B(n9578), .ZN(n9581)
         );
  INV_X1 U10844 ( .A(n9581), .ZN(n9583) );
  OAI211_X1 U10845 ( .C1(n9604), .C2(n9584), .A(n9583), .B(n9582), .ZN(
        P1_U3249) );
  INV_X1 U10846 ( .A(n9585), .ZN(n9598) );
  AOI21_X1 U10847 ( .B1(n9588), .B2(n9587), .A(n9586), .ZN(n9589) );
  NAND2_X1 U10848 ( .A1(n9590), .A2(n9589), .ZN(n9597) );
  AOI21_X1 U10849 ( .B1(n9593), .B2(n9592), .A(n9591), .ZN(n9594) );
  NAND2_X1 U10850 ( .A1(n9595), .A2(n9594), .ZN(n9596) );
  OAI211_X1 U10851 ( .C1(n9599), .C2(n9598), .A(n9597), .B(n9596), .ZN(n9600)
         );
  INV_X1 U10852 ( .A(n9600), .ZN(n9602) );
  OAI211_X1 U10853 ( .C1(n9604), .C2(n9603), .A(n9602), .B(n9601), .ZN(
        P1_U3254) );
  INV_X1 U10854 ( .A(n9605), .ZN(n9610) );
  AOI21_X1 U10855 ( .B1(n9607), .B2(n9606), .A(n4816), .ZN(n9608) );
  AOI211_X1 U10856 ( .C1(n9610), .C2(n9609), .A(n9754), .B(n9608), .ZN(n9614)
         );
  OAI22_X1 U10857 ( .A1(n9612), .A2(n9789), .B1(n9611), .B2(n9787), .ZN(n9613)
         );
  NOR2_X1 U10858 ( .A1(n9614), .A2(n9613), .ZN(n9780) );
  AOI222_X1 U10859 ( .A1(n9616), .A2(n9652), .B1(P1_REG2_REG_13__SCAN_IN), 
        .B2(n9634), .C1(n9651), .C2(n9615), .ZN(n9624) );
  XNOR2_X1 U10860 ( .A(n9618), .B(n9617), .ZN(n9785) );
  INV_X1 U10861 ( .A(n9619), .ZN(n9621) );
  OAI211_X1 U10862 ( .C1(n9621), .C2(n9782), .A(n9673), .B(n9620), .ZN(n9779)
         );
  INV_X1 U10863 ( .A(n9779), .ZN(n9622) );
  AOI22_X1 U10864 ( .A1(n9785), .A2(n9677), .B1(n9676), .B2(n9622), .ZN(n9623)
         );
  OAI211_X1 U10865 ( .C1(n9634), .C2(n9780), .A(n9624), .B(n9623), .ZN(
        P1_U3280) );
  XNOR2_X1 U10866 ( .A(n9625), .B(n9627), .ZN(n9763) );
  INV_X1 U10867 ( .A(n9626), .ZN(n9800) );
  XNOR2_X1 U10868 ( .A(n9628), .B(n9627), .ZN(n9632) );
  AOI22_X1 U10869 ( .A1(n9769), .A2(n9630), .B1(n9629), .B2(n9766), .ZN(n9631)
         );
  OAI21_X1 U10870 ( .B1(n9632), .B2(n9754), .A(n9631), .ZN(n9633) );
  AOI21_X1 U10871 ( .B1(n9763), .B2(n9800), .A(n9633), .ZN(n9760) );
  AOI222_X1 U10872 ( .A1(n9636), .A2(n9652), .B1(n9635), .B2(n9651), .C1(
        P1_REG2_REG_11__SCAN_IN), .C2(n9634), .ZN(n9642) );
  INV_X1 U10873 ( .A(n9637), .ZN(n9638) );
  OAI211_X1 U10874 ( .C1(n9759), .C2(n9639), .A(n9638), .B(n9673), .ZN(n9758)
         );
  INV_X1 U10875 ( .A(n9758), .ZN(n9640) );
  AOI22_X1 U10876 ( .A1(n9763), .A2(n9658), .B1(n9676), .B2(n9640), .ZN(n9641)
         );
  OAI211_X1 U10877 ( .C1(n9634), .C2(n9760), .A(n9642), .B(n9641), .ZN(
        P1_U3282) );
  XNOR2_X1 U10878 ( .A(n9643), .B(n4561), .ZN(n9727) );
  AOI21_X1 U10879 ( .B1(n4561), .B2(n9645), .A(n9644), .ZN(n9648) );
  AOI22_X1 U10880 ( .A1(n9769), .A2(n9739), .B1(n9646), .B2(n9766), .ZN(n9647)
         );
  OAI21_X1 U10881 ( .B1(n9648), .B2(n9754), .A(n9647), .ZN(n9649) );
  AOI21_X1 U10882 ( .B1(n9800), .B2(n9727), .A(n9649), .ZN(n9724) );
  AOI222_X1 U10883 ( .A1(n9653), .A2(n9652), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9634), .C1(n9651), .C2(n9650), .ZN(n9660) );
  INV_X1 U10884 ( .A(n9655), .ZN(n9656) );
  OAI211_X1 U10885 ( .C1(n9723), .C2(n4662), .A(n9656), .B(n9673), .ZN(n9722)
         );
  INV_X1 U10886 ( .A(n9722), .ZN(n9657) );
  AOI22_X1 U10887 ( .A1(n9727), .A2(n9658), .B1(n9676), .B2(n9657), .ZN(n9659)
         );
  OAI211_X1 U10888 ( .C1(n9666), .C2(n9724), .A(n9660), .B(n9659), .ZN(
        P1_U3286) );
  XNOR2_X1 U10889 ( .A(n9661), .B(n9670), .ZN(n9663) );
  AOI222_X1 U10890 ( .A1(n9777), .A2(n9663), .B1(n9662), .B2(n9769), .C1(n5779), .C2(n9766), .ZN(n9699) );
  NOR2_X1 U10891 ( .A1(n9664), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9665) );
  AOI21_X1 U10892 ( .B1(n9666), .B2(P1_REG2_REG_3__SCAN_IN), .A(n9665), .ZN(
        n9667) );
  OAI21_X1 U10893 ( .B1(n9668), .B2(n9698), .A(n9667), .ZN(n9669) );
  INV_X1 U10894 ( .A(n9669), .ZN(n9679) );
  XNOR2_X1 U10895 ( .A(n9671), .B(n9670), .ZN(n9702) );
  OAI211_X1 U10896 ( .C1(n9674), .C2(n9698), .A(n9673), .B(n9672), .ZN(n9697)
         );
  INV_X1 U10897 ( .A(n9697), .ZN(n9675) );
  AOI22_X1 U10898 ( .A1(n9702), .A2(n9677), .B1(n9676), .B2(n9675), .ZN(n9678)
         );
  OAI211_X1 U10899 ( .C1(n9634), .C2(n9699), .A(n9679), .B(n9678), .ZN(
        P1_U3290) );
  AND2_X1 U10900 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9680), .ZN(P1_U3294) );
  INV_X1 U10901 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U10902 ( .A1(n9681), .A2(n10225), .ZN(P1_U3295) );
  AND2_X1 U10903 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9680), .ZN(P1_U3296) );
  INV_X1 U10904 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10348) );
  NOR2_X1 U10905 ( .A1(n9681), .A2(n10348), .ZN(P1_U3297) );
  AND2_X1 U10906 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9680), .ZN(P1_U3298) );
  AND2_X1 U10907 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9680), .ZN(P1_U3299) );
  AND2_X1 U10908 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9680), .ZN(P1_U3300) );
  AND2_X1 U10909 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9680), .ZN(P1_U3301) );
  AND2_X1 U10910 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9680), .ZN(P1_U3302) );
  INV_X1 U10911 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10264) );
  NOR2_X1 U10912 ( .A1(n9681), .A2(n10264), .ZN(P1_U3303) );
  AND2_X1 U10913 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9680), .ZN(P1_U3304) );
  AND2_X1 U10914 ( .A1(n9680), .A2(P1_D_REG_20__SCAN_IN), .ZN(P1_U3305) );
  INV_X1 U10915 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10302) );
  NOR2_X1 U10916 ( .A1(n9681), .A2(n10302), .ZN(P1_U3306) );
  AND2_X1 U10917 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9680), .ZN(P1_U3307) );
  AND2_X1 U10918 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9680), .ZN(P1_U3308) );
  AND2_X1 U10919 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9680), .ZN(P1_U3309) );
  INV_X1 U10920 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10294) );
  NOR2_X1 U10921 ( .A1(n9681), .A2(n10294), .ZN(P1_U3310) );
  INV_X1 U10922 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10394) );
  NOR2_X1 U10923 ( .A1(n9681), .A2(n10394), .ZN(P1_U3311) );
  AND2_X1 U10924 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9680), .ZN(P1_U3312) );
  AND2_X1 U10925 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9680), .ZN(P1_U3313) );
  AND2_X1 U10926 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9680), .ZN(P1_U3314) );
  AND2_X1 U10927 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9680), .ZN(P1_U3315) );
  AND2_X1 U10928 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9680), .ZN(P1_U3316) );
  INV_X1 U10929 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10395) );
  NOR2_X1 U10930 ( .A1(n9681), .A2(n10395), .ZN(P1_U3317) );
  AND2_X1 U10931 ( .A1(n9680), .A2(P1_D_REG_7__SCAN_IN), .ZN(P1_U3318) );
  AND2_X1 U10932 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9680), .ZN(P1_U3319) );
  INV_X1 U10933 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10330) );
  NOR2_X1 U10934 ( .A1(n9681), .A2(n10330), .ZN(P1_U3320) );
  AND2_X1 U10935 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9680), .ZN(P1_U3321) );
  AND2_X1 U10936 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9680), .ZN(P1_U3322) );
  INV_X1 U10937 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10207) );
  NOR2_X1 U10938 ( .A1(n9681), .A2(n10207), .ZN(P1_U3323) );
  NAND2_X1 U10939 ( .A1(n9772), .A2(n9754), .ZN(n9685) );
  AOI222_X1 U10940 ( .A1(n9685), .A2(n9684), .B1(n9683), .B2(n9682), .C1(n6884), .C2(n9769), .ZN(n9803) );
  INV_X1 U10941 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9686) );
  AOI22_X1 U10942 ( .A1(n9802), .A2(n9803), .B1(n9686), .B2(n9801), .ZN(
        P1_U3453) );
  INV_X1 U10943 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9687) );
  AOI22_X1 U10944 ( .A1(n9802), .A2(n9688), .B1(n9687), .B2(n9801), .ZN(
        P1_U3456) );
  INV_X1 U10945 ( .A(n9689), .ZN(n9690) );
  OAI21_X1 U10946 ( .B1(n9691), .B2(n9781), .A(n9690), .ZN(n9694) );
  INV_X1 U10947 ( .A(n9692), .ZN(n9693) );
  AOI211_X1 U10948 ( .C1(n9784), .C2(n9695), .A(n9694), .B(n9693), .ZN(n9805)
         );
  INV_X1 U10949 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9696) );
  AOI22_X1 U10950 ( .A1(n9802), .A2(n9805), .B1(n9696), .B2(n9801), .ZN(
        P1_U3459) );
  OAI21_X1 U10951 ( .B1(n9698), .B2(n9781), .A(n9697), .ZN(n9701) );
  INV_X1 U10952 ( .A(n9699), .ZN(n9700) );
  AOI211_X1 U10953 ( .C1(n9784), .C2(n9702), .A(n9701), .B(n9700), .ZN(n9807)
         );
  INV_X1 U10954 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9703) );
  AOI22_X1 U10955 ( .A1(n9802), .A2(n9807), .B1(n9703), .B2(n9801), .ZN(
        P1_U3462) );
  OAI21_X1 U10956 ( .B1(n9705), .B2(n9781), .A(n9704), .ZN(n9706) );
  AOI21_X1 U10957 ( .B1(n9707), .B2(n9784), .A(n9706), .ZN(n9708) );
  AND2_X1 U10958 ( .A1(n9709), .A2(n9708), .ZN(n9808) );
  INV_X1 U10959 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9710) );
  AOI22_X1 U10960 ( .A1(n9802), .A2(n9808), .B1(n9710), .B2(n9801), .ZN(
        P1_U3465) );
  OAI211_X1 U10961 ( .C1(n9713), .C2(n9781), .A(n9712), .B(n9711), .ZN(n9714)
         );
  AOI21_X1 U10962 ( .B1(n9784), .B2(n9715), .A(n9714), .ZN(n9809) );
  INV_X1 U10963 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9716) );
  AOI22_X1 U10964 ( .A1(n9802), .A2(n9809), .B1(n9716), .B2(n9801), .ZN(
        P1_U3468) );
  OAI21_X1 U10965 ( .B1(n4789), .B2(n9781), .A(n9717), .ZN(n9719) );
  AOI211_X1 U10966 ( .C1(n9784), .C2(n9720), .A(n9719), .B(n9718), .ZN(n9810)
         );
  INV_X1 U10967 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9721) );
  AOI22_X1 U10968 ( .A1(n9802), .A2(n9810), .B1(n9721), .B2(n9801), .ZN(
        P1_U3471) );
  OAI21_X1 U10969 ( .B1(n9723), .B2(n9781), .A(n9722), .ZN(n9726) );
  INV_X1 U10970 ( .A(n9724), .ZN(n9725) );
  AOI211_X1 U10971 ( .C1(n9764), .C2(n9727), .A(n9726), .B(n9725), .ZN(n9812)
         );
  INV_X1 U10972 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9728) );
  AOI22_X1 U10973 ( .A1(n9802), .A2(n9812), .B1(n9728), .B2(n9801), .ZN(
        P1_U3474) );
  OAI22_X1 U10974 ( .A1(n9747), .A2(n9789), .B1(n9729), .B2(n9787), .ZN(n9731)
         );
  AOI211_X1 U10975 ( .C1(n9344), .C2(n9732), .A(n9731), .B(n9730), .ZN(n9734)
         );
  OAI211_X1 U10976 ( .C1(n9735), .C2(n9796), .A(n9734), .B(n9733), .ZN(n9736)
         );
  AOI21_X1 U10977 ( .B1(n9800), .B2(n9737), .A(n9736), .ZN(n9813) );
  INV_X1 U10978 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9738) );
  AOI22_X1 U10979 ( .A1(n9802), .A2(n9813), .B1(n9738), .B2(n9801), .ZN(
        P1_U3477) );
  AOI22_X1 U10980 ( .A1(n9740), .A2(n9344), .B1(n9766), .B2(n9739), .ZN(n9741)
         );
  OAI211_X1 U10981 ( .C1(n9743), .C2(n9772), .A(n9742), .B(n9741), .ZN(n9744)
         );
  AOI21_X1 U10982 ( .B1(n9777), .B2(n9745), .A(n9744), .ZN(n9815) );
  INV_X1 U10983 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9746) );
  AOI22_X1 U10984 ( .A1(n9802), .A2(n9815), .B1(n9746), .B2(n9801), .ZN(
        P1_U3480) );
  OAI22_X1 U10985 ( .A1(n9748), .A2(n9789), .B1(n9747), .B2(n9787), .ZN(n9750)
         );
  AOI211_X1 U10986 ( .C1(n9344), .C2(n9751), .A(n9750), .B(n9749), .ZN(n9752)
         );
  OAI21_X1 U10987 ( .B1(n9754), .B2(n9753), .A(n9752), .ZN(n9755) );
  AOI21_X1 U10988 ( .B1(n9756), .B2(n9784), .A(n9755), .ZN(n9817) );
  INV_X1 U10989 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9757) );
  AOI22_X1 U10990 ( .A1(n9802), .A2(n9817), .B1(n9757), .B2(n9801), .ZN(
        P1_U3483) );
  OAI21_X1 U10991 ( .B1(n9759), .B2(n9781), .A(n9758), .ZN(n9762) );
  INV_X1 U10992 ( .A(n9760), .ZN(n9761) );
  AOI211_X1 U10993 ( .C1(n9764), .C2(n9763), .A(n9762), .B(n9761), .ZN(n9818)
         );
  INV_X1 U10994 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9765) );
  AOI22_X1 U10995 ( .A1(n9802), .A2(n9818), .B1(n9765), .B2(n9801), .ZN(
        P1_U3486) );
  AOI22_X1 U10996 ( .A1(n9769), .A2(n9768), .B1(n9767), .B2(n9766), .ZN(n9770)
         );
  OAI211_X1 U10997 ( .C1(n4820), .C2(n9781), .A(n9771), .B(n9770), .ZN(n9775)
         );
  NOR2_X1 U10998 ( .A1(n9773), .A2(n9772), .ZN(n9774) );
  AOI211_X1 U10999 ( .C1(n9777), .C2(n9776), .A(n9775), .B(n9774), .ZN(n9820)
         );
  INV_X1 U11000 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U11001 ( .A1(n9802), .A2(n9820), .B1(n9778), .B2(n9801), .ZN(
        P1_U3489) );
  OAI211_X1 U11002 ( .C1(n9782), .C2(n9781), .A(n9780), .B(n9779), .ZN(n9783)
         );
  AOI21_X1 U11003 ( .B1(n9785), .B2(n9784), .A(n9783), .ZN(n9822) );
  INV_X1 U11004 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9786) );
  AOI22_X1 U11005 ( .A1(n9802), .A2(n9822), .B1(n9786), .B2(n9801), .ZN(
        P1_U3492) );
  INV_X1 U11006 ( .A(n9797), .ZN(n9799) );
  OAI22_X1 U11007 ( .A1(n9790), .A2(n9789), .B1(n9788), .B2(n9787), .ZN(n9792)
         );
  AOI211_X1 U11008 ( .C1(n9344), .C2(n9793), .A(n9792), .B(n9791), .ZN(n9795)
         );
  OAI211_X1 U11009 ( .C1(n9797), .C2(n9796), .A(n9795), .B(n9794), .ZN(n9798)
         );
  AOI21_X1 U11010 ( .B1(n9800), .B2(n9799), .A(n9798), .ZN(n9824) );
  INV_X1 U11011 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U11012 ( .A1(n9802), .A2(n9824), .B1(n10212), .B2(n9801), .ZN(
        P1_U3495) );
  AOI22_X1 U11013 ( .A1(n9825), .A2(n9803), .B1(n5770), .B2(n9823), .ZN(
        P1_U3522) );
  AOI22_X1 U11014 ( .A1(n9825), .A2(n9805), .B1(n9804), .B2(n9823), .ZN(
        P1_U3524) );
  INV_X1 U11015 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9806) );
  AOI22_X1 U11016 ( .A1(n9825), .A2(n9807), .B1(n9806), .B2(n9823), .ZN(
        P1_U3525) );
  INV_X1 U11017 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U11018 ( .A1(n9825), .A2(n9808), .B1(n10223), .B2(n9823), .ZN(
        P1_U3526) );
  AOI22_X1 U11019 ( .A1(n9825), .A2(n9809), .B1(n7081), .B2(n9823), .ZN(
        P1_U3527) );
  AOI22_X1 U11020 ( .A1(n9825), .A2(n9810), .B1(n7083), .B2(n9823), .ZN(
        P1_U3528) );
  INV_X1 U11021 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9811) );
  AOI22_X1 U11022 ( .A1(n9825), .A2(n9812), .B1(n9811), .B2(n9823), .ZN(
        P1_U3529) );
  INV_X1 U11023 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U11024 ( .A1(n9825), .A2(n9813), .B1(n10182), .B2(n9823), .ZN(
        P1_U3530) );
  INV_X1 U11025 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9814) );
  AOI22_X1 U11026 ( .A1(n9825), .A2(n9815), .B1(n9814), .B2(n9823), .ZN(
        P1_U3531) );
  INV_X1 U11027 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9816) );
  AOI22_X1 U11028 ( .A1(n9825), .A2(n9817), .B1(n9816), .B2(n9823), .ZN(
        P1_U3532) );
  AOI22_X1 U11029 ( .A1(n9825), .A2(n9818), .B1(n7091), .B2(n9823), .ZN(
        P1_U3533) );
  AOI22_X1 U11030 ( .A1(n9825), .A2(n9820), .B1(n9819), .B2(n9823), .ZN(
        P1_U3534) );
  AOI22_X1 U11031 ( .A1(n9825), .A2(n9822), .B1(n9821), .B2(n9823), .ZN(
        P1_U3535) );
  AOI22_X1 U11032 ( .A1(n9825), .A2(n9824), .B1(n10397), .B2(n9823), .ZN(
        P1_U3536) );
  INV_X1 U11033 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10084) );
  OR2_X1 U11034 ( .A1(n9897), .A2(n10084), .ZN(n9836) );
  XNOR2_X1 U11035 ( .A(n9826), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n9827) );
  NAND2_X1 U11036 ( .A1(n9974), .A2(n9827), .ZN(n9835) );
  NAND2_X1 U11037 ( .A1(n9828), .A2(n7189), .ZN(n9829) );
  AND2_X1 U11038 ( .A1(n9830), .A2(n9829), .ZN(n9831) );
  OR2_X1 U11039 ( .A1(n9980), .A2(n9831), .ZN(n9834) );
  NAND2_X1 U11040 ( .A1(n9964), .A2(n9832), .ZN(n9833) );
  AND4_X1 U11041 ( .A1(n9836), .A2(n9835), .A3(n9834), .A4(n9833), .ZN(n9841)
         );
  XOR2_X1 U11042 ( .A(n9838), .B(n9837), .Z(n9839) );
  NAND2_X1 U11043 ( .A1(n9973), .A2(n9839), .ZN(n9840) );
  OAI211_X1 U11044 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7183), .A(n9841), .B(
        n9840), .ZN(P2_U3183) );
  INV_X1 U11045 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9858) );
  OAI21_X1 U11046 ( .B1(n9842), .B2(P2_REG2_REG_3__SCAN_IN), .A(n9868), .ZN(
        n9843) );
  INV_X1 U11047 ( .A(n9843), .ZN(n9850) );
  XNOR2_X1 U11048 ( .A(n9844), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n9845) );
  NAND2_X1 U11049 ( .A1(n9974), .A2(n9845), .ZN(n9849) );
  AOI21_X1 U11050 ( .B1(n9964), .B2(n9847), .A(n9846), .ZN(n9848) );
  OAI211_X1 U11051 ( .C1(n9850), .C2(n9980), .A(n9849), .B(n9848), .ZN(n9851)
         );
  INV_X1 U11052 ( .A(n9851), .ZN(n9857) );
  OAI21_X1 U11053 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n9855) );
  NAND2_X1 U11054 ( .A1(n9855), .A2(n9973), .ZN(n9856) );
  OAI211_X1 U11055 ( .C1(n9858), .C2(n9897), .A(n9857), .B(n9856), .ZN(
        P2_U3185) );
  OAI21_X1 U11056 ( .B1(n9861), .B2(n9860), .A(n9859), .ZN(n9873) );
  OAI21_X1 U11057 ( .B1(n9864), .B2(n9863), .A(n9862), .ZN(n9872) );
  INV_X1 U11058 ( .A(n9865), .ZN(n9867) );
  NAND3_X1 U11059 ( .A1(n9868), .A2(n9867), .A3(n9866), .ZN(n9869) );
  AOI21_X1 U11060 ( .B1(n9870), .B2(n9869), .A(n9980), .ZN(n9871) );
  AOI211_X1 U11061 ( .C1(n9974), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9880)
         );
  AOI211_X1 U11062 ( .C1(n9877), .C2(n9876), .A(n9875), .B(n9874), .ZN(n9878)
         );
  INV_X1 U11063 ( .A(n9878), .ZN(n9879) );
  OAI211_X1 U11064 ( .C1(n9881), .C2(n9897), .A(n9880), .B(n9879), .ZN(
        P2_U3186) );
  OAI21_X1 U11065 ( .B1(n9883), .B2(P2_REG2_REG_5__SCAN_IN), .A(n9882), .ZN(
        n9884) );
  INV_X1 U11066 ( .A(n9884), .ZN(n9891) );
  XNOR2_X1 U11067 ( .A(n9885), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n9886) );
  NAND2_X1 U11068 ( .A1(n9974), .A2(n9886), .ZN(n9890) );
  AOI21_X1 U11069 ( .B1(n9964), .B2(n9888), .A(n9887), .ZN(n9889) );
  OAI211_X1 U11070 ( .C1(n9891), .C2(n9980), .A(n9890), .B(n9889), .ZN(n9892)
         );
  INV_X1 U11071 ( .A(n9892), .ZN(n9896) );
  XOR2_X1 U11072 ( .A(n9893), .B(n4595), .Z(n9894) );
  NAND2_X1 U11073 ( .A1(n9894), .A2(n9973), .ZN(n9895) );
  OAI211_X1 U11074 ( .C1(n9898), .C2(n9897), .A(n9896), .B(n9895), .ZN(
        P2_U3187) );
  AOI22_X1 U11075 ( .A1(n9966), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(n9899), .B2(
        n9964), .ZN(n9913) );
  OAI21_X1 U11076 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9901), .A(n9900), .ZN(
        n9906) );
  OAI21_X1 U11077 ( .B1(n9904), .B2(n9903), .A(n9902), .ZN(n9905) );
  AOI22_X1 U11078 ( .A1(n9906), .A2(n9974), .B1(n9973), .B2(n9905), .ZN(n9912)
         );
  AOI21_X1 U11079 ( .B1(n9908), .B2(n6266), .A(n9907), .ZN(n9909) );
  OR2_X1 U11080 ( .A1(n9909), .A2(n9980), .ZN(n9910) );
  NAND4_X1 U11081 ( .A1(n9913), .A2(n9912), .A3(n9911), .A4(n9910), .ZN(
        P2_U3195) );
  AOI22_X1 U11082 ( .A1(n9966), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(n9914), .B2(
        n9964), .ZN(n9930) );
  OAI21_X1 U11083 ( .B1(n9917), .B2(n9916), .A(n9915), .ZN(n9922) );
  OAI21_X1 U11084 ( .B1(n9920), .B2(n9919), .A(n9918), .ZN(n9921) );
  AOI22_X1 U11085 ( .A1(n9922), .A2(n9974), .B1(n9973), .B2(n9921), .ZN(n9929)
         );
  NAND2_X1 U11086 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n9928) );
  AOI21_X1 U11087 ( .B1(n9925), .B2(n9924), .A(n9923), .ZN(n9926) );
  OR2_X1 U11088 ( .A1(n9926), .A2(n9980), .ZN(n9927) );
  NAND4_X1 U11089 ( .A1(n9930), .A2(n9929), .A3(n9928), .A4(n9927), .ZN(
        P2_U3196) );
  AOI22_X1 U11090 ( .A1(n9966), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(n9931), .B2(
        n9964), .ZN(n9946) );
  OAI21_X1 U11091 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n9933), .A(n9932), .ZN(
        n9938) );
  OAI21_X1 U11092 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(n9937) );
  AOI22_X1 U11093 ( .A1(n9938), .A2(n9974), .B1(n9973), .B2(n9937), .ZN(n9945)
         );
  AOI21_X1 U11094 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(n9942) );
  OR2_X1 U11095 ( .A1(n9980), .A2(n9942), .ZN(n9943) );
  NAND4_X1 U11096 ( .A1(n9946), .A2(n9945), .A3(n9944), .A4(n9943), .ZN(
        P2_U3197) );
  AOI22_X1 U11097 ( .A1(n9966), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(n9947), .B2(
        n9964), .ZN(n9963) );
  OAI21_X1 U11098 ( .B1(n9950), .B2(n9949), .A(n9948), .ZN(n9955) );
  OAI21_X1 U11099 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n9954) );
  AOI22_X1 U11100 ( .A1(n9955), .A2(n9974), .B1(n9973), .B2(n9954), .ZN(n9962)
         );
  AOI21_X1 U11101 ( .B1(n9958), .B2(n9957), .A(n9956), .ZN(n9959) );
  OR2_X1 U11102 ( .A1(n9959), .A2(n9980), .ZN(n9960) );
  NAND4_X1 U11103 ( .A1(n9963), .A2(n9962), .A3(n9961), .A4(n9960), .ZN(
        P2_U3198) );
  AOI22_X1 U11104 ( .A1(n9966), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(n9965), .B2(
        n9964), .ZN(n9984) );
  OAI21_X1 U11105 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9968), .A(n9967), .ZN(
        n9975) );
  OAI21_X1 U11106 ( .B1(n9971), .B2(n9970), .A(n9969), .ZN(n9972) );
  AOI22_X1 U11107 ( .A1(n9975), .A2(n9974), .B1(n9973), .B2(n9972), .ZN(n9983)
         );
  NAND2_X1 U11108 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n9982) );
  AOI21_X1 U11109 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(n9979) );
  OR2_X1 U11110 ( .A1(n9980), .A2(n9979), .ZN(n9981) );
  NAND4_X1 U11111 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n9981), .ZN(
        P2_U3199) );
  OAI21_X1 U11112 ( .B1(n9986), .B2(n9990), .A(n9985), .ZN(n10016) );
  OAI22_X1 U11113 ( .A1(n9989), .A2(n9988), .B1(n10013), .B2(n9987), .ZN(
        n10001) );
  XNOR2_X1 U11114 ( .A(n9991), .B(n9990), .ZN(n9999) );
  INV_X1 U11115 ( .A(n9992), .ZN(n10012) );
  OAI22_X1 U11116 ( .A1(n9996), .A2(n9995), .B1(n9994), .B2(n9993), .ZN(n9997)
         );
  AOI21_X1 U11117 ( .B1(n10016), .B2(n10012), .A(n9997), .ZN(n9998) );
  OAI21_X1 U11118 ( .B1(n10000), .B2(n9999), .A(n9998), .ZN(n10014) );
  AOI211_X1 U11119 ( .C1(n10002), .C2(n10016), .A(n10001), .B(n10014), .ZN(
        n10003) );
  AOI22_X1 U11120 ( .A1(n10005), .A2(n10004), .B1(n10003), .B2(n4500), .ZN(
        P2_U3231) );
  INV_X1 U11121 ( .A(n10046), .ZN(n10017) );
  NAND2_X1 U11122 ( .A1(n10011), .A2(n10017), .ZN(n10006) );
  OAI21_X1 U11123 ( .B1(n10007), .B2(n10057), .A(n10006), .ZN(n10010) );
  INV_X1 U11124 ( .A(n10008), .ZN(n10009) );
  AOI211_X1 U11125 ( .C1(n10012), .C2(n10011), .A(n10010), .B(n10009), .ZN(
        n10066) );
  AOI22_X1 U11126 ( .A1(n10065), .A2(n6085), .B1(n10066), .B2(n10063), .ZN(
        P2_U3393) );
  NOR2_X1 U11127 ( .A1(n10013), .A2(n10057), .ZN(n10015) );
  AOI211_X1 U11128 ( .C1(n10017), .C2(n10016), .A(n10015), .B(n10014), .ZN(
        n10067) );
  AOI22_X1 U11129 ( .A1(n10065), .A2(n6102), .B1(n10067), .B2(n10063), .ZN(
        P2_U3396) );
  OAI21_X1 U11130 ( .B1(n10019), .B2(n10057), .A(n10018), .ZN(n10020) );
  AOI21_X1 U11131 ( .B1(n10021), .B2(n10030), .A(n10020), .ZN(n10069) );
  AOI22_X1 U11132 ( .A1(n10065), .A2(n6119), .B1(n10069), .B2(n10063), .ZN(
        P2_U3399) );
  NOR2_X1 U11133 ( .A1(n10022), .A2(n10057), .ZN(n10024) );
  AOI211_X1 U11134 ( .C1(n10030), .C2(n10025), .A(n10024), .B(n10023), .ZN(
        n10070) );
  AOI22_X1 U11135 ( .A1(n10065), .A2(n6137), .B1(n10070), .B2(n10063), .ZN(
        P2_U3402) );
  OAI22_X1 U11136 ( .A1(n10027), .A2(n10046), .B1(n10026), .B2(n10057), .ZN(
        n10028) );
  NOR2_X1 U11137 ( .A1(n10029), .A2(n10028), .ZN(n10071) );
  AOI22_X1 U11138 ( .A1(n10065), .A2(n6152), .B1(n10071), .B2(n10063), .ZN(
        P2_U3405) );
  AND2_X1 U11139 ( .A1(n10031), .A2(n10030), .ZN(n10035) );
  NOR2_X1 U11140 ( .A1(n10032), .A2(n10057), .ZN(n10033) );
  NOR3_X1 U11141 ( .A1(n10035), .A2(n10034), .A3(n10033), .ZN(n10072) );
  AOI22_X1 U11142 ( .A1(n10065), .A2(n6165), .B1(n10072), .B2(n10063), .ZN(
        P2_U3408) );
  OAI22_X1 U11143 ( .A1(n10037), .A2(n10046), .B1(n10036), .B2(n10057), .ZN(
        n10038) );
  NOR2_X1 U11144 ( .A1(n10039), .A2(n10038), .ZN(n10074) );
  AOI22_X1 U11145 ( .A1(n10065), .A2(n6187), .B1(n10074), .B2(n10063), .ZN(
        P2_U3411) );
  NOR2_X1 U11146 ( .A1(n10040), .A2(n10059), .ZN(n10043) );
  INV_X1 U11147 ( .A(n10041), .ZN(n10042) );
  AOI211_X1 U11148 ( .C1(n10055), .C2(n10044), .A(n10043), .B(n10042), .ZN(
        n10075) );
  AOI22_X1 U11149 ( .A1(n10065), .A2(n6197), .B1(n10075), .B2(n10063), .ZN(
        P2_U3414) );
  INV_X1 U11150 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10050) );
  OAI22_X1 U11151 ( .A1(n10047), .A2(n10046), .B1(n10045), .B2(n10057), .ZN(
        n10048) );
  NOR2_X1 U11152 ( .A1(n10049), .A2(n10048), .ZN(n10076) );
  AOI22_X1 U11153 ( .A1(n10065), .A2(n10050), .B1(n10076), .B2(n10063), .ZN(
        P2_U3420) );
  INV_X1 U11154 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10056) );
  NOR2_X1 U11155 ( .A1(n10051), .A2(n10059), .ZN(n10053) );
  AOI211_X1 U11156 ( .C1(n10055), .C2(n10054), .A(n10053), .B(n10052), .ZN(
        n10078) );
  AOI22_X1 U11157 ( .A1(n10065), .A2(n10056), .B1(n10078), .B2(n10063), .ZN(
        P2_U3423) );
  INV_X1 U11158 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10064) );
  OAI22_X1 U11159 ( .A1(n10060), .A2(n10059), .B1(n10058), .B2(n10057), .ZN(
        n10061) );
  NOR2_X1 U11160 ( .A1(n10062), .A2(n10061), .ZN(n10080) );
  AOI22_X1 U11161 ( .A1(n10065), .A2(n10064), .B1(n10080), .B2(n10063), .ZN(
        P2_U3426) );
  INV_X1 U11162 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10220) );
  AOI22_X1 U11163 ( .A1(n10081), .A2(n10066), .B1(n10220), .B2(n10079), .ZN(
        P2_U3460) );
  AOI22_X1 U11164 ( .A1(n10081), .A2(n10067), .B1(n6804), .B2(n10079), .ZN(
        P2_U3461) );
  INV_X1 U11165 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10068) );
  AOI22_X1 U11166 ( .A1(n10081), .A2(n10069), .B1(n10068), .B2(n10079), .ZN(
        P2_U3462) );
  AOI22_X1 U11167 ( .A1(n10081), .A2(n10070), .B1(n6839), .B2(n10079), .ZN(
        P2_U3463) );
  AOI22_X1 U11168 ( .A1(n10081), .A2(n10071), .B1(n6828), .B2(n10079), .ZN(
        P2_U3464) );
  AOI22_X1 U11169 ( .A1(n10081), .A2(n10072), .B1(n6916), .B2(n10079), .ZN(
        P2_U3465) );
  INV_X1 U11170 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U11171 ( .A1(n10081), .A2(n10074), .B1(n10073), .B2(n10079), .ZN(
        P2_U3466) );
  AOI22_X1 U11172 ( .A1(n10081), .A2(n10075), .B1(n7017), .B2(n10079), .ZN(
        P2_U3467) );
  AOI22_X1 U11173 ( .A1(n10081), .A2(n10076), .B1(n7434), .B2(n10079), .ZN(
        P2_U3469) );
  INV_X1 U11174 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10077) );
  AOI22_X1 U11175 ( .A1(n10081), .A2(n10078), .B1(n10077), .B2(n10079), .ZN(
        P2_U3470) );
  AOI22_X1 U11176 ( .A1(n10081), .A2(n10080), .B1(n7614), .B2(n10079), .ZN(
        P2_U3471) );
  NOR2_X1 U11177 ( .A1(n10083), .A2(n10082), .ZN(n10085) );
  XNOR2_X1 U11178 ( .A(n10085), .B(n10084), .ZN(ADD_1068_U5) );
  XOR2_X1 U11179 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11180 ( .A1(n10087), .A2(n10086), .ZN(n10088) );
  XOR2_X1 U11181 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10088), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11182 ( .A(n10090), .B(n10089), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11183 ( .A(n10092), .B(n10091), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11184 ( .A(n10094), .B(n10093), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11185 ( .A(n10096), .B(n10095), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11186 ( .A(n10098), .B(n10097), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11187 ( .A(n10100), .B(n10099), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11188 ( .A(n10102), .B(n10101), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11189 ( .A(n10104), .B(n10103), .ZN(ADD_1068_U63) );
  NAND2_X1 U11190 ( .A1(n10105), .A2(P2_D_REG_20__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U11191 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(keyinput238), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(keyinput138), .ZN(n10106) );
  OAI221_X1 U11192 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(keyinput238), .C1(
        P2_DATAO_REG_29__SCAN_IN), .C2(keyinput138), .A(n10106), .ZN(n10113)
         );
  AOI22_X1 U11193 ( .A1(P1_REG0_REG_6__SCAN_IN), .A2(keyinput162), .B1(SI_21_), 
        .B2(keyinput158), .ZN(n10107) );
  OAI221_X1 U11194 ( .B1(P1_REG0_REG_6__SCAN_IN), .B2(keyinput162), .C1(SI_21_), .C2(keyinput158), .A(n10107), .ZN(n10112) );
  AOI22_X1 U11195 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(keyinput188), .B1(
        P1_REG1_REG_29__SCAN_IN), .B2(keyinput214), .ZN(n10108) );
  OAI221_X1 U11196 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(keyinput188), .C1(
        P1_REG1_REG_29__SCAN_IN), .C2(keyinput214), .A(n10108), .ZN(n10111) );
  AOI22_X1 U11197 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(keyinput177), .B1(
        P1_IR_REG_24__SCAN_IN), .B2(keyinput174), .ZN(n10109) );
  OAI221_X1 U11198 ( .B1(P2_IR_REG_11__SCAN_IN), .B2(keyinput177), .C1(
        P1_IR_REG_24__SCAN_IN), .C2(keyinput174), .A(n10109), .ZN(n10110) );
  NOR4_X1 U11199 ( .A1(n10113), .A2(n10112), .A3(n10111), .A4(n10110), .ZN(
        n10141) );
  AOI22_X1 U11200 ( .A1(P1_REG0_REG_9__SCAN_IN), .A2(keyinput204), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput147), .ZN(n10114) );
  OAI221_X1 U11201 ( .B1(P1_REG0_REG_9__SCAN_IN), .B2(keyinput204), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput147), .A(n10114), .ZN(n10121) );
  AOI22_X1 U11202 ( .A1(P1_REG2_REG_30__SCAN_IN), .A2(keyinput172), .B1(SI_24_), .B2(keyinput132), .ZN(n10115) );
  OAI221_X1 U11203 ( .B1(P1_REG2_REG_30__SCAN_IN), .B2(keyinput172), .C1(
        SI_24_), .C2(keyinput132), .A(n10115), .ZN(n10120) );
  AOI22_X1 U11204 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(keyinput180), .B1(
        P1_REG3_REG_25__SCAN_IN), .B2(keyinput209), .ZN(n10116) );
  OAI221_X1 U11205 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(keyinput180), .C1(
        P1_REG3_REG_25__SCAN_IN), .C2(keyinput209), .A(n10116), .ZN(n10119) );
  AOI22_X1 U11206 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(keyinput206), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(keyinput139), .ZN(n10117) );
  OAI221_X1 U11207 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(keyinput206), .C1(
        P1_DATAO_REG_11__SCAN_IN), .C2(keyinput139), .A(n10117), .ZN(n10118)
         );
  NOR4_X1 U11208 ( .A1(n10121), .A2(n10120), .A3(n10119), .A4(n10118), .ZN(
        n10140) );
  AOI22_X1 U11209 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(keyinput170), .B1(
        P2_REG1_REG_20__SCAN_IN), .B2(keyinput134), .ZN(n10122) );
  OAI221_X1 U11210 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(keyinput170), .C1(
        P2_REG1_REG_20__SCAN_IN), .C2(keyinput134), .A(n10122), .ZN(n10129) );
  AOI22_X1 U11211 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput231), .B1(
        P1_D_REG_19__SCAN_IN), .B2(keyinput240), .ZN(n10123) );
  OAI221_X1 U11212 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput231), .C1(
        P1_D_REG_19__SCAN_IN), .C2(keyinput240), .A(n10123), .ZN(n10128) );
  AOI22_X1 U11213 ( .A1(P2_D_REG_2__SCAN_IN), .A2(keyinput178), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(keyinput217), .ZN(n10124) );
  OAI221_X1 U11214 ( .B1(P2_D_REG_2__SCAN_IN), .B2(keyinput178), .C1(
        P1_DATAO_REG_2__SCAN_IN), .C2(keyinput217), .A(n10124), .ZN(n10127) );
  AOI22_X1 U11215 ( .A1(P2_REG0_REG_6__SCAN_IN), .A2(keyinput182), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(keyinput142), .ZN(n10125) );
  OAI221_X1 U11216 ( .B1(P2_REG0_REG_6__SCAN_IN), .B2(keyinput182), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput142), .A(n10125), .ZN(n10126) );
  NOR4_X1 U11217 ( .A1(n10129), .A2(n10128), .A3(n10127), .A4(n10126), .ZN(
        n10139) );
  AOI22_X1 U11218 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(keyinput168), .B1(
        P2_D_REG_3__SCAN_IN), .B2(keyinput148), .ZN(n10130) );
  OAI221_X1 U11219 ( .B1(P1_DATAO_REG_29__SCAN_IN), .B2(keyinput168), .C1(
        P2_D_REG_3__SCAN_IN), .C2(keyinput148), .A(n10130), .ZN(n10137) );
  AOI22_X1 U11220 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(keyinput159), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput153), .ZN(n10131) );
  OAI221_X1 U11221 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(keyinput159), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput153), .A(n10131), .ZN(n10136) );
  AOI22_X1 U11222 ( .A1(P2_D_REG_0__SCAN_IN), .A2(keyinput175), .B1(
        P1_REG3_REG_12__SCAN_IN), .B2(keyinput160), .ZN(n10132) );
  OAI221_X1 U11223 ( .B1(P2_D_REG_0__SCAN_IN), .B2(keyinput175), .C1(
        P1_REG3_REG_12__SCAN_IN), .C2(keyinput160), .A(n10132), .ZN(n10135) );
  AOI22_X1 U11224 ( .A1(P1_REG0_REG_2__SCAN_IN), .A2(keyinput173), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput213), .ZN(n10133) );
  OAI221_X1 U11225 ( .B1(P1_REG0_REG_2__SCAN_IN), .B2(keyinput173), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput213), .A(n10133), .ZN(n10134)
         );
  NOR4_X1 U11226 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(n10134), .ZN(
        n10138) );
  NAND4_X1 U11227 ( .A1(n10141), .A2(n10140), .A3(n10139), .A4(n10138), .ZN(
        n10289) );
  AOI22_X1 U11228 ( .A1(P1_REG1_REG_26__SCAN_IN), .A2(keyinput254), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput247), .ZN(n10142) );
  OAI221_X1 U11229 ( .B1(P1_REG1_REG_26__SCAN_IN), .B2(keyinput254), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput247), .A(n10142), .ZN(n10149) );
  AOI22_X1 U11230 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput157), .B1(
        P1_D_REG_28__SCAN_IN), .B2(keyinput232), .ZN(n10143) );
  OAI221_X1 U11231 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput157), .C1(
        P1_D_REG_28__SCAN_IN), .C2(keyinput232), .A(n10143), .ZN(n10148) );
  AOI22_X1 U11232 ( .A1(P2_REG0_REG_8__SCAN_IN), .A2(keyinput143), .B1(
        P2_REG2_REG_16__SCAN_IN), .B2(keyinput197), .ZN(n10144) );
  OAI221_X1 U11233 ( .B1(P2_REG0_REG_8__SCAN_IN), .B2(keyinput143), .C1(
        P2_REG2_REG_16__SCAN_IN), .C2(keyinput197), .A(n10144), .ZN(n10147) );
  AOI22_X1 U11234 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(keyinput152), .B1(SI_22_), 
        .B2(keyinput215), .ZN(n10145) );
  OAI221_X1 U11235 ( .B1(P2_IR_REG_1__SCAN_IN), .B2(keyinput152), .C1(SI_22_), 
        .C2(keyinput215), .A(n10145), .ZN(n10146) );
  NOR4_X1 U11236 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10180) );
  AOI22_X1 U11237 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(keyinput140), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(keyinput130), .ZN(n10150) );
  OAI221_X1 U11238 ( .B1(P2_REG2_REG_25__SCAN_IN), .B2(keyinput140), .C1(
        P1_DATAO_REG_20__SCAN_IN), .C2(keyinput130), .A(n10150), .ZN(n10157)
         );
  AOI22_X1 U11239 ( .A1(P2_REG0_REG_2__SCAN_IN), .A2(keyinput189), .B1(
        P2_IR_REG_14__SCAN_IN), .B2(keyinput208), .ZN(n10151) );
  OAI221_X1 U11240 ( .B1(P2_REG0_REG_2__SCAN_IN), .B2(keyinput189), .C1(
        P2_IR_REG_14__SCAN_IN), .C2(keyinput208), .A(n10151), .ZN(n10156) );
  AOI22_X1 U11241 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(keyinput250), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(keyinput210), .ZN(n10152) );
  OAI221_X1 U11242 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(keyinput250), .C1(
        P1_REG3_REG_0__SCAN_IN), .C2(keyinput210), .A(n10152), .ZN(n10155) );
  AOI22_X1 U11243 ( .A1(P2_REG0_REG_31__SCAN_IN), .A2(keyinput227), .B1(
        P2_D_REG_8__SCAN_IN), .B2(keyinput233), .ZN(n10153) );
  OAI221_X1 U11244 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(keyinput227), .C1(
        P2_D_REG_8__SCAN_IN), .C2(keyinput233), .A(n10153), .ZN(n10154) );
  NOR4_X1 U11245 ( .A1(n10157), .A2(n10156), .A3(n10155), .A4(n10154), .ZN(
        n10179) );
  AOI22_X1 U11246 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(keyinput219), .B1(
        P1_REG0_REG_18__SCAN_IN), .B2(keyinput164), .ZN(n10158) );
  OAI221_X1 U11247 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(keyinput219), .C1(
        P1_REG0_REG_18__SCAN_IN), .C2(keyinput164), .A(n10158), .ZN(n10165) );
  AOI22_X1 U11248 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(keyinput145), .B1(
        P1_D_REG_7__SCAN_IN), .B2(keyinput165), .ZN(n10159) );
  OAI221_X1 U11249 ( .B1(P1_REG3_REG_13__SCAN_IN), .B2(keyinput145), .C1(
        P1_D_REG_7__SCAN_IN), .C2(keyinput165), .A(n10159), .ZN(n10164) );
  AOI22_X1 U11250 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput202), .B1(
        P1_REG2_REG_22__SCAN_IN), .B2(keyinput196), .ZN(n10160) );
  OAI221_X1 U11251 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput202), .C1(
        P1_REG2_REG_22__SCAN_IN), .C2(keyinput196), .A(n10160), .ZN(n10163) );
  AOI22_X1 U11252 ( .A1(P1_REG0_REG_7__SCAN_IN), .A2(keyinput185), .B1(
        P1_REG1_REG_20__SCAN_IN), .B2(keyinput251), .ZN(n10161) );
  OAI221_X1 U11253 ( .B1(P1_REG0_REG_7__SCAN_IN), .B2(keyinput185), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput251), .A(n10161), .ZN(n10162) );
  NOR4_X1 U11254 ( .A1(n10165), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        n10178) );
  AOI22_X1 U11255 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(keyinput226), .B1(
        P1_REG3_REG_8__SCAN_IN), .B2(keyinput198), .ZN(n10166) );
  OAI221_X1 U11256 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(keyinput226), .C1(
        P1_REG3_REG_8__SCAN_IN), .C2(keyinput198), .A(n10166), .ZN(n10176) );
  AOI22_X1 U11257 ( .A1(P1_D_REG_20__SCAN_IN), .A2(keyinput163), .B1(n10168), 
        .B2(keyinput141), .ZN(n10167) );
  OAI221_X1 U11258 ( .B1(P1_D_REG_20__SCAN_IN), .B2(keyinput163), .C1(n10168), 
        .C2(keyinput141), .A(n10167), .ZN(n10175) );
  INV_X1 U11259 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U11260 ( .A1(n10171), .A2(keyinput192), .B1(keyinput245), .B2(
        n10170), .ZN(n10169) );
  OAI221_X1 U11261 ( .B1(n10171), .B2(keyinput192), .C1(n10170), .C2(
        keyinput245), .A(n10169), .ZN(n10174) );
  INV_X1 U11262 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U11263 ( .A1(n10353), .A2(keyinput137), .B1(n10366), .B2(
        keyinput225), .ZN(n10172) );
  OAI221_X1 U11264 ( .B1(n10353), .B2(keyinput137), .C1(n10366), .C2(
        keyinput225), .A(n10172), .ZN(n10173) );
  NOR4_X1 U11265 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10177) );
  NAND4_X1 U11266 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10288) );
  INV_X1 U11267 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U11268 ( .A1(n10305), .A2(keyinput195), .B1(keyinput167), .B2(
        n10182), .ZN(n10181) );
  OAI221_X1 U11269 ( .B1(n10305), .B2(keyinput195), .C1(n10182), .C2(
        keyinput167), .A(n10181), .ZN(n10194) );
  AOI22_X1 U11270 ( .A1(n6121), .A2(keyinput150), .B1(n10184), .B2(keyinput154), .ZN(n10183) );
  OAI221_X1 U11271 ( .B1(n6121), .B2(keyinput150), .C1(n10184), .C2(
        keyinput154), .A(n10183), .ZN(n10193) );
  AOI22_X1 U11272 ( .A1(n10187), .A2(keyinput183), .B1(n10186), .B2(
        keyinput135), .ZN(n10185) );
  OAI221_X1 U11273 ( .B1(n10187), .B2(keyinput183), .C1(n10186), .C2(
        keyinput135), .A(n10185), .ZN(n10192) );
  XOR2_X1 U11274 ( .A(n10188), .B(keyinput156), .Z(n10190) );
  XNOR2_X1 U11275 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput224), .ZN(n10189)
         );
  NAND2_X1 U11276 ( .A1(n10190), .A2(n10189), .ZN(n10191) );
  NOR4_X1 U11277 ( .A1(n10194), .A2(n10193), .A3(n10192), .A4(n10191), .ZN(
        n10235) );
  AOI22_X1 U11278 ( .A1(n10196), .A2(keyinput190), .B1(keyinput223), .B2(
        n10315), .ZN(n10195) );
  OAI221_X1 U11279 ( .B1(n10196), .B2(keyinput190), .C1(n10315), .C2(
        keyinput223), .A(n10195), .ZN(n10205) );
  AOI22_X1 U11280 ( .A1(n10199), .A2(keyinput211), .B1(n10198), .B2(
        keyinput212), .ZN(n10197) );
  OAI221_X1 U11281 ( .B1(n10199), .B2(keyinput211), .C1(n10198), .C2(
        keyinput212), .A(n10197), .ZN(n10204) );
  AOI22_X1 U11282 ( .A1(n10335), .A2(keyinput205), .B1(n10394), .B2(
        keyinput136), .ZN(n10200) );
  OAI221_X1 U11283 ( .B1(n10335), .B2(keyinput205), .C1(n10394), .C2(
        keyinput136), .A(n10200), .ZN(n10203) );
  AOI22_X1 U11284 ( .A1(n6416), .A2(keyinput243), .B1(keyinput255), .B2(n6829), 
        .ZN(n10201) );
  OAI221_X1 U11285 ( .B1(n6416), .B2(keyinput243), .C1(n6829), .C2(keyinput255), .A(n10201), .ZN(n10202) );
  NOR4_X1 U11286 ( .A1(n10205), .A2(n10204), .A3(n10203), .A4(n10202), .ZN(
        n10234) );
  AOI22_X1 U11287 ( .A1(n10207), .A2(keyinput171), .B1(keyinput133), .B2(
        n10295), .ZN(n10206) );
  OAI221_X1 U11288 ( .B1(n10207), .B2(keyinput171), .C1(n10295), .C2(
        keyinput133), .A(n10206), .ZN(n10218) );
  AOI22_X1 U11289 ( .A1(n10304), .A2(keyinput253), .B1(keyinput241), .B2(
        n10209), .ZN(n10208) );
  OAI221_X1 U11290 ( .B1(n10304), .B2(keyinput253), .C1(n10209), .C2(
        keyinput241), .A(n10208), .ZN(n10217) );
  AOI22_X1 U11291 ( .A1(n10212), .A2(keyinput151), .B1(keyinput191), .B2(
        n10211), .ZN(n10210) );
  OAI221_X1 U11292 ( .B1(n10212), .B2(keyinput151), .C1(n10211), .C2(
        keyinput191), .A(n10210), .ZN(n10216) );
  XNOR2_X1 U11293 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput155), .ZN(n10214) );
  XNOR2_X1 U11294 ( .A(P1_REG3_REG_21__SCAN_IN), .B(keyinput242), .ZN(n10213)
         );
  NAND2_X1 U11295 ( .A1(n10214), .A2(n10213), .ZN(n10215) );
  NOR4_X1 U11296 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n10233) );
  INV_X1 U11297 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10221) );
  AOI22_X1 U11298 ( .A1(n10221), .A2(keyinput129), .B1(keyinput176), .B2(
        n10220), .ZN(n10219) );
  OAI221_X1 U11299 ( .B1(n10221), .B2(keyinput129), .C1(n10220), .C2(
        keyinput176), .A(n10219), .ZN(n10231) );
  INV_X1 U11300 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U11301 ( .A1(n10382), .A2(keyinput201), .B1(keyinput235), .B2(
        n10223), .ZN(n10222) );
  OAI221_X1 U11302 ( .B1(n10382), .B2(keyinput201), .C1(n10223), .C2(
        keyinput235), .A(n10222), .ZN(n10230) );
  AOI22_X1 U11303 ( .A1(n10225), .A2(keyinput229), .B1(keyinput166), .B2(
        n10378), .ZN(n10224) );
  OAI221_X1 U11304 ( .B1(n10225), .B2(keyinput229), .C1(n10378), .C2(
        keyinput166), .A(n10224), .ZN(n10229) );
  XNOR2_X1 U11305 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput246), .ZN(n10227) );
  XNOR2_X1 U11306 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput146), .ZN(n10226) );
  NAND2_X1 U11307 ( .A1(n10227), .A2(n10226), .ZN(n10228) );
  NOR4_X1 U11308 ( .A1(n10231), .A2(n10230), .A3(n10229), .A4(n10228), .ZN(
        n10232) );
  NAND4_X1 U11309 ( .A1(n10235), .A2(n10234), .A3(n10233), .A4(n10232), .ZN(
        n10287) );
  AOI22_X1 U11310 ( .A1(n10369), .A2(keyinput169), .B1(keyinput128), .B2(
        n10237), .ZN(n10236) );
  OAI221_X1 U11311 ( .B1(n10369), .B2(keyinput169), .C1(n10237), .C2(
        keyinput128), .A(n10236), .ZN(n10248) );
  INV_X1 U11312 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U11313 ( .A1(n10240), .A2(keyinput193), .B1(keyinput228), .B2(
        n10239), .ZN(n10238) );
  OAI221_X1 U11314 ( .B1(n10240), .B2(keyinput193), .C1(n10239), .C2(
        keyinput228), .A(n10238), .ZN(n10247) );
  AOI22_X1 U11315 ( .A1(n10242), .A2(keyinput187), .B1(keyinput248), .B2(n6725), .ZN(n10241) );
  OAI221_X1 U11316 ( .B1(n10242), .B2(keyinput187), .C1(n6725), .C2(
        keyinput248), .A(n10241), .ZN(n10246) );
  XNOR2_X1 U11317 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput161), .ZN(n10244) );
  XNOR2_X1 U11318 ( .A(SI_7_), .B(keyinput184), .ZN(n10243) );
  NAND2_X1 U11319 ( .A1(n10244), .A2(n10243), .ZN(n10245) );
  NOR4_X1 U11320 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10285) );
  INV_X1 U11321 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U11322 ( .A1(n10376), .A2(keyinput199), .B1(keyinput203), .B2(
        n10398), .ZN(n10249) );
  OAI221_X1 U11323 ( .B1(n10376), .B2(keyinput199), .C1(n10398), .C2(
        keyinput203), .A(n10249), .ZN(n10259) );
  AOI22_X1 U11324 ( .A1(n7615), .A2(keyinput249), .B1(n10251), .B2(keyinput149), .ZN(n10250) );
  OAI221_X1 U11325 ( .B1(n7615), .B2(keyinput249), .C1(n10251), .C2(
        keyinput149), .A(n10250), .ZN(n10258) );
  INV_X1 U11326 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U11327 ( .A1(n10253), .A2(keyinput207), .B1(n10390), .B2(
        keyinput220), .ZN(n10252) );
  OAI221_X1 U11328 ( .B1(n10253), .B2(keyinput207), .C1(n10390), .C2(
        keyinput220), .A(n10252), .ZN(n10257) );
  XNOR2_X1 U11329 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput216), .ZN(n10255)
         );
  XNOR2_X1 U11330 ( .A(SI_26_), .B(keyinput131), .ZN(n10254) );
  NAND2_X1 U11331 ( .A1(n10255), .A2(n10254), .ZN(n10256) );
  NOR4_X1 U11332 ( .A1(n10259), .A2(n10258), .A3(n10257), .A4(n10256), .ZN(
        n10284) );
  AOI22_X1 U11333 ( .A1(n6839), .A2(keyinput144), .B1(n10364), .B2(keyinput230), .ZN(n10260) );
  OAI221_X1 U11334 ( .B1(n6839), .B2(keyinput144), .C1(n10364), .C2(
        keyinput230), .A(n10260), .ZN(n10269) );
  AOI22_X1 U11335 ( .A1(n10392), .A2(keyinput186), .B1(n10262), .B2(
        keyinput218), .ZN(n10261) );
  OAI221_X1 U11336 ( .B1(n10392), .B2(keyinput186), .C1(n10262), .C2(
        keyinput218), .A(n10261), .ZN(n10268) );
  AOI22_X1 U11337 ( .A1(n10264), .A2(keyinput252), .B1(keyinput221), .B2(
        n10336), .ZN(n10263) );
  OAI221_X1 U11338 ( .B1(n10264), .B2(keyinput252), .C1(n10336), .C2(
        keyinput221), .A(n10263), .ZN(n10267) );
  AOI22_X1 U11339 ( .A1(n10330), .A2(keyinput239), .B1(keyinput200), .B2(
        n10397), .ZN(n10265) );
  OAI221_X1 U11340 ( .B1(n10330), .B2(keyinput239), .C1(n10397), .C2(
        keyinput200), .A(n10265), .ZN(n10266) );
  NOR4_X1 U11341 ( .A1(n10269), .A2(n10268), .A3(n10267), .A4(n10266), .ZN(
        n10283) );
  AOI22_X1 U11342 ( .A1(n10294), .A2(keyinput237), .B1(keyinput194), .B2(n8290), .ZN(n10270) );
  OAI221_X1 U11343 ( .B1(n10294), .B2(keyinput237), .C1(n8290), .C2(
        keyinput194), .A(n10270), .ZN(n10281) );
  AOI22_X1 U11344 ( .A1(n10395), .A2(keyinput234), .B1(keyinput244), .B2(
        n10272), .ZN(n10271) );
  OAI221_X1 U11345 ( .B1(n10395), .B2(keyinput234), .C1(n10272), .C2(
        keyinput244), .A(n10271), .ZN(n10280) );
  AOI22_X1 U11346 ( .A1(n10275), .A2(keyinput236), .B1(n10274), .B2(
        keyinput181), .ZN(n10273) );
  OAI221_X1 U11347 ( .B1(n10275), .B2(keyinput236), .C1(n10274), .C2(
        keyinput181), .A(n10273), .ZN(n10279) );
  INV_X1 U11348 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U11349 ( .A1(n10277), .A2(keyinput179), .B1(keyinput222), .B2(n6828), .ZN(n10276) );
  OAI221_X1 U11350 ( .B1(n10277), .B2(keyinput179), .C1(n6828), .C2(
        keyinput222), .A(n10276), .ZN(n10278) );
  NOR4_X1 U11351 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10282) );
  NAND4_X1 U11352 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10286) );
  NOR4_X1 U11353 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        n10484) );
  AOI22_X1 U11354 ( .A1(P2_D_REG_23__SCAN_IN), .A2(keyinput0), .B1(
        P1_REG3_REG_24__SCAN_IN), .B2(keyinput64), .ZN(n10290) );
  OAI221_X1 U11355 ( .B1(P2_D_REG_23__SCAN_IN), .B2(keyinput0), .C1(
        P1_REG3_REG_24__SCAN_IN), .C2(keyinput64), .A(n10290), .ZN(n10299) );
  AOI22_X1 U11356 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(keyinput94), .B1(
        P1_REG2_REG_19__SCAN_IN), .B2(keyinput103), .ZN(n10291) );
  OAI221_X1 U11357 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(keyinput94), .C1(
        P1_REG2_REG_19__SCAN_IN), .C2(keyinput103), .A(n10291), .ZN(n10298) );
  AOI22_X1 U11358 ( .A1(P2_D_REG_3__SCAN_IN), .A2(keyinput20), .B1(
        P1_REG0_REG_24__SCAN_IN), .B2(keyinput65), .ZN(n10292) );
  OAI221_X1 U11359 ( .B1(P2_D_REG_3__SCAN_IN), .B2(keyinput20), .C1(
        P1_REG0_REG_24__SCAN_IN), .C2(keyinput65), .A(n10292), .ZN(n10297) );
  AOI22_X1 U11360 ( .A1(n10295), .A2(keyinput5), .B1(n10294), .B2(keyinput109), 
        .ZN(n10293) );
  OAI221_X1 U11361 ( .B1(n10295), .B2(keyinput5), .C1(n10294), .C2(keyinput109), .A(n10293), .ZN(n10296) );
  NOR4_X1 U11362 ( .A1(n10299), .A2(n10298), .A3(n10297), .A4(n10296), .ZN(
        n10346) );
  AOI22_X1 U11363 ( .A1(n10302), .A2(keyinput112), .B1(keyinput40), .B2(n10301), .ZN(n10300) );
  OAI221_X1 U11364 ( .B1(n10302), .B2(keyinput112), .C1(n10301), .C2(
        keyinput40), .A(n10300), .ZN(n10312) );
  AOI22_X1 U11365 ( .A1(n10305), .A2(keyinput67), .B1(keyinput125), .B2(n10304), .ZN(n10303) );
  OAI221_X1 U11366 ( .B1(n10305), .B2(keyinput67), .C1(n10304), .C2(
        keyinput125), .A(n10303), .ZN(n10311) );
  XNOR2_X1 U11367 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput46), .ZN(n10309) );
  XNOR2_X1 U11368 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput96), .ZN(n10308) );
  XNOR2_X1 U11369 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput18), .ZN(n10307) );
  XNOR2_X1 U11370 ( .A(keyinput1), .B(P1_REG0_REG_16__SCAN_IN), .ZN(n10306) );
  NAND4_X1 U11371 ( .A1(n10309), .A2(n10308), .A3(n10307), .A4(n10306), .ZN(
        n10310) );
  NOR3_X1 U11372 ( .A1(n10312), .A2(n10311), .A3(n10310), .ZN(n10345) );
  AOI22_X1 U11373 ( .A1(n10315), .A2(keyinput95), .B1(n10314), .B2(keyinput114), .ZN(n10313) );
  OAI221_X1 U11374 ( .B1(n10315), .B2(keyinput95), .C1(n10314), .C2(
        keyinput114), .A(n10313), .ZN(n10328) );
  AOI22_X1 U11375 ( .A1(n10318), .A2(keyinput47), .B1(n10317), .B2(keyinput2), 
        .ZN(n10316) );
  OAI221_X1 U11376 ( .B1(n10318), .B2(keyinput47), .C1(n10317), .C2(keyinput2), 
        .A(n10316), .ZN(n10327) );
  AOI22_X1 U11377 ( .A1(n10321), .A2(keyinput81), .B1(n10320), .B2(keyinput56), 
        .ZN(n10319) );
  OAI221_X1 U11378 ( .B1(n10321), .B2(keyinput81), .C1(n10320), .C2(keyinput56), .A(n10319), .ZN(n10326) );
  XOR2_X1 U11379 ( .A(n10322), .B(keyinput110), .Z(n10324) );
  XNOR2_X1 U11380 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput49), .ZN(n10323) );
  NAND2_X1 U11381 ( .A1(n10324), .A2(n10323), .ZN(n10325) );
  NOR4_X1 U11382 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10344) );
  AOI22_X1 U11383 ( .A1(n10330), .A2(keyinput111), .B1(keyinput22), .B2(n6121), 
        .ZN(n10329) );
  OAI221_X1 U11384 ( .B1(n10330), .B2(keyinput111), .C1(n6121), .C2(keyinput22), .A(n10329), .ZN(n10342) );
  AOI22_X1 U11385 ( .A1(n10333), .A2(keyinput80), .B1(keyinput74), .B2(n10332), 
        .ZN(n10331) );
  OAI221_X1 U11386 ( .B1(n10333), .B2(keyinput80), .C1(n10332), .C2(keyinput74), .A(n10331), .ZN(n10341) );
  AOI22_X1 U11387 ( .A1(n10336), .A2(keyinput93), .B1(keyinput77), .B2(n10335), 
        .ZN(n10334) );
  OAI221_X1 U11388 ( .B1(n10336), .B2(keyinput93), .C1(n10335), .C2(keyinput77), .A(n10334), .ZN(n10340) );
  XNOR2_X1 U11389 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput25), .ZN(n10338) );
  XNOR2_X1 U11390 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput83), .ZN(n10337)
         );
  NAND2_X1 U11391 ( .A1(n10338), .A2(n10337), .ZN(n10339) );
  NOR4_X1 U11392 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10343) );
  NAND4_X1 U11393 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10483) );
  AOI22_X1 U11394 ( .A1(n10348), .A2(keyinput104), .B1(keyinput42), .B2(n7595), 
        .ZN(n10347) );
  OAI221_X1 U11395 ( .B1(n10348), .B2(keyinput104), .C1(n7595), .C2(keyinput42), .A(n10347), .ZN(n10359) );
  AOI22_X1 U11396 ( .A1(n10350), .A2(keyinput14), .B1(keyinput15), .B2(n6197), 
        .ZN(n10349) );
  OAI221_X1 U11397 ( .B1(n10350), .B2(keyinput14), .C1(n6197), .C2(keyinput15), 
        .A(n10349), .ZN(n10358) );
  AOI22_X1 U11398 ( .A1(n10353), .A2(keyinput9), .B1(n10352), .B2(keyinput6), 
        .ZN(n10351) );
  OAI221_X1 U11399 ( .B1(n10353), .B2(keyinput9), .C1(n10352), .C2(keyinput6), 
        .A(n10351), .ZN(n10357) );
  XNOR2_X1 U11400 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput27), .ZN(n10355) );
  XNOR2_X1 U11401 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(keyinput84), .ZN(n10354)
         );
  NAND2_X1 U11402 ( .A1(n10355), .A2(n10354), .ZN(n10356) );
  NOR4_X1 U11403 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n10406) );
  AOI22_X1 U11404 ( .A1(n10361), .A2(keyinput10), .B1(n5161), .B2(keyinput70), 
        .ZN(n10360) );
  OAI221_X1 U11405 ( .B1(n10361), .B2(keyinput10), .C1(n5161), .C2(keyinput70), 
        .A(n10360), .ZN(n10373) );
  AOI22_X1 U11406 ( .A1(n10364), .A2(keyinput102), .B1(n10363), .B2(keyinput11), .ZN(n10362) );
  OAI221_X1 U11407 ( .B1(n10364), .B2(keyinput102), .C1(n10363), .C2(
        keyinput11), .A(n10362), .ZN(n10372) );
  AOI22_X1 U11408 ( .A1(n10367), .A2(keyinput98), .B1(n10366), .B2(keyinput97), 
        .ZN(n10365) );
  OAI221_X1 U11409 ( .B1(n10367), .B2(keyinput98), .C1(n10366), .C2(keyinput97), .A(n10365), .ZN(n10371) );
  AOI22_X1 U11410 ( .A1(n6165), .A2(keyinput54), .B1(n10369), .B2(keyinput41), 
        .ZN(n10368) );
  OAI221_X1 U11411 ( .B1(n6165), .B2(keyinput54), .C1(n10369), .C2(keyinput41), 
        .A(n10368), .ZN(n10370) );
  NOR4_X1 U11412 ( .A1(n10373), .A2(n10372), .A3(n10371), .A4(n10370), .ZN(
        n10405) );
  INV_X1 U11413 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10375) );
  AOI22_X1 U11414 ( .A1(n10376), .A2(keyinput71), .B1(keyinput68), .B2(n10375), 
        .ZN(n10374) );
  OAI221_X1 U11415 ( .B1(n10376), .B2(keyinput71), .C1(n10375), .C2(keyinput68), .A(n10374), .ZN(n10388) );
  AOI22_X1 U11416 ( .A1(n10379), .A2(keyinput85), .B1(keyinput38), .B2(n10378), 
        .ZN(n10377) );
  OAI221_X1 U11417 ( .B1(n10379), .B2(keyinput85), .C1(n10378), .C2(keyinput38), .A(n10377), .ZN(n10387) );
  INV_X1 U11418 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U11419 ( .A1(n10382), .A2(keyinput73), .B1(keyinput36), .B2(n10381), 
        .ZN(n10380) );
  OAI221_X1 U11420 ( .B1(n10382), .B2(keyinput73), .C1(n10381), .C2(keyinput36), .A(n10380), .ZN(n10386) );
  XNOR2_X1 U11421 ( .A(P1_REG3_REG_0__SCAN_IN), .B(keyinput82), .ZN(n10384) );
  XNOR2_X1 U11422 ( .A(P2_B_REG_SCAN_IN), .B(keyinput29), .ZN(n10383) );
  NAND2_X1 U11423 ( .A1(n10384), .A2(n10383), .ZN(n10385) );
  NOR4_X1 U11424 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10404) );
  AOI22_X1 U11425 ( .A1(n6416), .A2(keyinput115), .B1(n10390), .B2(keyinput92), 
        .ZN(n10389) );
  OAI221_X1 U11426 ( .B1(n6416), .B2(keyinput115), .C1(n10390), .C2(keyinput92), .A(n10389), .ZN(n10402) );
  AOI22_X1 U11427 ( .A1(n6267), .A2(keyinput91), .B1(n10392), .B2(keyinput58), 
        .ZN(n10391) );
  OAI221_X1 U11428 ( .B1(n6267), .B2(keyinput91), .C1(n10392), .C2(keyinput58), 
        .A(n10391), .ZN(n10401) );
  AOI22_X1 U11429 ( .A1(n10395), .A2(keyinput106), .B1(keyinput8), .B2(n10394), 
        .ZN(n10393) );
  OAI221_X1 U11430 ( .B1(n10395), .B2(keyinput106), .C1(n10394), .C2(keyinput8), .A(n10393), .ZN(n10400) );
  AOI22_X1 U11431 ( .A1(n10398), .A2(keyinput75), .B1(n10397), .B2(keyinput72), 
        .ZN(n10396) );
  OAI221_X1 U11432 ( .B1(n10398), .B2(keyinput75), .C1(n10397), .C2(keyinput72), .A(n10396), .ZN(n10399) );
  NOR4_X1 U11433 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10403) );
  NAND4_X1 U11434 ( .A1(n10406), .A2(n10405), .A3(n10404), .A4(n10403), .ZN(
        n10482) );
  OAI22_X1 U11435 ( .A1(P1_D_REG_22__SCAN_IN), .A2(keyinput124), .B1(
        keyinput78), .B2(P1_DATAO_REG_31__SCAN_IN), .ZN(n10407) );
  AOI221_X1 U11436 ( .B1(P1_D_REG_22__SCAN_IN), .B2(keyinput124), .C1(
        P1_DATAO_REG_31__SCAN_IN), .C2(keyinput78), .A(n10407), .ZN(n10414) );
  OAI22_X1 U11437 ( .A1(P2_REG1_REG_23__SCAN_IN), .A2(keyinput63), .B1(
        P1_REG0_REG_30__SCAN_IN), .B2(keyinput79), .ZN(n10408) );
  AOI221_X1 U11438 ( .B1(P2_REG1_REG_23__SCAN_IN), .B2(keyinput63), .C1(
        keyinput79), .C2(P1_REG0_REG_30__SCAN_IN), .A(n10408), .ZN(n10413) );
  OAI22_X1 U11439 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(keyinput32), .B1(
        keyinput60), .B2(P1_ADDR_REG_10__SCAN_IN), .ZN(n10409) );
  AOI221_X1 U11440 ( .B1(P1_REG3_REG_12__SCAN_IN), .B2(keyinput32), .C1(
        P1_ADDR_REG_10__SCAN_IN), .C2(keyinput60), .A(n10409), .ZN(n10412) );
  OAI22_X1 U11441 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput19), .B1(
        P1_REG1_REG_26__SCAN_IN), .B2(keyinput126), .ZN(n10410) );
  AOI221_X1 U11442 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput19), .C1(
        keyinput126), .C2(P1_REG1_REG_26__SCAN_IN), .A(n10410), .ZN(n10411) );
  NAND4_X1 U11443 ( .A1(n10414), .A2(n10413), .A3(n10412), .A4(n10411), .ZN(
        n10442) );
  OAI22_X1 U11444 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(keyinput7), .B1(
        keyinput52), .B2(P1_REG3_REG_3__SCAN_IN), .ZN(n10415) );
  AOI221_X1 U11445 ( .B1(P1_DATAO_REG_7__SCAN_IN), .B2(keyinput7), .C1(
        P1_REG3_REG_3__SCAN_IN), .C2(keyinput52), .A(n10415), .ZN(n10422) );
  OAI22_X1 U11446 ( .A1(P1_REG1_REG_29__SCAN_IN), .A2(keyinput86), .B1(
        keyinput99), .B2(P2_REG0_REG_31__SCAN_IN), .ZN(n10416) );
  AOI221_X1 U11447 ( .B1(P1_REG1_REG_29__SCAN_IN), .B2(keyinput86), .C1(
        P2_REG0_REG_31__SCAN_IN), .C2(keyinput99), .A(n10416), .ZN(n10421) );
  OAI22_X1 U11448 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(keyinput12), .B1(
        keyinput113), .B2(P1_ADDR_REG_5__SCAN_IN), .ZN(n10417) );
  AOI221_X1 U11449 ( .B1(P2_REG2_REG_25__SCAN_IN), .B2(keyinput12), .C1(
        P1_ADDR_REG_5__SCAN_IN), .C2(keyinput113), .A(n10417), .ZN(n10420) );
  OAI22_X1 U11450 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(keyinput118), .B1(
        keyinput121), .B2(P2_REG2_REG_12__SCAN_IN), .ZN(n10418) );
  AOI221_X1 U11451 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(keyinput118), .C1(
        P2_REG2_REG_12__SCAN_IN), .C2(keyinput121), .A(n10418), .ZN(n10419) );
  NAND4_X1 U11452 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        n10441) );
  OAI22_X1 U11453 ( .A1(P1_REG0_REG_9__SCAN_IN), .A2(keyinput76), .B1(
        keyinput105), .B2(P2_D_REG_8__SCAN_IN), .ZN(n10423) );
  AOI221_X1 U11454 ( .B1(P1_REG0_REG_9__SCAN_IN), .B2(keyinput76), .C1(
        P2_D_REG_8__SCAN_IN), .C2(keyinput105), .A(n10423), .ZN(n10430) );
  OAI22_X1 U11455 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput43), .B1(
        P1_REG2_REG_15__SCAN_IN), .B2(keyinput116), .ZN(n10424) );
  AOI221_X1 U11456 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput43), .C1(
        keyinput116), .C2(P1_REG2_REG_15__SCAN_IN), .A(n10424), .ZN(n10429) );
  OAI22_X1 U11457 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(keyinput88), .B1(
        keyinput44), .B2(P1_REG2_REG_30__SCAN_IN), .ZN(n10425) );
  AOI221_X1 U11458 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(keyinput88), .C1(
        P1_REG2_REG_30__SCAN_IN), .C2(keyinput44), .A(n10425), .ZN(n10428) );
  OAI22_X1 U11459 ( .A1(P1_REG0_REG_6__SCAN_IN), .A2(keyinput34), .B1(
        P2_D_REG_30__SCAN_IN), .B2(keyinput108), .ZN(n10426) );
  AOI221_X1 U11460 ( .B1(P1_REG0_REG_6__SCAN_IN), .B2(keyinput34), .C1(
        keyinput108), .C2(P2_D_REG_30__SCAN_IN), .A(n10426), .ZN(n10427) );
  NAND4_X1 U11461 ( .A1(n10430), .A2(n10429), .A3(n10428), .A4(n10427), .ZN(
        n10440) );
  OAI22_X1 U11462 ( .A1(SI_22_), .A2(keyinput87), .B1(keyinput17), .B2(
        P1_REG3_REG_13__SCAN_IN), .ZN(n10431) );
  AOI221_X1 U11463 ( .B1(SI_22_), .B2(keyinput87), .C1(P1_REG3_REG_13__SCAN_IN), .C2(keyinput17), .A(n10431), .ZN(n10438) );
  OAI22_X1 U11464 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(keyinput24), .B1(keyinput55), .B2(P2_REG1_REG_21__SCAN_IN), .ZN(n10432) );
  AOI221_X1 U11465 ( .B1(P2_IR_REG_1__SCAN_IN), .B2(keyinput24), .C1(
        P2_REG1_REG_21__SCAN_IN), .C2(keyinput55), .A(n10432), .ZN(n10437) );
  OAI22_X1 U11466 ( .A1(P1_REG1_REG_20__SCAN_IN), .A2(keyinput123), .B1(
        keyinput16), .B2(P2_REG1_REG_4__SCAN_IN), .ZN(n10433) );
  AOI221_X1 U11467 ( .B1(P1_REG1_REG_20__SCAN_IN), .B2(keyinput123), .C1(
        P2_REG1_REG_4__SCAN_IN), .C2(keyinput16), .A(n10433), .ZN(n10436) );
  OAI22_X1 U11468 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput33), .B1(
        keyinput35), .B2(P1_D_REG_20__SCAN_IN), .ZN(n10434) );
  AOI221_X1 U11469 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput33), .C1(
        P1_D_REG_20__SCAN_IN), .C2(keyinput35), .A(n10434), .ZN(n10435) );
  NAND4_X1 U11470 ( .A1(n10438), .A2(n10437), .A3(n10436), .A4(n10435), .ZN(
        n10439) );
  NOR4_X1 U11471 ( .A1(n10442), .A2(n10441), .A3(n10440), .A4(n10439), .ZN(
        n10480) );
  OAI22_X1 U11472 ( .A1(P1_REG0_REG_15__SCAN_IN), .A2(keyinput28), .B1(
        keyinput13), .B2(P1_ADDR_REG_9__SCAN_IN), .ZN(n10443) );
  AOI221_X1 U11473 ( .B1(P1_REG0_REG_15__SCAN_IN), .B2(keyinput28), .C1(
        P1_ADDR_REG_9__SCAN_IN), .C2(keyinput13), .A(n10443), .ZN(n10450) );
  OAI22_X1 U11474 ( .A1(P1_D_REG_30__SCAN_IN), .A2(keyinput101), .B1(
        P2_D_REG_2__SCAN_IN), .B2(keyinput50), .ZN(n10444) );
  AOI221_X1 U11475 ( .B1(P1_D_REG_30__SCAN_IN), .B2(keyinput101), .C1(
        keyinput50), .C2(P2_D_REG_2__SCAN_IN), .A(n10444), .ZN(n10449) );
  OAI22_X1 U11476 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput21), .B1(
        keyinput39), .B2(P1_REG1_REG_8__SCAN_IN), .ZN(n10445) );
  AOI221_X1 U11477 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput21), .C1(
        P1_REG1_REG_8__SCAN_IN), .C2(keyinput39), .A(n10445), .ZN(n10448) );
  OAI22_X1 U11478 ( .A1(P1_D_REG_7__SCAN_IN), .A2(keyinput37), .B1(
        P1_REG2_REG_12__SCAN_IN), .B2(keyinput51), .ZN(n10446) );
  AOI221_X1 U11479 ( .B1(P1_D_REG_7__SCAN_IN), .B2(keyinput37), .C1(keyinput51), .C2(P1_REG2_REG_12__SCAN_IN), .A(n10446), .ZN(n10447) );
  NAND4_X1 U11480 ( .A1(n10450), .A2(n10449), .A3(n10448), .A4(n10447), .ZN(
        n10478) );
  OAI22_X1 U11481 ( .A1(P1_REG0_REG_14__SCAN_IN), .A2(keyinput23), .B1(
        keyinput48), .B2(P2_REG1_REG_1__SCAN_IN), .ZN(n10451) );
  AOI221_X1 U11482 ( .B1(P1_REG0_REG_14__SCAN_IN), .B2(keyinput23), .C1(
        P2_REG1_REG_1__SCAN_IN), .C2(keyinput48), .A(n10451), .ZN(n10458) );
  OAI22_X1 U11483 ( .A1(SI_21_), .A2(keyinput30), .B1(keyinput69), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n10452) );
  AOI221_X1 U11484 ( .B1(SI_21_), .B2(keyinput30), .C1(P2_REG2_REG_16__SCAN_IN), .C2(keyinput69), .A(n10452), .ZN(n10457) );
  OAI22_X1 U11485 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(keyinput26), .B1(
        keyinput62), .B2(P2_D_REG_9__SCAN_IN), .ZN(n10453) );
  AOI221_X1 U11486 ( .B1(P2_IR_REG_24__SCAN_IN), .B2(keyinput26), .C1(
        P2_D_REG_9__SCAN_IN), .C2(keyinput62), .A(n10453), .ZN(n10456) );
  OAI22_X1 U11487 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(keyinput89), .B1(
        keyinput120), .B2(P1_REG2_REG_31__SCAN_IN), .ZN(n10454) );
  AOI221_X1 U11488 ( .B1(P1_DATAO_REG_2__SCAN_IN), .B2(keyinput89), .C1(
        P1_REG2_REG_31__SCAN_IN), .C2(keyinput120), .A(n10454), .ZN(n10455) );
  NAND4_X1 U11489 ( .A1(n10458), .A2(n10457), .A3(n10456), .A4(n10455), .ZN(
        n10477) );
  OAI22_X1 U11490 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(keyinput122), .B1(
        P2_REG0_REG_2__SCAN_IN), .B2(keyinput61), .ZN(n10459) );
  AOI221_X1 U11491 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(keyinput122), .C1(
        keyinput61), .C2(P2_REG0_REG_2__SCAN_IN), .A(n10459), .ZN(n10466) );
  OAI22_X1 U11492 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput119), .B1(
        P1_REG0_REG_7__SCAN_IN), .B2(keyinput57), .ZN(n10460) );
  AOI221_X1 U11493 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput119), .C1(
        keyinput57), .C2(P1_REG0_REG_7__SCAN_IN), .A(n10460), .ZN(n10465) );
  OAI22_X1 U11494 ( .A1(P1_REG1_REG_24__SCAN_IN), .A2(keyinput117), .B1(
        keyinput66), .B2(P2_REG2_REG_31__SCAN_IN), .ZN(n10461) );
  AOI221_X1 U11495 ( .B1(P1_REG1_REG_24__SCAN_IN), .B2(keyinput117), .C1(
        P2_REG2_REG_31__SCAN_IN), .C2(keyinput66), .A(n10461), .ZN(n10464) );
  OAI22_X1 U11496 ( .A1(P1_REG1_REG_4__SCAN_IN), .A2(keyinput107), .B1(
        P1_REG0_REG_2__SCAN_IN), .B2(keyinput45), .ZN(n10462) );
  AOI221_X1 U11497 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(keyinput107), .C1(
        keyinput45), .C2(P1_REG0_REG_2__SCAN_IN), .A(n10462), .ZN(n10463) );
  NAND4_X1 U11498 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10476) );
  OAI22_X1 U11499 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput53), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput90), .ZN(n10467) );
  AOI221_X1 U11500 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput53), .C1(
        keyinput90), .C2(P2_DATAO_REG_14__SCAN_IN), .A(n10467), .ZN(n10474) );
  OAI22_X1 U11501 ( .A1(SI_26_), .A2(keyinput3), .B1(keyinput4), .B2(SI_24_), 
        .ZN(n10468) );
  AOI221_X1 U11502 ( .B1(SI_26_), .B2(keyinput3), .C1(SI_24_), .C2(keyinput4), 
        .A(n10468), .ZN(n10473) );
  OAI22_X1 U11503 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(keyinput31), .B1(
        P2_D_REG_6__SCAN_IN), .B2(keyinput59), .ZN(n10469) );
  AOI221_X1 U11504 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(keyinput31), .C1(
        keyinput59), .C2(P2_D_REG_6__SCAN_IN), .A(n10469), .ZN(n10472) );
  OAI22_X1 U11505 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(keyinput127), .B1(
        keyinput100), .B2(P2_ADDR_REG_15__SCAN_IN), .ZN(n10470) );
  AOI221_X1 U11506 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(keyinput127), .C1(
        P2_ADDR_REG_15__SCAN_IN), .C2(keyinput100), .A(n10470), .ZN(n10471) );
  NAND4_X1 U11507 ( .A1(n10474), .A2(n10473), .A3(n10472), .A4(n10471), .ZN(
        n10475) );
  NOR4_X1 U11508 ( .A1(n10478), .A2(n10477), .A3(n10476), .A4(n10475), .ZN(
        n10479) );
  NAND2_X1 U11509 ( .A1(n10480), .A2(n10479), .ZN(n10481) );
  NOR4_X1 U11510 ( .A1(n10484), .A2(n10483), .A3(n10482), .A4(n10481), .ZN(
        n10485) );
  XNOR2_X1 U11511 ( .A(n10486), .B(n10485), .ZN(P2_U3245) );
  XNOR2_X1 U11512 ( .A(n10488), .B(n10487), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11513 ( .A(n10490), .B(n10489), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11514 ( .A(n10492), .B(n10491), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11515 ( .A(n10494), .B(n10493), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11516 ( .A(n10496), .B(n10495), .ZN(ADD_1068_U48) );
  XOR2_X1 U11517 ( .A(n10498), .B(n10497), .Z(ADD_1068_U54) );
  XOR2_X1 U11518 ( .A(n10500), .B(n10499), .Z(ADD_1068_U53) );
  XNOR2_X1 U11519 ( .A(n10502), .B(n10501), .ZN(ADD_1068_U52) );
  NAND2_X2 U5222 ( .A1(n6707), .A2(n6680), .ZN(n8890) );
  CLKBUF_X1 U5006 ( .A(n7963), .Z(n4495) );
  CLKBUF_X1 U5008 ( .A(n6118), .Z(n7349) );
  NAND2_X1 U5026 ( .A1(n6070), .A2(n6021), .ZN(n6112) );
endmodule

