

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277;

  INV_X1 U4780 ( .A(n9899), .ZN(n9921) );
  NAND2_X1 U4781 ( .A1(n8636), .A2(n8635), .ZN(n4848) );
  NAND2_X1 U4782 ( .A1(n4591), .A2(n4589), .ZN(n7853) );
  CLKBUF_X2 U4783 ( .A(n6764), .Z(n4427) );
  NAND2_X1 U4784 ( .A1(n7662), .A2(n6628), .ZN(n5834) );
  NAND2_X1 U4785 ( .A1(n5170), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5208) );
  INV_X2 U4787 ( .A(n6727), .ZN(n4633) );
  NAND3_X1 U4788 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5130) );
  INV_X1 U4789 ( .A(n7684), .ZN(n6628) );
  INV_X1 U4790 ( .A(n8967), .ZN(n4457) );
  INV_X1 U4792 ( .A(n6526), .ZN(n6520) );
  NAND2_X1 U4793 ( .A1(n6737), .A2(n6736), .ZN(n8521) );
  NAND2_X1 U4794 ( .A1(n7833), .A2(n7684), .ZN(n6756) );
  INV_X1 U4795 ( .A(n8916), .ZN(n8965) );
  CLKBUF_X3 U4796 ( .A(n6100), .Z(n8087) );
  AOI21_X1 U4797 ( .B1(n9376), .B2(n7968), .A(n7967), .ZN(n9125) );
  NOR2_X1 U4798 ( .A1(n9389), .A2(n9631), .ZN(n9366) );
  NAND2_X1 U4799 ( .A1(n5228), .A2(n5227), .ZN(n8844) );
  CLKBUF_X3 U4800 ( .A(n5336), .Z(n6527) );
  NAND2_X1 U4801 ( .A1(n8576), .A2(n8581), .ZN(n8575) );
  INV_X2 U4802 ( .A(n6121), .ZN(n8085) );
  XNOR2_X1 U4803 ( .A(n4486), .B(n5263), .ZN(n6862) );
  NAND2_X1 U4804 ( .A1(n4299), .A2(n5101), .ZN(n8432) );
  AOI211_X1 U4805 ( .C1(n8777), .C2(n8670), .A(n8573), .B(n8572), .ZN(n8574)
         );
  INV_X1 U4806 ( .A(n9307), .ZN(n9126) );
  INV_X1 U4807 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5204) );
  CLKBUF_X3 U4808 ( .A(n5670), .Z(n5777) );
  OAI21_X2 U4809 ( .B1(n9886), .B2(n8175), .A(n7592), .ZN(n7748) );
  NAND2_X2 U4810 ( .A1(n7591), .A2(n7590), .ZN(n9886) );
  OAI21_X2 U4811 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10102), .ZN(n10100) );
  OAI21_X2 U4812 ( .B1(n5381), .B2(n4785), .A(n4783), .ZN(n5422) );
  INV_X2 U4813 ( .A(n7472), .ZN(n7012) );
  NOR2_X2 U4814 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5937) );
  AND3_X2 U4815 ( .A1(n4999), .A2(n5617), .A3(n4998), .ZN(n5001) );
  NOR2_X2 U4816 ( .A1(n4992), .A2(n4991), .ZN(n5617) );
  NAND2_X2 U4817 ( .A1(n7709), .A2(n7774), .ZN(n7730) );
  NOR2_X4 U4818 ( .A1(n7673), .A2(n8855), .ZN(n7709) );
  NAND2_X1 U4819 ( .A1(n6480), .A2(n8101), .ZN(n5990) );
  XNOR2_X2 U4820 ( .A(n5971), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6480) );
  NAND2_X2 U4821 ( .A1(n4848), .A2(n4846), .ZN(n8606) );
  XNOR2_X2 U4822 ( .A(n5082), .B(n4767), .ZN(n5081) );
  AND2_X2 U4823 ( .A1(n5062), .A2(n5063), .ZN(n5082) );
  NAND2_X2 U4824 ( .A1(n9477), .A2(n4324), .ZN(n9293) );
  AOI21_X2 U4825 ( .B1(n9489), .B2(n9289), .A(n9288), .ZN(n9477) );
  XNOR2_X2 U4826 ( .A(n5477), .B(n5476), .ZN(n7836) );
  NAND2_X2 U4828 ( .A1(n7853), .A2(n7854), .ZN(n7891) );
  NAND2_X2 U4829 ( .A1(n8435), .A2(n6987), .ZN(n6638) );
  INV_X2 U4830 ( .A(n5649), .ZN(n8435) );
  AOI21_X2 U4831 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7322), .A(n7317), .ZN(
        n7198) );
  AOI21_X2 U4832 ( .B1(n7117), .B2(n7115), .A(n7116), .ZN(n9193) );
  NOR2_X4 U4833 ( .A1(n5087), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5351) );
  XNOR2_X2 U4834 ( .A(n5241), .B(n5236), .ZN(n6849) );
  AOI21_X2 U4835 ( .B1(n4625), .B2(n6748), .A(n6607), .ZN(n6758) );
  XNOR2_X1 U4836 ( .A(n4595), .B(n5003), .ZN(n8267) );
  AOI21_X2 U4837 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10108), .ZN(n10107) );
  NAND2_X2 U4838 ( .A1(n7583), .A2(n7582), .ZN(n7581) );
  OAI21_X2 U4839 ( .B1(n7347), .B2(n4715), .A(n4712), .ZN(n7583) );
  BUF_X8 U4840 ( .A(n6807), .Z(n4277) );
  OAI22_X2 U4841 ( .A1(n8692), .A2(n4504), .B1(n5595), .B2(n4505), .ZN(n8633)
         );
  NAND2_X2 U4842 ( .A1(n8691), .A2(n8696), .ZN(n8692) );
  NOR2_X2 U4843 ( .A1(n9792), .A2(n10124), .ZN(n9794) );
  NAND2_X1 U4844 ( .A1(n4719), .A2(n4717), .ZN(n8308) );
  CLKBUF_X1 U4845 ( .A(n9400), .Z(n9401) );
  INV_X1 U4846 ( .A(n8501), .ZN(n8417) );
  NAND2_X1 U4847 ( .A1(n7845), .A2(n7844), .ZN(n7843) );
  NAND2_X1 U4848 ( .A1(n7766), .A2(n7765), .ZN(n7764) );
  NAND2_X1 U4849 ( .A1(n4511), .A2(n4509), .ZN(n7857) );
  NAND2_X1 U4850 ( .A1(n6365), .A2(n6364), .ZN(n9675) );
  INV_X1 U4851 ( .A(n10023), .ZN(n10019) );
  NAND2_X1 U4852 ( .A1(n4636), .A2(n4635), .ZN(n6625) );
  INV_X2 U4853 ( .A(n7538), .ZN(n7535) );
  INV_X1 U4854 ( .A(n9136), .ZN(n7428) );
  CLKBUF_X2 U4855 ( .A(n6008), .Z(n8961) );
  NAND2_X1 U4856 ( .A1(n5059), .A2(n4306), .ZN(n8434) );
  AND3_X1 U4857 ( .A1(n5092), .A2(n5091), .A3(n5090), .ZN(n10063) );
  INV_X2 U4858 ( .A(n8969), .ZN(n6008) );
  CLKBUF_X2 U4859 ( .A(n8067), .Z(n8054) );
  OR2_X1 U4860 ( .A1(n5263), .A2(n4793), .ZN(n4792) );
  OR2_X1 U4861 ( .A1(n5391), .A2(n5551), .ZN(n5392) );
  INV_X1 U4862 ( .A(n5962), .ZN(n8262) );
  MUX2_X1 U4863 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5929), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5930) );
  AND2_X1 U4864 ( .A1(n5351), .A2(n4886), .ZN(n4850) );
  NAND2_X1 U4865 ( .A1(n4516), .A2(n4515), .ZN(n4400) );
  NOR2_X1 U4866 ( .A1(n8395), .A2(n8396), .ZN(n8394) );
  AOI21_X1 U4867 ( .B1(n8751), .B2(n8750), .A(n4694), .ZN(n4693) );
  AOI21_X1 U4868 ( .B1(n5829), .B2(n10021), .A(n8388), .ZN(n8765) );
  NAND2_X1 U4869 ( .A1(n4863), .A2(n4337), .ZN(n8751) );
  NOR2_X1 U4870 ( .A1(n4604), .A2(n4399), .ZN(n4398) );
  OAI21_X1 U4871 ( .B1(n4957), .B2(n9309), .A(n4284), .ZN(n9375) );
  NOR4_X1 U4872 ( .A1(n8187), .A2(n9620), .A3(n9362), .A4(n8186), .ZN(n8190)
         );
  INV_X1 U4873 ( .A(n4913), .ZN(n4912) );
  NAND2_X1 U4874 ( .A1(n7905), .A2(n7904), .ZN(n7915) );
  NAND2_X1 U4875 ( .A1(n7843), .A2(n5713), .ZN(n7905) );
  NAND2_X1 U4876 ( .A1(n4622), .A2(n4394), .ZN(n8470) );
  NAND2_X1 U4877 ( .A1(n7857), .A2(n4869), .ZN(n8719) );
  OR2_X1 U4878 ( .A1(n9631), .A2(n9125), .ZN(n9340) );
  NAND2_X1 U4879 ( .A1(n7960), .A2(n7959), .ZN(n9631) );
  OR2_X2 U4880 ( .A1(n8654), .A2(n8802), .ZN(n4983) );
  NAND2_X1 U4881 ( .A1(n5585), .A2(n4513), .ZN(n4511) );
  NAND2_X1 U4882 ( .A1(n9402), .A2(n9306), .ZN(n9337) );
  NAND2_X1 U4883 ( .A1(n6400), .A2(n6399), .ZN(n9663) );
  NAND2_X1 U4884 ( .A1(n6381), .A2(n6380), .ZN(n9669) );
  NAND2_X1 U4885 ( .A1(n6419), .A2(n6418), .ZN(n9417) );
  NAND2_X1 U4886 ( .A1(n6324), .A2(n6323), .ZN(n9678) );
  CLKBUF_X2 U4887 ( .A(n9125), .Z(n4281) );
  XNOR2_X1 U4888 ( .A(n5439), .B(n5437), .ZN(n7680) );
  NAND2_X1 U4889 ( .A1(n7871), .A2(n4820), .ZN(n7926) );
  NAND2_X1 U4890 ( .A1(n5371), .A2(n5370), .ZN(n8805) );
  NAND2_X1 U4891 ( .A1(n6341), .A2(n6340), .ZN(n9510) );
  AND2_X1 U4892 ( .A1(n6491), .A2(n6490), .ZN(n9307) );
  AND2_X1 U4893 ( .A1(n7361), .A2(n5579), .ZN(n7618) );
  OR2_X1 U4894 ( .A1(n9701), .A2(n9020), .ZN(n9543) );
  NAND2_X1 U4895 ( .A1(n5354), .A2(n5353), .ZN(n8811) );
  NAND2_X1 U4896 ( .A1(n5312), .A2(n5311), .ZN(n8824) );
  NAND2_X1 U4897 ( .A1(n5292), .A2(n5291), .ZN(n8828) );
  NOR2_X1 U4898 ( .A1(n7822), .A2(n7821), .ZN(n7820) );
  NAND2_X1 U4899 ( .A1(n6253), .A2(n6252), .ZN(n9708) );
  NAND2_X1 U4900 ( .A1(n7637), .A2(n4621), .ZN(n7822) );
  AND2_X1 U4901 ( .A1(n4608), .A2(n4607), .ZN(n7490) );
  NAND2_X1 U4902 ( .A1(n5188), .A2(n5187), .ZN(n8855) );
  NAND2_X1 U4903 ( .A1(n6142), .A2(n6141), .ZN(n7653) );
  NAND2_X1 U4904 ( .A1(n5169), .A2(n5168), .ZN(n8860) );
  INV_X1 U4905 ( .A(n6366), .ZN(n5954) );
  INV_X1 U4906 ( .A(n7445), .ZN(n7562) );
  AND2_X1 U4907 ( .A1(n4616), .A2(n4374), .ZN(n7317) );
  INV_X1 U4908 ( .A(n7393), .ZN(n4635) );
  NAND2_X1 U4909 ( .A1(n4347), .A2(n5078), .ZN(n8433) );
  AOI21_X1 U4910 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n6931), .A(n6926), .ZN(
        n6892) );
  XNOR2_X1 U4911 ( .A(n5670), .B(n6987), .ZN(n7089) );
  NAND2_X1 U4912 ( .A1(n5125), .A2(n5124), .ZN(n7382) );
  NAND2_X1 U4913 ( .A1(n6770), .A2(n7012), .ZN(n6640) );
  NAND2_X1 U4914 ( .A1(n6104), .A2(n6103), .ZN(n7538) );
  AND2_X1 U4915 ( .A1(n6085), .A2(n6084), .ZN(n7445) );
  NAND4_X1 U4916 ( .A1(n6099), .A2(n6098), .A3(n6097), .A4(n6096), .ZN(n9136)
         );
  CLKBUF_X1 U4917 ( .A(n9938), .Z(n4433) );
  NAND2_X1 U4918 ( .A1(n8120), .A2(n7991), .ZN(n8168) );
  NAND2_X1 U4919 ( .A1(n10116), .A2(n10114), .ZN(n9789) );
  NAND2_X1 U4920 ( .A1(n5142), .A2(n5141), .ZN(n5158) );
  NAND2_X4 U4921 ( .A1(n8967), .A2(n5976), .ZN(n6047) );
  OR2_X1 U4922 ( .A1(n9138), .A2(n9836), .ZN(n8120) );
  NAND2_X2 U4923 ( .A1(n6792), .A2(n5992), .ZN(n8916) );
  INV_X2 U4924 ( .A(n10063), .ZN(n4278) );
  AND3_X2 U4925 ( .A1(n5048), .A2(n5047), .A3(n5046), .ZN(n7472) );
  NOR2_X1 U4926 ( .A1(n7277), .A2(n4319), .ZN(n7333) );
  AND3_X1 U4927 ( .A1(n6045), .A2(n6044), .A3(n6043), .ZN(n9836) );
  OAI211_X1 U4928 ( .C1(n6547), .C2(n5060), .A(n5073), .B(n4322), .ZN(n5663)
         );
  AND4_X1 U4929 ( .A1(n6079), .A2(n6078), .A3(n6077), .A4(n6076), .ZN(n7505)
         );
  NAND2_X2 U4930 ( .A1(n5951), .A2(n5969), .ZN(n8969) );
  NAND4_X1 U4931 ( .A1(n6060), .A2(n6059), .A3(n6058), .A4(n6057), .ZN(n9137)
         );
  CLKBUF_X1 U4932 ( .A(n5249), .Z(n6547) );
  NAND2_X1 U4933 ( .A1(n5006), .A2(n8267), .ZN(n5075) );
  NOR2_X1 U4934 ( .A1(n5249), .A2(n6809), .ZN(n4831) );
  BUF_X2 U4935 ( .A(n5074), .Z(n6526) );
  NAND4_X2 U4936 ( .A1(n5979), .A2(n5981), .A3(n5980), .A4(n4888), .ZN(n9140)
         );
  XNOR2_X1 U4937 ( .A(n5974), .B(n5973), .ZN(n6479) );
  CLKBUF_X1 U4938 ( .A(n5605), .Z(n6755) );
  OR2_X1 U4939 ( .A1(n6853), .A2(n4558), .ZN(n6040) );
  INV_X1 U4940 ( .A(n6238), .ZN(n6121) );
  OR2_X1 U4941 ( .A1(n5008), .A2(n8267), .ZN(n5058) );
  INV_X1 U4942 ( .A(n6002), .ZN(n6764) );
  NAND2_X1 U4943 ( .A1(n6458), .A2(n5950), .ZN(n5969) );
  AOI21_X1 U4944 ( .B1(n7295), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7290), .ZN(
        n7279) );
  OR2_X1 U4945 ( .A1(n6236), .A2(n7130), .ZN(n6254) );
  NAND2_X2 U4946 ( .A1(n5553), .A2(n5392), .ZN(n7558) );
  NAND2_X1 U4947 ( .A1(n5961), .A2(n5962), .ZN(n8067) );
  NAND2_X2 U4948 ( .A1(n8262), .A2(n5961), .ZN(n6238) );
  INV_X1 U4949 ( .A(n5851), .ZN(n4279) );
  INV_X1 U4950 ( .A(n6036), .ZN(n6442) );
  NAND2_X1 U4951 ( .A1(n5553), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4417) );
  NAND2_X1 U4952 ( .A1(n5391), .A2(n5551), .ZN(n5553) );
  NAND2_X1 U4953 ( .A1(n8240), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5002) );
  CLKBUF_X1 U4954 ( .A(n6492), .Z(n4426) );
  XNOR2_X1 U4955 ( .A(n5960), .B(n5959), .ZN(n9762) );
  NAND2_X1 U4956 ( .A1(n5549), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5391) );
  XNOR2_X1 U4957 ( .A(n5927), .B(n5957), .ZN(n6492) );
  NAND2_X1 U4958 ( .A1(n8254), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U4959 ( .A1(n4413), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5960) );
  OAI21_X1 U4960 ( .B1(n5631), .B2(n4885), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n4595) );
  NAND2_X1 U4961 ( .A1(n4967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5927) );
  NAND2_X2 U4962 ( .A1(n5061), .A2(P2_U3152), .ZN(n8894) );
  NOR2_X1 U4963 ( .A1(n10126), .A2(n4350), .ZN(n10131) );
  AND2_X1 U4964 ( .A1(n4965), .A2(n4377), .ZN(n4578) );
  NAND2_X1 U4965 ( .A1(n5987), .A2(n5986), .ZN(n6942) );
  BUF_X4 U4966 ( .A(n5104), .Z(n6807) );
  AND3_X1 U4967 ( .A1(n6023), .A2(n4751), .A3(n5924), .ZN(n6139) );
  CLKBUF_X1 U4968 ( .A(n5894), .Z(n7259) );
  AND2_X1 U4969 ( .A1(n5348), .A2(n4997), .ZN(n4998) );
  AND3_X1 U4970 ( .A1(n6081), .A2(n4646), .A3(n4645), .ZN(n4751) );
  INV_X4 U4971 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4972 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5625) );
  INV_X1 U4973 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5622) );
  NOR2_X1 U4974 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4990) );
  NOR2_X1 U4975 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4993) );
  NOR2_X1 U4976 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n4554) );
  INV_X2 U4977 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U4978 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4553) );
  NOR2_X1 U4979 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4552) );
  INV_X1 U4980 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6463) );
  NOR2_X1 U4981 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4994) );
  NAND2_X1 U4982 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10085) );
  NOR2_X1 U4983 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4548) );
  NOR2_X1 U4984 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4549) );
  NOR2_X1 U4985 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4550) );
  INV_X1 U4986 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5944) );
  NOR2_X1 U4987 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4995) );
  OAI21_X2 U4988 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10096), .ZN(n10094) );
  NAND2_X1 U4989 ( .A1(n5851), .A2(n5061), .ZN(n4280) );
  NAND2_X1 U4990 ( .A1(n5851), .A2(n5061), .ZN(n6549) );
  OR2_X1 U4991 ( .A1(n8620), .A2(n4855), .ZN(n4854) );
  AOI21_X2 U4992 ( .B1(n9432), .B2(n9301), .A(n4437), .ZN(n9416) );
  NAND2_X2 U4993 ( .A1(n4960), .A2(n4958), .ZN(n9432) );
  AOI21_X2 U4994 ( .B1(n9147), .B2(n9146), .A(n9145), .ZN(n9164) );
  NAND2_X1 U4995 ( .A1(n8646), .A2(n5605), .ZN(n6757) );
  NOR2_X2 U4996 ( .A1(n8728), .A2(n8824), .ZN(n8703) );
  NAND2_X2 U4997 ( .A1(n5854), .A2(n5016), .ZN(n4689) );
  AOI21_X2 U4998 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(n10275), .A(n10273), .ZN(
        n9795) );
  NAND3_X2 U4999 ( .A1(n4868), .A2(n4623), .A3(n5000), .ZN(n5087) );
  OAI21_X2 U5000 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10087), .ZN(n10119) );
  NOR3_X4 U5001 ( .A1(n4983), .A2(n4687), .A3(n8781), .ZN(n5606) );
  INV_X1 U5002 ( .A(n5476), .ZN(n4799) );
  NAND2_X1 U5003 ( .A1(n5408), .A2(n5407), .ZN(n5423) );
  NAND2_X1 U5004 ( .A1(n4839), .A2(n4834), .ZN(n4838) );
  AND2_X1 U5005 ( .A1(n4836), .A2(n8551), .ZN(n4834) );
  OR2_X1 U5006 ( .A1(n8762), .A2(n8250), .ZN(n6729) );
  OR2_X1 U5007 ( .A1(n8776), .A2(n8309), .ZN(n6612) );
  OR2_X1 U5008 ( .A1(n8786), .A2(n8281), .ZN(n6704) );
  NAND2_X1 U5009 ( .A1(n4410), .A2(n4338), .ZN(n8062) );
  NAND2_X1 U5010 ( .A1(n8044), .A2(n4411), .ZN(n4410) );
  OR2_X1 U5011 ( .A1(n9625), .A2(n8970), .ZN(n8151) );
  OR2_X1 U5012 ( .A1(n9636), .A2(n9307), .ZN(n9338) );
  AOI21_X1 U5013 ( .B1(n6510), .B2(n6509), .A(n4386), .ZN(n6561) );
  NAND2_X1 U5014 ( .A1(n5783), .A2(n5782), .ZN(n6510) );
  NOR2_X1 U5015 ( .A1(n7892), .A2(n4870), .ZN(n4869) );
  INV_X1 U5016 ( .A(n5586), .ZN(n4870) );
  OR2_X1 U5017 ( .A1(n8839), .A2(n8425), .ZN(n4512) );
  INV_X1 U5018 ( .A(n4828), .ZN(n4827) );
  OAI21_X1 U5019 ( .B1(n5298), .B2(n4829), .A(n6689), .ZN(n4828) );
  NAND2_X1 U5020 ( .A1(n5008), .A2(n5004), .ZN(n5074) );
  INV_X1 U5021 ( .A(n8267), .ZN(n5004) );
  AND2_X1 U5022 ( .A1(n6554), .A2(n6553), .ZN(n4837) );
  OR2_X1 U5023 ( .A1(n8755), .A2(n8416), .ZN(n6737) );
  OAI21_X2 U5024 ( .B1(n8606), .B2(n4602), .A(n4600), .ZN(n4839) );
  INV_X1 U5025 ( .A(n4603), .ZN(n4602) );
  AOI21_X1 U5026 ( .B1(n4603), .B2(n4601), .A(n4340), .ZN(n4600) );
  OR2_X1 U5027 ( .A1(n8811), .A2(n8382), .ZN(n6616) );
  AOI21_X1 U5028 ( .B1(n4827), .B2(n4829), .A(n4825), .ZN(n4824) );
  INV_X1 U5029 ( .A(n6690), .ZN(n4825) );
  NOR2_X1 U5030 ( .A1(n8839), .A2(n8844), .ZN(n4699) );
  NOR2_X1 U5031 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5015) );
  NAND2_X1 U5032 ( .A1(n4564), .A2(n8063), .ZN(n8095) );
  INV_X1 U5033 ( .A(n9762), .ZN(n5961) );
  NAND2_X1 U5034 ( .A1(n4539), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7962) );
  OR2_X1 U5035 ( .A1(n9417), .A2(n9303), .ZN(n9304) );
  NAND2_X1 U5036 ( .A1(n4900), .A2(n4898), .ZN(n4896) );
  INV_X1 U5037 ( .A(n9275), .ZN(n4934) );
  OR2_X1 U5038 ( .A1(n9708), .A2(n9057), .ZN(n9541) );
  OR2_X1 U5039 ( .A1(n9725), .A2(n7791), .ZN(n8013) );
  INV_X1 U5040 ( .A(n9140), .ZN(n6874) );
  INV_X1 U5041 ( .A(n6021), .ZN(n8089) );
  AND2_X1 U5042 ( .A1(n4918), .A2(n9334), .ZN(n4915) );
  NAND2_X1 U5043 ( .A1(n4527), .A2(n4528), .ZN(n5529) );
  AOI21_X1 U5044 ( .B1(n4530), .B2(n4529), .A(n4387), .ZN(n4528) );
  AND2_X1 U5045 ( .A1(n5423), .A2(n5410), .ZN(n5421) );
  XNOR2_X1 U5046 ( .A(n5365), .B(SI_17_), .ZN(n5364) );
  OAI21_X1 U5047 ( .B1(n5284), .B2(n4310), .A(n4517), .ZN(n5344) );
  INV_X1 U5048 ( .A(n4518), .ZN(n4517) );
  OAI21_X1 U5049 ( .B1(n4521), .B2(n4310), .A(n5322), .ZN(n4518) );
  NAND2_X1 U5050 ( .A1(n5262), .A2(n5245), .ZN(n5263) );
  AND2_X1 U5051 ( .A1(n4979), .A2(n5219), .ZN(n4488) );
  AND2_X1 U5052 ( .A1(n5216), .A2(n5217), .ZN(n4418) );
  OR2_X1 U5053 ( .A1(n5104), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5062) );
  NAND2_X1 U5054 ( .A1(n5449), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5469) );
  INV_X1 U5055 ( .A(n5450), .ZN(n5449) );
  NAND2_X1 U5056 ( .A1(n4705), .A2(n4704), .ZN(n4703) );
  INV_X1 U5057 ( .A(n8246), .ZN(n4704) );
  NAND2_X1 U5058 ( .A1(n5775), .A2(n8396), .ZN(n4705) );
  AOI21_X1 U5059 ( .B1(n8560), .B2(n5810), .A(n5486), .ZN(n8309) );
  OR2_X1 U5061 ( .A1(n7196), .A2(n4611), .ZN(n4608) );
  OR2_X1 U5062 ( .A1(n4815), .A2(n4323), .ZN(n4611) );
  NAND2_X1 U5063 ( .A1(n8511), .A2(n8510), .ZN(n8748) );
  NAND2_X1 U5064 ( .A1(n6739), .A2(n6740), .ZN(n8745) );
  AND2_X1 U5065 ( .A1(n4865), .A2(n8502), .ZN(n4864) );
  NAND2_X1 U5066 ( .A1(n4866), .A2(n8499), .ZN(n4865) );
  INV_X1 U5067 ( .A(n5603), .ZN(n4866) );
  NAND2_X1 U5068 ( .A1(n4500), .A2(n4873), .ZN(n5833) );
  AOI21_X1 U5069 ( .B1(n4874), .B2(n4876), .A(n4348), .ZN(n4873) );
  NAND2_X1 U5070 ( .A1(n8575), .A2(n4874), .ZN(n4500) );
  NAND2_X1 U5071 ( .A1(n8552), .A2(n8551), .ZN(n8550) );
  OR2_X1 U5072 ( .A1(n8579), .A2(n8564), .ZN(n4975) );
  AOI21_X1 U5073 ( .B1(n4853), .B2(n6598), .A(n5601), .ZN(n4852) );
  NOR2_X1 U5074 ( .A1(n8786), .A2(n5600), .ZN(n5601) );
  NOR2_X1 U5075 ( .A1(n8793), .A2(n8796), .ZN(n4688) );
  AOI21_X1 U5076 ( .B1(n4859), .B2(n4857), .A(n4336), .ZN(n4856) );
  NAND2_X1 U5077 ( .A1(n8606), .A2(n5436), .ZN(n8607) );
  OR2_X1 U5078 ( .A1(n8796), .A2(n8291), .ZN(n8605) );
  OR2_X1 U5079 ( .A1(n8828), .A2(n8404), .ZN(n6685) );
  NOR2_X1 U5080 ( .A1(n7854), .A2(n4510), .ZN(n4509) );
  INV_X1 U5081 ( .A(n4512), .ZN(n4510) );
  AOI21_X1 U5082 ( .B1(n4592), .B2(n4594), .A(n4590), .ZN(n4589) );
  INV_X1 U5083 ( .A(n6676), .ZN(n4590) );
  OR2_X1 U5084 ( .A1(n8844), .A2(n7908), .ZN(n6673) );
  NAND2_X1 U5085 ( .A1(n8850), .A2(n7847), .ZN(n6667) );
  NAND2_X1 U5086 ( .A1(n5514), .A2(n5513), .ZN(n8762) );
  NAND2_X1 U5087 ( .A1(n5468), .A2(n5467), .ZN(n8781) );
  NAND2_X1 U5088 ( .A1(n6516), .A2(n6515), .ZN(n6542) );
  OR2_X1 U5089 ( .A1(n6561), .A2(n6558), .ZN(n6515) );
  OR2_X1 U5090 ( .A1(n5044), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5071) );
  AND2_X1 U5091 ( .A1(n8156), .A2(n6906), .ZN(n9347) );
  NOR2_X1 U5092 ( .A1(n8076), .A2(n4562), .ZN(n4560) );
  AND2_X1 U5093 ( .A1(n5968), .A2(n5967), .ZN(n9298) );
  AND2_X1 U5094 ( .A1(n6409), .A2(n6408), .ZN(n9296) );
  AND2_X1 U5095 ( .A1(n6389), .A2(n6388), .ZN(n9070) );
  AND2_X1 U5096 ( .A1(n6304), .A2(n6303), .ZN(n9021) );
  INV_X1 U5097 ( .A(n6853), .ZN(n8068) );
  BUF_X1 U5098 ( .A(n6055), .Z(n6853) );
  NAND2_X1 U5099 ( .A1(n9762), .A2(n8262), .ZN(n6055) );
  AND2_X1 U5100 ( .A1(n4667), .A2(n4670), .ZN(n4666) );
  INV_X1 U5101 ( .A(n6908), .ZN(n4667) );
  XNOR2_X1 U5102 ( .A(n9243), .B(n4436), .ZN(n9253) );
  INV_X1 U5103 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4436) );
  OR2_X1 U5104 ( .A1(n9610), .A2(n9631), .ZN(n4654) );
  OR2_X1 U5105 ( .A1(n9614), .A2(n8978), .ZN(n8158) );
  NOR2_X1 U5106 ( .A1(n4912), .A2(n9339), .ZN(n4481) );
  NAND2_X1 U5107 ( .A1(n4494), .A2(n4908), .ZN(n4906) );
  AOI21_X1 U5108 ( .B1(n4940), .B2(n4942), .A(n4346), .ZN(n4937) );
  NOR2_X1 U5109 ( .A1(n4897), .A2(n9587), .ZN(n4489) );
  INV_X1 U5110 ( .A(n4898), .ZN(n4897) );
  NAND2_X1 U5111 ( .A1(n7784), .A2(n7783), .ZN(n4936) );
  OR2_X1 U5112 ( .A1(n9936), .A2(n6480), .ZN(n6870) );
  AND2_X1 U5113 ( .A1(n9759), .A2(n6796), .ZN(n7144) );
  NAND2_X1 U5114 ( .A1(n5941), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5971) );
  OR2_X1 U5115 ( .A1(n5104), .A2(n5039), .ZN(n5040) );
  NAND2_X1 U5116 ( .A1(n4577), .A2(n4576), .ZN(n4575) );
  AOI21_X1 U5117 ( .B1(n4574), .B2(n4573), .A(n4572), .ZN(n4571) );
  NOR2_X1 U5118 ( .A1(n8107), .A2(n8066), .ZN(n4576) );
  NAND2_X1 U5119 ( .A1(n6715), .A2(n4315), .ZN(n4643) );
  NOR2_X1 U5120 ( .A1(n8581), .A2(n4641), .ZN(n4640) );
  OAI21_X1 U5121 ( .B1(n6704), .B2(n4633), .A(n4321), .ZN(n4641) );
  AND2_X1 U5122 ( .A1(n8104), .A2(n8161), .ZN(n4408) );
  NOR2_X1 U5123 ( .A1(n6729), .A2(n4633), .ZN(n4811) );
  INV_X1 U5124 ( .A(n4734), .ZN(n4733) );
  NAND2_X1 U5125 ( .A1(n7956), .A2(n7955), .ZN(n8046) );
  NAND2_X1 U5126 ( .A1(n7954), .A2(n8066), .ZN(n7955) );
  NAND2_X1 U5127 ( .A1(n7951), .A2(n8097), .ZN(n7956) );
  OR2_X1 U5128 ( .A1(n7466), .A2(n7624), .ZN(n6651) );
  NOR2_X1 U5129 ( .A1(n4733), .A2(n8990), .ZN(n4732) );
  INV_X1 U5130 ( .A(n6322), .ZN(n4465) );
  OAI21_X1 U5131 ( .B1(n4733), .B2(n4730), .A(n8989), .ZN(n4729) );
  NAND2_X1 U5132 ( .A1(n4737), .A2(n4731), .ZN(n4730) );
  INV_X1 U5133 ( .A(n8990), .ZN(n4731) );
  NOR4_X1 U5134 ( .A1(n8178), .A2(n8177), .A3(n9891), .A4(n8176), .ZN(n8180)
         );
  NOR2_X1 U5135 ( .A1(n9587), .A2(n4423), .ZN(n4422) );
  NOR2_X1 U5136 ( .A1(n6438), .A2(n10218), .ZN(n4539) );
  AND2_X1 U5137 ( .A1(n9701), .A2(n9020), .ZN(n9317) );
  OR2_X1 U5138 ( .A1(n9818), .A2(n7744), .ZN(n7743) );
  NAND2_X1 U5139 ( .A1(n7596), .A2(n7653), .ZN(n8110) );
  OR2_X1 U5140 ( .A1(n7653), .A2(n7596), .ZN(n7978) );
  INV_X1 U5141 ( .A(n9437), .ZN(n4919) );
  NOR2_X1 U5142 ( .A1(n9433), .A2(n9663), .ZN(n4651) );
  INV_X1 U5143 ( .A(SI_15_), .ZN(n5305) );
  NOR2_X1 U5144 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5924) );
  INV_X1 U5145 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4646) );
  INV_X1 U5146 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4645) );
  OAI21_X1 U5147 ( .B1(n4277), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n4401), .ZN(
        n5161) );
  NAND2_X1 U5148 ( .A1(n4277), .A2(n6839), .ZN(n4401) );
  NAND2_X1 U5149 ( .A1(n8435), .A2(n5671), .ZN(n7088) );
  NAND2_X1 U5150 ( .A1(n4808), .A2(n4807), .ZN(n4806) );
  INV_X1 U5151 ( .A(n6735), .ZN(n4807) );
  AND2_X1 U5152 ( .A1(n7213), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4815) );
  INV_X1 U5153 ( .A(n4837), .ZN(n4584) );
  NOR2_X1 U5154 ( .A1(n8559), .A2(n4879), .ZN(n4878) );
  AND2_X1 U5155 ( .A1(n8596), .A2(n6714), .ZN(n4603) );
  NAND2_X1 U5156 ( .A1(n4688), .A2(n8594), .ZN(n4687) );
  OAI21_X1 U5157 ( .B1(n4871), .B2(n4507), .A(n5596), .ZN(n4506) );
  AND2_X1 U5158 ( .A1(n6616), .A2(n6696), .ZN(n4596) );
  NOR2_X1 U5159 ( .A1(n8686), .A2(n4872), .ZN(n4871) );
  INV_X1 U5160 ( .A(n5592), .ZN(n4872) );
  OR2_X1 U5161 ( .A1(n8824), .A2(n8324), .ZN(n6690) );
  NAND2_X1 U5162 ( .A1(n4699), .A2(n7866), .ZN(n4698) );
  NAND2_X1 U5163 ( .A1(n7462), .A2(n7382), .ZN(n6649) );
  NAND2_X1 U5164 ( .A1(n6620), .A2(n7234), .ZN(n10023) );
  AND2_X1 U5165 ( .A1(n10044), .A2(n5816), .ZN(n5831) );
  INV_X1 U5166 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4580) );
  INV_X1 U5167 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5389) );
  OR2_X1 U5168 ( .A1(n5285), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5286) );
  NOR2_X1 U5169 ( .A1(n5203), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5247) );
  INV_X1 U5170 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5000) );
  NOR2_X1 U5171 ( .A1(n7563), .A2(n7501), .ZN(n6108) );
  INV_X1 U5172 ( .A(n6231), .ZN(n4757) );
  OR2_X1 U5173 ( .A1(n9306), .A2(n8969), .ZN(n4456) );
  AOI21_X1 U5174 ( .B1(n7166), .B2(n4458), .A(n4314), .ZN(n4462) );
  INV_X1 U5175 ( .A(n6053), .ZN(n4458) );
  NOR2_X1 U5176 ( .A1(n6154), .A2(n7652), .ZN(n4470) );
  INV_X1 U5177 ( .A(n6137), .ZN(n4468) );
  NAND2_X1 U5178 ( .A1(n7036), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U5179 ( .A1(n4662), .A2(n4317), .ZN(n4661) );
  NAND2_X1 U5180 ( .A1(n9629), .A2(n9616), .ZN(n4655) );
  INV_X1 U5181 ( .A(n4539), .ZN(n6484) );
  OR2_X1 U5182 ( .A1(n6421), .A2(n6420), .ZN(n6438) );
  AOI21_X1 U5183 ( .B1(n4963), .B2(n4307), .A(n9297), .ZN(n4961) );
  NOR2_X1 U5184 ( .A1(n8994), .A2(n4547), .ZN(n4546) );
  NAND2_X1 U5185 ( .A1(n9328), .A2(n9292), .ZN(n4963) );
  AND2_X1 U5186 ( .A1(n9572), .A2(n9316), .ZN(n4902) );
  OR2_X1 U5187 ( .A1(n9717), .A2(n9056), .ZN(n8016) );
  AND2_X1 U5188 ( .A1(n7978), .A2(n8110), .ZN(n8175) );
  AND3_X1 U5189 ( .A1(n6067), .A2(n6066), .A3(n6065), .ZN(n7405) );
  NAND2_X1 U5190 ( .A1(n6479), .A2(n5990), .ZN(n6792) );
  INV_X1 U5191 ( .A(n6479), .ZN(n6781) );
  NAND2_X1 U5192 ( .A1(n4291), .A2(n4917), .ZN(n4916) );
  OR2_X1 U5193 ( .A1(n9433), .A2(n9298), .ZN(n9420) );
  NAND2_X1 U5194 ( .A1(n4917), .A2(n4919), .ZN(n9439) );
  NOR2_X1 U5195 ( .A1(n9450), .A2(n4649), .ZN(n9436) );
  INV_X1 U5196 ( .A(n4651), .ZN(n4649) );
  INV_X1 U5197 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5925) );
  AOI21_X1 U5198 ( .B1(n4356), .B2(n4798), .A(n4532), .ZN(n4531) );
  INV_X1 U5199 ( .A(n5478), .ZN(n4532) );
  INV_X1 U5200 ( .A(n5423), .ZN(n4533) );
  NAND2_X1 U5201 ( .A1(n4781), .A2(n4779), .ZN(n5424) );
  AOI21_X1 U5202 ( .B1(n4783), .B2(n4785), .A(n4780), .ZN(n4779) );
  INV_X1 U5203 ( .A(n5421), .ZN(n4780) );
  INV_X1 U5204 ( .A(n5442), .ZN(n4804) );
  AND2_X1 U5205 ( .A1(n5478), .A2(n5466), .ZN(n5476) );
  NAND2_X1 U5206 ( .A1(n5424), .A2(n5423), .ZN(n5439) );
  NAND2_X1 U5207 ( .A1(n4786), .A2(n5383), .ZN(n4785) );
  INV_X1 U5208 ( .A(n5405), .ZN(n4786) );
  INV_X1 U5209 ( .A(n4784), .ZN(n4783) );
  OAI21_X1 U5210 ( .B1(n4785), .B2(n5380), .A(n5404), .ZN(n4784) );
  NOR2_X1 U5211 ( .A1(n5303), .A2(n4522), .ZN(n4521) );
  INV_X1 U5212 ( .A(n5283), .ZN(n4522) );
  INV_X1 U5213 ( .A(n5299), .ZN(n5303) );
  NAND2_X1 U5214 ( .A1(n4787), .A2(n4788), .ZN(n5284) );
  AOI21_X1 U5215 ( .B1(n4790), .B2(n4792), .A(n4789), .ZN(n4788) );
  INV_X1 U5216 ( .A(n4981), .ZN(n4789) );
  OR2_X1 U5217 ( .A1(n6267), .A2(n4748), .ZN(n6249) );
  NOR2_X1 U5218 ( .A1(n5240), .A2(n4795), .ZN(n4794) );
  INV_X1 U5219 ( .A(n5236), .ZN(n5240) );
  XNOR2_X1 U5220 ( .A(n5237), .B(SI_11_), .ZN(n5236) );
  INV_X1 U5221 ( .A(n5217), .ZN(n4503) );
  NAND2_X1 U5222 ( .A1(n5084), .A2(n5083), .ZN(n5107) );
  INV_X1 U5223 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4644) );
  INV_X1 U5224 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5060) );
  OR2_X1 U5225 ( .A1(n5670), .A2(n7099), .ZN(n5653) );
  NOR2_X1 U5226 ( .A1(n8357), .A2(n4711), .ZN(n4710) );
  INV_X1 U5227 ( .A(n5753), .ZN(n4711) );
  NAND2_X1 U5228 ( .A1(n4442), .A2(n4441), .ZN(n5337) );
  NOR2_X1 U5229 ( .A1(n5315), .A2(n5314), .ZN(n4441) );
  INV_X1 U5230 ( .A(n5316), .ZN(n4442) );
  AND2_X1 U5231 ( .A1(n5813), .A2(n10044), .ZN(n5812) );
  OR2_X1 U5232 ( .A1(n8494), .A2(n8745), .ZN(n6566) );
  AND2_X1 U5233 ( .A1(n5457), .A2(n5456), .ZN(n8281) );
  AND3_X1 U5234 ( .A1(n5362), .A2(n5361), .A3(n5360), .ZN(n8382) );
  AND4_X1 U5235 ( .A1(n5281), .A2(n5280), .A3(n5279), .A4(n5278), .ZN(n8273)
         );
  NAND2_X1 U5236 ( .A1(n5053), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U5237 ( .A1(n7186), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4813) );
  NAND2_X1 U5238 ( .A1(n4620), .A2(n7306), .ZN(n4615) );
  NAND2_X1 U5239 ( .A1(n4816), .A2(n4617), .ZN(n4616) );
  NOR2_X1 U5240 ( .A1(n4619), .A2(n4285), .ZN(n4617) );
  INV_X1 U5241 ( .A(n7208), .ZN(n4612) );
  NOR2_X1 U5242 ( .A1(n7490), .A2(n5898), .ZN(n7639) );
  NAND2_X1 U5243 ( .A1(n7639), .A2(n7638), .ZN(n7637) );
  NOR2_X1 U5244 ( .A1(n7820), .A2(n4821), .ZN(n7872) );
  AND2_X1 U5245 ( .A1(n7826), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4821) );
  NAND2_X1 U5246 ( .A1(n7872), .A2(n7873), .ZN(n7871) );
  AND2_X1 U5247 ( .A1(n7929), .A2(n7928), .ZN(n7931) );
  NAND2_X1 U5248 ( .A1(n7925), .A2(n5903), .ZN(n5905) );
  XNOR2_X1 U5249 ( .A(n4606), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n5915) );
  NOR2_X1 U5250 ( .A1(n8482), .A2(n5910), .ZN(n4606) );
  NAND2_X1 U5251 ( .A1(n6519), .A2(n6518), .ZN(n8490) );
  OR2_X1 U5252 ( .A1(n5559), .A2(n5558), .ZN(n8508) );
  NAND2_X1 U5253 ( .A1(n8575), .A2(n4878), .ZN(n4877) );
  INV_X1 U5254 ( .A(n6598), .ZN(n8596) );
  NOR2_X1 U5255 ( .A1(n8627), .A2(n4847), .ZN(n4846) );
  INV_X1 U5256 ( .A(n6709), .ZN(n4847) );
  NAND2_X1 U5257 ( .A1(n5598), .A2(n4972), .ZN(n8620) );
  OR2_X1 U5258 ( .A1(n8638), .A2(n8380), .ZN(n4972) );
  OR2_X1 U5259 ( .A1(n8802), .A2(n8666), .ZN(n5597) );
  AND2_X1 U5260 ( .A1(n6707), .A2(n6709), .ZN(n8635) );
  AND2_X1 U5261 ( .A1(n8686), .A2(n6695), .ZN(n4849) );
  NAND2_X1 U5262 ( .A1(n4339), .A2(n4823), .ZN(n5343) );
  NAND2_X1 U5263 ( .A1(n8703), .A2(n8815), .ZN(n8705) );
  NOR2_X1 U5264 ( .A1(n7812), .A2(n4514), .ZN(n4513) );
  AND2_X1 U5265 ( .A1(n6678), .A2(n6676), .ZN(n7812) );
  NOR2_X1 U5266 ( .A1(n5235), .A2(n4844), .ZN(n4843) );
  INV_X1 U5267 ( .A(n6667), .ZN(n4844) );
  NAND2_X1 U5268 ( .A1(n7698), .A2(n7699), .ZN(n7697) );
  OR2_X1 U5269 ( .A1(n7668), .A2(n7669), .ZN(n7666) );
  AND4_X1 U5270 ( .A1(n5177), .A2(n5176), .A3(n5175), .A4(n5174), .ZN(n7691)
         );
  AND4_X1 U5271 ( .A1(n5215), .A2(n5214), .A3(n5213), .A4(n5212), .ZN(n7847)
         );
  INV_X1 U5272 ( .A(n5172), .ZN(n5170) );
  CLKBUF_X1 U5273 ( .A(n5648), .Z(n10033) );
  INV_X1 U5274 ( .A(n8768), .ZN(n8771) );
  NAND2_X1 U5275 ( .A1(n8769), .A2(n8840), .ZN(n8770) );
  NAND2_X1 U5276 ( .A1(n4499), .A2(n5205), .ZN(n8850) );
  NAND2_X1 U5277 ( .A1(n6840), .A2(n5787), .ZN(n4499) );
  AND2_X1 U5278 ( .A1(n10033), .A2(n7662), .ZN(n8861) );
  AND2_X1 U5279 ( .A1(n5633), .A2(n5637), .ZN(n10042) );
  OR2_X1 U5280 ( .A1(n5638), .A2(n5630), .ZN(n5633) );
  NAND2_X1 U5281 ( .A1(n5015), .A2(n4886), .ZN(n4885) );
  NAND2_X1 U5282 ( .A1(n5624), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5636) );
  CLKBUF_X1 U5283 ( .A(n5625), .Z(n5626) );
  INV_X1 U5284 ( .A(n5549), .ZN(n5552) );
  INV_X1 U5285 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5551) );
  OR2_X1 U5286 ( .A1(n5165), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5332) );
  OR2_X1 U5287 ( .A1(n5332), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5203) );
  CLKBUF_X1 U5288 ( .A(n5087), .Z(n5088) );
  OR2_X1 U5289 ( .A1(n9080), .A2(n4756), .ZN(n4475) );
  NAND2_X1 U5290 ( .A1(n5955), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6421) );
  INV_X1 U5291 ( .A(n6403), .ZN(n5955) );
  INV_X1 U5292 ( .A(n4311), .ZN(n4766) );
  AND2_X1 U5293 ( .A1(n6434), .A2(n6433), .ZN(n6454) );
  NAND2_X1 U5294 ( .A1(n6159), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6199) );
  AND2_X1 U5295 ( .A1(n8101), .A2(n9471), .ZN(n6497) );
  NAND2_X1 U5296 ( .A1(n4766), .A2(n4293), .ZN(n4765) );
  NAND2_X1 U5297 ( .A1(n5953), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U5298 ( .A1(n8208), .A2(n9124), .ZN(n4537) );
  INV_X1 U5299 ( .A(n8232), .ZN(n8187) );
  AND2_X1 U5300 ( .A1(n8075), .A2(n8074), .ZN(n8978) );
  OR2_X1 U5301 ( .A1(n9103), .A2(n8054), .ZN(n6491) );
  AND2_X1 U5302 ( .A1(n6349), .A2(n6348), .ZN(n9285) );
  CLKBUF_X1 U5303 ( .A(n6036), .Z(n8069) );
  OR2_X1 U5304 ( .A1(n8067), .A2(n7022), .ZN(n6016) );
  INV_X1 U5305 ( .A(n4892), .ZN(n4891) );
  OAI21_X1 U5306 ( .B1(n6238), .B2(n6006), .A(n5997), .ZN(n4892) );
  INV_X1 U5307 ( .A(n4890), .ZN(n4889) );
  OAI22_X1 U5308 ( .A1(n8067), .A2(n7542), .B1(n6055), .B2(n5996), .ZN(n4890)
         );
  AOI21_X1 U5309 ( .B1(n6932), .B2(n6968), .A(n4354), .ZN(n4670) );
  OR2_X1 U5310 ( .A1(n7516), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4662) );
  XNOR2_X1 U5311 ( .A(n4661), .B(n9860), .ZN(n9864) );
  NAND2_X1 U5312 ( .A1(n4747), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U5313 ( .A1(n5935), .A2(n4749), .ZN(n4747) );
  NAND2_X1 U5314 ( .A1(n4535), .A2(n4534), .ZN(n9352) );
  INV_X1 U5315 ( .A(n4655), .ZN(n4535) );
  NOR2_X1 U5316 ( .A1(n9389), .A2(n9631), .ZN(n4534) );
  NAND2_X1 U5317 ( .A1(n8065), .A2(n8064), .ZN(n9614) );
  OAI211_X1 U5318 ( .C1(n9620), .C2(n4318), .A(n4923), .B(n9349), .ZN(n4922)
         );
  AOI21_X1 U5319 ( .B1(n9348), .B2(n9347), .A(n9346), .ZN(n9349) );
  NAND2_X1 U5320 ( .A1(n4924), .A2(n9620), .ZN(n4923) );
  NOR2_X1 U5321 ( .A1(n9362), .A2(n9908), .ZN(n4926) );
  NAND2_X1 U5322 ( .A1(n4904), .A2(n9329), .ZN(n4903) );
  INV_X1 U5323 ( .A(n9337), .ZN(n4914) );
  NOR2_X1 U5324 ( .A1(n8159), .A2(n9339), .ZN(n9393) );
  INV_X1 U5325 ( .A(n9338), .ZN(n8159) );
  AND2_X1 U5326 ( .A1(n9433), .A2(n9300), .ZN(n4437) );
  NOR2_X1 U5327 ( .A1(n9450), .A2(n9663), .ZN(n9256) );
  INV_X1 U5328 ( .A(n9326), .ZN(n4909) );
  NAND2_X1 U5329 ( .A1(n4911), .A2(n8163), .ZN(n4910) );
  OR2_X1 U5330 ( .A1(n9675), .A2(n9291), .ZN(n9292) );
  OR2_X1 U5331 ( .A1(n4964), .A2(n4963), .ZN(n4962) );
  INV_X1 U5332 ( .A(n9293), .ZN(n4964) );
  AND2_X1 U5333 ( .A1(n8163), .A2(n9326), .ZN(n9479) );
  AND2_X1 U5334 ( .A1(n9678), .A2(n9287), .ZN(n9288) );
  AND2_X1 U5335 ( .A1(n9544), .A2(n4287), .ZN(n4944) );
  NAND2_X1 U5336 ( .A1(n4357), .A2(n4287), .ZN(n4943) );
  INV_X1 U5337 ( .A(n4943), .ZN(n4942) );
  INV_X1 U5338 ( .A(n4941), .ZN(n4940) );
  OAI21_X1 U5339 ( .B1(n4944), .B2(n4942), .A(n9513), .ZN(n4941) );
  NAND2_X1 U5340 ( .A1(n4290), .A2(n4335), .ZN(n4898) );
  NOR2_X1 U5341 ( .A1(n4327), .A2(n4932), .ZN(n4931) );
  AND2_X1 U5342 ( .A1(n9541), .A2(n8165), .ZN(n9572) );
  NAND2_X1 U5343 ( .A1(n9315), .A2(n9314), .ZN(n9590) );
  NAND2_X1 U5344 ( .A1(n4894), .A2(n4498), .ZN(n9313) );
  NOR2_X1 U5345 ( .A1(n7792), .A2(n4893), .ZN(n4498) );
  INV_X1 U5346 ( .A(n8006), .ZN(n4893) );
  NAND2_X1 U5347 ( .A1(n7790), .A2(n8013), .ZN(n4894) );
  AND4_X1 U5348 ( .A1(n6205), .A2(n6204), .A3(n6203), .A4(n6202), .ZN(n7791)
         );
  INV_X1 U5349 ( .A(n9347), .ZN(n9102) );
  INV_X1 U5350 ( .A(n6497), .ZN(n8226) );
  CLKBUF_X1 U5351 ( .A(n6874), .Z(n4446) );
  NAND2_X1 U5352 ( .A1(n6871), .A2(n6799), .ZN(n7416) );
  OR2_X1 U5353 ( .A1(n6873), .A2(n6497), .ZN(n7145) );
  OAI21_X1 U5354 ( .B1(n8256), .B2(n8089), .A(n8088), .ZN(n9604) );
  NAND2_X1 U5355 ( .A1(n8081), .A2(n8080), .ZN(n9610) );
  INV_X1 U5356 ( .A(n9618), .ZN(n4526) );
  AND2_X1 U5357 ( .A1(n6870), .A2(n6869), .ZN(n7147) );
  NAND2_X1 U5358 ( .A1(n6479), .A2(n7681), .ZN(n7149) );
  AND2_X1 U5359 ( .A1(n9772), .A2(n6466), .ZN(n5950) );
  INV_X1 U5360 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5959) );
  AND2_X1 U5361 ( .A1(n4971), .A2(n4966), .ZN(n4965) );
  INV_X1 U5362 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4966) );
  XNOR2_X1 U5363 ( .A(n5786), .B(n6512), .ZN(n8890) );
  XNOR2_X1 U5364 ( .A(n5512), .B(n5511), .ZN(n8898) );
  NAND2_X1 U5365 ( .A1(n5506), .A2(n5531), .ZN(n5512) );
  OR2_X1 U5366 ( .A1(n5529), .A2(n5527), .ZN(n5506) );
  NAND2_X1 U5367 ( .A1(n5944), .A2(n6463), .ZN(n4474) );
  NAND2_X1 U5368 ( .A1(n4745), .A2(n4743), .ZN(n5942) );
  AOI21_X1 U5369 ( .B1(n5939), .B2(n4744), .A(n4748), .ZN(n4743) );
  AND2_X1 U5370 ( .A1(n4748), .A2(n4746), .ZN(n4744) );
  OAI211_X1 U5371 ( .C1(n5935), .C2(n4748), .A(n5939), .B(n4742), .ZN(n5975)
         );
  OR2_X1 U5372 ( .A1(n4749), .A2(n4748), .ZN(n4742) );
  NAND2_X1 U5373 ( .A1(n4782), .A2(n5383), .ZN(n5406) );
  NAND2_X1 U5374 ( .A1(n5381), .A2(n5380), .ZN(n4782) );
  NAND2_X1 U5375 ( .A1(n4796), .A2(n5345), .ZN(n5363) );
  OAI21_X1 U5376 ( .B1(n5222), .B2(n4792), .A(n4790), .ZN(n5282) );
  OR2_X1 U5377 ( .A1(n6063), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6101) );
  NAND3_X1 U5378 ( .A1(n4776), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4777) );
  NAND3_X1 U5379 ( .A1(n4775), .A2(n4774), .A3(n4773), .ZN(n4778) );
  INV_X1 U5380 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4776) );
  INV_X1 U5381 ( .A(n4716), .ZN(n4715) );
  AOI21_X1 U5382 ( .B1(n4716), .B2(n4714), .A(n4713), .ZN(n4712) );
  INV_X1 U5383 ( .A(n5691), .ZN(n4713) );
  AND4_X1 U5384 ( .A1(n5234), .A2(n5233), .A3(n5232), .A4(n5231), .ZN(n7908)
         );
  NAND2_X1 U5385 ( .A1(n5252), .A2(n5251), .ZN(n8839) );
  AOI21_X1 U5386 ( .B1(n5769), .B2(n5770), .A(n4718), .ZN(n4717) );
  NOR2_X1 U5387 ( .A1(n8346), .A2(n8347), .ZN(n4718) );
  INV_X1 U5388 ( .A(n8815), .ZN(n8709) );
  AND2_X1 U5389 ( .A1(n5112), .A2(n5111), .ZN(n7393) );
  OR2_X1 U5390 ( .A1(n8392), .A2(n8563), .ZN(n8383) );
  AND2_X1 U5391 ( .A1(n5434), .A2(n5433), .ZN(n8371) );
  NAND2_X1 U5392 ( .A1(n5412), .A2(n5411), .ZN(n8796) );
  AND4_X1 U5393 ( .A1(n5296), .A2(n5295), .A3(n5294), .A4(n5293), .ZN(n8404)
         );
  AND2_X1 U5394 ( .A1(n5475), .A2(n5474), .ZN(n8564) );
  NAND2_X1 U5395 ( .A1(n5448), .A2(n5447), .ZN(n8786) );
  AND4_X1 U5396 ( .A1(n5261), .A2(n5260), .A3(n5259), .A4(n5258), .ZN(n7919)
         );
  OR2_X1 U5397 ( .A1(n8392), .A2(n8336), .ZN(n8381) );
  AND2_X1 U5398 ( .A1(n8762), .A2(n8411), .ZN(n4449) );
  INV_X1 U5399 ( .A(n8394), .ZN(n4451) );
  INV_X1 U5400 ( .A(n8389), .ZN(n8409) );
  INV_X1 U5401 ( .A(n8300), .ZN(n8411) );
  INV_X1 U5402 ( .A(n6759), .ZN(n4769) );
  AND2_X1 U5403 ( .A1(n6756), .A2(n6757), .ZN(n4770) );
  OAI21_X1 U5404 ( .B1(n7100), .B2(n6582), .A(n7839), .ZN(n6583) );
  INV_X1 U5405 ( .A(n8564), .ZN(n8598) );
  NAND2_X1 U5406 ( .A1(n7926), .A2(n7927), .ZN(n7925) );
  AND2_X1 U5407 ( .A1(n5911), .A2(n5913), .ZN(n8487) );
  OAI21_X1 U5408 ( .B1(n8256), .B2(n6549), .A(n6548), .ZN(n8737) );
  NAND2_X1 U5409 ( .A1(n6564), .A2(n6563), .ZN(n8746) );
  NAND2_X1 U5410 ( .A1(n8498), .A2(n10021), .ZN(n4822) );
  OAI21_X1 U5411 ( .B1(n5604), .B2(n4867), .A(n4864), .ZN(n8522) );
  NAND2_X1 U5412 ( .A1(n4588), .A2(n6557), .ZN(n8518) );
  OAI21_X1 U5413 ( .B1(n5826), .B2(n5525), .A(n6726), .ZN(n5548) );
  OR2_X1 U5414 ( .A1(n5249), .A2(n6808), .ZN(n5047) );
  OR2_X1 U5415 ( .A1(n4280), .A2(n6811), .ZN(n5048) );
  AND2_X1 U5416 ( .A1(n10029), .A2(n5836), .ZN(n8727) );
  NAND2_X2 U5417 ( .A1(n7178), .A2(n10041), .ZN(n10029) );
  AND2_X1 U5418 ( .A1(n10029), .A2(n10027), .ZN(n8531) );
  AND2_X1 U5419 ( .A1(n7889), .A2(n8900), .ZN(n10046) );
  OAI21_X1 U5420 ( .B1(n6457), .B2(n4761), .A(n4759), .ZN(n8960) );
  AOI21_X1 U5421 ( .B1(n4762), .B2(n4760), .A(n4383), .ZN(n4759) );
  INV_X1 U5422 ( .A(n4762), .ZN(n4761) );
  INV_X1 U5423 ( .A(n4313), .ZN(n4760) );
  AND2_X1 U5424 ( .A1(n6503), .A2(n9935), .ZN(n9837) );
  INV_X1 U5425 ( .A(n8970), .ZN(n9348) );
  INV_X1 U5426 ( .A(n9286), .ZN(n9287) );
  INV_X1 U5427 ( .A(n9021), .ZN(n9284) );
  INV_X1 U5428 ( .A(n9020), .ZN(n9279) );
  INV_X1 U5429 ( .A(n8008), .ZN(n9274) );
  OR2_X1 U5430 ( .A1(n8067), .A2(n7450), .ZN(n5979) );
  NAND2_X1 U5431 ( .A1(n4435), .A2(n4678), .ZN(n4677) );
  OR2_X1 U5432 ( .A1(n9250), .A2(n9249), .ZN(n4678) );
  NAND2_X1 U5433 ( .A1(n9253), .A2(n9879), .ZN(n4435) );
  OAI21_X1 U5434 ( .B1(n9253), .B2(n9252), .A(n9251), .ZN(n4674) );
  XNOR2_X1 U5435 ( .A(n9264), .B(n4305), .ZN(n9607) );
  AOI21_X1 U5436 ( .B1(n9401), .B2(n4947), .A(n4349), .ZN(n9361) );
  NOR2_X1 U5437 ( .A1(n4950), .A2(n4948), .ZN(n4947) );
  NAND2_X1 U5438 ( .A1(n4936), .A2(n7785), .ZN(n7786) );
  CLKBUF_X1 U5439 ( .A(n5991), .Z(n9444) );
  NAND2_X1 U5440 ( .A1(n6795), .A2(n9935), .ZN(n9814) );
  INV_X1 U5441 ( .A(n6870), .ZN(n6795) );
  AND2_X1 U5442 ( .A1(n6468), .A2(n6467), .ZN(n9759) );
  NAND2_X1 U5443 ( .A1(n9787), .A2(n4402), .ZN(n10116) );
  INV_X1 U5444 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n4402) );
  NOR2_X1 U5445 ( .A1(n10107), .A2(n10106), .ZN(n10105) );
  NAND2_X1 U5446 ( .A1(n10100), .A2(n10101), .ZN(n10099) );
  NAND2_X1 U5447 ( .A1(n10091), .A2(n10092), .ZN(n10090) );
  NAND2_X1 U5448 ( .A1(n4637), .A2(n4632), .ZN(n6634) );
  NAND2_X1 U5449 ( .A1(n6621), .A2(n6727), .ZN(n4637) );
  INV_X1 U5450 ( .A(n8179), .ZN(n4572) );
  AND2_X1 U5451 ( .A1(n7985), .A2(n8066), .ZN(n4573) );
  AOI21_X1 U5452 ( .B1(n4631), .B2(n4332), .A(n4630), .ZN(n4629) );
  NAND2_X1 U5453 ( .A1(n6698), .A2(n6699), .ZN(n4630) );
  AND2_X1 U5454 ( .A1(n9541), .A2(n8066), .ZN(n4567) );
  NAND2_X1 U5455 ( .A1(n8012), .A2(n4569), .ZN(n4568) );
  NOR2_X1 U5456 ( .A1(n4570), .A2(n8066), .ZN(n4569) );
  INV_X1 U5457 ( .A(n8165), .ZN(n4570) );
  AND2_X1 U5458 ( .A1(n8559), .A2(n6720), .ZN(n4638) );
  NAND2_X1 U5459 ( .A1(n8179), .A2(n9810), .ZN(n4423) );
  NAND3_X1 U5460 ( .A1(n8042), .A2(n8040), .A3(n8041), .ZN(n4557) );
  OR3_X1 U5461 ( .A1(n8146), .A2(n8198), .A3(n8033), .ZN(n8042) );
  NOR2_X1 U5462 ( .A1(n7999), .A2(n7990), .ZN(n8125) );
  OAI21_X1 U5463 ( .B1(n4624), .B2(n4325), .A(n4810), .ZN(n4809) );
  AND2_X1 U5464 ( .A1(n6737), .A2(n6732), .ZN(n4810) );
  AND2_X1 U5465 ( .A1(n8559), .A2(n4295), .ZN(n4836) );
  INV_X1 U5466 ( .A(n6704), .ZN(n4835) );
  INV_X1 U5467 ( .A(n5436), .ZN(n4601) );
  INV_X1 U5468 ( .A(n6685), .ZN(n4829) );
  NAND2_X1 U5469 ( .A1(n8434), .A2(n10035), .ZN(n6620) );
  NOR2_X1 U5470 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5348) );
  INV_X1 U5471 ( .A(n4412), .ZN(n4411) );
  OAI21_X1 U5472 ( .B1(n8046), .B2(n8045), .A(n9380), .ZN(n4412) );
  NAND2_X1 U5473 ( .A1(n7743), .A2(n9805), .ZN(n7983) );
  NAND2_X1 U5474 ( .A1(n5385), .A2(n5384), .ZN(n5404) );
  INV_X1 U5475 ( .A(SI_19_), .ZN(n5384) );
  INV_X1 U5476 ( .A(n5302), .ZN(n4519) );
  INV_X1 U5477 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5326) );
  INV_X1 U5478 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5325) );
  INV_X1 U5479 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5264) );
  OAI21_X1 U5480 ( .B1(n4277), .B2(n4431), .A(n4430), .ZN(n5140) );
  INV_X1 U5481 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4431) );
  NAND2_X1 U5482 ( .A1(n4276), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4430) );
  INV_X1 U5483 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5103) );
  INV_X1 U5485 ( .A(n5777), .ZN(n5790) );
  XNOR2_X1 U5486 ( .A(n7472), .B(n5670), .ZN(n5659) );
  INV_X1 U5487 ( .A(n6570), .ZN(n6572) );
  AND2_X2 U5488 ( .A1(n6752), .A2(n5648), .ZN(n5651) );
  NOR2_X1 U5489 ( .A1(n8762), .A2(n8769), .ZN(n4683) );
  NOR2_X1 U5490 ( .A1(n6733), .A2(n4682), .ZN(n4681) );
  INV_X1 U5491 ( .A(n4683), .ZN(n4682) );
  INV_X1 U5492 ( .A(n4875), .ZN(n4874) );
  OAI21_X1 U5493 ( .B1(n4878), .B2(n4876), .A(n4880), .ZN(n4875) );
  INV_X1 U5494 ( .A(n4289), .ZN(n4876) );
  NAND2_X1 U5495 ( .A1(n6598), .A2(n4859), .ZN(n4855) );
  INV_X1 U5496 ( .A(n4856), .ZN(n4853) );
  NOR2_X1 U5497 ( .A1(n5397), .A2(n5396), .ZN(n4439) );
  INV_X1 U5498 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5357) );
  OR2_X1 U5499 ( .A1(n5358), .A2(n5357), .ZN(n5374) );
  AND2_X1 U5500 ( .A1(n4840), .A2(n4593), .ZN(n4592) );
  NOR2_X1 U5501 ( .A1(n4845), .A2(n4841), .ZN(n4840) );
  NAND2_X1 U5502 ( .A1(n4843), .A2(n7702), .ZN(n4593) );
  INV_X1 U5503 ( .A(n6673), .ZN(n4841) );
  INV_X1 U5504 ( .A(n4843), .ZN(n4594) );
  INV_X1 U5505 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5254) );
  OR2_X1 U5506 ( .A1(n5255), .A2(n5254), .ZN(n5276) );
  NAND2_X1 U5507 ( .A1(n4634), .A2(n4278), .ZN(n6617) );
  NAND2_X1 U5508 ( .A1(n5018), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5567) );
  INV_X1 U5509 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U5510 ( .A1(n4701), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5623) );
  XNOR2_X1 U5511 ( .A(n4605), .B(P2_IR_REG_1__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U5512 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4605) );
  OAI22_X1 U5513 ( .A1(n4756), .A2(n6228), .B1(n9053), .B2(n9052), .ZN(n4755)
         );
  AND2_X1 U5514 ( .A1(n6363), .A2(n4308), .ZN(n4738) );
  NAND2_X1 U5515 ( .A1(n6138), .A2(n6137), .ZN(n4471) );
  INV_X1 U5516 ( .A(n4729), .ZN(n4728) );
  INV_X1 U5517 ( .A(n4732), .ZN(n4466) );
  NOR2_X1 U5518 ( .A1(n6198), .A2(n4541), .ZN(n4540) );
  NAND2_X1 U5519 ( .A1(n4475), .A2(n4298), .ZN(n9014) );
  NAND2_X1 U5520 ( .A1(n4420), .A2(n4419), .ZN(n8182) );
  NOR2_X1 U5521 ( .A1(n9571), .A2(n4421), .ZN(n4420) );
  NOR2_X1 U5522 ( .A1(n4562), .A2(n8077), .ZN(n4561) );
  INV_X1 U5523 ( .A(n8208), .ZN(n4562) );
  OR2_X1 U5524 ( .A1(n6853), .A2(n4559), .ZN(n6079) );
  OR2_X1 U5525 ( .A1(n6969), .A2(n6889), .ZN(n6970) );
  AND2_X1 U5526 ( .A1(n6233), .A2(n6232), .ZN(n6267) );
  AND2_X1 U5527 ( .A1(n9362), .A2(n4286), .ZN(n4924) );
  INV_X1 U5528 ( .A(n4908), .ZN(n4904) );
  NOR2_X1 U5529 ( .A1(n9022), .A2(n4544), .ZN(n4543) );
  INV_X1 U5530 ( .A(n6282), .ZN(n5953) );
  AND2_X1 U5531 ( .A1(n9540), .A2(n4657), .ZN(n4656) );
  INV_X1 U5532 ( .A(n4935), .ZN(n4932) );
  NOR2_X1 U5533 ( .A1(n9701), .A2(n9708), .ZN(n4657) );
  AND2_X1 U5534 ( .A1(n8017), .A2(n8016), .ZN(n9312) );
  NOR2_X1 U5535 ( .A1(n7653), .A2(n7589), .ZN(n4653) );
  NOR2_X1 U5536 ( .A1(n6161), .A2(n6160), .ZN(n6159) );
  OR2_X1 U5537 ( .A1(n8004), .A2(n9889), .ZN(n7735) );
  AND2_X1 U5538 ( .A1(n7440), .A2(n7437), .ZN(n7427) );
  NAND2_X1 U5539 ( .A1(n7412), .A2(n4288), .ZN(n4648) );
  OAI21_X1 U5540 ( .B1(n7454), .B2(n9140), .A(n6872), .ZN(n8118) );
  NAND2_X1 U5541 ( .A1(n9311), .A2(n4955), .ZN(n4954) );
  INV_X1 U5542 ( .A(n9309), .ZN(n4955) );
  NAND2_X1 U5543 ( .A1(n9419), .A2(n4651), .ZN(n4650) );
  NOR2_X2 U5544 ( .A1(n9491), .A2(n9675), .ZN(n9482) );
  NAND2_X1 U5545 ( .A1(n7402), .A2(n8117), .ZN(n8169) );
  INV_X1 U5546 ( .A(n8101), .ZN(n8216) );
  NAND2_X1 U5547 ( .A1(n5535), .A2(n5534), .ZN(n5783) );
  OR2_X1 U5548 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  OR2_X1 U5549 ( .A1(n5529), .A2(n5528), .ZN(n5535) );
  NOR3_X1 U5550 ( .A1(n5936), .A2(P1_IR_REG_9__SCAN_IN), .A3(
        P1_IR_REG_19__SCAN_IN), .ZN(n4741) );
  NOR2_X1 U5551 ( .A1(n5936), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n4749) );
  INV_X1 U5552 ( .A(n5379), .ZN(n5380) );
  XNOR2_X1 U5553 ( .A(n5382), .B(SI_18_), .ZN(n5379) );
  XNOR2_X1 U5554 ( .A(n5300), .B(SI_14_), .ZN(n5299) );
  NAND2_X1 U5555 ( .A1(n5265), .A2(n10216), .ZN(n5283) );
  INV_X1 U5556 ( .A(n5239), .ZN(n4793) );
  INV_X1 U5557 ( .A(n4791), .ZN(n4790) );
  OAI21_X1 U5558 ( .B1(n4794), .B2(n4792), .A(n5262), .ZN(n4791) );
  NAND2_X1 U5559 ( .A1(n5935), .A2(n5934), .ZN(n6194) );
  INV_X1 U5560 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5933) );
  INV_X1 U5561 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6081) );
  XNOR2_X1 U5562 ( .A(n5114), .B(SI_5_), .ZN(n5116) );
  INV_X1 U5563 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4773) );
  INV_X1 U5564 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4775) );
  INV_X1 U5565 ( .A(SI_13_), .ZN(n10216) );
  OR2_X1 U5566 ( .A1(n8270), .A2(n8271), .ZN(n8316) );
  INV_X1 U5567 ( .A(n7346), .ZN(n4714) );
  NAND2_X1 U5568 ( .A1(n4722), .A2(n4721), .ZN(n4720) );
  INV_X1 U5569 ( .A(n5769), .ZN(n4721) );
  OR2_X1 U5570 ( .A1(n4320), .A2(n4723), .ZN(n4722) );
  NAND2_X1 U5571 ( .A1(n4440), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5358) );
  INV_X1 U5572 ( .A(n5337), .ZN(n4440) );
  OR2_X1 U5573 ( .A1(n4404), .A2(n5770), .ZN(n8279) );
  NAND2_X1 U5574 ( .A1(n4404), .A2(n5770), .ZN(n8343) );
  BUF_X1 U5575 ( .A(n8287), .Z(n4447) );
  NAND2_X1 U5576 ( .A1(n8297), .A2(n4709), .ZN(n4708) );
  INV_X1 U5577 ( .A(n5758), .ZN(n4709) );
  CLKBUF_X1 U5578 ( .A(n7088), .Z(n4416) );
  NAND2_X1 U5579 ( .A1(n5275), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5316) );
  INV_X1 U5580 ( .A(n5276), .ZN(n5275) );
  INV_X1 U5581 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5314) );
  NOR2_X1 U5582 ( .A1(n4627), .A2(n6749), .ZN(n4626) );
  NOR2_X1 U5583 ( .A1(n6738), .A2(n8745), .ZN(n4805) );
  AND2_X1 U5584 ( .A1(n5547), .A2(n5546), .ZN(n8501) );
  AND2_X1 U5585 ( .A1(n5420), .A2(n5419), .ZN(n8291) );
  OR2_X1 U5586 ( .A1(n5147), .A2(n7250), .ZN(n5077) );
  OR2_X1 U5587 ( .A1(n5074), .A2(n5858), .ZN(n5027) );
  OR2_X1 U5588 ( .A1(n5074), .A2(n5005), .ZN(n5013) );
  NOR2_X1 U5589 ( .A1(n7256), .A2(n7257), .ZN(n7255) );
  OR2_X1 U5590 ( .A1(n7196), .A2(n4323), .ZN(n4613) );
  OR2_X1 U5591 ( .A1(n5900), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4621) );
  AND2_X1 U5592 ( .A1(n5247), .A2(n5246), .ZN(n5269) );
  NOR2_X1 U5593 ( .A1(n8457), .A2(n8456), .ZN(n8455) );
  AND2_X1 U5594 ( .A1(n8470), .A2(n4814), .ZN(n5909) );
  NAND2_X1 U5595 ( .A1(n5908), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4814) );
  NAND2_X1 U5596 ( .A1(n8523), .A2(n7940), .ZN(n8510) );
  OAI21_X1 U5597 ( .B1(n4838), .B2(n4585), .A(n4582), .ZN(n8494) );
  AOI21_X1 U5598 ( .B1(n4586), .B2(n4584), .A(n4583), .ZN(n4582) );
  INV_X1 U5599 ( .A(n6737), .ZN(n4583) );
  AND2_X1 U5600 ( .A1(n5560), .A2(n8508), .ZN(n8525) );
  AND2_X1 U5601 ( .A1(n8541), .A2(n4679), .ZN(n8523) );
  AND2_X1 U5602 ( .A1(n4681), .A2(n4680), .ZN(n4679) );
  NAND2_X1 U5603 ( .A1(n4838), .A2(n4837), .ZN(n4588) );
  AND2_X1 U5604 ( .A1(n5524), .A2(n5523), .ZN(n8250) );
  NAND2_X1 U5605 ( .A1(n8762), .A2(n8250), .ZN(n6726) );
  NAND2_X1 U5606 ( .A1(n8541), .A2(n4681), .ZN(n8524) );
  NAND2_X1 U5607 ( .A1(n8541), .A2(n8545), .ZN(n8542) );
  AND2_X1 U5608 ( .A1(n5499), .A2(n5482), .ZN(n8560) );
  NAND2_X1 U5609 ( .A1(n4439), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5427) );
  OR2_X1 U5610 ( .A1(n5427), .A2(n8299), .ZN(n5450) );
  NOR2_X1 U5611 ( .A1(n4983), .A2(n8796), .ZN(n8621) );
  NAND2_X1 U5612 ( .A1(n4508), .A2(n5594), .ZN(n4504) );
  INV_X1 U5613 ( .A(n4506), .ZN(n4505) );
  NAND2_X1 U5614 ( .A1(n5372), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5397) );
  INV_X1 U5615 ( .A(n5374), .ZN(n5372) );
  INV_X1 U5616 ( .A(n4439), .ZN(n5413) );
  OR2_X1 U5617 ( .A1(n4849), .A2(n4599), .ZN(n4598) );
  INV_X1 U5618 ( .A(n6616), .ZN(n4599) );
  CLKBUF_X1 U5619 ( .A(n8692), .Z(n4403) );
  NAND2_X1 U5620 ( .A1(n4403), .A2(n4871), .ZN(n8684) );
  NOR2_X2 U5621 ( .A1(n8705), .A2(n8811), .ZN(n8677) );
  NAND2_X1 U5622 ( .A1(n4696), .A2(n7899), .ZN(n4695) );
  INV_X1 U5623 ( .A(n4698), .ZN(n4696) );
  NOR2_X1 U5624 ( .A1(n7730), .A2(n4697), .ZN(n7861) );
  INV_X1 U5625 ( .A(n4699), .ZN(n4697) );
  NAND2_X1 U5626 ( .A1(n5210), .A2(n5209), .ZN(n5229) );
  INV_X1 U5627 ( .A(n5208), .ZN(n5210) );
  AOI21_X1 U5628 ( .B1(n5583), .B2(n7669), .A(n4343), .ZN(n4882) );
  NAND2_X1 U5629 ( .A1(n5148), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5172) );
  INV_X1 U5630 ( .A(n5150), .ZN(n5148) );
  NOR2_X1 U5631 ( .A1(n7363), .A2(n8860), .ZN(n4438) );
  AND2_X1 U5632 ( .A1(n6654), .A2(n6655), .ZN(n7623) );
  INV_X1 U5633 ( .A(n5576), .ZN(n5577) );
  OR2_X1 U5634 ( .A1(n7238), .A2(n4635), .ZN(n7376) );
  NOR2_X2 U5635 ( .A1(n7376), .A2(n7382), .ZN(n7377) );
  AND2_X1 U5636 ( .A1(n5663), .A2(n4306), .ZN(n4581) );
  OR2_X1 U5637 ( .A1(n5845), .A2(n5890), .ZN(n8336) );
  NAND2_X1 U5638 ( .A1(n6617), .A2(n7054), .ZN(n7235) );
  CLKBUF_X1 U5639 ( .A(n6588), .Z(n6995) );
  AND2_X1 U5640 ( .A1(n10042), .A2(n10140), .ZN(n5640) );
  NAND2_X1 U5641 ( .A1(n5604), .A2(n4864), .ZN(n4863) );
  NAND2_X1 U5642 ( .A1(n4864), .A2(n4867), .ZN(n4862) );
  NAND2_X1 U5643 ( .A1(n8749), .A2(n8747), .ZN(n4694) );
  INV_X1 U5644 ( .A(n4822), .ZN(n4399) );
  NAND2_X1 U5645 ( .A1(n8748), .A2(n8497), .ZN(n4604) );
  NOR2_X1 U5646 ( .A1(n6603), .A2(n8849), .ZN(n4515) );
  NAND2_X1 U5647 ( .A1(n8595), .A2(n6704), .ZN(n8582) );
  AND2_X1 U5648 ( .A1(n5335), .A2(n5334), .ZN(n8815) );
  INV_X1 U5649 ( .A(n8861), .ZN(n8816) );
  NOR2_X1 U5650 ( .A1(n5639), .A2(n5793), .ZN(n5643) );
  XNOR2_X1 U5651 ( .A(n5632), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5637) );
  XNOR2_X1 U5652 ( .A(n5621), .B(P2_IR_REG_25__SCAN_IN), .ZN(n5638) );
  CLKBUF_X1 U5653 ( .A(n5617), .Z(n5618) );
  XNOR2_X1 U5654 ( .A(n5623), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5605) );
  OR2_X1 U5655 ( .A1(n5332), .A2(n5331), .ZN(n5620) );
  AND2_X1 U5656 ( .A1(n5290), .A2(n5309), .ZN(n5902) );
  NOR2_X2 U5657 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4868) );
  AND2_X2 U5658 ( .A1(n5045), .A2(n5071), .ZN(n7186) );
  AND2_X1 U5659 ( .A1(n4460), .A2(n6110), .ZN(n4459) );
  OR2_X1 U5660 ( .A1(n7166), .A2(n4314), .ZN(n4460) );
  INV_X1 U5661 ( .A(n6113), .ZN(n6109) );
  NOR2_X1 U5662 ( .A1(n4763), .A2(n9099), .ZN(n4762) );
  INV_X1 U5663 ( .A(n4765), .ZN(n4763) );
  AND2_X1 U5664 ( .A1(n4754), .A2(n4477), .ZN(n4476) );
  NAND2_X1 U5665 ( .A1(n4479), .A2(n4478), .ZN(n4477) );
  INV_X1 U5666 ( .A(n4755), .ZN(n4754) );
  INV_X1 U5667 ( .A(n6212), .ZN(n4478) );
  NAND2_X1 U5668 ( .A1(n5954), .A2(n4304), .ZN(n6403) );
  OR2_X1 U5669 ( .A1(n6342), .A2(n9094), .ZN(n6344) );
  INV_X1 U5670 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7656) );
  AOI21_X1 U5671 ( .B1(n4738), .B2(n4736), .A(n4735), .ZN(n4734) );
  INV_X1 U5672 ( .A(n9045), .ZN(n4735) );
  INV_X1 U5673 ( .A(n6355), .ZN(n4736) );
  INV_X1 U5674 ( .A(n4738), .ZN(n4737) );
  INV_X1 U5675 ( .A(n7166), .ZN(n4463) );
  NAND2_X1 U5676 ( .A1(n6311), .A2(n6275), .ZN(n9026) );
  NAND2_X1 U5677 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6092) );
  NAND2_X1 U5678 ( .A1(n4471), .A2(n6153), .ZN(n7649) );
  OR2_X1 U5679 ( .A1(n4471), .A2(n6153), .ZN(n7650) );
  NAND2_X1 U5680 ( .A1(n6154), .A2(n7652), .ZN(n4469) );
  NAND2_X1 U5681 ( .A1(n9030), .A2(n6322), .ZN(n8943) );
  NAND2_X1 U5682 ( .A1(n4758), .A2(n6228), .ZN(n8999) );
  NOR2_X1 U5683 ( .A1(n9083), .A2(n4725), .ZN(n4724) );
  INV_X1 U5684 ( .A(n6193), .ZN(n4725) );
  NAND2_X1 U5685 ( .A1(n7776), .A2(n7775), .ZN(n4726) );
  NAND2_X1 U5686 ( .A1(n6159), .A2(n4540), .ZN(n6218) );
  NAND2_X1 U5687 ( .A1(n6011), .A2(n8965), .ZN(n6012) );
  AND2_X1 U5688 ( .A1(n5995), .A2(n5994), .ZN(n6948) );
  OR2_X1 U5689 ( .A1(n6047), .A2(n4446), .ZN(n5995) );
  OAI22_X1 U5690 ( .A1(n6952), .A2(n8969), .B1(n4433), .B2(n4457), .ZN(n6028)
         );
  AND2_X1 U5691 ( .A1(n8943), .A2(n8944), .ZN(n9090) );
  OR2_X1 U5692 ( .A1(n6254), .A2(n8927), .ZN(n6282) );
  AND2_X1 U5693 ( .A1(n9014), .A2(n9013), .ZN(n9113) );
  AND2_X1 U5694 ( .A1(n8091), .A2(n8090), .ZN(n8189) );
  AOI21_X1 U5695 ( .B1(n8150), .B2(n4443), .A(n8206), .ZN(n8152) );
  AND2_X1 U5696 ( .A1(n9380), .A2(n9338), .ZN(n4443) );
  OR3_X1 U5697 ( .A1(n9336), .A2(n9335), .A3(n8148), .ZN(n8149) );
  AND2_X1 U5698 ( .A1(n8060), .A2(n8059), .ZN(n8970) );
  OR2_X1 U5699 ( .A1(n8979), .A2(n8054), .ZN(n8060) );
  AND2_X1 U5700 ( .A1(n6428), .A2(n6427), .ZN(n9302) );
  AND2_X1 U5701 ( .A1(n6330), .A2(n6329), .ZN(n9286) );
  AND3_X1 U5702 ( .A1(n6289), .A2(n6288), .A3(n6287), .ZN(n9020) );
  INV_X1 U5703 ( .A(n8054), .ZN(n7968) );
  AND4_X1 U5704 ( .A1(n6242), .A2(n6241), .A3(n6240), .A4(n6239), .ZN(n8008)
         );
  AND4_X1 U5705 ( .A1(n6223), .A2(n6222), .A3(n6221), .A4(n6220), .ZN(n9056)
         );
  AND4_X1 U5706 ( .A1(n6185), .A2(n6184), .A3(n6183), .A4(n6182), .ZN(n7744)
         );
  AND4_X1 U5707 ( .A1(n6148), .A2(n6147), .A3(n6146), .A4(n6145), .ZN(n7596)
         );
  AND4_X1 U5708 ( .A1(n6128), .A2(n6127), .A3(n6126), .A4(n6125), .ZN(n7441)
         );
  NAND2_X1 U5709 ( .A1(n6970), .A2(n6971), .ZN(n6928) );
  NAND2_X1 U5710 ( .A1(n6966), .A2(n6932), .ZN(n4668) );
  OAI21_X1 U5711 ( .B1(n4665), .B2(n4666), .A(n4664), .ZN(n9142) );
  INV_X1 U5712 ( .A(n4671), .ZN(n4665) );
  NAND2_X1 U5713 ( .A1(n4434), .A2(n4384), .ZN(n9209) );
  INV_X1 U5714 ( .A(n7513), .ZN(n4434) );
  NOR2_X1 U5715 ( .A1(n7522), .A2(n7521), .ZN(n9199) );
  NOR2_X1 U5716 ( .A1(n4661), .A2(n9204), .ZN(n4660) );
  INV_X1 U5717 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9022) );
  AND2_X1 U5718 ( .A1(n9366), .A2(n9629), .ZN(n9367) );
  NAND2_X1 U5719 ( .A1(n4951), .A2(n8061), .ZN(n4950) );
  INV_X1 U5720 ( .A(n4954), .ZN(n4951) );
  INV_X1 U5721 ( .A(n9403), .ZN(n4948) );
  AND2_X1 U5722 ( .A1(n8052), .A2(n7963), .ZN(n9376) );
  OR2_X1 U5723 ( .A1(n9309), .A2(n4358), .ZN(n4956) );
  NAND2_X1 U5724 ( .A1(n9400), .A2(n9403), .ZN(n4957) );
  AND2_X1 U5725 ( .A1(n6484), .A2(n6439), .ZN(n9409) );
  AND2_X1 U5726 ( .A1(n6437), .A2(n6436), .ZN(n9407) );
  AOI21_X1 U5727 ( .B1(n4961), .B2(n4959), .A(n4355), .ZN(n4958) );
  INV_X1 U5728 ( .A(n4307), .ZN(n4959) );
  NAND2_X1 U5729 ( .A1(n5954), .A2(n4546), .ZN(n6401) );
  OR2_X1 U5730 ( .A1(n6344), .A2(n8954), .ZN(n6366) );
  AOI21_X1 U5731 ( .B1(n4353), .B2(n4492), .A(n4490), .ZN(n9497) );
  NOR2_X1 U5732 ( .A1(n9322), .A2(n4491), .ZN(n4490) );
  INV_X1 U5733 ( .A(n9323), .ZN(n4491) );
  AND2_X1 U5734 ( .A1(n8162), .A2(n9324), .ZN(n9496) );
  NAND2_X1 U5735 ( .A1(n5953), .A2(n4543), .ZN(n6298) );
  AND2_X1 U5736 ( .A1(n9594), .A2(n4656), .ZN(n9536) );
  NAND2_X1 U5737 ( .A1(n9594), .A2(n4657), .ZN(n9559) );
  NAND2_X1 U5738 ( .A1(n9590), .A2(n4902), .ZN(n9542) );
  NAND2_X1 U5739 ( .A1(n4933), .A2(n4935), .ZN(n9552) );
  NAND2_X1 U5740 ( .A1(n9594), .A2(n9581), .ZN(n9577) );
  AND4_X1 U5741 ( .A1(n6166), .A2(n6165), .A3(n6164), .A4(n6163), .ZN(n7778)
         );
  NOR2_X1 U5742 ( .A1(n9810), .A2(n4929), .ZN(n4928) );
  INV_X1 U5743 ( .A(n7750), .ZN(n4929) );
  NAND2_X1 U5744 ( .A1(n7414), .A2(n4653), .ZN(n9901) );
  AND2_X1 U5745 ( .A1(n7414), .A2(n4300), .ZN(n9816) );
  OR2_X1 U5746 ( .A1(n6143), .A2(n7656), .ZN(n6161) );
  INV_X1 U5747 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6160) );
  AND2_X1 U5748 ( .A1(n9888), .A2(n8109), .ZN(n9887) );
  AND2_X1 U5749 ( .A1(n8175), .A2(n8109), .ZN(n9889) );
  INV_X1 U5750 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6122) );
  OR2_X1 U5751 ( .A1(n6123), .A2(n6122), .ZN(n6143) );
  AND2_X1 U5752 ( .A1(n7535), .A2(n7445), .ZN(n4647) );
  NAND2_X1 U5753 ( .A1(n9135), .A2(n7445), .ZN(n7986) );
  NAND2_X1 U5754 ( .A1(n4536), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6094) );
  INV_X1 U5755 ( .A(n6092), .ZN(n4536) );
  NAND2_X1 U5756 ( .A1(n5952), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6123) );
  INV_X1 U5757 ( .A(n6094), .ZN(n5952) );
  NOR2_X1 U5758 ( .A1(n4648), .A2(n7538), .ZN(n7533) );
  AOI21_X1 U5759 ( .B1(n7994), .B2(n7604), .A(n7404), .ZN(n9907) );
  NAND2_X1 U5760 ( .A1(n7402), .A2(n7403), .ZN(n7994) );
  NAND2_X1 U5761 ( .A1(n6779), .A2(n6780), .ZN(n7403) );
  AND2_X1 U5762 ( .A1(n8118), .A2(n8116), .ZN(n6779) );
  NOR2_X1 U5763 ( .A1(n7158), .A2(n7541), .ZN(n7151) );
  OR2_X1 U5764 ( .A1(n9615), .A2(n9977), .ZN(n4523) );
  NOR2_X1 U5765 ( .A1(n4309), .A2(n4525), .ZN(n4524) );
  NAND2_X1 U5766 ( .A1(n4916), .A2(n4915), .ZN(n9404) );
  NAND2_X1 U5767 ( .A1(n4916), .A2(n9334), .ZN(n9421) );
  INV_X1 U5768 ( .A(n9256), .ZN(n9451) );
  OR2_X1 U5769 ( .A1(n8066), .A2(n8216), .ZN(n9936) );
  INV_X1 U5770 ( .A(n9977), .ZN(n9986) );
  NAND2_X1 U5771 ( .A1(n7412), .A2(n9836), .ZN(n9915) );
  OR2_X1 U5772 ( .A1(n7149), .A2(n8216), .ZN(n9977) );
  AND2_X1 U5773 ( .A1(n7145), .A2(n6798), .ZN(n6871) );
  XNOR2_X1 U5774 ( .A(n6542), .B(n6517), .ZN(n8079) );
  XNOR2_X1 U5775 ( .A(n6561), .B(n6560), .ZN(n8265) );
  XNOR2_X1 U5776 ( .A(n5783), .B(n5782), .ZN(n8895) );
  XNOR2_X1 U5777 ( .A(n5529), .B(n5527), .ZN(n8901) );
  OAI21_X1 U5778 ( .B1(n5424), .B2(n4529), .A(n4531), .ZN(n5490) );
  NAND2_X1 U5779 ( .A1(n4797), .A2(n4800), .ZN(n5477) );
  NAND2_X1 U5780 ( .A1(n5439), .A2(n4803), .ZN(n4797) );
  OAI21_X1 U5781 ( .B1(n5439), .B2(n5438), .A(n5442), .ZN(n5460) );
  OR2_X1 U5782 ( .A1(n6276), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U5783 ( .A1(n4520), .A2(n5302), .ZN(n5324) );
  NAND2_X1 U5784 ( .A1(n5284), .A2(n4521), .ZN(n4520) );
  NAND2_X1 U5785 ( .A1(n4487), .A2(n5239), .ZN(n4486) );
  NAND2_X1 U5786 ( .A1(n5222), .A2(n4794), .ZN(n4487) );
  XNOR2_X1 U5787 ( .A(n5202), .B(n4979), .ZN(n6840) );
  XNOR2_X1 U5788 ( .A(n5195), .B(n5194), .ZN(n6842) );
  INV_X1 U5789 ( .A(SI_3_), .ZN(n4767) );
  OAI22_X1 U5790 ( .A1(n6022), .A2(n4663), .B1(P1_IR_REG_31__SCAN_IN), .B2(
        P1_IR_REG_2__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U5791 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4663) );
  AND2_X1 U5792 ( .A1(n4753), .A2(n4752), .ZN(n6022) );
  NOR2_X1 U5793 ( .A1(n10111), .A2(n9790), .ZN(n9791) );
  INV_X1 U5794 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10184) );
  AND2_X1 U5796 ( .A1(n7460), .A2(n5685), .ZN(n4716) );
  AND2_X1 U5797 ( .A1(n7345), .A2(n5685), .ZN(n7461) );
  AND4_X1 U5798 ( .A1(n5321), .A2(n5320), .A3(n5319), .A4(n5318), .ZN(n8324)
         );
  AND4_X1 U5799 ( .A1(n5193), .A2(n5192), .A3(n5191), .A4(n5190), .ZN(n7767)
         );
  NAND2_X1 U5800 ( .A1(n4707), .A2(n5758), .ZN(n8298) );
  NAND2_X1 U5801 ( .A1(n4447), .A2(n4710), .ZN(n4707) );
  NAND2_X1 U5802 ( .A1(n4691), .A2(n4690), .ZN(n7099) );
  NAND2_X1 U5803 ( .A1(n4689), .A2(n4329), .ZN(n4691) );
  NAND2_X1 U5804 ( .A1(n5851), .A2(n8905), .ZN(n4690) );
  NAND2_X1 U5805 ( .A1(n4447), .A2(n5753), .ZN(n8358) );
  NAND2_X1 U5806 ( .A1(n5272), .A2(n5271), .ZN(n8833) );
  CLKBUF_X1 U5807 ( .A(n7347), .Z(n4429) );
  NAND2_X1 U5808 ( .A1(n5505), .A2(n5504), .ZN(n8571) );
  INV_X2 U5809 ( .A(P2_U3966), .ZN(n8436) );
  OAI21_X1 U5810 ( .B1(n7186), .B2(P2_REG2_REG_2__SCAN_IN), .A(n4813), .ZN(
        n7184) );
  NOR2_X1 U5811 ( .A1(n7184), .A2(n7185), .ZN(n7183) );
  AOI21_X1 U5812 ( .B1(n7259), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7255), .ZN(
        n7185) );
  NOR2_X1 U5813 ( .A1(n7183), .A2(n4812), .ZN(n7292) );
  INV_X1 U5814 ( .A(n4813), .ZN(n4812) );
  NOR2_X1 U5815 ( .A1(n4618), .A2(n4285), .ZN(n7307) );
  NOR2_X1 U5816 ( .A1(n7307), .A2(n7306), .ZN(n7305) );
  NAND2_X1 U5817 ( .A1(n4616), .A2(n4615), .ZN(n7319) );
  INV_X1 U5818 ( .A(n7318), .ZN(n4614) );
  AND2_X1 U5819 ( .A1(n4613), .A2(n4612), .ZN(n7207) );
  NOR2_X1 U5820 ( .A1(n7491), .A2(n4610), .ZN(n4607) );
  NAND2_X1 U5821 ( .A1(n4608), .A2(n4609), .ZN(n7492) );
  OR2_X1 U5822 ( .A1(n7870), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4820) );
  XNOR2_X1 U5823 ( .A(n5905), .B(n5904), .ZN(n8439) );
  NOR2_X1 U5824 ( .A1(n10012), .A2(n5913), .ZN(n10008) );
  OAI21_X1 U5825 ( .B1(n10044), .B2(n7839), .A(n5918), .ZN(n8480) );
  XNOR2_X1 U5826 ( .A(n5909), .B(n7486), .ZN(n8483) );
  NOR2_X1 U5827 ( .A1(n8483), .A2(n5378), .ZN(n8482) );
  OAI21_X1 U5828 ( .B1(n5915), .B2(n10012), .A(n4819), .ZN(n4818) );
  AOI21_X1 U5829 ( .B1(n5912), .B2(n10007), .A(n8487), .ZN(n4819) );
  INV_X1 U5830 ( .A(n8490), .ZN(n8743) );
  INV_X1 U5831 ( .A(n4877), .ZN(n8557) );
  INV_X1 U5832 ( .A(n8781), .ZN(n8579) );
  AND2_X1 U5833 ( .A1(n8600), .A2(n8599), .ZN(n8789) );
  AND2_X1 U5834 ( .A1(n8607), .A2(n6714), .ZN(n8597) );
  INV_X1 U5835 ( .A(n4688), .ZN(n4686) );
  NAND2_X1 U5836 ( .A1(n4851), .A2(n4856), .ZN(n8589) );
  OR2_X1 U5837 ( .A1(n8620), .A2(n4858), .ZN(n4851) );
  AND2_X1 U5838 ( .A1(n4860), .A2(n4861), .ZN(n8604) );
  NAND2_X1 U5839 ( .A1(n8620), .A2(n8627), .ZN(n4860) );
  NAND2_X1 U5840 ( .A1(n4848), .A2(n6709), .ZN(n8626) );
  NAND2_X1 U5841 ( .A1(n5395), .A2(n5394), .ZN(n8802) );
  NAND2_X1 U5842 ( .A1(n5343), .A2(n4849), .ZN(n8675) );
  NAND2_X1 U5843 ( .A1(n7891), .A2(n5298), .ZN(n4826) );
  NAND2_X1 U5844 ( .A1(n4511), .A2(n4512), .ZN(n7855) );
  NAND2_X1 U5845 ( .A1(n4842), .A2(n6673), .ZN(n7806) );
  NAND2_X1 U5846 ( .A1(n7697), .A2(n4843), .ZN(n4842) );
  NAND2_X1 U5847 ( .A1(n7697), .A2(n6667), .ZN(n7726) );
  NAND2_X1 U5848 ( .A1(n7666), .A2(n5583), .ZN(n7701) );
  INV_X1 U5849 ( .A(n8727), .ZN(n8681) );
  INV_X2 U5850 ( .A(n10029), .ZN(n10031) );
  AND2_X1 U5851 ( .A1(n8757), .A2(n8756), .ZN(n8758) );
  AOI21_X1 U5852 ( .B1(n8532), .B2(n10074), .A(n4397), .ZN(n4988) );
  INV_X1 U5853 ( .A(n5609), .ZN(n4397) );
  INV_X1 U5854 ( .A(n8766), .ZN(n8775) );
  AOI21_X1 U5855 ( .B1(n8773), .B2(n10074), .A(n8772), .ZN(n8774) );
  NAND2_X1 U5856 ( .A1(n8771), .A2(n8770), .ZN(n8772) );
  AND2_X1 U5857 ( .A1(n5846), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10050) );
  OAI211_X1 U5858 ( .C1(n6546), .C2(n6545), .A(n6544), .B(n6543), .ZN(n8256)
         );
  OR2_X1 U5859 ( .A1(n6542), .A2(n6537), .ZN(n6544) );
  INV_X1 U5860 ( .A(n4885), .ZN(n4883) );
  INV_X1 U5861 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7887) );
  XNOR2_X1 U5862 ( .A(n5629), .B(n5628), .ZN(n7889) );
  NAND2_X1 U5863 ( .A1(n5627), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5629) );
  INV_X1 U5864 ( .A(n6754), .ZN(n7839) );
  INV_X1 U5865 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7835) );
  INV_X1 U5866 ( .A(n5605), .ZN(n7833) );
  INV_X1 U5867 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U5868 ( .A1(n5554), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5556) );
  INV_X1 U5869 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7663) );
  INV_X1 U5870 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7559) );
  INV_X1 U5871 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7086) );
  INV_X1 U5872 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6879) );
  INV_X1 U5873 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10220) );
  INV_X1 U5874 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6852) );
  AND2_X1 U5875 ( .A1(n5167), .A2(n5203), .ZN(n7201) );
  XNOR2_X1 U5876 ( .A(n5110), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7336) );
  CLKBUF_X1 U5877 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n4407) );
  NAND2_X1 U5878 ( .A1(n8050), .A2(n8049), .ZN(n9625) );
  NOR2_X1 U5879 ( .A1(n8960), .A2(n8959), .ZN(n8988) );
  OAI22_X1 U5880 ( .A1(n4446), .A2(n8969), .B1(n7454), .B2(n4457), .ZN(n5993)
         );
  NAND2_X1 U5881 ( .A1(n4727), .A2(n4734), .ZN(n8993) );
  OR2_X1 U5882 ( .A1(n8943), .A2(n4737), .ZN(n4727) );
  NAND2_X1 U5883 ( .A1(n9080), .A2(n6212), .ZN(n9001) );
  INV_X1 U5884 ( .A(n8907), .ZN(n4445) );
  AOI21_X1 U5885 ( .B1(n6457), .B2(n6456), .A(n4766), .ZN(n8907) );
  NAND2_X1 U5886 ( .A1(n4740), .A2(n7650), .ZN(n7717) );
  NAND2_X1 U5887 ( .A1(n7649), .A2(n7652), .ZN(n4740) );
  NAND2_X1 U5888 ( .A1(n4739), .A2(n6363), .ZN(n9047) );
  NAND2_X1 U5889 ( .A1(n8943), .A2(n6355), .ZN(n4739) );
  NAND2_X1 U5890 ( .A1(n8999), .A2(n6231), .ZN(n9055) );
  NAND2_X1 U5891 ( .A1(n6235), .A2(n6234), .ZN(n9712) );
  INV_X1 U5892 ( .A(n9106), .ZN(n9832) );
  NAND2_X1 U5893 ( .A1(n4726), .A2(n6193), .ZN(n9082) );
  INV_X1 U5894 ( .A(n9510), .ZN(n9685) );
  INV_X1 U5895 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9094) );
  INV_X1 U5896 ( .A(n9110), .ZN(n9838) );
  INV_X1 U5897 ( .A(n9842), .ZN(n9104) );
  NAND2_X1 U5898 ( .A1(n4764), .A2(n4765), .ZN(n9101) );
  NAND2_X1 U5899 ( .A1(n7949), .A2(n7948), .ZN(n9636) );
  AND2_X1 U5900 ( .A1(n9837), .A2(n9726), .ZN(n9121) );
  AND2_X1 U5901 ( .A1(n8099), .A2(n8100), .ZN(n8234) );
  INV_X1 U5902 ( .A(n9302), .ZN(n9303) );
  INV_X1 U5903 ( .A(n9298), .ZN(n9300) );
  INV_X1 U5904 ( .A(n7791), .ZN(n9130) );
  INV_X1 U5905 ( .A(n7744), .ZN(n9131) );
  CLKBUF_X1 U5906 ( .A(n6778), .Z(n9139) );
  OR2_X1 U5907 ( .A1(n6966), .A2(n6968), .ZN(n4669) );
  NAND2_X1 U5908 ( .A1(n4668), .A2(n4670), .ZN(n6909) );
  AOI21_X1 U5909 ( .B1(n7032), .B2(n9160), .A(n9157), .ZN(n9172) );
  OR2_X1 U5910 ( .A1(n6914), .A2(n6896), .ZN(n9249) );
  AND2_X1 U5911 ( .A1(n7108), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4659) );
  AND2_X1 U5912 ( .A1(n7110), .A2(n7109), .ZN(n7124) );
  NOR2_X1 U5913 ( .A1(n7124), .A2(n4658), .ZN(n9186) );
  NOR2_X1 U5914 ( .A1(n7132), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4658) );
  NAND2_X1 U5915 ( .A1(n9186), .A2(n9185), .ZN(n9184) );
  AOI21_X1 U5916 ( .B1(n9184), .B2(n7126), .A(n7127), .ZN(n7513) );
  INV_X1 U5917 ( .A(n4662), .ZN(n9211) );
  OAI21_X1 U5918 ( .B1(n9266), .B2(n9265), .A(n4305), .ZN(n9613) );
  NAND2_X1 U5919 ( .A1(n4927), .A2(n4926), .ZN(n4925) );
  INV_X1 U5920 ( .A(n4922), .ZN(n4921) );
  AND2_X1 U5921 ( .A1(n9383), .A2(n9382), .ZN(n9634) );
  INV_X1 U5922 ( .A(n4485), .ZN(n9394) );
  INV_X1 U5923 ( .A(n9636), .ZN(n7952) );
  INV_X1 U5924 ( .A(n9407), .ZN(n9402) );
  NAND2_X1 U5925 ( .A1(n4906), .A2(n4905), .ZN(n9456) );
  AOI21_X1 U5926 ( .B1(n4908), .B2(n9327), .A(n4907), .ZN(n4905) );
  AND2_X1 U5927 ( .A1(n4962), .A2(n4307), .ZN(n9449) );
  NAND2_X1 U5928 ( .A1(n4910), .A2(n4908), .ZN(n9465) );
  INV_X1 U5929 ( .A(n4962), .ZN(n9462) );
  CLKBUF_X1 U5930 ( .A(n9477), .Z(n9478) );
  NAND2_X1 U5931 ( .A1(n4939), .A2(n4943), .ZN(n9514) );
  NAND2_X1 U5932 ( .A1(n9533), .A2(n4944), .ZN(n4939) );
  OAI21_X1 U5933 ( .B1(n9533), .B2(n4942), .A(n4940), .ZN(n9515) );
  NAND2_X1 U5934 ( .A1(n4492), .A2(n4334), .ZN(n9504) );
  NAND2_X1 U5935 ( .A1(n6297), .A2(n6296), .ZN(n9530) );
  INV_X1 U5936 ( .A(n9283), .ZN(n4945) );
  NAND2_X1 U5937 ( .A1(n9533), .A2(n9544), .ZN(n4946) );
  NAND2_X1 U5938 ( .A1(n4895), .A2(n4898), .ZN(n9520) );
  NAND2_X1 U5939 ( .A1(n9590), .A2(n4899), .ZN(n4895) );
  NOR2_X1 U5940 ( .A1(n4901), .A2(n8011), .ZN(n9573) );
  INV_X1 U5941 ( .A(n9590), .ZN(n4901) );
  NAND2_X1 U5942 ( .A1(n4894), .A2(n8006), .ZN(n7793) );
  CLKBUF_X1 U5943 ( .A(n7748), .Z(n7593) );
  OR2_X1 U5944 ( .A1(n9603), .A2(n6800), .ZN(n9899) );
  OR2_X1 U5945 ( .A1(n9603), .A2(n6801), .ZN(n9527) );
  INV_X1 U5946 ( .A(n9527), .ZN(n9919) );
  AND2_X2 U5947 ( .A1(n7147), .A2(n7146), .ZN(n10006) );
  OR2_X1 U5948 ( .A1(n4495), .A2(n4432), .ZN(n9737) );
  INV_X1 U5949 ( .A(n9932), .ZN(n9933) );
  OR2_X1 U5950 ( .A1(n6868), .A2(n8225), .ZN(n9934) );
  AND2_X1 U5951 ( .A1(n5969), .A2(n6465), .ZN(n9935) );
  AND2_X1 U5952 ( .A1(n4965), .A2(n5957), .ZN(n4579) );
  NAND2_X1 U5953 ( .A1(n5946), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U5954 ( .A1(n4473), .A2(n4472), .ZN(n5946) );
  AOI21_X1 U5955 ( .B1(n4283), .B2(n4474), .A(P1_IR_REG_25__SCAN_IN), .ZN(
        n4472) );
  XNOR2_X1 U5956 ( .A(n5948), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9772) );
  INV_X1 U5957 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7885) );
  INV_X1 U5958 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U5959 ( .A1(n5972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5974) );
  INV_X1 U5960 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7682) );
  INV_X1 U5961 ( .A(n6480), .ZN(n7681) );
  INV_X1 U5962 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7648) );
  XNOR2_X1 U5963 ( .A(n5942), .B(n5940), .ZN(n8101) );
  INV_X1 U5964 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7561) );
  INV_X1 U5965 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7084) );
  INV_X1 U5966 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6880) );
  INV_X1 U5967 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6866) );
  INV_X1 U5968 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6850) );
  INV_X1 U5969 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6848) );
  INV_X1 U5970 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6845) );
  XNOR2_X1 U5971 ( .A(n6102), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6931) );
  XNOR2_X1 U5972 ( .A(n5043), .B(n5042), .ZN(n6811) );
  INV_X2 U5973 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10185) );
  NOR2_X1 U5974 ( .A1(n10129), .A2(n4351), .ZN(n10133) );
  NOR2_X1 U5975 ( .A1(n10113), .A2(n10112), .ZN(n10111) );
  NOR2_X1 U5976 ( .A1(n10122), .A2(n9797), .ZN(n10110) );
  NOR2_X1 U5977 ( .A1(n10105), .A2(n4396), .ZN(n10104) );
  NAND2_X1 U5978 ( .A1(n10104), .A2(n10103), .ZN(n10102) );
  NAND2_X1 U5979 ( .A1(n7878), .A2(n4453), .ZN(n4452) );
  INV_X1 U5980 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n4453) );
  NAND2_X1 U5981 ( .A1(n8454), .A2(n4455), .ZN(n4454) );
  AND2_X1 U5982 ( .A1(n8253), .A2(n4388), .ZN(n4414) );
  NAND2_X1 U5983 ( .A1(n8248), .A2(n7842), .ZN(n4415) );
  NAND2_X1 U5984 ( .A1(n7581), .A2(n5697), .ZN(n7688) );
  AOI21_X1 U5985 ( .B1(n4451), .B2(n4450), .A(n4448), .ZN(n8398) );
  OR2_X1 U5986 ( .A1(n8397), .A2(n4449), .ZN(n4448) );
  AOI21_X1 U5987 ( .B1(n8395), .B2(n8396), .A(n8413), .ZN(n4450) );
  AOI21_X1 U5988 ( .B1(n6758), .B2(n4395), .A(n4769), .ZN(n4768) );
  NAND2_X1 U5989 ( .A1(n4772), .A2(n4326), .ZN(n4771) );
  NAND2_X1 U5990 ( .A1(n5923), .A2(n4817), .ZN(P2_U3264) );
  INV_X1 U5991 ( .A(n5922), .ZN(n5923) );
  NAND2_X1 U5992 ( .A1(n4818), .A2(n8646), .ZN(n4817) );
  OAI21_X1 U5993 ( .B1(n5921), .B2(n8646), .A(n5920), .ZN(n5922) );
  AND2_X1 U5994 ( .A1(n4822), .A2(n8497), .ZN(n8517) );
  AOI21_X1 U5995 ( .B1(n9874), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9254), .ZN(
        n4675) );
  NAND2_X1 U5996 ( .A1(n4677), .A2(n9471), .ZN(n4676) );
  MUX2_X1 U5997 ( .A(n9608), .B(n9732), .S(n10006), .Z(n9609) );
  MUX2_X1 U5998 ( .A(n9733), .B(n9732), .S(n9995), .Z(n9734) );
  INV_X1 U5999 ( .A(n10116), .ZN(n10115) );
  AND2_X1 U6000 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4342), .ZN(n4283) );
  AND2_X1 U6001 ( .A1(n4956), .A2(n9308), .ZN(n4284) );
  INV_X1 U6002 ( .A(n8551), .ZN(n4880) );
  AND2_X1 U6003 ( .A1(n6663), .A2(n6658), .ZN(n7669) );
  INV_X1 U6004 ( .A(n4798), .ZN(n4529) );
  NAND2_X1 U6005 ( .A1(n4312), .A2(n4889), .ZN(n6872) );
  INV_X1 U6006 ( .A(n9836), .ZN(n7612) );
  AND2_X1 U6007 ( .A1(n7336), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4285) );
  INV_X1 U6008 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5934) );
  INV_X1 U6009 ( .A(n5770), .ZN(n4723) );
  INV_X1 U6010 ( .A(n8627), .ZN(n4857) );
  AND2_X1 U6011 ( .A1(n9341), .A2(n9553), .ZN(n4286) );
  OR2_X1 U6012 ( .A1(n9530), .A2(n9284), .ZN(n4287) );
  AND2_X1 U6013 ( .A1(n9836), .A2(n7405), .ZN(n4288) );
  OR2_X1 U6014 ( .A1(n8776), .A2(n5602), .ZN(n4289) );
  AND2_X1 U6015 ( .A1(n9320), .A2(n9319), .ZN(n4290) );
  AND2_X1 U6016 ( .A1(n4919), .A2(n9333), .ZN(n4291) );
  AND2_X1 U6017 ( .A1(n9323), .A2(n9321), .ZN(n4292) );
  NAND2_X1 U6018 ( .A1(n8908), .A2(n8909), .ZN(n4293) );
  OR2_X1 U6019 ( .A1(n8208), .A2(n8097), .ZN(n4294) );
  OR2_X1 U6020 ( .A1(n8579), .A2(n8598), .ZN(n4295) );
  OR2_X1 U6021 ( .A1(n9631), .A2(n9310), .ZN(n4296) );
  AND2_X1 U6022 ( .A1(n8796), .A2(n8419), .ZN(n5599) );
  OR2_X1 U6023 ( .A1(n4983), .A2(n4686), .ZN(n4297) );
  AND2_X1 U6024 ( .A1(n4476), .A2(n4366), .ZN(n4298) );
  AND2_X1 U6025 ( .A1(n6616), .A2(n6614), .ZN(n8686) );
  INV_X1 U6026 ( .A(n8433), .ZN(n4634) );
  AND3_X1 U6027 ( .A1(n5100), .A2(n5098), .A3(n5099), .ZN(n4299) );
  AND2_X1 U6028 ( .A1(n4653), .A2(n4652), .ZN(n4300) );
  AND2_X1 U6029 ( .A1(n9628), .A2(n4361), .ZN(n4301) );
  AND2_X1 U6030 ( .A1(n5698), .A2(n5697), .ZN(n4302) );
  AND2_X1 U6031 ( .A1(n4883), .A2(n5003), .ZN(n4303) );
  AND2_X1 U6032 ( .A1(n4531), .A2(n5487), .ZN(n4530) );
  AND2_X1 U6033 ( .A1(n4546), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n4304) );
  INV_X1 U6034 ( .A(n9850), .ZN(n9879) );
  OR3_X1 U6035 ( .A1(n9389), .A2(n4654), .A3(n4655), .ZN(n4305) );
  NAND2_X1 U6037 ( .A1(n7562), .A2(n7505), .ZN(n7996) );
  AND3_X1 U6038 ( .A1(n5057), .A2(n5056), .A3(n5055), .ZN(n4306) );
  NAND2_X1 U6039 ( .A1(n9669), .A2(n9294), .ZN(n4307) );
  XNOR2_X1 U6040 ( .A(n6733), .B(n8501), .ZN(n8499) );
  INV_X1 U6041 ( .A(n8499), .ZN(n4867) );
  OR2_X1 U6042 ( .A1(n8437), .A2(n10052), .ZN(n6589) );
  NAND2_X1 U6043 ( .A1(n6376), .A2(n6377), .ZN(n4308) );
  NOR3_X1 U6044 ( .A1(n9620), .A2(n9991), .A3(n9619), .ZN(n4309) );
  AOI21_X1 U6045 ( .B1(n4800), .B2(n4802), .A(n4799), .ZN(n4798) );
  OR2_X1 U6046 ( .A1(n5323), .A2(n4519), .ZN(n4310) );
  XNOR2_X1 U6047 ( .A(n8906), .B(n8908), .ZN(n4311) );
  INV_X1 U6048 ( .A(n7792), .ZN(n8181) );
  INV_X1 U6049 ( .A(n4494), .ZN(n4911) );
  NAND2_X1 U6050 ( .A1(n9325), .A2(n9324), .ZN(n4494) );
  AND2_X1 U6051 ( .A1(n4891), .A2(n7541), .ZN(n4312) );
  INV_X1 U6052 ( .A(n9364), .ZN(n4496) );
  AND2_X1 U6053 ( .A1(n6456), .A2(n4293), .ZN(n4313) );
  AND2_X1 U6054 ( .A1(n6073), .A2(n6072), .ZN(n4314) );
  INV_X1 U6055 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4746) );
  AND2_X1 U6056 ( .A1(n9636), .A2(n9307), .ZN(n9339) );
  NAND2_X1 U6057 ( .A1(n4823), .A2(n4824), .ZN(n8695) );
  NAND2_X1 U6058 ( .A1(n8684), .A2(n5594), .ZN(n8653) );
  NAND2_X1 U6059 ( .A1(n4826), .A2(n6685), .ZN(n8715) );
  INV_X1 U6060 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U6061 ( .A1(n8151), .A2(n9341), .ZN(n9362) );
  AND3_X1 U6062 ( .A1(n6716), .A2(n6727), .A3(n6714), .ZN(n4315) );
  AND2_X1 U6063 ( .A1(n4877), .A2(n4289), .ZN(n4316) );
  OR2_X1 U6064 ( .A1(n9210), .A2(n9209), .ZN(n4317) );
  INV_X1 U6065 ( .A(n9329), .ZN(n4907) );
  INV_X1 U6066 ( .A(n9438), .ZN(n4917) );
  INV_X1 U6067 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6068 ( .A1(n8158), .A2(n8209), .ZN(n9620) );
  INV_X1 U6069 ( .A(n9620), .ZN(n4927) );
  NAND2_X1 U6070 ( .A1(n4403), .A2(n5592), .ZN(n8683) );
  OR2_X1 U6071 ( .A1(n9341), .A2(n9908), .ZN(n4318) );
  XNOR2_X1 U6072 ( .A(n8781), .B(n8564), .ZN(n8581) );
  AND2_X1 U6073 ( .A1(n7282), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4319) );
  AND2_X1 U6074 ( .A1(n8346), .A2(n8347), .ZN(n4320) );
  NAND2_X1 U6075 ( .A1(n5343), .A2(n6695), .ZN(n8672) );
  OR2_X1 U6076 ( .A1(n6716), .A2(n6727), .ZN(n4321) );
  OR2_X1 U6077 ( .A1(n6549), .A2(n6814), .ZN(n4322) );
  AND2_X1 U6078 ( .A1(n7201), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4323) );
  NAND2_X1 U6079 ( .A1(n8607), .A2(n4603), .ZN(n8595) );
  OR2_X1 U6080 ( .A1(n9486), .A2(n9290), .ZN(n4324) );
  NOR2_X2 U6081 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5347) );
  OR2_X1 U6082 ( .A1(n4811), .A2(n8499), .ZN(n4325) );
  AND2_X1 U6083 ( .A1(n6750), .A2(n7839), .ZN(n4326) );
  NAND2_X1 U6084 ( .A1(n5542), .A2(n5541), .ZN(n6733) );
  NAND2_X1 U6085 ( .A1(n5480), .A2(n5479), .ZN(n8776) );
  OR2_X1 U6086 ( .A1(n8023), .A2(n9317), .ZN(n9551) );
  INV_X1 U6087 ( .A(n9551), .ZN(n4419) );
  NAND2_X1 U6088 ( .A1(n5497), .A2(n5496), .ZN(n8769) );
  NOR2_X1 U6089 ( .A1(n9701), .A2(n9279), .ZN(n4327) );
  AND2_X1 U6090 ( .A1(n4910), .A2(n9326), .ZN(n4328) );
  AND2_X1 U6091 ( .A1(n5019), .A2(n4407), .ZN(n4329) );
  AND3_X1 U6092 ( .A1(n4526), .A2(n4524), .A3(n4523), .ZN(n4330) );
  AND2_X1 U6093 ( .A1(n9530), .A2(n9284), .ZN(n4331) );
  AND2_X1 U6094 ( .A1(n6697), .A2(n8686), .ZN(n4332) );
  NOR2_X1 U6095 ( .A1(n8617), .A2(n8371), .ZN(n4333) );
  INV_X1 U6096 ( .A(n8786), .ZN(n8594) );
  AND2_X1 U6097 ( .A1(n4896), .A2(n9321), .ZN(n4334) );
  INV_X1 U6098 ( .A(n4859), .ZN(n4858) );
  NOR2_X1 U6099 ( .A1(n5599), .A2(n4333), .ZN(n4859) );
  NAND2_X1 U6100 ( .A1(n8541), .A2(n4683), .ZN(n4684) );
  NAND3_X1 U6101 ( .A1(n9318), .A2(n9541), .A3(n9543), .ZN(n4335) );
  INV_X1 U6102 ( .A(n4801), .ZN(n4800) );
  OAI21_X1 U6103 ( .B1(n5437), .B2(n4802), .A(n5458), .ZN(n4801) );
  INV_X1 U6104 ( .A(n5594), .ZN(n4507) );
  INV_X1 U6105 ( .A(n7405), .ZN(n9920) );
  AND2_X1 U6106 ( .A1(n8617), .A2(n8371), .ZN(n4336) );
  AND2_X1 U6107 ( .A1(n6685), .A2(n6686), .ZN(n7892) );
  AND2_X1 U6108 ( .A1(n4862), .A2(n8521), .ZN(n4337) );
  AND2_X1 U6109 ( .A1(n8048), .A2(n8047), .ZN(n4338) );
  INV_X1 U6110 ( .A(n5595), .ZN(n4508) );
  AND2_X1 U6111 ( .A1(n4824), .A2(n6696), .ZN(n4339) );
  OR2_X1 U6112 ( .A1(n8581), .A2(n4835), .ZN(n4340) );
  AND2_X1 U6113 ( .A1(n9340), .A2(n8103), .ZN(n9380) );
  NAND2_X1 U6114 ( .A1(n4291), .A2(n9337), .ZN(n4341) );
  INV_X1 U6115 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U6116 ( .A1(n5944), .A2(n4748), .ZN(n4342) );
  AND2_X1 U6117 ( .A1(n6682), .A2(n7890), .ZN(n7854) );
  INV_X1 U6118 ( .A(n9127), .ZN(n9306) );
  NAND2_X1 U6119 ( .A1(n6445), .A2(n6444), .ZN(n9127) );
  AND2_X1 U6120 ( .A1(n8850), .A2(n8427), .ZN(n4343) );
  NOR2_X1 U6121 ( .A1(n5746), .A2(n8378), .ZN(n4344) );
  NOR2_X1 U6122 ( .A1(n5738), .A2(n8331), .ZN(n4345) );
  NOR2_X1 U6123 ( .A1(n9685), .A2(n9285), .ZN(n4346) );
  INV_X1 U6124 ( .A(n4685), .ZN(n8590) );
  NOR2_X1 U6125 ( .A1(n4983), .A2(n4687), .ZN(n4685) );
  INV_X1 U6126 ( .A(n4610), .ZN(n4609) );
  NOR2_X1 U6127 ( .A1(n4612), .A2(n4815), .ZN(n4610) );
  AND3_X1 U6128 ( .A1(n5077), .A2(n5076), .A3(n5079), .ZN(n4347) );
  NOR2_X1 U6129 ( .A1(n7962), .A2(n7961), .ZN(n4538) );
  NOR2_X1 U6130 ( .A1(n8769), .A2(n8571), .ZN(n4348) );
  NOR2_X1 U6131 ( .A1(n4952), .A2(n9362), .ZN(n4349) );
  AND2_X1 U6132 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n4350) );
  AND2_X1 U6133 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n4351) );
  NOR2_X1 U6134 ( .A1(n4907), .A2(n9327), .ZN(n4352) );
  AND2_X1 U6135 ( .A1(n4896), .A2(n4292), .ZN(n4353) );
  AND2_X1 U6136 ( .A1(n4672), .A2(n6095), .ZN(n4354) );
  AND2_X1 U6137 ( .A1(n5426), .A2(n5425), .ZN(n8617) );
  INV_X1 U6138 ( .A(n8617), .ZN(n8793) );
  NOR2_X1 U6139 ( .A1(n9454), .A2(n9296), .ZN(n4355) );
  XNOR2_X1 U6140 ( .A(n8769), .B(n8571), .ZN(n8551) );
  OR2_X1 U6141 ( .A1(n4801), .A2(n4533), .ZN(n4356) );
  OR2_X1 U6142 ( .A1(n9283), .A2(n4331), .ZN(n4357) );
  OR2_X1 U6143 ( .A1(n9402), .A2(n9127), .ZN(n4358) );
  INV_X1 U6144 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5945) );
  INV_X1 U6145 ( .A(n4620), .ZN(n4619) );
  OR2_X1 U6146 ( .A1(n8455), .A2(n5907), .ZN(n4622) );
  INV_X1 U6147 ( .A(n4900), .ZN(n4899) );
  NAND2_X1 U6148 ( .A1(n4290), .A2(n4902), .ZN(n4900) );
  AND2_X1 U6149 ( .A1(n6728), .A2(n6727), .ZN(n4359) );
  AND2_X1 U6150 ( .A1(n6932), .A2(n4671), .ZN(n4360) );
  OR2_X1 U6151 ( .A1(n9629), .A2(n9617), .ZN(n4361) );
  AND2_X1 U6152 ( .A1(n4824), .A2(n4596), .ZN(n4362) );
  AND2_X1 U6153 ( .A1(n4710), .A2(n8297), .ZN(n4363) );
  AND3_X1 U6154 ( .A1(n6712), .A2(n6704), .A3(n4633), .ZN(n4364) );
  AND2_X1 U6155 ( .A1(n4946), .A2(n4945), .ZN(n4365) );
  NAND2_X1 U6156 ( .A1(n8924), .A2(n6291), .ZN(n4366) );
  AND2_X1 U6157 ( .A1(n8247), .A2(n8246), .ZN(n4367) );
  AND2_X1 U6158 ( .A1(n4352), .A2(n9324), .ZN(n4368) );
  AND2_X1 U6159 ( .A1(n5364), .A2(n5345), .ZN(n4369) );
  AND2_X1 U6160 ( .A1(n4540), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n4370) );
  AND2_X1 U6161 ( .A1(n9407), .A2(n9127), .ZN(n9336) );
  INV_X1 U6162 ( .A(n9336), .ZN(n8202) );
  NOR2_X1 U6163 ( .A1(n4470), .A2(n4468), .ZN(n4371) );
  NOR2_X1 U6164 ( .A1(n9278), .A2(n4934), .ZN(n4372) );
  AND2_X1 U6165 ( .A1(n8063), .A2(n4561), .ZN(n4373) );
  INV_X1 U6166 ( .A(n9540), .ZN(n9697) );
  AND2_X1 U6167 ( .A1(n6270), .A2(n6269), .ZN(n9540) );
  AND2_X1 U6168 ( .A1(n9419), .A2(n9303), .ZN(n9335) );
  INV_X1 U6169 ( .A(n9335), .ZN(n4918) );
  AND2_X1 U6170 ( .A1(n4615), .A2(n4614), .ZN(n4374) );
  AND2_X1 U6171 ( .A1(n4970), .A2(n5555), .ZN(n4375) );
  INV_X1 U6172 ( .A(n8559), .ZN(n8568) );
  AND2_X1 U6173 ( .A1(n6612), .A2(n6613), .ZN(n8559) );
  AND2_X1 U6174 ( .A1(n7792), .A2(n7785), .ZN(n4376) );
  AND2_X1 U6175 ( .A1(n5957), .A2(n5959), .ZN(n4377) );
  INV_X1 U6176 ( .A(n4953), .ZN(n4952) );
  OAI21_X1 U6177 ( .B1(n4284), .B2(n9380), .A(n4296), .ZN(n4953) );
  AND2_X1 U6178 ( .A1(n8026), .A2(n8025), .ZN(n4378) );
  AND2_X1 U6179 ( .A1(n6694), .A2(n6692), .ZN(n4379) );
  AND2_X1 U6180 ( .A1(n6171), .A2(n4469), .ZN(n4380) );
  INV_X1 U6181 ( .A(n4756), .ZN(n4479) );
  OR2_X1 U6182 ( .A1(n6247), .A2(n4757), .ZN(n4756) );
  AND2_X1 U6183 ( .A1(n4300), .A2(n7777), .ZN(n4381) );
  INV_X1 U6184 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4748) );
  INV_X1 U6185 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4886) );
  OR2_X1 U6186 ( .A1(n4311), .A2(n6454), .ZN(n4382) );
  INV_X1 U6187 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4752) );
  INV_X1 U6188 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4753) );
  NAND2_X1 U6189 ( .A1(n5789), .A2(n5788), .ZN(n8755) );
  INV_X1 U6190 ( .A(n8755), .ZN(n4680) );
  NAND2_X1 U6191 ( .A1(n9814), .A2(n7416), .ZN(n9583) );
  NAND2_X1 U6192 ( .A1(n5812), .A2(n5799), .ZN(n8413) );
  INV_X1 U6193 ( .A(n8413), .ZN(n7842) );
  NOR2_X1 U6194 ( .A1(n7730), .A2(n4698), .ZN(n7862) );
  NAND2_X1 U6195 ( .A1(n7857), .A2(n5586), .ZN(n7900) );
  NAND2_X1 U6196 ( .A1(n9276), .A2(n9275), .ZN(n9570) );
  XNOR2_X1 U6197 ( .A(n5947), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U6198 ( .A1(n4429), .A2(n7346), .ZN(n7345) );
  AND2_X1 U6199 ( .A1(n8915), .A2(n8914), .ZN(n4383) );
  NAND2_X1 U6200 ( .A1(n7345), .A2(n4716), .ZN(n7459) );
  INV_X1 U6201 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n4541) );
  INV_X1 U6202 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n4542) );
  OR2_X1 U6203 ( .A1(n7514), .A2(n7515), .ZN(n4384) );
  AND2_X1 U6204 ( .A1(n4930), .A2(n7750), .ZN(n4385) );
  INV_X1 U6205 ( .A(n4803), .ZN(n4802) );
  NOR2_X1 U6206 ( .A1(n5459), .A2(n4804), .ZN(n4803) );
  AND3_X1 U6207 ( .A1(n9594), .A2(n4656), .A3(n9690), .ZN(n9508) );
  NOR2_X1 U6208 ( .A1(n6513), .A2(n6512), .ZN(n4386) );
  NOR2_X1 U6209 ( .A1(n7730), .A2(n8844), .ZN(n4700) );
  AND2_X1 U6210 ( .A1(n5489), .A2(SI_24_), .ZN(n4387) );
  OR2_X1 U6211 ( .A1(n8535), .A2(n8300), .ZN(n4388) );
  AND2_X1 U6212 ( .A1(n4543), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n4389) );
  INV_X1 U6213 ( .A(n5599), .ZN(n4861) );
  INV_X1 U6214 ( .A(n8432), .ZN(n4636) );
  AND2_X1 U6215 ( .A1(n7414), .A2(n7413), .ZN(n4390) );
  INV_X1 U6216 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n4547) );
  NAND2_X1 U6217 ( .A1(n6054), .A2(n6053), .ZN(n7165) );
  NAND2_X1 U6218 ( .A1(n6479), .A2(n9444), .ZN(n8066) );
  INV_X1 U6219 ( .A(n7749), .ZN(n4652) );
  AND2_X1 U6220 ( .A1(n4669), .A2(n6932), .ZN(n4391) );
  AND2_X1 U6221 ( .A1(n10034), .A2(n10035), .ZN(n4392) );
  INV_X1 U6222 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n4544) );
  INV_X1 U6223 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n4545) );
  AND2_X1 U6224 ( .A1(n6279), .A2(n6278), .ZN(n9860) );
  AND2_X1 U6225 ( .A1(n4668), .A2(n4666), .ZN(n4393) );
  OR2_X1 U6226 ( .A1(n7333), .A2(n7332), .ZN(n4816) );
  INV_X1 U6227 ( .A(n4816), .ZN(n4618) );
  INV_X1 U6228 ( .A(n5991), .ZN(n9471) );
  XOR2_X1 U6229 ( .A(n5908), .B(P2_REG2_REG_17__SCAN_IN), .Z(n4394) );
  AND2_X1 U6230 ( .A1(n7839), .A2(n4770), .ZN(n4395) );
  AND2_X1 U6231 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4396) );
  INV_X1 U6232 ( .A(n4407), .ZN(n4692) );
  INV_X1 U6233 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n4455) );
  INV_X1 U6234 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4558) );
  INV_X1 U6235 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n4559) );
  NAND2_X1 U6236 ( .A1(n8633), .A2(n5597), .ZN(n5598) );
  INV_X1 U6237 ( .A(n7009), .ZN(n7005) );
  NAND3_X1 U6238 ( .A1(n4400), .A2(n4693), .A3(n4398), .ZN(n8869) );
  AOI21_X2 U6239 ( .B1(n8377), .B2(n5747), .A(n4344), .ZN(n8290) );
  NAND2_X1 U6240 ( .A1(n7245), .A2(n5675), .ZN(n7396) );
  NOR2_X1 U6241 ( .A1(n4702), .A2(n5781), .ZN(n5806) );
  NAND3_X1 U6242 ( .A1(n6756), .A2(n6757), .A3(n7684), .ZN(n5647) );
  NAND2_X1 U6243 ( .A1(n4881), .A2(n4882), .ZN(n7725) );
  NAND2_X1 U6244 ( .A1(n5578), .A2(n5577), .ZN(n7361) );
  NAND2_X1 U6245 ( .A1(n4425), .A2(n5591), .ZN(n8691) );
  NAND2_X1 U6246 ( .A1(n7617), .A2(n5581), .ZN(n7668) );
  NAND2_X1 U6247 ( .A1(n6777), .A2(n4428), .ZN(n7402) );
  OAI21_X1 U6248 ( .B1(n5181), .B2(n4503), .A(n5194), .ZN(n4502) );
  NAND2_X1 U6249 ( .A1(n9360), .A2(n9362), .ZN(n9622) );
  NAND2_X1 U6250 ( .A1(n9586), .A2(n9273), .ZN(n9276) );
  NAND2_X1 U6251 ( .A1(n4579), .A2(n5926), .ZN(n4413) );
  AND2_X2 U6252 ( .A1(n4887), .A2(n6139), .ZN(n5926) );
  NAND2_X1 U6253 ( .A1(n9804), .A2(n7752), .ZN(n7784) );
  NAND3_X2 U6254 ( .A1(n5984), .A2(n5989), .A3(n5983), .ZN(n7158) );
  NAND2_X1 U6255 ( .A1(n10099), .A2(n4452), .ZN(n10097) );
  NAND2_X1 U6256 ( .A1(n10090), .A2(n4454), .ZN(n10088) );
  OAI21_X1 U6257 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9801), .A(n10118), .ZN(
        n9803) );
  OAI21_X1 U6258 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10093), .ZN(n10091) );
  NAND2_X1 U6259 ( .A1(n6994), .A2(n5652), .ZN(n7103) );
  NAND2_X1 U6260 ( .A1(n5771), .A2(n4720), .ZN(n4719) );
  NAND2_X1 U6261 ( .A1(n7247), .A2(n7246), .ZN(n7245) );
  NAND4_X1 U6262 ( .A1(n5013), .A2(n5012), .A3(n5011), .A4(n5010), .ZN(n6590)
         );
  NAND2_X1 U6263 ( .A1(n7426), .A2(n7425), .ZN(n7436) );
  NAND2_X1 U6264 ( .A1(n7618), .A2(n5580), .ZN(n7617) );
  INV_X1 U6265 ( .A(n8767), .ZN(n8773) );
  NAND2_X1 U6266 ( .A1(n8775), .A2(n8774), .ZN(n8872) );
  OAI22_X2 U6267 ( .A1(n5772), .A2(n8306), .B1(n8305), .B2(n8308), .ZN(n8395)
         );
  NAND2_X1 U6268 ( .A1(n5768), .A2(n5767), .ZN(n5771) );
  NAND2_X1 U6269 ( .A1(n6766), .A2(n6768), .ZN(n6767) );
  NAND2_X1 U6270 ( .A1(n5680), .A2(n5679), .ZN(n7394) );
  NAND2_X1 U6271 ( .A1(n4405), .A2(n7091), .ZN(n6766) );
  NAND3_X1 U6272 ( .A1(n4406), .A2(n5658), .A3(n7090), .ZN(n4405) );
  NAND2_X1 U6273 ( .A1(n5653), .A2(n7103), .ZN(n6982) );
  NAND2_X1 U6274 ( .A1(n5655), .A2(n7089), .ZN(n4406) );
  NAND2_X1 U6275 ( .A1(n4392), .A2(n10063), .ZN(n7238) );
  AOI21_X2 U6276 ( .B1(n8330), .B2(n5727), .A(n4345), .ZN(n8377) );
  INV_X2 U6277 ( .A(n5851), .ZN(n5393) );
  NAND2_X1 U6278 ( .A1(n4409), .A2(n4408), .ZN(n8032) );
  NAND2_X1 U6279 ( .A1(n8034), .A2(n8031), .ZN(n4409) );
  OR3_X2 U6280 ( .A1(n8234), .A2(n8235), .A3(n8233), .ZN(n8236) );
  NAND2_X1 U6281 ( .A1(n4575), .A2(n4571), .ZN(n8019) );
  NAND2_X1 U6282 ( .A1(n4557), .A2(n4918), .ZN(n4555) );
  NAND2_X1 U6283 ( .A1(n8022), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U6284 ( .A1(n4565), .A2(n4378), .ZN(n8028) );
  NAND2_X1 U6285 ( .A1(n8005), .A2(n8131), .ZN(n4577) );
  OAI21_X1 U6286 ( .B1(n8095), .B2(n4537), .A(n8215), .ZN(n8098) );
  NAND2_X1 U6287 ( .A1(n7748), .A2(n7747), .ZN(n4930) );
  INV_X1 U6288 ( .A(n8174), .ZN(n9913) );
  OAI21_X1 U6289 ( .B1(n4415), .B2(n4367), .A(n4414), .ZN(P2_U3216) );
  XNOR2_X2 U6290 ( .A(n4417), .B(n5550), .ZN(n7662) );
  NAND2_X1 U6291 ( .A1(n5218), .A2(n4418), .ZN(n5220) );
  NAND2_X1 U6292 ( .A1(n5182), .A2(n5181), .ZN(n5218) );
  NAND3_X1 U6293 ( .A1(n8181), .A2(n4422), .A3(n8180), .ZN(n4421) );
  NAND3_X1 U6294 ( .A1(n5572), .A2(n7235), .A3(n4424), .ZN(n7231) );
  NAND2_X1 U6295 ( .A1(n10019), .A2(n7229), .ZN(n4424) );
  NAND2_X1 U6296 ( .A1(n8719), .A2(n5588), .ZN(n4425) );
  INV_X1 U6297 ( .A(n8751), .ZN(n4516) );
  NAND2_X1 U6298 ( .A1(n5654), .A2(n6982), .ZN(n5655) );
  NAND2_X1 U6299 ( .A1(n5552), .A2(n4375), .ZN(n4701) );
  NOR2_X1 U6300 ( .A1(n4957), .A2(n4954), .ZN(n4949) );
  NAND4_X2 U6301 ( .A1(n6040), .A2(n6039), .A3(n6038), .A4(n6037), .ZN(n9138)
         );
  NAND2_X1 U6302 ( .A1(n6789), .A2(n7148), .ZN(n6791) );
  OR2_X1 U6303 ( .A1(n6238), .A2(n6884), .ZN(n6018) );
  NAND2_X1 U6304 ( .A1(n9276), .A2(n4372), .ZN(n4933) );
  INV_X4 U6305 ( .A(n8089), .ZN(n8078) );
  NAND2_X1 U6306 ( .A1(n7996), .A2(n7986), .ZN(n7440) );
  AOI21_X2 U6307 ( .B1(n8935), .B2(n8933), .A(n8932), .ZN(n9039) );
  OAI211_X1 U6308 ( .C1(n4466), .C2(n9030), .A(n4464), .B(n4728), .ZN(n6413)
         );
  NOR2_X1 U6309 ( .A1(n4949), .A2(n4953), .ZN(n9360) );
  NAND3_X2 U6310 ( .A1(n6027), .A2(n6025), .A3(n6026), .ZN(n4428) );
  INV_X1 U6311 ( .A(n4428), .ZN(n9938) );
  NAND2_X1 U6312 ( .A1(n5001), .A2(n5351), .ZN(n5631) );
  NAND2_X1 U6313 ( .A1(n9365), .A2(n9553), .ZN(n4497) );
  NAND2_X1 U6314 ( .A1(n4301), .A2(n9627), .ZN(n4432) );
  OAI21_X1 U6315 ( .B1(n4915), .B2(n4914), .A(n8202), .ZN(n4913) );
  NAND2_X1 U6316 ( .A1(n4341), .A2(n4912), .ZN(n4484) );
  NAND2_X1 U6317 ( .A1(n4930), .A2(n4928), .ZN(n9804) );
  NAND2_X1 U6318 ( .A1(n7420), .A2(n8169), .ZN(n7422) );
  NAND2_X1 U6319 ( .A1(n6791), .A2(n6790), .ZN(n7420) );
  AND2_X2 U6320 ( .A1(n6002), .A2(n4277), .ZN(n6021) );
  NAND2_X2 U6321 ( .A1(n6492), .A2(n9258), .ZN(n6002) );
  NAND2_X1 U6322 ( .A1(n9293), .A2(n4961), .ZN(n4960) );
  AOI21_X1 U6323 ( .B1(n9864), .B2(P1_REG2_REG_15__SCAN_IN), .A(n4660), .ZN(
        n9212) );
  NOR2_X1 U6324 ( .A1(n7107), .A2(n4659), .ZN(n7110) );
  INV_X1 U6325 ( .A(n5926), .ZN(n5943) );
  NAND2_X1 U6326 ( .A1(n5926), .A2(n4971), .ZN(n5928) );
  NAND2_X1 U6327 ( .A1(n6703), .A2(n4364), .ZN(n4642) );
  NAND2_X1 U6328 ( .A1(n4639), .A2(n4638), .ZN(n6721) );
  INV_X1 U6329 ( .A(n6758), .ZN(n4772) );
  AOI21_X1 U6330 ( .B1(n4806), .B2(n4805), .A(n4628), .ZN(n4627) );
  INV_X1 U6331 ( .A(n4629), .ZN(n6706) );
  NAND2_X1 U6332 ( .A1(n4809), .A2(n6736), .ZN(n4808) );
  NAND2_X1 U6333 ( .A1(n6693), .A2(n4379), .ZN(n4631) );
  INV_X1 U6334 ( .A(n4626), .ZN(n4625) );
  AOI21_X1 U6335 ( .B1(n6725), .B2(n6726), .A(n4359), .ZN(n4624) );
  OR2_X2 U6336 ( .A1(n6609), .A2(n6755), .ZN(n6727) );
  INV_X1 U6337 ( .A(n4438), .ZN(n7673) );
  XNOR2_X1 U6338 ( .A(n8489), .B(n7941), .ZN(n8739) );
  NOR2_X4 U6339 ( .A1(n8577), .A2(n8776), .ZN(n8541) );
  NAND2_X1 U6340 ( .A1(n4830), .A2(n4833), .ZN(n5028) );
  NOR2_X1 U6341 ( .A1(n8394), .A2(n5776), .ZN(n8247) );
  NAND2_X1 U6342 ( .A1(n4850), .A2(n5001), .ZN(n5018) );
  NOR2_X1 U6343 ( .A1(n4832), .A2(n4831), .ZN(n4830) );
  NAND2_X1 U6344 ( .A1(n5128), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5150) );
  NAND2_X1 U6345 ( .A1(n5498), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5517) );
  INV_X1 U6346 ( .A(n4586), .ZN(n4585) );
  INV_X1 U6347 ( .A(n6557), .ZN(n4587) );
  XNOR2_X2 U6348 ( .A(n5559), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U6349 ( .A1(n5158), .A2(n5157), .ZN(n5182) );
  OR3_X2 U6350 ( .A1(n8140), .A2(n8139), .A3(n8138), .ZN(n8191) );
  NAND2_X1 U6351 ( .A1(n4444), .A2(n9838), .ZN(n6505) );
  OAI21_X1 U6352 ( .B1(n9037), .B2(n4382), .A(n4445), .ZN(n4444) );
  NAND2_X1 U6353 ( .A1(n5344), .A2(n4980), .ZN(n4796) );
  NAND2_X1 U6354 ( .A1(n4674), .A2(n9444), .ZN(n4673) );
  NOR2_X1 U6355 ( .A1(n9630), .A2(n9991), .ZN(n4495) );
  AND3_X2 U6356 ( .A1(n4753), .A2(n4752), .A3(n4644), .ZN(n6023) );
  NAND2_X1 U6357 ( .A1(n4938), .A2(n4937), .ZN(n9489) );
  NAND2_X1 U6358 ( .A1(n5138), .A2(n5139), .ZN(n5142) );
  NAND2_X2 U6359 ( .A1(n6158), .A2(n6157), .ZN(n7749) );
  NOR2_X1 U6360 ( .A1(n10241), .A2(n10125), .ZN(n10124) );
  NOR2_X1 U6361 ( .A1(n10201), .A2(n10123), .ZN(n10122) );
  NOR2_X1 U6362 ( .A1(n9794), .A2(n9793), .ZN(n10273) );
  OAI22_X1 U6363 ( .A1(n7606), .A2(n8969), .B1(n7405), .B2(n4457), .ZN(n6068)
         );
  OAI22_X1 U6364 ( .A1(n6785), .A2(n8969), .B1(n9836), .B2(n4457), .ZN(n6046)
         );
  OAI22_X1 U6365 ( .A1(n7428), .A2(n8969), .B1(n7535), .B2(n4457), .ZN(n6105)
         );
  OAI22_X1 U6366 ( .A1(n9540), .A2(n4457), .B1(n8969), .B2(n9033), .ZN(n6274)
         );
  OAI21_X1 U6367 ( .B1(n9407), .B2(n4457), .A(n4456), .ZN(n6446) );
  OAI22_X1 U6368 ( .A1(n9454), .A2(n4457), .B1(n8969), .B2(n9296), .ZN(n6411)
         );
  OAI22_X1 U6369 ( .A1(n9378), .A2(n4457), .B1(n8969), .B2(n4281), .ZN(n8917)
         );
  NAND2_X1 U6370 ( .A1(n4461), .A2(n4459), .ZN(n6116) );
  NAND2_X1 U6371 ( .A1(n6054), .A2(n4462), .ZN(n4461) );
  OAI21_X1 U6372 ( .B1(n6054), .B2(n4463), .A(n4462), .ZN(n7502) );
  NAND2_X1 U6373 ( .A1(n4732), .A2(n4465), .ZN(n4464) );
  NOR2_X1 U6374 ( .A1(n6413), .A2(n6412), .ZN(n9067) );
  NAND2_X1 U6375 ( .A1(n6138), .A2(n4371), .ZN(n4467) );
  NAND2_X1 U6376 ( .A1(n4467), .A2(n4380), .ZN(n7715) );
  OAI21_X1 U6377 ( .B1(n5943), .B2(n4474), .A(n4283), .ZN(n5948) );
  NAND2_X1 U6378 ( .A1(n5943), .A2(n4283), .ZN(n4473) );
  OAI21_X1 U6379 ( .B1(n5943), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U6380 ( .A1(n4475), .A2(n4476), .ZN(n8926) );
  NAND3_X1 U6381 ( .A1(n4482), .A2(n4480), .A3(n9338), .ZN(n9381) );
  NAND2_X1 U6382 ( .A1(n4484), .A2(n4481), .ZN(n4480) );
  NAND2_X1 U6383 ( .A1(n4483), .A2(n4484), .ZN(n4482) );
  NOR2_X1 U6384 ( .A1(n9438), .A2(n9339), .ZN(n4483) );
  OAI21_X1 U6385 ( .B1(n9438), .B2(n4341), .A(n4912), .ZN(n4485) );
  NAND2_X2 U6386 ( .A1(n5220), .A2(n4488), .ZN(n5222) );
  NAND2_X1 U6387 ( .A1(n9315), .A2(n4489), .ZN(n4492) );
  NAND2_X1 U6388 ( .A1(n9325), .A2(n4368), .ZN(n4493) );
  NAND3_X1 U6389 ( .A1(n4493), .A2(n9330), .A3(n4903), .ZN(n9332) );
  XNOR2_X1 U6390 ( .A(n4911), .B(n9479), .ZN(n9481) );
  AND2_X2 U6391 ( .A1(n4497), .A2(n4496), .ZN(n9627) );
  NAND3_X1 U6392 ( .A1(n7741), .A2(n8106), .A3(n7742), .ZN(n7790) );
  NAND2_X2 U6393 ( .A1(n5833), .A2(n6587), .ZN(n5604) );
  OAI21_X1 U6394 ( .B1(n5182), .B2(n4503), .A(n4501), .ZN(n5196) );
  INV_X1 U6395 ( .A(n4502), .ZN(n4501) );
  NAND2_X1 U6396 ( .A1(n5218), .A2(n5217), .ZN(n5195) );
  NAND2_X1 U6397 ( .A1(n5585), .A2(n5584), .ZN(n7813) );
  INV_X1 U6398 ( .A(n5584), .ZN(n4514) );
  NAND2_X1 U6399 ( .A1(n5284), .A2(n5283), .ZN(n5304) );
  NAND3_X1 U6400 ( .A1(n9624), .A2(n9623), .A3(n4330), .ZN(n9736) );
  NOR2_X1 U6401 ( .A1(n9616), .A2(n9617), .ZN(n4525) );
  NAND2_X1 U6402 ( .A1(n5424), .A2(n4530), .ZN(n4527) );
  INV_X1 U6403 ( .A(n4538), .ZN(n8052) );
  NAND2_X1 U6404 ( .A1(n6159), .A2(n4370), .ZN(n6236) );
  NAND2_X1 U6405 ( .A1(n5953), .A2(n4389), .ZN(n6342) );
  NAND2_X1 U6406 ( .A1(n5954), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6382) );
  NAND4_X1 U6407 ( .A1(n4550), .A2(n4549), .A3(n4548), .A4(n6213), .ZN(n5936)
         );
  NOR2_X1 U6408 ( .A1(n5936), .A2(n4551), .ZN(n4887) );
  NAND4_X1 U6409 ( .A1(n5937), .A2(n4554), .A3(n4553), .A4(n4552), .ZN(n4551)
         );
  NAND3_X1 U6410 ( .A1(n8043), .A2(n4556), .A3(n4555), .ZN(n8044) );
  NAND3_X1 U6411 ( .A1(n8039), .A2(n9420), .A3(n4918), .ZN(n4556) );
  AOI21_X1 U6412 ( .B1(n4564), .B2(n4373), .A(n4560), .ZN(n4563) );
  NAND2_X1 U6413 ( .A1(n4563), .A2(n4294), .ZN(n8094) );
  NAND2_X1 U6414 ( .A1(n8062), .A2(n8061), .ZN(n4564) );
  NAND3_X1 U6415 ( .A1(n4568), .A2(n4419), .A3(n4566), .ZN(n4565) );
  NAND3_X1 U6416 ( .A1(n7982), .A2(n8110), .A3(n7981), .ZN(n4574) );
  NAND2_X1 U6417 ( .A1(n5926), .A2(n4578), .ZN(n8254) );
  NAND2_X1 U6418 ( .A1(n5926), .A2(n4965), .ZN(n4967) );
  NAND4_X1 U6419 ( .A1(n5550), .A2(n5622), .A3(n5625), .A4(n4580), .ZN(n4991)
         );
  INV_X2 U6420 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U6421 ( .A1(n5059), .A2(n4581), .ZN(n7234) );
  NOR2_X2 U6422 ( .A1(n8521), .A2(n4587), .ZN(n4586) );
  XNOR2_X1 U6423 ( .A(n8494), .B(n8745), .ZN(n8498) );
  NAND2_X1 U6424 ( .A1(n7698), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U6425 ( .A1(n4823), .A2(n4362), .ZN(n4597) );
  NAND2_X1 U6426 ( .A1(n4597), .A2(n4598), .ZN(n8662) );
  MUX2_X1 U6427 ( .A(n5895), .B(P2_REG2_REG_1__SCAN_IN), .S(n5894), .Z(n7256)
         );
  INV_X1 U6428 ( .A(n4613), .ZN(n7209) );
  NAND2_X1 U6429 ( .A1(n7310), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4620) );
  NOR2_X1 U6430 ( .A1(n4623), .A2(n5204), .ZN(n5044) );
  NAND2_X1 U6431 ( .A1(n4868), .A2(n4623), .ZN(n5085) );
  NOR2_X4 U6432 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4623) );
  NAND3_X1 U6433 ( .A1(n6742), .A2(n6741), .A3(n6743), .ZN(n4628) );
  NAND3_X1 U6434 ( .A1(n6625), .A2(n6617), .A3(n4633), .ZN(n4632) );
  NAND3_X1 U6435 ( .A1(n4643), .A2(n4642), .A3(n4640), .ZN(n4639) );
  INV_X2 U6436 ( .A(n7150), .ZN(n7541) );
  MUX2_X1 U6437 ( .A(n6919), .B(n9776), .S(n6002), .Z(n7150) );
  NAND3_X1 U6438 ( .A1(n7412), .A2(n4288), .A3(n4647), .ZN(n7415) );
  INV_X1 U6439 ( .A(n4648), .ZN(n9916) );
  OR2_X2 U6440 ( .A1(n9450), .A2(n4650), .ZN(n9418) );
  NAND2_X1 U6441 ( .A1(n4381), .A2(n7414), .ZN(n7755) );
  NAND2_X1 U6442 ( .A1(n6966), .A2(n4360), .ZN(n4664) );
  INV_X1 U6443 ( .A(n6931), .ZN(n4672) );
  NAND3_X1 U6444 ( .A1(n4676), .A2(n4675), .A3(n4673), .ZN(P1_U3260) );
  INV_X1 U6445 ( .A(n4684), .ZN(n5835) );
  NAND2_X2 U6446 ( .A1(n4689), .A2(n5019), .ZN(n5851) );
  OR2_X2 U6447 ( .A1(n5567), .A2(n5566), .ZN(n5854) );
  OR2_X2 U6448 ( .A1(n7730), .A2(n4695), .ZN(n8728) );
  INV_X1 U6449 ( .A(n4700), .ZN(n7808) );
  NAND2_X1 U6450 ( .A1(n5552), .A2(n4970), .ZN(n5554) );
  AND2_X2 U6451 ( .A1(n7686), .A2(n5703), .ZN(n7766) );
  NAND2_X1 U6452 ( .A1(n7581), .A2(n4302), .ZN(n7686) );
  INV_X1 U6453 ( .A(n5388), .ZN(n5390) );
  NAND2_X1 U6454 ( .A1(n5350), .A2(n5351), .ZN(n5388) );
  AOI21_X2 U6455 ( .B1(n8395), .B2(n5775), .A(n4703), .ZN(n4702) );
  NAND2_X1 U6456 ( .A1(n8287), .A2(n4363), .ZN(n4706) );
  NAND2_X1 U6457 ( .A1(n4706), .A2(n4708), .ZN(n8365) );
  INV_X1 U6458 ( .A(n5651), .ZN(n5652) );
  NAND2_X1 U6459 ( .A1(n4726), .A2(n4724), .ZN(n9080) );
  NAND3_X1 U6460 ( .A1(n5935), .A2(n5939), .A3(n4741), .ZN(n4745) );
  AND2_X1 U6461 ( .A1(n5924), .A2(n5933), .ZN(n4750) );
  NAND3_X1 U6462 ( .A1(n4751), .A2(n4750), .A3(n6023), .ZN(n6155) );
  INV_X1 U6463 ( .A(n9001), .ZN(n4758) );
  NAND2_X1 U6464 ( .A1(n6457), .A2(n4313), .ZN(n4764) );
  NAND3_X1 U6465 ( .A1(n4771), .A2(n4768), .A3(n6760), .ZN(P2_U3244) );
  INV_X2 U6466 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4774) );
  NAND2_X4 U6467 ( .A1(n4778), .A2(n4777), .ZN(n5104) );
  NAND2_X1 U6468 ( .A1(n5381), .A2(n4783), .ZN(n4781) );
  NAND2_X1 U6469 ( .A1(n5222), .A2(n4790), .ZN(n4787) );
  NAND2_X1 U6470 ( .A1(n5222), .A2(n5221), .ZN(n5241) );
  INV_X1 U6471 ( .A(n5221), .ZN(n4795) );
  NAND2_X1 U6472 ( .A1(n4796), .A2(n4369), .ZN(n5368) );
  NAND2_X1 U6473 ( .A1(n7891), .A2(n4827), .ZN(n4823) );
  INV_X2 U6474 ( .A(n5028), .ZN(n6987) );
  NOR2_X1 U6475 ( .A1(n4280), .A2(n6816), .ZN(n4832) );
  NAND2_X1 U6476 ( .A1(n4279), .A2(n7259), .ZN(n4833) );
  NAND2_X2 U6477 ( .A1(n5851), .A2(n4277), .ZN(n5249) );
  NAND2_X1 U6478 ( .A1(n4839), .A2(n4836), .ZN(n8565) );
  NAND2_X1 U6479 ( .A1(n4839), .A2(n4295), .ZN(n8567) );
  INV_X1 U6480 ( .A(n6678), .ZN(n4845) );
  AND2_X2 U6481 ( .A1(n4854), .A2(n4852), .ZN(n8576) );
  NAND2_X1 U6482 ( .A1(n5604), .A2(n5603), .ZN(n8500) );
  NAND2_X1 U6483 ( .A1(n8575), .A2(n4975), .ZN(n8558) );
  INV_X1 U6484 ( .A(n4975), .ZN(n4879) );
  NAND2_X1 U6485 ( .A1(n7668), .A2(n5583), .ZN(n4881) );
  INV_X1 U6486 ( .A(n5631), .ZN(n4884) );
  NAND2_X1 U6487 ( .A1(n4884), .A2(n4303), .ZN(n8240) );
  OR2_X1 U6488 ( .A1(n6238), .A2(n7162), .ZN(n4888) );
  NAND2_X1 U6489 ( .A1(n4891), .A2(n4889), .ZN(n6788) );
  NOR2_X2 U6490 ( .A1(n9328), .A2(n4909), .ZN(n4908) );
  OAI211_X1 U6491 ( .C1(n9363), .C2(n4925), .A(n4921), .B(n4920), .ZN(n9618)
         );
  NAND3_X1 U6492 ( .A1(n9363), .A2(n4286), .A3(n9620), .ZN(n4920) );
  NAND2_X1 U6493 ( .A1(n4933), .A2(n4931), .ZN(n9281) );
  OR2_X1 U6494 ( .A1(n9708), .A2(n9277), .ZN(n4935) );
  NAND2_X1 U6495 ( .A1(n4936), .A2(n4376), .ZN(n9272) );
  NAND2_X1 U6496 ( .A1(n9533), .A2(n4940), .ZN(n4938) );
  AND2_X1 U6497 ( .A1(n4957), .A2(n4358), .ZN(n9387) );
  NAND2_X1 U6498 ( .A1(n9293), .A2(n9292), .ZN(n9463) );
  AND2_X1 U6499 ( .A1(n8764), .A2(n8763), .ZN(n4977) );
  CLKBUF_X1 U6500 ( .A(n6982), .Z(n6983) );
  INV_X1 U6501 ( .A(n6155), .ZN(n5935) );
  NAND2_X1 U6502 ( .A1(n8765), .A2(n4977), .ZN(n8871) );
  OR2_X1 U6503 ( .A1(n8760), .A2(n8849), .ZN(n8764) );
  INV_X1 U6504 ( .A(n5990), .ZN(n5951) );
  AND2_X1 U6505 ( .A1(n8330), .A2(n8268), .ZN(n8270) );
  NAND2_X1 U6506 ( .A1(n5644), .A2(n10082), .ZN(n5642) );
  NAND2_X1 U6507 ( .A1(n8540), .A2(n4988), .ZN(n5644) );
  NAND2_X1 U6508 ( .A1(n8565), .A2(n6612), .ZN(n8552) );
  AND2_X1 U6509 ( .A1(n6629), .A2(n6638), .ZN(n7008) );
  INV_X1 U6510 ( .A(n7415), .ZN(n7414) );
  OR2_X1 U6511 ( .A1(n8585), .A2(n5147), .ZN(n5475) );
  OR2_X1 U6512 ( .A1(n5837), .A2(n5147), .ZN(n5524) );
  INV_X1 U6513 ( .A(n5147), .ZN(n5810) );
  OR2_X1 U6514 ( .A1(n8547), .A2(n5147), .ZN(n5505) );
  NAND2_X1 U6515 ( .A1(n9352), .A2(n9351), .ZN(n9615) );
  NAND2_X1 U6516 ( .A1(n7757), .A2(n7756), .ZN(n7799) );
  INV_X1 U6517 ( .A(n7755), .ZN(n7757) );
  NOR2_X1 U6518 ( .A1(n5806), .A2(n5805), .ZN(n5824) );
  OR2_X1 U6519 ( .A1(n5075), .A2(n5007), .ZN(n5012) );
  INV_X1 U6520 ( .A(n7611), .ZN(n7412) );
  INV_X1 U6521 ( .A(n9417), .ZN(n9419) );
  NAND2_X1 U6522 ( .A1(n9388), .A2(n7952), .ZN(n9389) );
  CLKBUF_X1 U6523 ( .A(n7052), .Z(n7358) );
  NAND2_X2 U6524 ( .A1(n9281), .A2(n9280), .ZN(n9533) );
  NAND2_X1 U6525 ( .A1(n5028), .A2(n5649), .ZN(n6639) );
  BUF_X4 U6526 ( .A(n5058), .Z(n5147) );
  INV_X1 U6527 ( .A(n4702), .ZN(n8248) );
  INV_X1 U6528 ( .A(n5008), .ZN(n5006) );
  AND2_X1 U6529 ( .A1(n9619), .A2(n9971), .ZN(n4968) );
  NAND2_X1 U6530 ( .A1(n9622), .A2(n9619), .ZN(n4969) );
  AND2_X1 U6531 ( .A1(n5551), .A2(n5550), .ZN(n4970) );
  AND2_X2 U6532 ( .A1(n5643), .A2(n5832), .ZN(n10076) );
  AND2_X2 U6533 ( .A1(n5643), .A2(n5794), .ZN(n10082) );
  AND2_X1 U6534 ( .A1(n6481), .A2(n8226), .ZN(n9726) );
  INV_X1 U6535 ( .A(n10070), .ZN(n10032) );
  AND4_X1 U6536 ( .A1(n5945), .A2(n5944), .A3(n6463), .A4(n5925), .ZN(n4971)
         );
  INV_X1 U6537 ( .A(n8371), .ZN(n8628) );
  NAND2_X1 U6538 ( .A1(n4927), .A2(n9971), .ZN(n4973) );
  OR2_X1 U6539 ( .A1(n9135), .A2(n7562), .ZN(n4974) );
  OR2_X1 U6540 ( .A1(n9419), .A2(n9302), .ZN(n4976) );
  INV_X1 U6541 ( .A(n8309), .ZN(n5602) );
  INV_X1 U6542 ( .A(n8281), .ZN(n5600) );
  INV_X1 U6543 ( .A(n9810), .ZN(n7751) );
  NAND2_X1 U6544 ( .A1(n6590), .A2(n7099), .ZN(n5650) );
  INV_X1 U6545 ( .A(n9725), .ZN(n7756) );
  OR2_X1 U6546 ( .A1(n8765), .A2(n10031), .ZN(n4978) );
  AND2_X1 U6547 ( .A1(n5221), .A2(n5201), .ZN(n4979) );
  AND2_X1 U6548 ( .A1(n5345), .A2(n5330), .ZN(n4980) );
  NAND2_X1 U6549 ( .A1(n6783), .A2(n6782), .ZN(n9553) );
  INV_X1 U6550 ( .A(n9553), .ZN(n9908) );
  AND2_X1 U6551 ( .A1(n5283), .A2(n5267), .ZN(n4981) );
  AND2_X1 U6552 ( .A1(n6699), .A2(n6705), .ZN(n4982) );
  INV_X1 U6553 ( .A(n7623), .ZN(n5580) );
  AND2_X1 U6554 ( .A1(n6450), .A2(n6448), .ZN(n4984) );
  AND2_X1 U6555 ( .A1(n7357), .A2(n7359), .ZN(n4985) );
  INV_X1 U6556 ( .A(n5606), .ZN(n8577) );
  OR2_X1 U6557 ( .A1(n6611), .A2(n6567), .ZN(n4986) );
  AND2_X1 U6558 ( .A1(n6572), .A2(n6571), .ZN(n4987) );
  OR2_X1 U6559 ( .A1(n9641), .A2(n8938), .ZN(n4989) );
  INV_X1 U6560 ( .A(n7589), .ZN(n7413) );
  NAND2_X1 U6561 ( .A1(n9337), .A2(n7952), .ZN(n7953) );
  NAND2_X1 U6562 ( .A1(n9338), .A2(n7953), .ZN(n7954) );
  INV_X1 U6563 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4997) );
  INV_X1 U6564 ( .A(n6982), .ZN(n5656) );
  NAND2_X1 U6565 ( .A1(n6575), .A2(n6611), .ZN(n6571) );
  NAND2_X1 U6566 ( .A1(n6617), .A2(n7234), .ZN(n6627) );
  INV_X1 U6567 ( .A(n7892), .ZN(n5587) );
  OR2_X1 U6568 ( .A1(n6447), .A2(n8935), .ZN(n6448) );
  AND2_X1 U6569 ( .A1(n7429), .A2(n4974), .ZN(n7430) );
  INV_X1 U6570 ( .A(n9343), .ZN(n9344) );
  INV_X1 U6571 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5940) );
  AND2_X1 U6572 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5209) );
  INV_X1 U6573 ( .A(n6756), .ZN(n5648) );
  INV_X1 U6574 ( .A(n7397), .ZN(n5679) );
  NAND2_X1 U6575 ( .A1(n7934), .A2(n5901), .ZN(n5903) );
  INV_X1 U6576 ( .A(n8523), .ZN(n8509) );
  INV_X1 U6577 ( .A(n7669), .ZN(n5582) );
  INV_X1 U6578 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5143) );
  INV_X1 U6579 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U6580 ( .A1(n7737), .A2(n7736), .ZN(n7742) );
  OR2_X1 U6581 ( .A1(n5527), .A2(n5533), .ZN(n5528) );
  INV_X1 U6582 ( .A(SI_23_), .ZN(n5463) );
  INV_X1 U6583 ( .A(SI_20_), .ZN(n5407) );
  INV_X1 U6584 ( .A(SI_16_), .ZN(n5327) );
  INV_X1 U6585 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6213) );
  AND2_X1 U6586 ( .A1(n5180), .A2(n5179), .ZN(n5181) );
  NAND2_X1 U6587 ( .A1(n5104), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5102) );
  INV_X1 U6588 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5315) );
  AND2_X1 U6589 ( .A1(n7495), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5898) );
  AND2_X1 U6590 ( .A1(n8460), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U6591 ( .A1(n6729), .A2(n6726), .ZN(n6587) );
  OR2_X1 U6592 ( .A1(n8839), .A2(n7919), .ZN(n6678) );
  NOR2_X1 U6593 ( .A1(n6109), .A2(n6108), .ZN(n6110) );
  INV_X1 U6594 ( .A(n7718), .ZN(n6171) );
  INV_X1 U6595 ( .A(n9002), .ZN(n6228) );
  INV_X1 U6596 ( .A(n9587), .ZN(n9314) );
  NAND2_X1 U6597 ( .A1(n5328), .A2(n5327), .ZN(n5345) );
  NAND2_X1 U6598 ( .A1(n5306), .A2(n5305), .ZN(n5322) );
  NAND2_X1 U6599 ( .A1(n5243), .A2(n5242), .ZN(n5262) );
  NAND2_X1 U6600 ( .A1(n5104), .A2(n6812), .ZN(n5063) );
  INV_X1 U6601 ( .A(n8666), .ZN(n8380) );
  INV_X1 U6602 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U6603 ( .A1(n8439), .A2(n8725), .ZN(n8438) );
  INV_X1 U6604 ( .A(n7374), .ZN(n7371) );
  OR2_X1 U6605 ( .A1(n7178), .A2(n8646), .ZN(n8512) );
  NAND2_X1 U6606 ( .A1(n8755), .A2(n10032), .ZN(n8756) );
  AND2_X1 U6607 ( .A1(n10033), .A2(n5608), .ZN(n8840) );
  INV_X1 U6608 ( .A(n8663), .ZN(n8563) );
  INV_X1 U6609 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8241) );
  OAI21_X1 U6610 ( .B1(n5620), .B2(n5619), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5621) );
  INV_X1 U6611 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8927) );
  OR2_X1 U6612 ( .A1(n9407), .A2(n9617), .ZN(n9641) );
  NOR2_X1 U6613 ( .A1(n6417), .A2(n6452), .ZN(n8932) );
  NAND2_X1 U6614 ( .A1(n6781), .A2(n6480), .ZN(n6873) );
  NAND2_X1 U6615 ( .A1(n6121), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6147) );
  INV_X1 U6616 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7130) );
  INV_X1 U6617 ( .A(n9388), .ZN(n9406) );
  NAND2_X1 U6618 ( .A1(n8202), .A2(n9337), .ZN(n9403) );
  OR2_X1 U6619 ( .A1(n6873), .A2(n6906), .ZN(n9260) );
  INV_X1 U6620 ( .A(n9814), .ZN(n9924) );
  INV_X1 U6621 ( .A(n9934), .ZN(n6799) );
  AND2_X1 U6622 ( .A1(n6508), .A2(n5540), .ZN(n5782) );
  INV_X1 U6623 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5973) );
  OR3_X1 U6624 ( .A1(n7889), .A2(n8900), .A3(n8902), .ZN(n5847) );
  AND2_X1 U6625 ( .A1(n5820), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8389) );
  INV_X1 U6626 ( .A(n6583), .ZN(n6584) );
  INV_X1 U6627 ( .A(n10008), .ZN(n8481) );
  AND2_X1 U6628 ( .A1(n5855), .A2(n8897), .ZN(n10007) );
  OAI21_X1 U6629 ( .B1(n8760), .B2(n8734), .A(n5841), .ZN(n5842) );
  AND2_X1 U6630 ( .A1(n5916), .A2(n5890), .ZN(n8663) );
  INV_X1 U6631 ( .A(n8336), .ZN(n8665) );
  NOR2_X1 U6632 ( .A1(n10046), .A2(n5640), .ZN(n5794) );
  INV_X1 U6633 ( .A(n8840), .ZN(n10070) );
  AND2_X1 U6634 ( .A1(n8693), .A2(n8866), .ZN(n8849) );
  INV_X1 U6635 ( .A(n8849), .ZN(n10074) );
  AND2_X1 U6636 ( .A1(n5847), .A2(n10050), .ZN(n10044) );
  AND2_X1 U6637 ( .A1(n8973), .A2(n8958), .ZN(n8959) );
  INV_X1 U6638 ( .A(n9260), .ZN(n9116) );
  OR2_X1 U6639 ( .A1(n5969), .A2(n6762), .ZN(n6882) );
  INV_X1 U6640 ( .A(n9861), .ZN(n9871) );
  INV_X1 U6641 ( .A(n9249), .ZN(n9878) );
  NOR2_X1 U6642 ( .A1(n9252), .A2(n6906), .ZN(n9861) );
  AND2_X1 U6643 ( .A1(n7145), .A2(n7144), .ZN(n7146) );
  OR2_X1 U6644 ( .A1(n9622), .A2(n4973), .ZN(n9624) );
  INV_X1 U6645 ( .A(n9971), .ZN(n9991) );
  NAND2_X1 U6646 ( .A1(n7796), .A2(n9936), .ZN(n9971) );
  XNOR2_X1 U6647 ( .A(n5949), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6466) );
  INV_X1 U6648 ( .A(n8480), .ZN(n10009) );
  INV_X1 U6649 ( .A(n6733), .ZN(n8535) );
  INV_X1 U6650 ( .A(n5822), .ZN(n5823) );
  AND2_X1 U6651 ( .A1(n5796), .A2(n10041), .ZN(n8300) );
  INV_X1 U6652 ( .A(n8291), .ZN(n8419) );
  INV_X1 U6653 ( .A(n10007), .ZN(n10011) );
  INV_X1 U6654 ( .A(n8487), .ZN(n10010) );
  AOI21_X1 U6655 ( .B1(n5570), .B2(n10021), .A(n5569), .ZN(n8540) );
  AND3_X1 U6656 ( .A1(n8700), .A2(n8699), .A3(n8698), .ZN(n8822) );
  INV_X1 U6657 ( .A(n8531), .ZN(n8734) );
  NAND2_X1 U6658 ( .A1(n10044), .A2(n5795), .ZN(n10041) );
  NAND2_X1 U6659 ( .A1(n10080), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5641) );
  INV_X1 U6660 ( .A(n10082), .ZN(n10080) );
  NAND2_X1 U6661 ( .A1(n10075), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5645) );
  INV_X1 U6662 ( .A(n10076), .ZN(n10075) );
  NAND2_X1 U6663 ( .A1(n10044), .A2(n10043), .ZN(n10047) );
  INV_X1 U6664 ( .A(n5637), .ZN(n8900) );
  INV_X1 U6665 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7387) );
  INV_X1 U6666 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U6667 ( .A1(n6499), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9842) );
  INV_X1 U6668 ( .A(n9530), .ZN(n9690) );
  INV_X1 U6669 ( .A(n9121), .ZN(n9098) );
  OR2_X1 U6670 ( .A1(n6482), .A2(n9726), .ZN(n9110) );
  INV_X1 U6671 ( .A(n9070), .ZN(n9294) );
  OR2_X1 U6672 ( .A1(n6882), .A2(P1_U3084), .ZN(n9129) );
  INV_X1 U6673 ( .A(n7505), .ZN(n9135) );
  INV_X1 U6674 ( .A(n9874), .ZN(n9241) );
  OR2_X1 U6675 ( .A1(n9925), .A2(n7433), .ZN(n9585) );
  INV_X1 U6676 ( .A(n9583), .ZN(n9603) );
  INV_X1 U6677 ( .A(n10006), .ZN(n10004) );
  OR3_X1 U6678 ( .A1(n9689), .A2(n9688), .A3(n9687), .ZN(n9747) );
  INV_X1 U6679 ( .A(n9995), .ZN(n9993) );
  AND2_X2 U6680 ( .A1(n7147), .A2(n6871), .ZN(n9995) );
  AND2_X1 U6681 ( .A1(n9935), .A2(n9931), .ZN(n9932) );
  INV_X1 U6682 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7388) );
  INV_X1 U6683 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6865) );
  INV_X1 U6684 ( .A(n9771), .ZN(n7832) );
  NOR2_X1 U6685 ( .A1(n10110), .A2(n10109), .ZN(n10108) );
  AND2_X1 U6686 ( .A1(n5844), .A2(n10050), .ZN(P2_U3966) );
  NAND2_X1 U6687 ( .A1(n4978), .A2(n5843), .ZN(P2_U3270) );
  INV_X2 U6688 ( .A(n9129), .ZN(P1_U4006) );
  INV_X2 U6689 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5628) );
  NAND3_X1 U6690 ( .A1(n5347), .A2(n4990), .A3(n5628), .ZN(n4992) );
  NOR2_X1 U6691 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n4996) );
  NAND4_X1 U6692 ( .A1(n4996), .A2(n4995), .A3(n4994), .A4(n4993), .ZN(n5331)
         );
  INV_X1 U6693 ( .A(n5331), .ZN(n4999) );
  XNOR2_X2 U6694 ( .A(n5002), .B(n8241), .ZN(n5008) );
  INV_X1 U6695 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5005) );
  INV_X1 U6696 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5007) );
  AND2_X2 U6697 ( .A1(n5008), .A2(n8267), .ZN(n5126) );
  NAND2_X1 U6698 ( .A1(n5126), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5011) );
  INV_X1 U6699 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5009) );
  OR2_X1 U6700 ( .A1(n5058), .A2(n5009), .ZN(n5010) );
  NAND2_X1 U6701 ( .A1(n5061), .A2(SI_0_), .ZN(n5014) );
  XNOR2_X1 U6702 ( .A(n5014), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8905) );
  INV_X1 U6703 ( .A(n5015), .ZN(n5016) );
  INV_X1 U6704 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5017) );
  NAND3_X1 U6705 ( .A1(n5018), .A2(P2_IR_REG_31__SCAN_IN), .A3(n5017), .ZN(
        n5019) );
  INV_X1 U6706 ( .A(n7099), .ZN(n10052) );
  NAND2_X1 U6707 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5036) );
  AND2_X1 U6708 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n5030) );
  NAND2_X1 U6709 ( .A1(n5104), .A2(n5030), .ZN(n6000) );
  OAI21_X1 U6710 ( .B1(n5104), .B2(n5036), .A(n6000), .ZN(n5021) );
  INV_X1 U6711 ( .A(SI_1_), .ZN(n5020) );
  XNOR2_X1 U6712 ( .A(n5021), .B(n5020), .ZN(n5023) );
  MUX2_X1 U6713 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5104), .Z(n5022) );
  XNOR2_X1 U6714 ( .A(n5023), .B(n5022), .ZN(n6816) );
  INV_X1 U6715 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6809) );
  INV_X1 U6716 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U6717 ( .A1(n5126), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5026) );
  INV_X1 U6718 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7263) );
  OR2_X1 U6719 ( .A1(n5058), .A2(n7263), .ZN(n5025) );
  INV_X1 U6720 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5895) );
  OR2_X1 U6721 ( .A1(n5075), .A2(n5895), .ZN(n5024) );
  AND4_X2 U6722 ( .A1(n5027), .A2(n5026), .A3(n5025), .A4(n5024), .ZN(n5649)
         );
  NAND2_X1 U6723 ( .A1(n6589), .A2(n6639), .ZN(n6629) );
  NAND2_X1 U6724 ( .A1(n5126), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5052) );
  INV_X1 U6725 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5857) );
  OR2_X1 U6726 ( .A1(n5074), .A2(n5857), .ZN(n5051) );
  INV_X1 U6727 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5029) );
  OR2_X1 U6728 ( .A1(n5058), .A2(n5029), .ZN(n5050) );
  INV_X1 U6729 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5896) );
  OR2_X1 U6730 ( .A1(n5075), .A2(n5896), .ZN(n5049) );
  AND4_X1 U6731 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(n6770)
         );
  NOR2_X1 U6732 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5033) );
  INV_X1 U6733 ( .A(n5030), .ZN(n5032) );
  NAND2_X1 U6734 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5031) );
  OAI21_X1 U6735 ( .B1(n5033), .B2(n5032), .A(n5031), .ZN(n5034) );
  NAND2_X1 U6736 ( .A1(n5104), .A2(n5034), .ZN(n5041) );
  NOR2_X1 U6737 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6738 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5035) );
  OAI21_X1 U6739 ( .B1(n5037), .B2(n5036), .A(n5035), .ZN(n5038) );
  INV_X1 U6740 ( .A(n5038), .ZN(n5039) );
  NAND2_X1 U6741 ( .A1(n5041), .A2(n5040), .ZN(n5066) );
  INV_X1 U6742 ( .A(SI_2_), .ZN(n5064) );
  XNOR2_X1 U6743 ( .A(n5066), .B(n5064), .ZN(n5043) );
  MUX2_X1 U6744 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n5061), .Z(n5042) );
  INV_X1 U6745 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U6746 ( .A1(n5044), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U6747 ( .A1(n4279), .A2(n7186), .ZN(n5046) );
  NAND4_X1 U6748 ( .A1(n5052), .A2(n5051), .A3(n5050), .A4(n5049), .ZN(n5657)
         );
  NAND2_X1 U6749 ( .A1(n5657), .A2(n7472), .ZN(n6630) );
  AND2_X1 U6750 ( .A1(n6640), .A2(n6630), .ZN(n7009) );
  NAND2_X1 U6751 ( .A1(n7008), .A2(n7009), .ZN(n7007) );
  NAND2_X1 U6752 ( .A1(n7007), .A2(n6640), .ZN(n10018) );
  INV_X1 U6753 ( .A(n5074), .ZN(n5053) );
  INV_X1 U6754 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5054) );
  OR2_X1 U6755 ( .A1(n5075), .A2(n5054), .ZN(n5056) );
  NAND2_X1 U6756 ( .A1(n5126), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5055) );
  OR2_X1 U6757 ( .A1(n5147), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5059) );
  INV_X1 U6758 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6812) );
  INV_X2 U6759 ( .A(n5104), .ZN(n5061) );
  NAND2_X1 U6760 ( .A1(n5104), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5065) );
  OAI211_X1 U6761 ( .C1(n5104), .C2(n6808), .A(n5065), .B(n5064), .ZN(n5067)
         );
  NAND2_X1 U6762 ( .A1(n5067), .A2(n5066), .ZN(n5070) );
  INV_X1 U6763 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U6764 ( .A1(n5104), .A2(n6810), .ZN(n5068) );
  OAI211_X1 U6765 ( .C1(n5104), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5068), .B(
        SI_2_), .ZN(n5069) );
  NAND2_X1 U6766 ( .A1(n5070), .A2(n5069), .ZN(n5080) );
  XNOR2_X1 U6767 ( .A(n5081), .B(n5080), .ZN(n6814) );
  NAND2_X1 U6768 ( .A1(n5071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5072) );
  XNOR2_X2 U6769 ( .A(n5072), .B(P2_IR_REG_3__SCAN_IN), .ZN(n7295) );
  NAND2_X1 U6770 ( .A1(n5393), .A2(n7295), .ZN(n5073) );
  INV_X1 U6771 ( .A(n5663), .ZN(n10035) );
  NAND2_X1 U6772 ( .A1(n10018), .A2(n10019), .ZN(n7233) );
  NAND2_X1 U6773 ( .A1(n5126), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5079) );
  INV_X1 U6774 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5865) );
  OR2_X1 U6775 ( .A1(n6526), .A2(n5865), .ZN(n5078) );
  XNOR2_X1 U6776 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7250) );
  INV_X1 U6777 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7239) );
  OR2_X1 U6778 ( .A1(n5336), .A2(n7239), .ZN(n5076) );
  INV_X4 U6779 ( .A(n6549), .ZN(n5787) );
  NAND2_X1 U6780 ( .A1(n5081), .A2(n5080), .ZN(n5084) );
  NAND2_X1 U6781 ( .A1(n5082), .A2(SI_3_), .ZN(n5083) );
  MUX2_X1 U6782 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5104), .Z(n5108) );
  XNOR2_X1 U6783 ( .A(n5108), .B(SI_4_), .ZN(n5105) );
  XNOR2_X1 U6784 ( .A(n5107), .B(n5105), .ZN(n6817) );
  NAND2_X1 U6785 ( .A1(n5787), .A2(n6817), .ZN(n5092) );
  INV_X4 U6786 ( .A(n5249), .ZN(n6562) );
  NAND2_X1 U6787 ( .A1(n6562), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5091) );
  NAND2_X1 U6788 ( .A1(n5085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5086) );
  MUX2_X1 U6789 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5086), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5089) );
  AND2_X1 U6790 ( .A1(n5089), .A2(n5088), .ZN(n7282) );
  NAND2_X1 U6791 ( .A1(n5393), .A2(n7282), .ZN(n5090) );
  INV_X1 U6792 ( .A(n6627), .ZN(n5093) );
  NAND2_X1 U6793 ( .A1(n7233), .A2(n5093), .ZN(n7055) );
  NAND2_X1 U6794 ( .A1(n5126), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5101) );
  INV_X1 U6795 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5868) );
  OR2_X1 U6796 ( .A1(n6526), .A2(n5868), .ZN(n5100) );
  INV_X1 U6797 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6798 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5094) );
  NAND2_X1 U6799 ( .A1(n5095), .A2(n5094), .ZN(n5096) );
  NAND2_X1 U6800 ( .A1(n5130), .A2(n5096), .ZN(n7390) );
  OR2_X1 U6801 ( .A1(n5147), .A2(n7390), .ZN(n5099) );
  INV_X1 U6802 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5097) );
  OR2_X1 U6803 ( .A1(n5336), .A2(n5097), .ZN(n5098) );
  OAI21_X1 U6804 ( .B1(n5104), .B2(n5103), .A(n5102), .ZN(n5114) );
  INV_X1 U6805 ( .A(n5105), .ZN(n5106) );
  NAND2_X1 U6806 ( .A1(n5107), .A2(n5106), .ZN(n5122) );
  NAND2_X1 U6807 ( .A1(n5108), .A2(SI_4_), .ZN(n5115) );
  NAND2_X1 U6808 ( .A1(n5122), .A2(n5115), .ZN(n5109) );
  XNOR2_X1 U6809 ( .A(n5116), .B(n5109), .ZN(n6821) );
  NAND2_X1 U6810 ( .A1(n6821), .A2(n5787), .ZN(n5112) );
  NAND2_X1 U6811 ( .A1(n5088), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5110) );
  AOI22_X1 U6812 ( .A1(n6562), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n5393), .B2(
        n7336), .ZN(n5111) );
  NAND2_X1 U6813 ( .A1(n8432), .A2(n7393), .ZN(n6618) );
  NAND2_X1 U6814 ( .A1(n8433), .A2(n10063), .ZN(n7054) );
  AND2_X1 U6815 ( .A1(n6618), .A2(n7054), .ZN(n6621) );
  NAND2_X1 U6816 ( .A1(n7055), .A2(n6621), .ZN(n5113) );
  NAND2_X1 U6817 ( .A1(n5113), .A2(n6625), .ZN(n7370) );
  NAND2_X1 U6818 ( .A1(n5114), .A2(SI_5_), .ZN(n5117) );
  AND2_X1 U6819 ( .A1(n5115), .A2(n5117), .ZN(n5121) );
  INV_X1 U6820 ( .A(n5116), .ZN(n5119) );
  INV_X1 U6821 ( .A(n5117), .ZN(n5118) );
  NOR2_X1 U6822 ( .A1(n5119), .A2(n5118), .ZN(n5120) );
  AOI21_X2 U6823 ( .B1(n5122), .B2(n5121), .A(n5120), .ZN(n5139) );
  XNOR2_X1 U6824 ( .A(n5140), .B(SI_6_), .ZN(n5137) );
  XNOR2_X1 U6825 ( .A(n5139), .B(n5137), .ZN(n6080) );
  NAND2_X1 U6826 ( .A1(n6080), .A2(n5787), .ZN(n5125) );
  OR2_X1 U6827 ( .A1(n5351), .A2(n5204), .ZN(n5123) );
  XNOR2_X1 U6828 ( .A(n5123), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7310) );
  AOI22_X1 U6829 ( .A1(n6562), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5393), .B2(
        n7310), .ZN(n5124) );
  INV_X1 U6830 ( .A(n7382), .ZN(n10071) );
  NAND2_X1 U6831 ( .A1(n5126), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5136) );
  INV_X1 U6832 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5127) );
  OR2_X1 U6833 ( .A1(n6526), .A2(n5127), .ZN(n5135) );
  INV_X1 U6834 ( .A(n5130), .ZN(n5128) );
  INV_X1 U6835 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6836 ( .A1(n5130), .A2(n5129), .ZN(n5131) );
  NAND2_X1 U6837 ( .A1(n5150), .A2(n5131), .ZN(n7380) );
  OR2_X1 U6838 ( .A1(n5147), .A2(n7380), .ZN(n5134) );
  INV_X1 U6839 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5132) );
  OR2_X1 U6840 ( .A1(n5336), .A2(n5132), .ZN(n5133) );
  NAND4_X1 U6841 ( .A1(n5136), .A2(n5135), .A3(n5134), .A4(n5133), .ZN(n8431)
         );
  NAND2_X1 U6842 ( .A1(n10071), .A2(n8431), .ZN(n6644) );
  INV_X1 U6843 ( .A(n8431), .ZN(n7462) );
  NAND2_X1 U6844 ( .A1(n6644), .A2(n6649), .ZN(n7374) );
  NAND2_X1 U6845 ( .A1(n7370), .A2(n7371), .ZN(n7369) );
  NAND2_X1 U6846 ( .A1(n7369), .A2(n6649), .ZN(n7355) );
  INV_X1 U6847 ( .A(n5137), .ZN(n5138) );
  NAND2_X1 U6848 ( .A1(n5140), .A2(SI_6_), .ZN(n5141) );
  MUX2_X1 U6849 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4277), .Z(n5159) );
  XNOR2_X1 U6850 ( .A(n5159), .B(SI_7_), .ZN(n5156) );
  XNOR2_X1 U6851 ( .A(n5158), .B(n5156), .ZN(n6829) );
  NAND2_X1 U6852 ( .A1(n6829), .A2(n5787), .ZN(n5146) );
  NAND2_X1 U6853 ( .A1(n5351), .A2(n5143), .ZN(n5165) );
  NAND2_X1 U6854 ( .A1(n5165), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5144) );
  XNOR2_X1 U6855 ( .A(n5144), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7322) );
  AOI22_X1 U6856 ( .A1(n6562), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5393), .B2(
        n7322), .ZN(n5145) );
  NAND2_X1 U6857 ( .A1(n5146), .A2(n5145), .ZN(n7466) );
  NAND2_X1 U6858 ( .A1(n6520), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5155) );
  INV_X1 U6859 ( .A(n5126), .ZN(n5274) );
  INV_X1 U6860 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10176) );
  OR2_X1 U6861 ( .A1(n5274), .A2(n10176), .ZN(n5154) );
  INV_X1 U6862 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6863 ( .A1(n5150), .A2(n5149), .ZN(n5151) );
  NAND2_X1 U6864 ( .A1(n5172), .A2(n5151), .ZN(n7463) );
  OR2_X1 U6865 ( .A1(n5147), .A2(n7463), .ZN(n5153) );
  INV_X1 U6866 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7364) );
  OR2_X1 U6867 ( .A1(n6527), .A2(n7364), .ZN(n5152) );
  AND4_X2 U6868 ( .A1(n5155), .A2(n5154), .A3(n5153), .A4(n5152), .ZN(n7624)
         );
  NAND2_X1 U6869 ( .A1(n7466), .A2(n7624), .ZN(n6650) );
  NAND2_X1 U6870 ( .A1(n6651), .A2(n6650), .ZN(n5574) );
  INV_X1 U6871 ( .A(n5574), .ZN(n7360) );
  NAND2_X1 U6872 ( .A1(n7355), .A2(n7360), .ZN(n7354) );
  NAND2_X1 U6873 ( .A1(n7354), .A2(n6650), .ZN(n7622) );
  INV_X1 U6874 ( .A(n5156), .ZN(n5157) );
  NAND2_X1 U6875 ( .A1(n5159), .A2(SI_7_), .ZN(n5179) );
  NAND2_X1 U6876 ( .A1(n5182), .A2(n5179), .ZN(n5164) );
  INV_X1 U6877 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6839) );
  INV_X1 U6878 ( .A(SI_8_), .ZN(n5160) );
  NAND2_X1 U6879 ( .A1(n5161), .A2(n5160), .ZN(n5217) );
  INV_X1 U6880 ( .A(n5161), .ZN(n5162) );
  NAND2_X1 U6881 ( .A1(n5162), .A2(SI_8_), .ZN(n5163) );
  NAND2_X1 U6882 ( .A1(n5217), .A2(n5163), .ZN(n5178) );
  XNOR2_X1 U6883 ( .A(n5178), .B(n5164), .ZN(n6834) );
  NAND2_X1 U6884 ( .A1(n6834), .A2(n5787), .ZN(n5169) );
  NAND2_X1 U6885 ( .A1(n5332), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5166) );
  MUX2_X1 U6886 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5166), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5167) );
  AOI22_X1 U6887 ( .A1(n6562), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5393), .B2(
        n7201), .ZN(n5168) );
  NAND2_X1 U6888 ( .A1(n6520), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5177) );
  INV_X1 U6889 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10231) );
  OR2_X1 U6890 ( .A1(n5274), .A2(n10231), .ZN(n5176) );
  INV_X1 U6891 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6892 ( .A1(n5172), .A2(n5171), .ZN(n5173) );
  NAND2_X1 U6893 ( .A1(n5208), .A2(n5173), .ZN(n7630) );
  OR2_X1 U6894 ( .A1(n5147), .A2(n7630), .ZN(n5175) );
  INV_X1 U6895 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7628) );
  OR2_X1 U6896 ( .A1(n6527), .A2(n7628), .ZN(n5174) );
  OR2_X1 U6897 ( .A1(n8860), .A2(n7691), .ZN(n6654) );
  NAND2_X1 U6898 ( .A1(n8860), .A2(n7691), .ZN(n6655) );
  NAND2_X1 U6899 ( .A1(n7622), .A2(n7623), .ZN(n7621) );
  NAND2_X1 U6900 ( .A1(n7621), .A2(n6655), .ZN(n7665) );
  INV_X1 U6901 ( .A(n5178), .ZN(n5180) );
  MUX2_X1 U6902 ( .A(n6844), .B(n6845), .S(n4277), .Z(n5184) );
  INV_X1 U6903 ( .A(SI_9_), .ZN(n5183) );
  NAND2_X1 U6904 ( .A1(n5184), .A2(n5183), .ZN(n5216) );
  INV_X1 U6905 ( .A(n5184), .ZN(n5185) );
  NAND2_X1 U6906 ( .A1(n5185), .A2(SI_9_), .ZN(n5219) );
  AND2_X1 U6907 ( .A1(n5216), .A2(n5219), .ZN(n5194) );
  NAND2_X1 U6908 ( .A1(n6842), .A2(n5787), .ZN(n5188) );
  NAND2_X1 U6909 ( .A1(n5203), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5186) );
  XNOR2_X1 U6910 ( .A(n5186), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7213) );
  AOI22_X1 U6911 ( .A1(n6562), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5393), .B2(
        n7213), .ZN(n5187) );
  NAND2_X1 U6912 ( .A1(n6524), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5193) );
  INV_X1 U6913 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5873) );
  OR2_X1 U6914 ( .A1(n6526), .A2(n5873), .ZN(n5192) );
  INV_X1 U6915 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5207) );
  XNOR2_X1 U6916 ( .A(n5208), .B(n5207), .ZN(n7692) );
  OR2_X1 U6917 ( .A1(n5147), .A2(n7692), .ZN(n5191) );
  INV_X1 U6918 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5189) );
  OR2_X1 U6919 ( .A1(n6527), .A2(n5189), .ZN(n5190) );
  OR2_X1 U6920 ( .A1(n8855), .A2(n7767), .ZN(n6663) );
  NAND2_X1 U6921 ( .A1(n8855), .A2(n7767), .ZN(n6658) );
  NAND2_X1 U6922 ( .A1(n7665), .A2(n7669), .ZN(n7664) );
  NAND2_X1 U6923 ( .A1(n7664), .A2(n6658), .ZN(n7698) );
  NAND2_X1 U6924 ( .A1(n5196), .A2(n5216), .ZN(n5202) );
  INV_X1 U6925 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5197) );
  MUX2_X1 U6926 ( .A(n5197), .B(n6848), .S(n4277), .Z(n5199) );
  INV_X1 U6927 ( .A(SI_10_), .ZN(n5198) );
  NAND2_X1 U6928 ( .A1(n5199), .A2(n5198), .ZN(n5221) );
  INV_X1 U6929 ( .A(n5199), .ZN(n5200) );
  NAND2_X1 U6930 ( .A1(n5200), .A2(SI_10_), .ZN(n5201) );
  OR2_X1 U6931 ( .A1(n5247), .A2(n5204), .ZN(n5224) );
  XNOR2_X1 U6932 ( .A(n5224), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7495) );
  AOI22_X1 U6933 ( .A1(n7495), .A2(n5393), .B1(n6562), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6934 ( .A1(n6520), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5215) );
  INV_X1 U6935 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10213) );
  OR2_X1 U6936 ( .A1(n5274), .A2(n10213), .ZN(n5214) );
  INV_X1 U6937 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5206) );
  OAI21_X1 U6938 ( .B1(n5208), .B2(n5207), .A(n5206), .ZN(n5211) );
  NAND2_X1 U6939 ( .A1(n5211), .A2(n5229), .ZN(n7768) );
  OR2_X1 U6940 ( .A1(n5147), .A2(n7768), .ZN(n5213) );
  INV_X1 U6941 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7707) );
  OR2_X1 U6942 ( .A1(n6527), .A2(n7707), .ZN(n5212) );
  OR2_X1 U6943 ( .A1(n8850), .A2(n7847), .ZN(n6665) );
  NAND2_X1 U6944 ( .A1(n6665), .A2(n6667), .ZN(n7702) );
  INV_X1 U6945 ( .A(n7702), .ZN(n7699) );
  MUX2_X1 U6946 ( .A(n6852), .B(n6850), .S(n4277), .Z(n5237) );
  NAND2_X1 U6947 ( .A1(n6849), .A2(n5787), .ZN(n5228) );
  INV_X1 U6948 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U6949 ( .A1(n5224), .A2(n5223), .ZN(n5225) );
  NAND2_X1 U6950 ( .A1(n5225), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5226) );
  XNOR2_X1 U6951 ( .A(n5226), .B(P2_IR_REG_11__SCAN_IN), .ZN(n5900) );
  AOI22_X1 U6952 ( .A1(n5900), .A2(n5393), .B1(n6562), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6953 ( .A1(n5126), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5234) );
  INV_X1 U6954 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5874) );
  OR2_X1 U6955 ( .A1(n6526), .A2(n5874), .ZN(n5233) );
  OR2_X2 U6956 ( .A1(n5229), .A2(n7846), .ZN(n5255) );
  NAND2_X1 U6957 ( .A1(n5229), .A2(n7846), .ZN(n5230) );
  NAND2_X1 U6958 ( .A1(n5255), .A2(n5230), .ZN(n7848) );
  OR2_X1 U6959 ( .A1(n5147), .A2(n7848), .ZN(n5232) );
  INV_X1 U6960 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7729) );
  OR2_X1 U6961 ( .A1(n6527), .A2(n7729), .ZN(n5231) );
  NAND2_X1 U6962 ( .A1(n8844), .A2(n7908), .ZN(n6675) );
  INV_X1 U6963 ( .A(n6675), .ZN(n5235) );
  INV_X1 U6964 ( .A(n5237), .ZN(n5238) );
  NAND2_X1 U6965 ( .A1(n5238), .A2(SI_11_), .ZN(n5239) );
  MUX2_X1 U6966 ( .A(n10220), .B(n6865), .S(n4276), .Z(n5243) );
  INV_X1 U6967 ( .A(SI_12_), .ZN(n5242) );
  INV_X1 U6968 ( .A(n5243), .ZN(n5244) );
  NAND2_X1 U6969 ( .A1(n5244), .A2(SI_12_), .ZN(n5245) );
  NAND2_X1 U6970 ( .A1(n6862), .A2(n5787), .ZN(n5252) );
  NOR2_X1 U6971 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5246) );
  OR2_X1 U6972 ( .A1(n5269), .A2(n5204), .ZN(n5248) );
  XNOR2_X1 U6973 ( .A(n5248), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7826) );
  NOR2_X1 U6974 ( .A1(n6547), .A2(n10220), .ZN(n5250) );
  AOI21_X1 U6975 ( .B1(n7826), .B2(n5393), .A(n5250), .ZN(n5251) );
  NAND2_X1 U6976 ( .A1(n6520), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5261) );
  INV_X1 U6977 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5253) );
  OR2_X1 U6978 ( .A1(n6527), .A2(n5253), .ZN(n5260) );
  NAND2_X1 U6979 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  NAND2_X1 U6980 ( .A1(n5276), .A2(n5256), .ZN(n7909) );
  OR2_X1 U6981 ( .A1(n5147), .A2(n7909), .ZN(n5259) );
  INV_X1 U6982 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5257) );
  OR2_X1 U6983 ( .A1(n5274), .A2(n5257), .ZN(n5258) );
  NAND2_X1 U6984 ( .A1(n8839), .A2(n7919), .ZN(n6676) );
  MUX2_X1 U6985 ( .A(n5264), .B(n6866), .S(n4277), .Z(n5265) );
  INV_X1 U6986 ( .A(n5265), .ZN(n5266) );
  NAND2_X1 U6987 ( .A1(n5266), .A2(SI_13_), .ZN(n5267) );
  XNOR2_X1 U6988 ( .A(n5282), .B(n4981), .ZN(n6860) );
  NAND2_X1 U6989 ( .A1(n6860), .A2(n5787), .ZN(n5272) );
  INV_X1 U6990 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6991 ( .A1(n5269), .A2(n5268), .ZN(n5285) );
  NAND2_X1 U6992 ( .A1(n5285), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5270) );
  XNOR2_X1 U6993 ( .A(n5270), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7870) );
  AOI22_X1 U6994 ( .A1(n7870), .A2(n5393), .B1(n6562), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6995 ( .A1(n6520), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5281) );
  INV_X1 U6996 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n5273) );
  OR2_X1 U6997 ( .A1(n5274), .A2(n5273), .ZN(n5280) );
  INV_X1 U6998 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U6999 ( .A1(n5276), .A2(n10245), .ZN(n5277) );
  NAND2_X1 U7000 ( .A1(n5316), .A2(n5277), .ZN(n7920) );
  OR2_X1 U7001 ( .A1(n5147), .A2(n7920), .ZN(n5279) );
  INV_X1 U7002 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5892) );
  OR2_X1 U7003 ( .A1(n6527), .A2(n5892), .ZN(n5278) );
  OR2_X1 U7004 ( .A1(n8833), .A2(n8273), .ZN(n6682) );
  NAND2_X1 U7005 ( .A1(n8833), .A2(n8273), .ZN(n7890) );
  MUX2_X1 U7006 ( .A(n6879), .B(n6880), .S(n4277), .Z(n5300) );
  XNOR2_X1 U7007 ( .A(n5304), .B(n5299), .ZN(n6878) );
  NAND2_X1 U7008 ( .A1(n6878), .A2(n5787), .ZN(n5292) );
  NAND2_X1 U7009 ( .A1(n5286), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5289) );
  INV_X1 U7010 ( .A(n5289), .ZN(n5287) );
  NAND2_X1 U7011 ( .A1(n5287), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5290) );
  INV_X1 U7012 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U7013 ( .A1(n5289), .A2(n5288), .ZN(n5309) );
  AOI22_X1 U7014 ( .A1(n5902), .A2(n5393), .B1(n6562), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U7015 ( .A1(n6524), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5296) );
  INV_X1 U7016 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5879) );
  OR2_X1 U7017 ( .A1(n6526), .A2(n5879), .ZN(n5295) );
  INV_X1 U7018 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5901) );
  OR2_X1 U7019 ( .A1(n6527), .A2(n5901), .ZN(n5294) );
  XNOR2_X1 U7020 ( .A(n5316), .B(n5315), .ZN(n8274) );
  OR2_X1 U7021 ( .A1(n5147), .A2(n8274), .ZN(n5293) );
  NAND2_X1 U7022 ( .A1(n8828), .A2(n8404), .ZN(n6686) );
  INV_X1 U7023 ( .A(n7890), .ZN(n5297) );
  NOR2_X1 U7024 ( .A1(n5587), .A2(n5297), .ZN(n5298) );
  INV_X1 U7025 ( .A(n5300), .ZN(n5301) );
  NAND2_X1 U7026 ( .A1(n5301), .A2(SI_14_), .ZN(n5302) );
  MUX2_X1 U7027 ( .A(n7086), .B(n7084), .S(n4277), .Z(n5306) );
  INV_X1 U7028 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U7029 ( .A1(n5307), .A2(SI_15_), .ZN(n5308) );
  NAND2_X1 U7030 ( .A1(n5322), .A2(n5308), .ZN(n5323) );
  XNOR2_X1 U7031 ( .A(n5324), .B(n5323), .ZN(n7083) );
  NAND2_X1 U7032 ( .A1(n7083), .A2(n5787), .ZN(n5312) );
  NAND2_X1 U7033 ( .A1(n5309), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5310) );
  XNOR2_X1 U7034 ( .A(n5310), .B(P2_IR_REG_15__SCAN_IN), .ZN(n5904) );
  AOI22_X1 U7035 ( .A1(n5904), .A2(n5393), .B1(n6562), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U7036 ( .A1(n6524), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5321) );
  INV_X1 U7037 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5313) );
  OR2_X1 U7038 ( .A1(n6526), .A2(n5313), .ZN(n5320) );
  INV_X1 U7039 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8725) );
  OR2_X1 U7040 ( .A1(n6527), .A2(n8725), .ZN(n5319) );
  OAI21_X1 U7041 ( .B1(n5316), .B2(n5315), .A(n5314), .ZN(n5317) );
  NAND2_X1 U7042 ( .A1(n5317), .A2(n5337), .ZN(n8724) );
  OR2_X1 U7043 ( .A1(n5147), .A2(n8724), .ZN(n5318) );
  NAND2_X1 U7044 ( .A1(n8824), .A2(n8324), .ZN(n6691) );
  NAND2_X1 U7045 ( .A1(n6690), .A2(n6691), .ZN(n8721) );
  INV_X1 U7046 ( .A(n8721), .ZN(n6689) );
  MUX2_X1 U7047 ( .A(n5326), .B(n5325), .S(n4277), .Z(n5328) );
  INV_X1 U7048 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U7049 ( .A1(n5329), .A2(SI_16_), .ZN(n5330) );
  XNOR2_X1 U7050 ( .A(n5344), .B(n4980), .ZN(n7174) );
  NAND2_X1 U7051 ( .A1(n7174), .A2(n5787), .ZN(n5335) );
  NAND2_X1 U7052 ( .A1(n5620), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5333) );
  XNOR2_X1 U7053 ( .A(n5333), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8460) );
  AOI22_X1 U7054 ( .A1(n6562), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5393), .B2(
        n8460), .ZN(n5334) );
  INV_X1 U7055 ( .A(n5336), .ZN(n5561) );
  NAND2_X1 U7056 ( .A1(n5561), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U7057 ( .A1(n6524), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5341) );
  INV_X1 U7058 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n5882) );
  OR2_X1 U7059 ( .A1(n6526), .A2(n5882), .ZN(n5340) );
  INV_X1 U7060 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U7061 ( .A1(n5337), .A2(n8452), .ZN(n5338) );
  NAND2_X1 U7062 ( .A1(n5358), .A2(n5338), .ZN(n8706) );
  OR2_X1 U7063 ( .A1(n5147), .A2(n8706), .ZN(n5339) );
  NAND4_X1 U7064 ( .A1(n5342), .A2(n5341), .A3(n5340), .A4(n5339), .ZN(n8421)
         );
  NAND2_X1 U7065 ( .A1(n8815), .A2(n8421), .ZN(n6696) );
  INV_X1 U7066 ( .A(n8421), .ZN(n8335) );
  NAND2_X1 U7067 ( .A1(n8709), .A2(n8335), .ZN(n6695) );
  MUX2_X1 U7068 ( .A(n7387), .B(n7388), .S(n4277), .Z(n5365) );
  XNOR2_X1 U7069 ( .A(n5363), .B(n5364), .ZN(n7386) );
  NAND2_X1 U7070 ( .A1(n7386), .A2(n5787), .ZN(n5354) );
  OAI21_X1 U7071 ( .B1(n5620), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5346) );
  MUX2_X1 U7072 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5346), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5352) );
  NAND2_X1 U7073 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  NOR2_X1 U7074 ( .A1(n5331), .A2(n5349), .ZN(n5350) );
  NAND2_X1 U7075 ( .A1(n5352), .A2(n5388), .ZN(n8473) );
  INV_X1 U7076 ( .A(n8473), .ZN(n5908) );
  AOI22_X1 U7077 ( .A1(n5908), .A2(n5393), .B1(n6562), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U7078 ( .A1(n6520), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U7079 ( .A1(n5126), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5355) );
  AND2_X1 U7080 ( .A1(n5356), .A2(n5355), .ZN(n5362) );
  NAND2_X1 U7081 ( .A1(n5358), .A2(n5357), .ZN(n5359) );
  AND2_X1 U7082 ( .A1(n5374), .A2(n5359), .ZN(n8679) );
  NAND2_X1 U7083 ( .A1(n8679), .A2(n5810), .ZN(n5361) );
  NAND2_X1 U7084 ( .A1(n5561), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U7085 ( .A1(n8811), .A2(n8382), .ZN(n6614) );
  INV_X1 U7086 ( .A(n5365), .ZN(n5366) );
  NAND2_X1 U7087 ( .A1(n5366), .A2(SI_17_), .ZN(n5367) );
  NAND2_X1 U7088 ( .A1(n5368), .A2(n5367), .ZN(n5381) );
  MUX2_X1 U7089 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4277), .Z(n5382) );
  XNOR2_X1 U7090 ( .A(n5381), .B(n5379), .ZN(n7485) );
  NAND2_X1 U7091 ( .A1(n7485), .A2(n5787), .ZN(n5371) );
  NAND2_X1 U7092 ( .A1(n5388), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5369) );
  XNOR2_X1 U7093 ( .A(n5369), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8486) );
  AOI22_X1 U7094 ( .A1(n6562), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5393), .B2(
        n8486), .ZN(n5370) );
  INV_X1 U7095 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5378) );
  INV_X1 U7096 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U7097 ( .A1(n5374), .A2(n5373), .ZN(n5375) );
  NAND2_X1 U7098 ( .A1(n5397), .A2(n5375), .ZN(n8657) );
  OR2_X1 U7099 ( .A1(n8657), .A2(n5147), .ZN(n5377) );
  AOI22_X1 U7100 ( .A1(n5126), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n6520), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n5376) );
  OAI211_X1 U7101 ( .C1(n6527), .C2(n5378), .A(n5377), .B(n5376), .ZN(n8420)
         );
  INV_X1 U7102 ( .A(n8420), .ZN(n8337) );
  OR2_X1 U7103 ( .A1(n8805), .A2(n8337), .ZN(n6699) );
  NAND2_X1 U7104 ( .A1(n8805), .A2(n8337), .ZN(n6705) );
  NAND2_X1 U7105 ( .A1(n8662), .A2(n4982), .ZN(n8661) );
  NAND2_X1 U7106 ( .A1(n8661), .A2(n6705), .ZN(n8636) );
  NAND2_X1 U7107 ( .A1(n5382), .A2(SI_18_), .ZN(n5383) );
  MUX2_X1 U7108 ( .A(n7559), .B(n7561), .S(n4277), .Z(n5385) );
  INV_X1 U7109 ( .A(n5385), .ZN(n5386) );
  NAND2_X1 U7110 ( .A1(n5386), .A2(SI_19_), .ZN(n5387) );
  NAND2_X1 U7111 ( .A1(n5404), .A2(n5387), .ZN(n5405) );
  XNOR2_X1 U7112 ( .A(n5406), .B(n5405), .ZN(n7557) );
  NAND2_X1 U7113 ( .A1(n7557), .A2(n5787), .ZN(n5395) );
  NAND2_X1 U7114 ( .A1(n5390), .A2(n5389), .ZN(n5549) );
  INV_X4 U7115 ( .A(n7558), .ZN(n8646) );
  AOI22_X1 U7116 ( .A1(n6562), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8646), .B2(
        n5393), .ZN(n5394) );
  INV_X1 U7117 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U7118 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  NAND2_X1 U7119 ( .A1(n5413), .A2(n5398), .ZN(n8648) );
  OR2_X1 U7120 ( .A1(n8648), .A2(n5147), .ZN(n5403) );
  INV_X1 U7121 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7122 ( .A1(n6524), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5400) );
  NAND2_X1 U7123 ( .A1(n5561), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5399) );
  OAI211_X1 U7124 ( .C1(n6526), .C2(n5888), .A(n5400), .B(n5399), .ZN(n5401)
         );
  INV_X1 U7125 ( .A(n5401), .ZN(n5402) );
  NAND2_X1 U7126 ( .A1(n5403), .A2(n5402), .ZN(n8666) );
  OR2_X1 U7127 ( .A1(n8802), .A2(n8380), .ZN(n6707) );
  NAND2_X1 U7128 ( .A1(n8802), .A2(n8380), .ZN(n6709) );
  MUX2_X1 U7129 ( .A(n7663), .B(n7648), .S(n4277), .Z(n5408) );
  INV_X1 U7130 ( .A(n5408), .ZN(n5409) );
  NAND2_X1 U7131 ( .A1(n5409), .A2(SI_20_), .ZN(n5410) );
  XNOR2_X1 U7132 ( .A(n5422), .B(n5421), .ZN(n7647) );
  NAND2_X1 U7133 ( .A1(n7647), .A2(n5787), .ZN(n5412) );
  NAND2_X1 U7134 ( .A1(n6562), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5411) );
  INV_X1 U7135 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U7136 ( .A1(n5413), .A2(n10232), .ZN(n5414) );
  NAND2_X1 U7137 ( .A1(n5427), .A2(n5414), .ZN(n8622) );
  OR2_X1 U7138 ( .A1(n8622), .A2(n5147), .ZN(n5420) );
  INV_X1 U7139 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U7140 ( .A1(n6520), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U7141 ( .A1(n6524), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5415) );
  OAI211_X1 U7142 ( .C1(n6527), .C2(n5417), .A(n5416), .B(n5415), .ZN(n5418)
         );
  INV_X1 U7143 ( .A(n5418), .ZN(n5419) );
  NAND2_X1 U7144 ( .A1(n8796), .A2(n8291), .ZN(n6710) );
  NAND2_X1 U7145 ( .A1(n8605), .A2(n6710), .ZN(n8627) );
  MUX2_X1 U7146 ( .A(n7685), .B(n7682), .S(n4277), .Z(n5440) );
  XNOR2_X1 U7147 ( .A(n5440), .B(SI_21_), .ZN(n5437) );
  NAND2_X1 U7148 ( .A1(n7680), .A2(n5787), .ZN(n5426) );
  NAND2_X1 U7149 ( .A1(n6562), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5425) );
  INV_X1 U7150 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8299) );
  NAND2_X1 U7151 ( .A1(n5427), .A2(n8299), .ZN(n5428) );
  AND2_X1 U7152 ( .A1(n5450), .A2(n5428), .ZN(n8614) );
  NAND2_X1 U7153 ( .A1(n8614), .A2(n5810), .ZN(n5434) );
  INV_X1 U7154 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U7155 ( .A1(n6520), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U7156 ( .A1(n6524), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5429) );
  OAI211_X1 U7157 ( .C1(n5431), .C2(n6527), .A(n5430), .B(n5429), .ZN(n5432)
         );
  INV_X1 U7158 ( .A(n5432), .ZN(n5433) );
  OR2_X1 U7159 ( .A1(n8793), .A2(n8371), .ZN(n6712) );
  NAND2_X1 U7160 ( .A1(n8793), .A2(n8371), .ZN(n6714) );
  NAND2_X1 U7161 ( .A1(n6712), .A2(n6714), .ZN(n8610) );
  INV_X1 U7162 ( .A(n8605), .ZN(n5435) );
  NOR2_X1 U7163 ( .A1(n8610), .A2(n5435), .ZN(n5436) );
  INV_X1 U7164 ( .A(n5437), .ZN(n5438) );
  INV_X1 U7165 ( .A(n5440), .ZN(n5441) );
  NAND2_X1 U7166 ( .A1(n5441), .A2(SI_21_), .ZN(n5442) );
  MUX2_X1 U7167 ( .A(n7835), .B(n7831), .S(n4277), .Z(n5444) );
  INV_X1 U7168 ( .A(SI_22_), .ZN(n5443) );
  NAND2_X1 U7169 ( .A1(n5444), .A2(n5443), .ZN(n5458) );
  INV_X1 U7170 ( .A(n5444), .ZN(n5445) );
  NAND2_X1 U7171 ( .A1(n5445), .A2(SI_22_), .ZN(n5446) );
  NAND2_X1 U7172 ( .A1(n5458), .A2(n5446), .ZN(n5459) );
  XNOR2_X1 U7173 ( .A(n5460), .B(n5459), .ZN(n7830) );
  NAND2_X1 U7174 ( .A1(n7830), .A2(n5787), .ZN(n5448) );
  NAND2_X1 U7175 ( .A1(n6562), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5447) );
  INV_X1 U7176 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U7177 ( .A1(n5450), .A2(n8370), .ZN(n5451) );
  NAND2_X1 U7178 ( .A1(n5469), .A2(n5451), .ZN(n8591) );
  OR2_X1 U7179 ( .A1(n8591), .A2(n5147), .ZN(n5457) );
  INV_X1 U7180 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U7181 ( .A1(n6520), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U7182 ( .A1(n6524), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5452) );
  OAI211_X1 U7183 ( .C1(n6527), .C2(n5454), .A(n5453), .B(n5452), .ZN(n5455)
         );
  INV_X1 U7184 ( .A(n5455), .ZN(n5456) );
  NAND2_X1 U7185 ( .A1(n8786), .A2(n8281), .ZN(n6716) );
  NAND2_X1 U7186 ( .A1(n6704), .A2(n6716), .ZN(n6598) );
  INV_X1 U7187 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5462) );
  INV_X1 U7188 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5461) );
  MUX2_X1 U7189 ( .A(n5462), .B(n5461), .S(n4277), .Z(n5464) );
  NAND2_X1 U7190 ( .A1(n5464), .A2(n5463), .ZN(n5478) );
  INV_X1 U7191 ( .A(n5464), .ZN(n5465) );
  NAND2_X1 U7192 ( .A1(n5465), .A2(SI_23_), .ZN(n5466) );
  NAND2_X1 U7193 ( .A1(n7836), .A2(n5787), .ZN(n5468) );
  NAND2_X1 U7194 ( .A1(n6562), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5467) );
  INV_X1 U7195 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8282) );
  OR2_X2 U7196 ( .A1(n5469), .A2(n8282), .ZN(n5481) );
  NAND2_X1 U7197 ( .A1(n5469), .A2(n8282), .ZN(n5470) );
  NAND2_X1 U7198 ( .A1(n5481), .A2(n5470), .ZN(n8585) );
  INV_X1 U7199 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U7200 ( .A1(n6520), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U7201 ( .A1(n5126), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5471) );
  OAI211_X1 U7202 ( .C1(n6527), .C2(n8578), .A(n5472), .B(n5471), .ZN(n5473)
         );
  INV_X1 U7203 ( .A(n5473), .ZN(n5474) );
  MUX2_X1 U7204 ( .A(n7887), .B(n7885), .S(n4277), .Z(n5488) );
  XNOR2_X1 U7205 ( .A(n5488), .B(SI_24_), .ZN(n5487) );
  XNOR2_X1 U7206 ( .A(n5490), .B(n5487), .ZN(n7884) );
  NAND2_X1 U7207 ( .A1(n7884), .A2(n5787), .ZN(n5480) );
  NAND2_X1 U7208 ( .A1(n6562), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5479) );
  INV_X1 U7209 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8350) );
  OR2_X2 U7210 ( .A1(n5481), .A2(n8350), .ZN(n5499) );
  NAND2_X1 U7211 ( .A1(n5481), .A2(n8350), .ZN(n5482) );
  INV_X1 U7212 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U7213 ( .A1(n6520), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7214 ( .A1(n6524), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5483) );
  OAI211_X1 U7215 ( .C1(n5485), .C2(n6527), .A(n5484), .B(n5483), .ZN(n5486)
         );
  NAND2_X1 U7216 ( .A1(n8776), .A2(n8309), .ZN(n6613) );
  INV_X1 U7217 ( .A(n5488), .ZN(n5489) );
  INV_X1 U7218 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8903) );
  INV_X1 U7219 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5491) );
  MUX2_X1 U7220 ( .A(n8903), .B(n5491), .S(n4277), .Z(n5493) );
  INV_X1 U7221 ( .A(SI_25_), .ZN(n5492) );
  NAND2_X1 U7222 ( .A1(n5493), .A2(n5492), .ZN(n5531) );
  INV_X1 U7223 ( .A(n5493), .ZN(n5494) );
  NAND2_X1 U7224 ( .A1(n5494), .A2(SI_25_), .ZN(n5495) );
  NAND2_X1 U7225 ( .A1(n5531), .A2(n5495), .ZN(n5527) );
  NAND2_X1 U7226 ( .A1(n8901), .A2(n5787), .ZN(n5497) );
  NAND2_X1 U7227 ( .A1(n6562), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5496) );
  INV_X1 U7228 ( .A(n5499), .ZN(n5498) );
  INV_X1 U7229 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U7230 ( .A1(n5499), .A2(n8310), .ZN(n5500) );
  NAND2_X1 U7231 ( .A1(n5517), .A2(n5500), .ZN(n8547) );
  INV_X1 U7232 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U7233 ( .A1(n6524), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U7234 ( .A1(n6520), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5501) );
  OAI211_X1 U7235 ( .C1(n8546), .C2(n6527), .A(n5502), .B(n5501), .ZN(n5503)
         );
  INV_X1 U7236 ( .A(n5503), .ZN(n5504) );
  INV_X1 U7237 ( .A(n8571), .ZN(n8352) );
  OR2_X1 U7238 ( .A1(n8769), .A2(n8352), .ZN(n6551) );
  NAND2_X1 U7239 ( .A1(n8550), .A2(n6551), .ZN(n5826) );
  INV_X1 U7240 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8899) );
  INV_X1 U7241 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5507) );
  MUX2_X1 U7242 ( .A(n8899), .B(n5507), .S(n4277), .Z(n5509) );
  INV_X1 U7243 ( .A(SI_26_), .ZN(n5508) );
  NAND2_X1 U7244 ( .A1(n5509), .A2(n5508), .ZN(n5530) );
  INV_X1 U7245 ( .A(n5509), .ZN(n5510) );
  NAND2_X1 U7246 ( .A1(n5510), .A2(SI_26_), .ZN(n5526) );
  AND2_X1 U7247 ( .A1(n5530), .A2(n5526), .ZN(n5511) );
  NAND2_X1 U7248 ( .A1(n8898), .A2(n5787), .ZN(n5514) );
  NAND2_X1 U7249 ( .A1(n6562), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5513) );
  INV_X1 U7250 ( .A(n5517), .ZN(n5515) );
  NAND2_X2 U7251 ( .A1(n5515), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5559) );
  INV_X1 U7252 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7253 ( .A1(n5517), .A2(n5516), .ZN(n5518) );
  NAND2_X1 U7254 ( .A1(n5559), .A2(n5518), .ZN(n5837) );
  INV_X1 U7255 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7256 ( .A1(n6524), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7257 ( .A1(n6520), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5519) );
  OAI211_X1 U7258 ( .C1(n5521), .C2(n6527), .A(n5520), .B(n5519), .ZN(n5522)
         );
  INV_X1 U7259 ( .A(n5522), .ZN(n5523) );
  INV_X1 U7260 ( .A(n6729), .ZN(n5525) );
  INV_X1 U7261 ( .A(n5526), .ZN(n5533) );
  AND2_X1 U7262 ( .A1(n5531), .A2(n5530), .ZN(n5532) );
  INV_X1 U7263 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8896) );
  INV_X1 U7264 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5536) );
  MUX2_X1 U7265 ( .A(n8896), .B(n5536), .S(n4277), .Z(n5538) );
  INV_X1 U7266 ( .A(SI_27_), .ZN(n5537) );
  NAND2_X1 U7267 ( .A1(n5538), .A2(n5537), .ZN(n6508) );
  INV_X1 U7268 ( .A(n5538), .ZN(n5539) );
  NAND2_X1 U7269 ( .A1(n5539), .A2(SI_27_), .ZN(n5540) );
  NAND2_X1 U7270 ( .A1(n8895), .A2(n5787), .ZN(n5542) );
  NAND2_X1 U7271 ( .A1(n6562), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7272 ( .A1(n8533), .A2(n5810), .ZN(n5547) );
  INV_X1 U7273 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10162) );
  NAND2_X1 U7274 ( .A1(n6524), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7275 ( .A1(n5561), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5543) );
  OAI211_X1 U7276 ( .C1(n6526), .C2(n10162), .A(n5544), .B(n5543), .ZN(n5545)
         );
  INV_X1 U7277 ( .A(n5545), .ZN(n5546) );
  XNOR2_X1 U7278 ( .A(n5548), .B(n4867), .ZN(n5570) );
  INV_X1 U7279 ( .A(n7662), .ZN(n6607) );
  XNOR2_X2 U7280 ( .A(n5556), .B(n5555), .ZN(n7684) );
  NAND2_X1 U7281 ( .A1(n6607), .A2(n6628), .ZN(n6581) );
  NAND2_X2 U7282 ( .A1(n6757), .A2(n6581), .ZN(n10021) );
  INV_X1 U7283 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8249) );
  INV_X1 U7284 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5557) );
  OAI21_X1 U7285 ( .B1(n5559), .B2(n8249), .A(n5557), .ZN(n5560) );
  NAND2_X1 U7286 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5558) );
  INV_X1 U7287 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7288 ( .A1(n6524), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7289 ( .A1(n5561), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5562) );
  OAI211_X1 U7290 ( .C1(n5564), .C2(n6526), .A(n5563), .B(n5562), .ZN(n5565)
         );
  AOI21_X2 U7291 ( .B1(n8525), .B2(n5810), .A(n5565), .ZN(n8416) );
  NAND2_X1 U7292 ( .A1(n6755), .A2(n6628), .ZN(n5845) );
  NAND2_X1 U7293 ( .A1(n5567), .A2(n5566), .ZN(n5853) );
  NAND2_X1 U7294 ( .A1(n5853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5568) );
  XNOR2_X1 U7295 ( .A(n5568), .B(P2_IR_REG_28__SCAN_IN), .ZN(n5890) );
  INV_X1 U7296 ( .A(n5845), .ZN(n5916) );
  OAI22_X1 U7297 ( .A1(n8416), .A2(n8336), .B1(n8250), .B2(n8563), .ZN(n5569)
         );
  NAND2_X1 U7298 ( .A1(n6639), .A2(n6638), .ZN(n6588) );
  NAND2_X1 U7299 ( .A1(n6588), .A2(n5650), .ZN(n6991) );
  NAND2_X1 U7300 ( .A1(n5649), .A2(n6987), .ZN(n5571) );
  NAND2_X1 U7301 ( .A1(n6991), .A2(n5571), .ZN(n7006) );
  NAND2_X1 U7302 ( .A1(n7006), .A2(n7005), .ZN(n7004) );
  OR2_X1 U7303 ( .A1(n5657), .A2(n7012), .ZN(n7228) );
  OR2_X1 U7304 ( .A1(n8434), .A2(n5663), .ZN(n7229) );
  NAND3_X1 U7305 ( .A1(n7004), .A2(n7228), .A3(n7229), .ZN(n5572) );
  NAND2_X1 U7306 ( .A1(n4634), .A2(n10063), .ZN(n5573) );
  NAND2_X1 U7307 ( .A1(n7231), .A2(n5573), .ZN(n7051) );
  NAND2_X1 U7308 ( .A1(n6625), .A2(n6618), .ZN(n7056) );
  NAND2_X1 U7309 ( .A1(n7051), .A2(n7056), .ZN(n7052) );
  OR2_X1 U7310 ( .A1(n8432), .A2(n4635), .ZN(n7357) );
  OR2_X1 U7311 ( .A1(n8431), .A2(n7382), .ZN(n7359) );
  NAND2_X1 U7312 ( .A1(n7052), .A2(n4985), .ZN(n5578) );
  INV_X1 U7313 ( .A(n7359), .ZN(n5575) );
  OAI21_X1 U7314 ( .B1(n5575), .B2(n7374), .A(n5574), .ZN(n5576) );
  INV_X1 U7315 ( .A(n7624), .ZN(n8430) );
  OR2_X1 U7316 ( .A1(n7466), .A2(n8430), .ZN(n5579) );
  INV_X1 U7317 ( .A(n7691), .ZN(n8429) );
  NAND2_X1 U7318 ( .A1(n8860), .A2(n8429), .ZN(n5581) );
  INV_X1 U7319 ( .A(n7767), .ZN(n8428) );
  OR2_X1 U7320 ( .A1(n8855), .A2(n8428), .ZN(n7700) );
  AND2_X1 U7321 ( .A1(n7702), .A2(n7700), .ZN(n5583) );
  INV_X1 U7322 ( .A(n7847), .ZN(n8427) );
  NAND2_X1 U7323 ( .A1(n6673), .A2(n6675), .ZN(n7727) );
  NAND2_X1 U7324 ( .A1(n7725), .A2(n7727), .ZN(n5585) );
  INV_X1 U7325 ( .A(n7908), .ZN(n8426) );
  NAND2_X1 U7326 ( .A1(n8844), .A2(n8426), .ZN(n5584) );
  INV_X1 U7327 ( .A(n7919), .ZN(n8425) );
  INV_X1 U7328 ( .A(n8273), .ZN(n8424) );
  NAND2_X1 U7329 ( .A1(n8833), .A2(n8424), .ZN(n5586) );
  INV_X1 U7330 ( .A(n8404), .ZN(n8423) );
  OR2_X1 U7331 ( .A1(n8828), .A2(n8423), .ZN(n8718) );
  INV_X1 U7332 ( .A(n8324), .ZN(n8422) );
  OR2_X1 U7333 ( .A1(n8824), .A2(n8422), .ZN(n5589) );
  AND2_X1 U7334 ( .A1(n8718), .A2(n5589), .ZN(n5588) );
  INV_X1 U7335 ( .A(n5589), .ZN(n5590) );
  OR2_X1 U7336 ( .A1(n5590), .A2(n8721), .ZN(n5591) );
  NAND2_X1 U7337 ( .A1(n6696), .A2(n6695), .ZN(n8696) );
  NAND2_X1 U7338 ( .A1(n8709), .A2(n8421), .ZN(n5592) );
  INV_X1 U7339 ( .A(n8686), .ZN(n5593) );
  INV_X1 U7340 ( .A(n8382), .ZN(n8664) );
  OR2_X1 U7341 ( .A1(n8811), .A2(n8664), .ZN(n5594) );
  NAND2_X1 U7342 ( .A1(n8805), .A2(n8420), .ZN(n5596) );
  NOR2_X1 U7343 ( .A1(n8805), .A2(n8420), .ZN(n5595) );
  INV_X1 U7344 ( .A(n8802), .ZN(n8638) );
  INV_X1 U7345 ( .A(n8776), .ZN(n8562) );
  INV_X1 U7346 ( .A(n8762), .ZN(n5839) );
  NAND2_X1 U7347 ( .A1(n5839), .A2(n8250), .ZN(n5603) );
  XNOR2_X1 U7348 ( .A(n8500), .B(n8499), .ZN(n8532) );
  XNOR2_X1 U7349 ( .A(n6755), .B(n5834), .ZN(n8642) );
  NAND2_X1 U7350 ( .A1(n8642), .A2(n7558), .ZN(n8693) );
  NAND3_X1 U7351 ( .A1(n7833), .A2(n8646), .A3(n7662), .ZN(n8866) );
  INV_X1 U7352 ( .A(n8769), .ZN(n8545) );
  NAND2_X1 U7353 ( .A1(n6987), .A2(n10052), .ZN(n7011) );
  NOR2_X2 U7354 ( .A1(n7011), .A2(n7012), .ZN(n10034) );
  INV_X1 U7355 ( .A(n7466), .ZN(n7549) );
  NAND2_X1 U7356 ( .A1(n7377), .A2(n7549), .ZN(n7363) );
  INV_X1 U7357 ( .A(n8850), .ZN(n7774) );
  INV_X1 U7358 ( .A(n8833), .ZN(n7866) );
  INV_X1 U7359 ( .A(n8828), .ZN(n7899) );
  INV_X1 U7360 ( .A(n8805), .ZN(n8660) );
  NAND2_X1 U7361 ( .A1(n8677), .A2(n8660), .ZN(n8654) );
  INV_X1 U7362 ( .A(n8524), .ZN(n5607) );
  AOI21_X1 U7363 ( .B1(n6733), .B2(n4684), .A(n5607), .ZN(n8537) );
  INV_X1 U7365 ( .A(n6752), .ZN(n5608) );
  AOI22_X1 U7366 ( .A1(n8537), .A2(n8861), .B1(n8840), .B2(n6733), .ZN(n5609)
         );
  NOR4_X1 U7367 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5613) );
  NOR4_X1 U7368 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5612) );
  NOR4_X1 U7369 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5611) );
  NOR4_X1 U7370 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n5610) );
  NAND4_X1 U7371 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n5635)
         );
  NOR2_X1 U7372 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .ZN(
        n10148) );
  NOR4_X1 U7373 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n5616) );
  NOR4_X1 U7374 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5615) );
  NOR4_X1 U7375 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5614) );
  NAND4_X1 U7376 ( .A1(n10148), .A2(n5616), .A3(n5615), .A4(n5614), .ZN(n5634)
         );
  INV_X1 U7377 ( .A(n5618), .ZN(n5619) );
  NAND2_X1 U7378 ( .A1(n5623), .A2(n5622), .ZN(n5624) );
  NAND2_X1 U7379 ( .A1(n5636), .A2(n5626), .ZN(n5627) );
  INV_X1 U7380 ( .A(P2_B_REG_SCAN_IN), .ZN(n7943) );
  XNOR2_X1 U7381 ( .A(n7889), .B(n7943), .ZN(n5630) );
  NAND2_X1 U7382 ( .A1(n5631), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5632) );
  OAI21_X1 U7383 ( .B1(n5635), .B2(n5634), .A(n10042), .ZN(n5792) );
  INV_X1 U7384 ( .A(n5638), .ZN(n8902) );
  XNOR2_X1 U7385 ( .A(n5626), .B(n5636), .ZN(n5846) );
  OR2_X1 U7386 ( .A1(n5845), .A2(n6752), .ZN(n5816) );
  NAND2_X1 U7387 ( .A1(n8861), .A2(n8646), .ZN(n5814) );
  NAND3_X1 U7388 ( .A1(n5792), .A2(n5831), .A3(n5814), .ZN(n5639) );
  INV_X1 U7389 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10048) );
  NOR2_X1 U7390 ( .A1(n5638), .A2(n5637), .ZN(n10049) );
  AOI21_X1 U7391 ( .B1(n10042), .B2(n10048), .A(n10049), .ZN(n5793) );
  INV_X1 U7392 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10140) );
  NAND2_X1 U7393 ( .A1(n5642), .A2(n5641), .ZN(P2_U3547) );
  INV_X1 U7394 ( .A(n5794), .ZN(n5832) );
  NAND2_X1 U7395 ( .A1(n5644), .A2(n10076), .ZN(n5646) );
  NAND2_X1 U7396 ( .A1(n5646), .A2(n5645), .ZN(P2_U3515) );
  NAND2_X2 U7397 ( .A1(n5647), .A2(n5834), .ZN(n5670) );
  XNOR2_X1 U7398 ( .A(n8776), .B(n5790), .ZN(n8346) );
  OR2_X1 U7399 ( .A1(n8309), .A2(n7100), .ZN(n8347) );
  INV_X2 U7400 ( .A(n5651), .ZN(n5671) );
  INV_X1 U7401 ( .A(n7088), .ZN(n5654) );
  INV_X1 U7402 ( .A(n5650), .ZN(n6994) );
  NAND2_X1 U7403 ( .A1(n5656), .A2(n7088), .ZN(n5658) );
  NAND2_X1 U7404 ( .A1(n5657), .A2(n5671), .ZN(n5660) );
  NAND2_X1 U7405 ( .A1(n5659), .A2(n5660), .ZN(n7090) );
  INV_X1 U7406 ( .A(n5659), .ZN(n5662) );
  INV_X1 U7407 ( .A(n5660), .ZN(n5661) );
  NAND2_X1 U7408 ( .A1(n5662), .A2(n5661), .ZN(n7091) );
  XNOR2_X1 U7409 ( .A(n5663), .B(n5670), .ZN(n5664) );
  AND2_X1 U7410 ( .A1(n8434), .A2(n5671), .ZN(n5665) );
  NAND2_X1 U7411 ( .A1(n5664), .A2(n5665), .ZN(n5669) );
  INV_X1 U7412 ( .A(n5664), .ZN(n5667) );
  INV_X1 U7413 ( .A(n5665), .ZN(n5666) );
  NAND2_X1 U7414 ( .A1(n5667), .A2(n5666), .ZN(n5668) );
  AND2_X1 U7415 ( .A1(n5669), .A2(n5668), .ZN(n6768) );
  AND2_X2 U7416 ( .A1(n6767), .A2(n5669), .ZN(n7247) );
  XNOR2_X1 U7417 ( .A(n5670), .B(n4278), .ZN(n5672) );
  NAND2_X1 U7418 ( .A1(n8433), .A2(n5671), .ZN(n5673) );
  XNOR2_X1 U7419 ( .A(n5672), .B(n5673), .ZN(n7246) );
  INV_X1 U7420 ( .A(n5672), .ZN(n5674) );
  NAND2_X1 U7421 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  INV_X1 U7422 ( .A(n7396), .ZN(n5680) );
  XNOR2_X1 U7423 ( .A(n5777), .B(n7393), .ZN(n5677) );
  NAND2_X1 U7424 ( .A1(n8432), .A2(n5671), .ZN(n5676) );
  OR2_X1 U7425 ( .A1(n5677), .A2(n5676), .ZN(n5681) );
  NAND2_X1 U7426 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  NAND2_X1 U7427 ( .A1(n5681), .A2(n5678), .ZN(n7397) );
  AND2_X2 U7428 ( .A1(n7394), .A2(n5681), .ZN(n7347) );
  XNOR2_X1 U7429 ( .A(n7382), .B(n5777), .ZN(n5684) );
  NAND2_X1 U7430 ( .A1(n8431), .A2(n5671), .ZN(n5682) );
  XNOR2_X1 U7431 ( .A(n5684), .B(n5682), .ZN(n7346) );
  INV_X1 U7432 ( .A(n5682), .ZN(n5683) );
  OR2_X1 U7433 ( .A1(n5684), .A2(n5683), .ZN(n5685) );
  XNOR2_X1 U7434 ( .A(n7466), .B(n5777), .ZN(n5686) );
  NOR2_X1 U7435 ( .A1(n7624), .A2(n7100), .ZN(n5687) );
  NAND2_X1 U7436 ( .A1(n5686), .A2(n5687), .ZN(n5691) );
  INV_X1 U7437 ( .A(n5686), .ZN(n5689) );
  INV_X1 U7438 ( .A(n5687), .ZN(n5688) );
  NAND2_X1 U7439 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  AND2_X1 U7440 ( .A1(n5691), .A2(n5690), .ZN(n7460) );
  XNOR2_X1 U7441 ( .A(n8860), .B(n5777), .ZN(n5692) );
  NOR2_X1 U7442 ( .A1(n7691), .A2(n7100), .ZN(n5693) );
  NAND2_X1 U7443 ( .A1(n5692), .A2(n5693), .ZN(n5697) );
  INV_X1 U7444 ( .A(n5692), .ZN(n5695) );
  INV_X1 U7445 ( .A(n5693), .ZN(n5694) );
  NAND2_X1 U7446 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  AND2_X1 U7447 ( .A1(n5697), .A2(n5696), .ZN(n7582) );
  XNOR2_X1 U7448 ( .A(n8855), .B(n5777), .ZN(n5699) );
  NOR2_X1 U7449 ( .A1(n7767), .A2(n7100), .ZN(n5700) );
  XNOR2_X1 U7450 ( .A(n5699), .B(n5700), .ZN(n7689) );
  INV_X1 U7451 ( .A(n7689), .ZN(n5698) );
  INV_X1 U7452 ( .A(n5699), .ZN(n5702) );
  INV_X1 U7453 ( .A(n5700), .ZN(n5701) );
  NAND2_X1 U7454 ( .A1(n5702), .A2(n5701), .ZN(n5703) );
  XNOR2_X1 U7455 ( .A(n8850), .B(n5777), .ZN(n5704) );
  NOR2_X1 U7456 ( .A1(n7847), .A2(n7100), .ZN(n5705) );
  NAND2_X1 U7457 ( .A1(n5704), .A2(n5705), .ZN(n5709) );
  INV_X1 U7458 ( .A(n5704), .ZN(n5707) );
  INV_X1 U7459 ( .A(n5705), .ZN(n5706) );
  NAND2_X1 U7460 ( .A1(n5707), .A2(n5706), .ZN(n5708) );
  AND2_X1 U7461 ( .A1(n5709), .A2(n5708), .ZN(n7765) );
  NAND2_X1 U7462 ( .A1(n7764), .A2(n5709), .ZN(n7845) );
  XNOR2_X1 U7463 ( .A(n8844), .B(n5790), .ZN(n5710) );
  NOR2_X1 U7464 ( .A1(n7908), .A2(n7100), .ZN(n5711) );
  XNOR2_X1 U7465 ( .A(n5710), .B(n5711), .ZN(n7844) );
  INV_X1 U7466 ( .A(n5710), .ZN(n5712) );
  NAND2_X1 U7467 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  XNOR2_X1 U7468 ( .A(n8839), .B(n5790), .ZN(n5714) );
  OR2_X1 U7469 ( .A1(n7919), .A2(n7100), .ZN(n5715) );
  NAND2_X1 U7470 ( .A1(n5714), .A2(n5715), .ZN(n7904) );
  INV_X1 U7471 ( .A(n5714), .ZN(n5717) );
  INV_X1 U7472 ( .A(n5715), .ZN(n5716) );
  NAND2_X1 U7473 ( .A1(n5717), .A2(n5716), .ZN(n7914) );
  XNOR2_X1 U7474 ( .A(n8833), .B(n5790), .ZN(n5722) );
  INV_X1 U7475 ( .A(n5722), .ZN(n5718) );
  NOR2_X1 U7476 ( .A1(n8273), .A2(n7100), .ZN(n5721) );
  NAND2_X1 U7477 ( .A1(n5718), .A2(n5721), .ZN(n5720) );
  AND2_X1 U7478 ( .A1(n7914), .A2(n5720), .ZN(n5719) );
  NAND2_X1 U7479 ( .A1(n7915), .A2(n5719), .ZN(n8330) );
  INV_X1 U7480 ( .A(n5720), .ZN(n5723) );
  XNOR2_X1 U7481 ( .A(n5722), .B(n5721), .ZN(n7916) );
  OR2_X1 U7482 ( .A1(n5723), .A2(n7916), .ZN(n8268) );
  XNOR2_X1 U7483 ( .A(n8815), .B(n5777), .ZN(n8321) );
  NAND2_X1 U7484 ( .A1(n8421), .A2(n5652), .ZN(n8320) );
  XNOR2_X1 U7485 ( .A(n8824), .B(n5777), .ZN(n5731) );
  NOR2_X1 U7486 ( .A1(n8324), .A2(n7100), .ZN(n8319) );
  XNOR2_X1 U7487 ( .A(n8828), .B(n5777), .ZN(n5729) );
  INV_X1 U7488 ( .A(n5729), .ZN(n5725) );
  NOR2_X1 U7489 ( .A1(n8404), .A2(n7100), .ZN(n5728) );
  INV_X1 U7490 ( .A(n5728), .ZN(n5724) );
  NAND2_X1 U7491 ( .A1(n5725), .A2(n5724), .ZN(n8315) );
  OAI21_X1 U7492 ( .B1(n5731), .B2(n8319), .A(n8315), .ZN(n5726) );
  AOI21_X1 U7493 ( .B1(n8321), .B2(n8320), .A(n5726), .ZN(n5730) );
  AND2_X1 U7494 ( .A1(n8268), .A2(n5730), .ZN(n8329) );
  XNOR2_X1 U7495 ( .A(n8811), .B(n5777), .ZN(n5741) );
  NAND2_X1 U7496 ( .A1(n8664), .A2(n5671), .ZN(n5739) );
  XNOR2_X1 U7497 ( .A(n5741), .B(n5739), .ZN(n8333) );
  AND2_X1 U7498 ( .A1(n8329), .A2(n8333), .ZN(n5727) );
  INV_X1 U7499 ( .A(n8333), .ZN(n5738) );
  XNOR2_X1 U7500 ( .A(n5729), .B(n5728), .ZN(n8271) );
  AND2_X1 U7501 ( .A1(n5730), .A2(n8271), .ZN(n5737) );
  INV_X1 U7502 ( .A(n8321), .ZN(n5734) );
  INV_X1 U7503 ( .A(n5731), .ZN(n8317) );
  INV_X1 U7504 ( .A(n8319), .ZN(n8402) );
  OAI21_X1 U7505 ( .B1(n8317), .B2(n8402), .A(n8320), .ZN(n5733) );
  NOR2_X1 U7506 ( .A1(n8402), .A2(n8320), .ZN(n5732) );
  AOI22_X1 U7507 ( .A1(n5734), .A2(n5733), .B1(n5732), .B2(n5731), .ZN(n5735)
         );
  INV_X1 U7508 ( .A(n5735), .ZN(n5736) );
  NOR2_X1 U7509 ( .A1(n5737), .A2(n5736), .ZN(n8331) );
  INV_X1 U7510 ( .A(n5739), .ZN(n5740) );
  NAND2_X1 U7511 ( .A1(n5741), .A2(n5740), .ZN(n8376) );
  XNOR2_X1 U7512 ( .A(n8805), .B(n5777), .ZN(n5745) );
  NAND2_X1 U7513 ( .A1(n8420), .A2(n5652), .ZN(n5744) );
  INV_X1 U7514 ( .A(n5744), .ZN(n5742) );
  NAND2_X1 U7515 ( .A1(n5745), .A2(n5742), .ZN(n5743) );
  AND2_X1 U7516 ( .A1(n8376), .A2(n5743), .ZN(n5747) );
  INV_X1 U7517 ( .A(n5743), .ZN(n5746) );
  XNOR2_X1 U7518 ( .A(n5745), .B(n5744), .ZN(n8378) );
  XNOR2_X1 U7519 ( .A(n8802), .B(n5790), .ZN(n5748) );
  NAND2_X1 U7520 ( .A1(n8666), .A2(n5671), .ZN(n5749) );
  NAND2_X1 U7521 ( .A1(n5748), .A2(n5749), .ZN(n5753) );
  INV_X1 U7522 ( .A(n5748), .ZN(n5751) );
  INV_X1 U7523 ( .A(n5749), .ZN(n5750) );
  NAND2_X1 U7524 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  NAND2_X1 U7525 ( .A1(n5753), .A2(n5752), .ZN(n8289) );
  OR2_X2 U7526 ( .A1(n8290), .A2(n8289), .ZN(n8287) );
  XNOR2_X1 U7527 ( .A(n8796), .B(n5790), .ZN(n5754) );
  NAND2_X1 U7528 ( .A1(n8419), .A2(n5671), .ZN(n5755) );
  XNOR2_X1 U7529 ( .A(n5754), .B(n5755), .ZN(n8357) );
  INV_X1 U7530 ( .A(n5754), .ZN(n5757) );
  INV_X1 U7531 ( .A(n5755), .ZN(n5756) );
  NAND2_X1 U7532 ( .A1(n5757), .A2(n5756), .ZN(n5758) );
  XNOR2_X1 U7533 ( .A(n8617), .B(n5777), .ZN(n5760) );
  NOR2_X1 U7534 ( .A1(n8371), .A2(n7100), .ZN(n5761) );
  XNOR2_X1 U7535 ( .A(n5760), .B(n5761), .ZN(n8297) );
  XNOR2_X1 U7536 ( .A(n8786), .B(n5790), .ZN(n8367) );
  NAND2_X1 U7537 ( .A1(n5600), .A2(n5652), .ZN(n8366) );
  NAND2_X1 U7538 ( .A1(n8367), .A2(n8366), .ZN(n5759) );
  NAND2_X1 U7539 ( .A1(n8365), .A2(n5759), .ZN(n5768) );
  INV_X1 U7540 ( .A(n5760), .ZN(n5763) );
  NAND2_X1 U7541 ( .A1(n5763), .A2(n5761), .ZN(n8363) );
  NAND2_X1 U7542 ( .A1(n8363), .A2(n8366), .ZN(n5766) );
  INV_X1 U7543 ( .A(n8367), .ZN(n5765) );
  INV_X1 U7544 ( .A(n5761), .ZN(n5762) );
  NOR2_X1 U7545 ( .A1(n8281), .A2(n5762), .ZN(n5764) );
  AOI22_X1 U7546 ( .A1(n5766), .A2(n5765), .B1(n5764), .B2(n5763), .ZN(n5767)
         );
  XNOR2_X1 U7547 ( .A(n8781), .B(n5777), .ZN(n5770) );
  NAND2_X1 U7548 ( .A1(n8598), .A2(n5671), .ZN(n8344) );
  AOI21_X1 U7549 ( .B1(n8346), .B2(n8309), .A(n8344), .ZN(n5769) );
  XNOR2_X1 U7550 ( .A(n8769), .B(n5777), .ZN(n8305) );
  AND2_X2 U7551 ( .A1(n8308), .A2(n8305), .ZN(n5772) );
  NOR2_X1 U7552 ( .A1(n8352), .A2(n7100), .ZN(n8306) );
  XNOR2_X1 U7553 ( .A(n8762), .B(n5777), .ZN(n5774) );
  NOR2_X1 U7554 ( .A1(n8250), .A2(n7100), .ZN(n5773) );
  NAND2_X1 U7555 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  OAI21_X1 U7556 ( .B1(n5774), .B2(n5773), .A(n5775), .ZN(n8396) );
  INV_X1 U7557 ( .A(n5775), .ZN(n5776) );
  XNOR2_X1 U7558 ( .A(n6733), .B(n5777), .ZN(n5779) );
  NOR2_X1 U7559 ( .A1(n8501), .A2(n7100), .ZN(n5778) );
  NAND2_X1 U7560 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  OAI21_X1 U7561 ( .B1(n5779), .B2(n5778), .A(n5780), .ZN(n8246) );
  INV_X1 U7562 ( .A(n5780), .ZN(n5781) );
  NAND2_X1 U7563 ( .A1(n6510), .A2(n6508), .ZN(n5786) );
  INV_X1 U7564 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5785) );
  INV_X1 U7565 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5784) );
  MUX2_X1 U7566 ( .A(n5785), .B(n5784), .S(n4277), .Z(n6507) );
  XNOR2_X1 U7567 ( .A(n6507), .B(SI_28_), .ZN(n6512) );
  NAND2_X1 U7568 ( .A1(n8890), .A2(n5787), .ZN(n5789) );
  NAND2_X1 U7569 ( .A1(n6562), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5788) );
  OR2_X1 U7570 ( .A1(n8416), .A2(n7100), .ZN(n5791) );
  XNOR2_X1 U7571 ( .A(n5791), .B(n5790), .ZN(n5804) );
  AND2_X1 U7572 ( .A1(n5793), .A2(n5792), .ZN(n5830) );
  AND2_X1 U7573 ( .A1(n5794), .A2(n5830), .ZN(n5813) );
  AND2_X1 U7574 ( .A1(n10033), .A2(n6607), .ZN(n5836) );
  NAND2_X1 U7575 ( .A1(n5812), .A2(n5836), .ZN(n5796) );
  INV_X1 U7576 ( .A(n5814), .ZN(n5795) );
  NAND3_X1 U7577 ( .A1(n8755), .A2(n5804), .A3(n8300), .ZN(n5797) );
  OAI21_X1 U7578 ( .B1(n8755), .B2(n5804), .A(n5797), .ZN(n5798) );
  NAND2_X1 U7579 ( .A1(n5806), .A2(n5798), .ZN(n5802) );
  NAND2_X1 U7580 ( .A1(n8755), .A2(n8411), .ZN(n5800) );
  NOR2_X1 U7581 ( .A1(n10032), .A2(n5916), .ZN(n5799) );
  NAND2_X1 U7582 ( .A1(n5800), .A2(n8413), .ZN(n5801) );
  NAND2_X1 U7583 ( .A1(n5802), .A2(n5801), .ZN(n5825) );
  NOR3_X1 U7584 ( .A1(n4680), .A2(n5804), .A3(n8411), .ZN(n5803) );
  AOI21_X1 U7585 ( .B1(n5804), .B2(n4680), .A(n5803), .ZN(n5805) );
  INV_X1 U7586 ( .A(n8508), .ZN(n5811) );
  INV_X1 U7587 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U7588 ( .A1(n6520), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U7589 ( .A1(n6524), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5807) );
  OAI211_X1 U7590 ( .C1(n8507), .C2(n6527), .A(n5808), .B(n5807), .ZN(n5809)
         );
  AOI21_X1 U7591 ( .B1(n5811), .B2(n5810), .A(n5809), .ZN(n6565) );
  INV_X1 U7592 ( .A(n6565), .ZN(n8415) );
  AOI22_X1 U7593 ( .A1(n8417), .A2(n8663), .B1(n8415), .B2(n8665), .ZN(n8519)
         );
  NAND2_X1 U7594 ( .A1(n5812), .A2(n6752), .ZN(n8392) );
  INV_X1 U7595 ( .A(n5813), .ZN(n5815) );
  NAND2_X1 U7596 ( .A1(n5815), .A2(n5814), .ZN(n5818) );
  AND2_X1 U7597 ( .A1(n5847), .A2(n5816), .ZN(n5817) );
  NAND2_X1 U7598 ( .A1(n5818), .A2(n5817), .ZN(n6985) );
  INV_X1 U7599 ( .A(n5846), .ZN(n5819) );
  OR2_X1 U7600 ( .A1(n6985), .A2(n5819), .ZN(n5820) );
  AOI22_X1 U7601 ( .A1(n8525), .A2(n8389), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5821) );
  OAI21_X1 U7602 ( .B1(n8519), .B2(n8392), .A(n5821), .ZN(n5822) );
  OAI21_X1 U7603 ( .B1(n5825), .B2(n5824), .A(n5823), .ZN(P2_U3222) );
  XNOR2_X1 U7604 ( .A(n5826), .B(n6587), .ZN(n5829) );
  OR2_X1 U7605 ( .A1(n8501), .A2(n8336), .ZN(n5828) );
  NAND2_X1 U7606 ( .A1(n8571), .A2(n8663), .ZN(n5827) );
  NAND2_X1 U7607 ( .A1(n5828), .A2(n5827), .ZN(n8388) );
  NAND3_X1 U7608 ( .A1(n5832), .A2(n5831), .A3(n5830), .ZN(n7178) );
  XOR2_X1 U7609 ( .A(n5833), .B(n6587), .Z(n8760) );
  OR2_X1 U7610 ( .A1(n5834), .A2(n7558), .ZN(n7619) );
  NAND2_X1 U7611 ( .A1(n8693), .A2(n7619), .ZN(n10027) );
  AOI211_X1 U7612 ( .C1(n8762), .C2(n8542), .A(n8816), .B(n5835), .ZN(n8761)
         );
  NOR2_X1 U7613 ( .A1(n10031), .A2(n8646), .ZN(n8689) );
  INV_X1 U7614 ( .A(n5837), .ZN(n8390) );
  INV_X1 U7615 ( .A(n10041), .ZN(n8678) );
  AOI22_X1 U7616 ( .A1(n8390), .A2(n8678), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n10031), .ZN(n5838) );
  OAI21_X1 U7617 ( .B1(n5839), .B2(n8681), .A(n5838), .ZN(n5840) );
  AOI21_X1 U7618 ( .B1(n8761), .B2(n8689), .A(n5840), .ZN(n5841) );
  INV_X1 U7619 ( .A(n5842), .ZN(n5843) );
  INV_X1 U7620 ( .A(n5847), .ZN(n5844) );
  NAND2_X1 U7621 ( .A1(n10044), .A2(n5845), .ZN(n5850) );
  NAND2_X1 U7622 ( .A1(n5890), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8893) );
  OR2_X1 U7623 ( .A1(n5846), .A2(P2_U3152), .ZN(n6754) );
  OAI21_X1 U7624 ( .B1(n5847), .B2(n8893), .A(n6754), .ZN(n5848) );
  INV_X1 U7625 ( .A(n5848), .ZN(n5849) );
  NAND2_X1 U7626 ( .A1(n5850), .A2(n5849), .ZN(n5852) );
  NAND2_X1 U7627 ( .A1(n5852), .A2(n5851), .ZN(n5889) );
  INV_X1 U7628 ( .A(n5889), .ZN(n5855) );
  NAND2_X1 U7629 ( .A1(n5854), .A2(n5853), .ZN(n8897) );
  INV_X1 U7630 ( .A(n8486), .ZN(n7486) );
  INV_X1 U7631 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n5886) );
  XNOR2_X1 U7632 ( .A(n8473), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8463) );
  INV_X1 U7633 ( .A(n8460), .ZN(n5883) );
  XNOR2_X1 U7634 ( .A(n8460), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8450) );
  INV_X1 U7635 ( .A(n5902), .ZN(n7934) );
  OR2_X1 U7636 ( .A1(n7870), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7637 ( .A1(n7870), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5856) );
  AND2_X1 U7638 ( .A1(n5878), .A2(n5856), .ZN(n7877) );
  INV_X1 U7639 ( .A(n7826), .ZN(n6863) );
  INV_X1 U7640 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7641 ( .A1(n6863), .A2(n5875), .ZN(n5877) );
  MUX2_X1 U7642 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5857), .S(n7186), .Z(n5862)
         );
  MUX2_X1 U7643 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n5858), .S(n7259), .Z(n5860)
         );
  AND2_X1 U7644 ( .A1(n4407), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7645 ( .A1(n5860), .A2(n5859), .ZN(n7261) );
  NAND2_X1 U7646 ( .A1(n7259), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7187) );
  NAND2_X1 U7647 ( .A1(n7261), .A2(n7187), .ZN(n5861) );
  NAND2_X1 U7648 ( .A1(n5862), .A2(n5861), .ZN(n7190) );
  NAND2_X1 U7649 ( .A1(n7186), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7650 ( .A1(n7190), .A2(n5863), .ZN(n7285) );
  INV_X1 U7651 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5864) );
  MUX2_X1 U7652 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n5864), .S(n7295), .Z(n7286)
         );
  NAND2_X1 U7653 ( .A1(n7285), .A2(n7286), .ZN(n7284) );
  NAND2_X1 U7654 ( .A1(n7295), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7271) );
  NAND2_X1 U7655 ( .A1(n7284), .A2(n7271), .ZN(n5867) );
  MUX2_X1 U7656 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n5865), .S(n7282), .Z(n5866)
         );
  NAND2_X1 U7657 ( .A1(n5867), .A2(n5866), .ZN(n7326) );
  NAND2_X1 U7658 ( .A1(n7282), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7325) );
  NAND2_X1 U7659 ( .A1(n7326), .A2(n7325), .ZN(n5870) );
  MUX2_X1 U7660 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n5868), .S(n7336), .Z(n5869)
         );
  NAND2_X1 U7661 ( .A1(n5870), .A2(n5869), .ZN(n7328) );
  NAND2_X1 U7662 ( .A1(n7336), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7299) );
  MUX2_X1 U7663 ( .A(n5127), .B(P2_REG1_REG_6__SCAN_IN), .S(n7310), .Z(n7298)
         );
  AOI21_X1 U7664 ( .B1(n7328), .B2(n7299), .A(n7298), .ZN(n7297) );
  AND2_X1 U7665 ( .A1(n7310), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5871) );
  NOR2_X1 U7666 ( .A1(n7297), .A2(n5871), .ZN(n7313) );
  XNOR2_X1 U7667 ( .A(n7322), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n7312) );
  INV_X1 U7668 ( .A(n7322), .ZN(n6830) );
  INV_X1 U7669 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5872) );
  OAI22_X1 U7670 ( .A1(n7313), .A2(n7312), .B1(n6830), .B2(n5872), .ZN(n7200)
         );
  XOR2_X1 U7671 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7201), .Z(n7199) );
  AOI22_X1 U7672 ( .A1(n7200), .A2(n7199), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n7201), .ZN(n7211) );
  XNOR2_X1 U7673 ( .A(n7213), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7210) );
  INV_X1 U7674 ( .A(n7213), .ZN(n6843) );
  OAI22_X1 U7675 ( .A1(n7211), .A2(n7210), .B1(n5873), .B2(n6843), .ZN(n7494)
         );
  XOR2_X1 U7676 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7495), .Z(n7493) );
  AOI22_X1 U7677 ( .A1(n7494), .A2(n7493), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7495), .ZN(n7636) );
  XNOR2_X1 U7678 ( .A(n5900), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n7635) );
  INV_X1 U7679 ( .A(n5900), .ZN(n7641) );
  OAI22_X1 U7680 ( .A1(n7636), .A2(n7635), .B1(n5874), .B2(n7641), .ZN(n7819)
         );
  OAI21_X1 U7681 ( .B1(n6863), .B2(n5875), .A(n5877), .ZN(n7818) );
  NOR2_X1 U7682 ( .A1(n7819), .A2(n7818), .ZN(n7817) );
  INV_X1 U7683 ( .A(n7817), .ZN(n5876) );
  NAND2_X1 U7684 ( .A1(n5877), .A2(n5876), .ZN(n7876) );
  NAND2_X1 U7685 ( .A1(n7877), .A2(n7876), .ZN(n7875) );
  NAND2_X1 U7686 ( .A1(n7875), .A2(n5878), .ZN(n7929) );
  XNOR2_X1 U7687 ( .A(n5902), .B(n5879), .ZN(n7928) );
  AOI21_X1 U7688 ( .B1(n7934), .B2(n5879), .A(n7931), .ZN(n5880) );
  NAND2_X1 U7689 ( .A1(n5904), .A2(n5880), .ZN(n5881) );
  INV_X1 U7690 ( .A(n5904), .ZN(n8445) );
  XNOR2_X1 U7691 ( .A(n8445), .B(n5880), .ZN(n8442) );
  NAND2_X1 U7692 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8442), .ZN(n8441) );
  NAND2_X1 U7693 ( .A1(n5881), .A2(n8441), .ZN(n8451) );
  NOR2_X1 U7694 ( .A1(n8450), .A2(n8451), .ZN(n8449) );
  AOI21_X1 U7695 ( .B1(n5883), .B2(n5882), .A(n8449), .ZN(n8464) );
  AND2_X1 U7696 ( .A1(n8463), .A2(n8464), .ZN(n8465) );
  INV_X1 U7697 ( .A(n8465), .ZN(n5885) );
  NAND2_X1 U7698 ( .A1(n5908), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7699 ( .A1(n5885), .A2(n5884), .ZN(n8475) );
  AOI22_X1 U7700 ( .A1(n8486), .A2(n5886), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n7486), .ZN(n8474) );
  NOR2_X1 U7701 ( .A1(n8475), .A2(n8474), .ZN(n8477) );
  AOI21_X1 U7702 ( .B1(n7486), .B2(n5886), .A(n8477), .ZN(n5887) );
  XNOR2_X1 U7703 ( .A(n5888), .B(n5887), .ZN(n5914) );
  INV_X1 U7704 ( .A(n5914), .ZN(n5912) );
  NAND2_X1 U7705 ( .A1(n5889), .A2(n8436), .ZN(n5911) );
  INV_X1 U7706 ( .A(n5890), .ZN(n5913) );
  NAND2_X1 U7707 ( .A1(n8460), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5891) );
  OAI21_X1 U7708 ( .B1(n8460), .B2(P2_REG2_REG_16__SCAN_IN), .A(n5891), .ZN(
        n8456) );
  XNOR2_X1 U7709 ( .A(n7870), .B(n5892), .ZN(n7873) );
  NAND2_X1 U7710 ( .A1(n7826), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5893) );
  OAI21_X1 U7711 ( .B1(n7826), .B2(P2_REG2_REG_12__SCAN_IN), .A(n5893), .ZN(
        n7821) );
  NAND2_X1 U7712 ( .A1(n4407), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7257) );
  XNOR2_X1 U7713 ( .A(n7295), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n7291) );
  NOR2_X1 U7714 ( .A1(n7292), .A2(n7291), .ZN(n7290) );
  XNOR2_X1 U7715 ( .A(n7282), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7278) );
  NOR2_X1 U7716 ( .A1(n7279), .A2(n7278), .ZN(n7277) );
  XNOR2_X1 U7717 ( .A(n7336), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n7332) );
  XNOR2_X1 U7718 ( .A(n7310), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7306) );
  XNOR2_X1 U7719 ( .A(n7322), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n7318) );
  MUX2_X1 U7720 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7628), .S(n7201), .Z(n5897)
         );
  INV_X1 U7721 ( .A(n5897), .ZN(n7197) );
  NOR2_X1 U7722 ( .A1(n7198), .A2(n7197), .ZN(n7196) );
  XNOR2_X1 U7723 ( .A(n7213), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n7208) );
  XNOR2_X1 U7724 ( .A(n7495), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7491) );
  MUX2_X1 U7725 ( .A(n7729), .B(P2_REG2_REG_11__SCAN_IN), .S(n5900), .Z(n5899)
         );
  INV_X1 U7726 ( .A(n5899), .ZN(n7638) );
  XNOR2_X1 U7727 ( .A(n5902), .B(n5901), .ZN(n7927) );
  NAND2_X1 U7728 ( .A1(n8445), .A2(n5905), .ZN(n5906) );
  NAND2_X1 U7729 ( .A1(n8438), .A2(n5906), .ZN(n8457) );
  NOR2_X1 U7730 ( .A1(n5909), .A2(n7486), .ZN(n5910) );
  INV_X1 U7731 ( .A(n8897), .ZN(n6751) );
  NAND2_X1 U7732 ( .A1(n5911), .A2(n6751), .ZN(n10012) );
  AOI22_X1 U7733 ( .A1(n5915), .A2(n10008), .B1(n10007), .B2(n5914), .ZN(n5921) );
  NAND2_X1 U7734 ( .A1(n10044), .A2(n5916), .ZN(n5917) );
  NAND2_X1 U7735 ( .A1(n5917), .A2(n5851), .ZN(n5918) );
  NAND2_X1 U7736 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8293) );
  OAI21_X1 U7737 ( .B1(n8480), .B2(n4774), .A(n8293), .ZN(n5919) );
  INV_X1 U7738 ( .A(n5919), .ZN(n5920) );
  NAND2_X1 U7739 ( .A1(n5928), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5929) );
  NAND2_X2 U7740 ( .A1(n5930), .A2(n4967), .ZN(n9258) );
  NAND2_X1 U7741 ( .A1(n7836), .A2(n8078), .ZN(n5932) );
  AND2_X2 U7742 ( .A1(n6002), .A2(n5061), .ZN(n6100) );
  NAND2_X1 U7743 ( .A1(n8087), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5931) );
  NAND2_X2 U7744 ( .A1(n5932), .A2(n5931), .ZN(n9433) );
  INV_X1 U7745 ( .A(n5937), .ZN(n5938) );
  NAND2_X1 U7746 ( .A1(n5938), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7747 ( .A1(n5942), .A2(n5940), .ZN(n5941) );
  INV_X1 U7748 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8954) );
  INV_X1 U7749 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9071) );
  INV_X1 U7750 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U7751 ( .A1(n6403), .A2(n8937), .ZN(n5956) );
  NAND2_X1 U7752 ( .A1(n6421), .A2(n5956), .ZN(n9441) );
  XNOR2_X2 U7753 ( .A(n5958), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5962) );
  OR2_X1 U7754 ( .A1(n9441), .A2(n8054), .ZN(n5968) );
  INV_X1 U7755 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7756 ( .A1(n4282), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5964) );
  AND2_X2 U7757 ( .A1(n5962), .A2(n9762), .ZN(n6036) );
  NAND2_X1 U7758 ( .A1(n8069), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5963) );
  OAI211_X1 U7759 ( .C1(n8085), .C2(n5965), .A(n5964), .B(n5963), .ZN(n5966)
         );
  INV_X1 U7760 ( .A(n5966), .ZN(n5967) );
  AND2_X4 U7761 ( .A1(n5990), .A2(n5969), .ZN(n8967) );
  INV_X1 U7762 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7763 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  XNOR2_X1 U7764 ( .A(n5975), .B(n4746), .ZN(n5991) );
  NAND2_X1 U7765 ( .A1(n6479), .A2(n6497), .ZN(n5976) );
  NOR2_X1 U7766 ( .A1(n9298), .A2(n6047), .ZN(n5977) );
  AOI21_X1 U7767 ( .B1(n9433), .B2(n8961), .A(n5977), .ZN(n8935) );
  INV_X1 U7768 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5978) );
  OR2_X1 U7769 ( .A1(n6055), .A2(n5978), .ZN(n5981) );
  NAND2_X1 U7770 ( .A1(n6036), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5980) );
  INV_X1 U7771 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7450) );
  INV_X1 U7772 ( .A(n6816), .ZN(n5982) );
  NAND2_X1 U7773 ( .A1(n6021), .A2(n5982), .ZN(n5984) );
  NAND2_X1 U7774 ( .A1(n6100), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7775 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5985) );
  MUX2_X1 U7776 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5985), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5987) );
  INV_X1 U7777 ( .A(n6022), .ZN(n5986) );
  INV_X1 U7778 ( .A(n6942), .ZN(n5988) );
  NAND2_X1 U7779 ( .A1(n6764), .A2(n5988), .ZN(n5989) );
  INV_X2 U7780 ( .A(n7158), .ZN(n7454) );
  NAND2_X1 U7781 ( .A1(n5990), .A2(n9444), .ZN(n5992) );
  XNOR2_X1 U7782 ( .A(n5993), .B(n8916), .ZN(n6950) );
  NAND2_X1 U7783 ( .A1(n6008), .A2(n7158), .ZN(n5994) );
  INV_X1 U7784 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7542) );
  INV_X1 U7785 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7786 ( .A1(n6036), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5997) );
  INV_X1 U7787 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5996) );
  INV_X1 U7788 ( .A(n6788), .ZN(n6953) );
  OR2_X1 U7789 ( .A1(n6047), .A2(n6953), .ZN(n6005) );
  INV_X1 U7790 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6919) );
  INV_X1 U7791 ( .A(SI_0_), .ZN(n5999) );
  INV_X1 U7792 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5998) );
  OAI21_X1 U7793 ( .B1(n5061), .B2(n5999), .A(n5998), .ZN(n6001) );
  NAND2_X1 U7794 ( .A1(n6001), .A2(n6000), .ZN(n9776) );
  OAI22_X1 U7795 ( .A1(n8969), .A2(n7150), .B1(n6919), .B2(n5969), .ZN(n6003)
         );
  INV_X1 U7796 ( .A(n6003), .ZN(n6004) );
  AND2_X1 U7797 ( .A1(n6005), .A2(n6004), .ZN(n6961) );
  NOR2_X1 U7798 ( .A1(n5969), .A2(n6006), .ZN(n6007) );
  AOI21_X1 U7799 ( .B1(n8967), .B2(n7541), .A(n6007), .ZN(n6010) );
  NAND2_X1 U7800 ( .A1(n6008), .A2(n6788), .ZN(n6009) );
  NAND2_X1 U7801 ( .A1(n6010), .A2(n6009), .ZN(n6960) );
  NAND2_X1 U7802 ( .A1(n6961), .A2(n6960), .ZN(n6959) );
  INV_X1 U7803 ( .A(n6960), .ZN(n6011) );
  NAND2_X1 U7804 ( .A1(n6959), .A2(n6012), .ZN(n6949) );
  OAI21_X1 U7805 ( .B1(n6950), .B2(n6948), .A(n6949), .ZN(n6014) );
  NAND2_X1 U7806 ( .A1(n6950), .A2(n6948), .ZN(n6013) );
  NAND2_X1 U7807 ( .A1(n6014), .A2(n6013), .ZN(n7020) );
  NAND2_X1 U7808 ( .A1(n6036), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6019) );
  INV_X1 U7809 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6884) );
  INV_X1 U7810 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6015) );
  OR2_X1 U7811 ( .A1(n6055), .A2(n6015), .ZN(n6017) );
  INV_X1 U7812 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7022) );
  NAND4_X1 U7813 ( .A1(n6019), .A2(n6016), .A3(n6017), .A4(n6018), .ZN(n6778)
         );
  INV_X1 U7814 ( .A(n9139), .ZN(n6952) );
  INV_X1 U7815 ( .A(n6811), .ZN(n6020) );
  NAND2_X1 U7816 ( .A1(n6021), .A2(n6020), .ZN(n6027) );
  NAND2_X1 U7817 ( .A1(n6100), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6026) );
  NOR2_X1 U7818 ( .A1(n6024), .A2(n6023), .ZN(n9847) );
  NAND2_X1 U7819 ( .A1(n6764), .A2(n9847), .ZN(n6025) );
  XNOR2_X1 U7820 ( .A(n6028), .B(n8916), .ZN(n6033) );
  OR2_X1 U7821 ( .A1(n6047), .A2(n6952), .ZN(n6030) );
  NAND2_X1 U7822 ( .A1(n6008), .A2(n4428), .ZN(n6029) );
  NAND2_X1 U7823 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  XNOR2_X1 U7824 ( .A(n6033), .B(n6031), .ZN(n7019) );
  NAND2_X1 U7825 ( .A1(n7020), .A2(n7019), .ZN(n6035) );
  INV_X1 U7826 ( .A(n6031), .ZN(n6032) );
  NAND2_X1 U7827 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  NAND2_X1 U7828 ( .A1(n6035), .A2(n6034), .ZN(n9835) );
  INV_X1 U7829 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6885) );
  OR2_X1 U7830 ( .A1(n6238), .A2(n6885), .ZN(n6039) );
  INV_X1 U7831 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6902) );
  OR2_X1 U7832 ( .A1(n6442), .A2(n6902), .ZN(n6038) );
  OR2_X1 U7833 ( .A1(n8067), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6037) );
  INV_X1 U7834 ( .A(n9138), .ZN(n6785) );
  INV_X1 U7835 ( .A(n6814), .ZN(n6041) );
  NAND2_X1 U7836 ( .A1(n6021), .A2(n6041), .ZN(n6045) );
  NAND2_X1 U7837 ( .A1(n6100), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6044) );
  OR2_X1 U7838 ( .A1(n6023), .A2(n4748), .ZN(n6042) );
  XNOR2_X1 U7839 ( .A(n6042), .B(P1_IR_REG_3__SCAN_IN), .ZN(n7072) );
  NAND2_X1 U7840 ( .A1(n6764), .A2(n7072), .ZN(n6043) );
  XNOR2_X1 U7841 ( .A(n6046), .B(n8916), .ZN(n6052) );
  OR2_X1 U7842 ( .A1(n6047), .A2(n6785), .ZN(n6049) );
  NAND2_X1 U7843 ( .A1(n6008), .A2(n7612), .ZN(n6048) );
  NAND2_X1 U7844 ( .A1(n6049), .A2(n6048), .ZN(n6050) );
  XNOR2_X1 U7845 ( .A(n6052), .B(n6050), .ZN(n9834) );
  NAND2_X1 U7846 ( .A1(n9835), .A2(n9834), .ZN(n6054) );
  INV_X1 U7847 ( .A(n6050), .ZN(n6051) );
  NAND2_X1 U7848 ( .A1(n6052), .A2(n6051), .ZN(n6053) );
  NAND2_X1 U7849 ( .A1(n6121), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6060) );
  INV_X1 U7850 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6903) );
  OR2_X1 U7851 ( .A1(n6442), .A2(n6903), .ZN(n6059) );
  OAI21_X1 U7852 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6092), .ZN(n9922) );
  OR2_X1 U7853 ( .A1(n8067), .A2(n9922), .ZN(n6058) );
  INV_X1 U7854 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6056) );
  OR2_X1 U7855 ( .A1(n6055), .A2(n6056), .ZN(n6057) );
  INV_X1 U7856 ( .A(n9137), .ZN(n7606) );
  NAND2_X1 U7857 ( .A1(n6021), .A2(n6817), .ZN(n6067) );
  NAND2_X1 U7858 ( .A1(n6100), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6066) );
  INV_X1 U7859 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7860 ( .A1(n6023), .A2(n6061), .ZN(n6063) );
  NAND2_X1 U7861 ( .A1(n6063), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6062) );
  MUX2_X1 U7862 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6062), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n6064) );
  AND2_X1 U7863 ( .A1(n6064), .A2(n6101), .ZN(n6905) );
  NAND2_X1 U7864 ( .A1(n6764), .A2(n6905), .ZN(n6065) );
  XNOR2_X1 U7865 ( .A(n6068), .B(n8916), .ZN(n6073) );
  OR2_X1 U7866 ( .A1(n6047), .A2(n7606), .ZN(n6070) );
  NAND2_X1 U7867 ( .A1(n6008), .A2(n9920), .ZN(n6069) );
  NAND2_X1 U7868 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  XNOR2_X1 U7869 ( .A(n6073), .B(n6071), .ZN(n7166) );
  INV_X1 U7870 ( .A(n6071), .ZN(n6072) );
  INV_X1 U7871 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6074) );
  OR2_X1 U7872 ( .A1(n6238), .A2(n6074), .ZN(n6078) );
  INV_X1 U7873 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7575) );
  NAND2_X1 U7874 ( .A1(n6094), .A2(n7575), .ZN(n6075) );
  NAND2_X1 U7875 ( .A1(n6123), .A2(n6075), .ZN(n7574) );
  OR2_X1 U7876 ( .A1(n8067), .A2(n7574), .ZN(n6077) );
  INV_X1 U7877 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7444) );
  OR2_X1 U7878 ( .A1(n6442), .A2(n7444), .ZN(n6076) );
  NAND2_X1 U7879 ( .A1(n6080), .A2(n6021), .ZN(n6085) );
  INV_X1 U7880 ( .A(n6101), .ZN(n6082) );
  NAND2_X1 U7881 ( .A1(n6082), .A2(n6081), .ZN(n6117) );
  NAND2_X1 U7882 ( .A1(n6117), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6083) );
  XNOR2_X1 U7883 ( .A(n6083), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7036) );
  AOI22_X1 U7884 ( .A1(n6100), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6764), .B2(
        n7036), .ZN(n6084) );
  NAND2_X1 U7885 ( .A1(n8967), .A2(n7562), .ZN(n6086) );
  OAI21_X1 U7886 ( .B1(n7505), .B2(n8969), .A(n6086), .ZN(n6087) );
  XNOR2_X1 U7887 ( .A(n6087), .B(n8965), .ZN(n7565) );
  OR2_X1 U7888 ( .A1(n6047), .A2(n7505), .ZN(n6089) );
  NAND2_X1 U7889 ( .A1(n6008), .A2(n7562), .ZN(n6088) );
  NAND2_X1 U7890 ( .A1(n6089), .A2(n6088), .ZN(n6111) );
  NAND2_X1 U7891 ( .A1(n7565), .A2(n6111), .ZN(n6113) );
  NAND2_X1 U7892 ( .A1(n4282), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6099) );
  INV_X1 U7893 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6090) );
  OR2_X1 U7894 ( .A1(n8085), .A2(n6090), .ZN(n6098) );
  INV_X1 U7895 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7896 ( .A1(n6092), .A2(n6091), .ZN(n6093) );
  NAND2_X1 U7897 ( .A1(n6094), .A2(n6093), .ZN(n7532) );
  OR2_X1 U7898 ( .A1(n8054), .A2(n7532), .ZN(n6097) );
  INV_X1 U7899 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6095) );
  OR2_X1 U7900 ( .A1(n6442), .A2(n6095), .ZN(n6096) );
  NAND2_X1 U7901 ( .A1(n6101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6102) );
  AOI22_X1 U7902 ( .A1(n8087), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n4427), .B2(
        n6931), .ZN(n6104) );
  NAND2_X1 U7903 ( .A1(n6821), .A2(n8078), .ZN(n6103) );
  XNOR2_X1 U7904 ( .A(n6105), .B(n8916), .ZN(n7563) );
  OR2_X1 U7905 ( .A1(n6047), .A2(n7428), .ZN(n6107) );
  NAND2_X1 U7906 ( .A1(n6008), .A2(n7538), .ZN(n6106) );
  AND2_X1 U7907 ( .A1(n6107), .A2(n6106), .ZN(n7501) );
  AND2_X1 U7908 ( .A1(n7563), .A2(n7501), .ZN(n6114) );
  INV_X1 U7909 ( .A(n6111), .ZN(n7564) );
  INV_X1 U7910 ( .A(n7565), .ZN(n6112) );
  AOI22_X1 U7911 ( .A1(n6114), .A2(n6113), .B1(n7564), .B2(n6112), .ZN(n6115)
         );
  NAND2_X1 U7912 ( .A1(n6116), .A2(n6115), .ZN(n7478) );
  NAND2_X1 U7913 ( .A1(n6829), .A2(n8078), .ZN(n6120) );
  OAI21_X1 U7914 ( .B1(n6117), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6118) );
  XNOR2_X1 U7915 ( .A(n6118), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9143) );
  AOI22_X1 U7916 ( .A1(n8087), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6764), .B2(
        n9143), .ZN(n6119) );
  NAND2_X1 U7917 ( .A1(n6120), .A2(n6119), .ZN(n7589) );
  NAND2_X1 U7918 ( .A1(n7589), .A2(n8967), .ZN(n6130) );
  NAND2_X1 U7919 ( .A1(n4282), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6128) );
  INV_X1 U7920 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7037) );
  OR2_X1 U7921 ( .A1(n8085), .A2(n7037), .ZN(n6127) );
  NAND2_X1 U7922 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  NAND2_X1 U7923 ( .A1(n6143), .A2(n6124), .ZN(n7481) );
  OR2_X1 U7924 ( .A1(n8054), .A2(n7481), .ZN(n6126) );
  INV_X1 U7925 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7417) );
  OR2_X1 U7926 ( .A1(n6442), .A2(n7417), .ZN(n6125) );
  OR2_X1 U7927 ( .A1(n7441), .A2(n8969), .ZN(n6129) );
  NAND2_X1 U7928 ( .A1(n6130), .A2(n6129), .ZN(n6131) );
  XNOR2_X1 U7929 ( .A(n6131), .B(n8916), .ZN(n6136) );
  NAND2_X1 U7930 ( .A1(n7589), .A2(n8961), .ZN(n6133) );
  OR2_X1 U7931 ( .A1(n6047), .A2(n7441), .ZN(n6132) );
  NAND2_X1 U7932 ( .A1(n6133), .A2(n6132), .ZN(n6134) );
  XNOR2_X1 U7933 ( .A(n6136), .B(n6134), .ZN(n7477) );
  NAND2_X1 U7934 ( .A1(n7478), .A2(n7477), .ZN(n6138) );
  INV_X1 U7935 ( .A(n6134), .ZN(n6135) );
  NAND2_X1 U7936 ( .A1(n6136), .A2(n6135), .ZN(n6137) );
  NAND2_X1 U7937 ( .A1(n6834), .A2(n8078), .ZN(n6142) );
  OR2_X1 U7938 ( .A1(n6139), .A2(n4748), .ZN(n6140) );
  XNOR2_X1 U7939 ( .A(n6140), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7040) );
  AOI22_X1 U7940 ( .A1(n8087), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4427), .B2(
        n7040), .ZN(n6141) );
  NAND2_X1 U7941 ( .A1(n4282), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7942 ( .A1(n6143), .A2(n7656), .ZN(n6144) );
  NAND2_X1 U7943 ( .A1(n6161), .A2(n6144), .ZN(n9896) );
  OR2_X1 U7944 ( .A1(n8054), .A2(n9896), .ZN(n6146) );
  INV_X1 U7945 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7032) );
  OR2_X1 U7946 ( .A1(n6442), .A2(n7032), .ZN(n6145) );
  NOR2_X1 U7947 ( .A1(n6047), .A2(n7596), .ZN(n6149) );
  AOI21_X1 U7948 ( .B1(n7653), .B2(n6008), .A(n6149), .ZN(n6153) );
  NAND2_X1 U7949 ( .A1(n7653), .A2(n8967), .ZN(n6151) );
  OR2_X1 U7950 ( .A1(n7596), .A2(n8969), .ZN(n6150) );
  NAND2_X1 U7951 ( .A1(n6151), .A2(n6150), .ZN(n6152) );
  XNOR2_X1 U7952 ( .A(n6152), .B(n8965), .ZN(n7652) );
  INV_X1 U7953 ( .A(n6153), .ZN(n6154) );
  NAND2_X1 U7954 ( .A1(n6842), .A2(n8078), .ZN(n6158) );
  NAND2_X1 U7955 ( .A1(n6155), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6156) );
  XNOR2_X1 U7956 ( .A(n6156), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7042) );
  AOI22_X1 U7957 ( .A1(n8087), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4427), .B2(
        n7042), .ZN(n6157) );
  NAND2_X1 U7958 ( .A1(n7749), .A2(n8967), .ZN(n6168) );
  NAND2_X1 U7959 ( .A1(n4282), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6166) );
  INV_X1 U7960 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7041) );
  OR2_X1 U7961 ( .A1(n8085), .A2(n7041), .ZN(n6165) );
  INV_X1 U7962 ( .A(n6159), .ZN(n6178) );
  NAND2_X1 U7963 ( .A1(n6161), .A2(n6160), .ZN(n6162) );
  NAND2_X1 U7964 ( .A1(n6178), .A2(n6162), .ZN(n7721) );
  OR2_X1 U7965 ( .A1(n8054), .A2(n7721), .ZN(n6164) );
  INV_X1 U7966 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7598) );
  OR2_X1 U7967 ( .A1(n6442), .A2(n7598), .ZN(n6163) );
  OR2_X1 U7968 ( .A1(n7778), .A2(n8969), .ZN(n6167) );
  NAND2_X1 U7969 ( .A1(n6168), .A2(n6167), .ZN(n6169) );
  XNOR2_X1 U7970 ( .A(n6169), .B(n8916), .ZN(n6173) );
  NOR2_X1 U7971 ( .A1(n6047), .A2(n7778), .ZN(n6170) );
  AOI21_X1 U7972 ( .B1(n7749), .B2(n6008), .A(n6170), .ZN(n6172) );
  XNOR2_X1 U7973 ( .A(n6173), .B(n6172), .ZN(n7718) );
  NAND2_X1 U7974 ( .A1(n6173), .A2(n6172), .ZN(n6174) );
  NAND2_X1 U7975 ( .A1(n7715), .A2(n6174), .ZN(n7776) );
  NAND2_X1 U7976 ( .A1(n6840), .A2(n8078), .ZN(n6177) );
  NAND2_X1 U7977 ( .A1(n6194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6175) );
  XNOR2_X1 U7978 ( .A(n6175), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7108) );
  AOI22_X1 U7979 ( .A1(n8087), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4427), .B2(
        n7108), .ZN(n6176) );
  NAND2_X2 U7980 ( .A1(n6177), .A2(n6176), .ZN(n9818) );
  NAND2_X1 U7981 ( .A1(n9818), .A2(n8967), .ZN(n6187) );
  NAND2_X1 U7982 ( .A1(n4282), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7983 ( .A1(n6178), .A2(n4541), .ZN(n6179) );
  NAND2_X1 U7984 ( .A1(n6199), .A2(n6179), .ZN(n9813) );
  OR2_X1 U7985 ( .A1(n8054), .A2(n9813), .ZN(n6184) );
  INV_X1 U7986 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6180) );
  OR2_X1 U7987 ( .A1(n8085), .A2(n6180), .ZN(n6183) );
  INV_X1 U7988 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6181) );
  OR2_X1 U7989 ( .A1(n6442), .A2(n6181), .ZN(n6182) );
  OR2_X1 U7990 ( .A1(n7744), .A2(n8969), .ZN(n6186) );
  NAND2_X1 U7991 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  XNOR2_X1 U7992 ( .A(n6188), .B(n8965), .ZN(n6190) );
  NOR2_X1 U7993 ( .A1(n6047), .A2(n7744), .ZN(n6189) );
  AOI21_X1 U7994 ( .B1(n9818), .B2(n6008), .A(n6189), .ZN(n6191) );
  XNOR2_X1 U7995 ( .A(n6190), .B(n6191), .ZN(n7775) );
  INV_X1 U7996 ( .A(n6190), .ZN(n6192) );
  NAND2_X1 U7997 ( .A1(n6192), .A2(n6191), .ZN(n6193) );
  NAND2_X1 U7998 ( .A1(n6849), .A2(n8078), .ZN(n6197) );
  NOR2_X1 U7999 ( .A1(n6194), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6214) );
  OR2_X1 U8000 ( .A1(n6214), .A2(n4748), .ZN(n6195) );
  XNOR2_X1 U8001 ( .A(n6195), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7132) );
  AOI22_X1 U8002 ( .A1(n8087), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4427), .B2(
        n7132), .ZN(n6196) );
  NAND2_X2 U8003 ( .A1(n6197), .A2(n6196), .ZN(n9725) );
  NAND2_X1 U8004 ( .A1(n9725), .A2(n8967), .ZN(n6207) );
  NAND2_X1 U8005 ( .A1(n4282), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6205) );
  INV_X1 U8006 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7114) );
  OR2_X1 U8007 ( .A1(n6238), .A2(n7114), .ZN(n6204) );
  NAND2_X1 U8008 ( .A1(n6199), .A2(n6198), .ZN(n6200) );
  NAND2_X1 U8009 ( .A1(n6218), .A2(n6200), .ZN(n9079) );
  OR2_X1 U8010 ( .A1(n8054), .A2(n9079), .ZN(n6203) );
  INV_X1 U8011 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6201) );
  OR2_X1 U8012 ( .A1(n6442), .A2(n6201), .ZN(n6202) );
  OR2_X1 U8013 ( .A1(n7791), .A2(n8969), .ZN(n6206) );
  NAND2_X1 U8014 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  XNOR2_X1 U8015 ( .A(n6208), .B(n8916), .ZN(n6211) );
  NOR2_X1 U8016 ( .A1(n6047), .A2(n7791), .ZN(n6209) );
  AOI21_X1 U8017 ( .B1(n9725), .B2(n6008), .A(n6209), .ZN(n6210) );
  XNOR2_X1 U8018 ( .A(n6211), .B(n6210), .ZN(n9083) );
  OR2_X1 U8019 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  NAND2_X1 U8020 ( .A1(n6862), .A2(n8078), .ZN(n6217) );
  AND2_X1 U8021 ( .A1(n6214), .A2(n6213), .ZN(n6233) );
  OR2_X1 U8022 ( .A1(n6233), .A2(n4748), .ZN(n6215) );
  XNOR2_X1 U8023 ( .A(n6215), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7133) );
  AOI22_X1 U8024 ( .A1(n8087), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7133), .B2(
        n4427), .ZN(n6216) );
  NAND2_X2 U8025 ( .A1(n6217), .A2(n6216), .ZN(n9717) );
  NAND2_X1 U8026 ( .A1(n9717), .A2(n8967), .ZN(n6225) );
  NAND2_X1 U8027 ( .A1(n6121), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6223) );
  INV_X1 U8028 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9754) );
  OR2_X1 U8029 ( .A1(n6853), .A2(n9754), .ZN(n6222) );
  NAND2_X1 U8030 ( .A1(n6218), .A2(n4542), .ZN(n6219) );
  NAND2_X1 U8031 ( .A1(n6236), .A2(n6219), .ZN(n9006) );
  OR2_X1 U8032 ( .A1(n8054), .A2(n9006), .ZN(n6221) );
  INV_X1 U8033 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7797) );
  OR2_X1 U8034 ( .A1(n6442), .A2(n7797), .ZN(n6220) );
  OR2_X1 U8035 ( .A1(n9056), .A2(n8969), .ZN(n6224) );
  NAND2_X1 U8036 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  XNOR2_X1 U8037 ( .A(n6226), .B(n8916), .ZN(n6230) );
  NOR2_X1 U8038 ( .A1(n6047), .A2(n9056), .ZN(n6227) );
  AOI21_X1 U8039 ( .B1(n9717), .B2(n8961), .A(n6227), .ZN(n6229) );
  XNOR2_X1 U8040 ( .A(n6230), .B(n6229), .ZN(n9002) );
  NAND2_X1 U8041 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  NAND2_X1 U8042 ( .A1(n6860), .A2(n8078), .ZN(n6235) );
  INV_X1 U8043 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6232) );
  XNOR2_X1 U8044 ( .A(n6249), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7136) );
  AOI22_X1 U8045 ( .A1(n7136), .A2(n4427), .B1(n8087), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U8046 ( .A1(n9712), .A2(n8967), .ZN(n6244) );
  NAND2_X1 U8047 ( .A1(n4282), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U8048 ( .A1(n6236), .A2(n7130), .ZN(n6237) );
  NAND2_X1 U8049 ( .A1(n6254), .A2(n6237), .ZN(n9596) );
  OR2_X1 U8050 ( .A1(n9596), .A2(n8054), .ZN(n6241) );
  INV_X1 U8051 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7135) );
  OR2_X1 U8052 ( .A1(n6238), .A2(n7135), .ZN(n6240) );
  INV_X1 U8053 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7515) );
  OR2_X1 U8054 ( .A1(n6442), .A2(n7515), .ZN(n6239) );
  NAND2_X1 U8055 ( .A1(n9274), .A2(n8961), .ZN(n6243) );
  NAND2_X1 U8056 ( .A1(n6244), .A2(n6243), .ZN(n6245) );
  XNOR2_X1 U8057 ( .A(n6245), .B(n8916), .ZN(n9053) );
  NOR2_X1 U8058 ( .A1(n6047), .A2(n8008), .ZN(n6246) );
  AOI21_X1 U8059 ( .B1(n9712), .B2(n8961), .A(n6246), .ZN(n9052) );
  AND2_X1 U8060 ( .A1(n9053), .A2(n9052), .ZN(n6247) );
  NAND2_X1 U8061 ( .A1(n6878), .A2(n8078), .ZN(n6253) );
  INV_X1 U8062 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U8063 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  NAND2_X1 U8064 ( .A1(n6250), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6251) );
  XNOR2_X1 U8065 ( .A(n6251), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9210) );
  AOI22_X1 U8066 ( .A1(n9210), .A2(n4427), .B1(n8087), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U8067 ( .A1(n9708), .A2(n8967), .ZN(n6261) );
  NAND2_X1 U8068 ( .A1(n6254), .A2(n8927), .ZN(n6255) );
  AND2_X1 U8069 ( .A1(n6282), .A2(n6255), .ZN(n9578) );
  NAND2_X1 U8070 ( .A1(n9578), .A2(n7968), .ZN(n6259) );
  NAND2_X1 U8071 ( .A1(n8069), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6258) );
  INV_X1 U8072 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10248) );
  OR2_X1 U8073 ( .A1(n6853), .A2(n10248), .ZN(n6257) );
  INV_X1 U8074 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10135) );
  OR2_X1 U8075 ( .A1(n8085), .A2(n10135), .ZN(n6256) );
  NAND4_X1 U8076 ( .A1(n6259), .A2(n6258), .A3(n6257), .A4(n6256), .ZN(n9277)
         );
  NAND2_X1 U8077 ( .A1(n6008), .A2(n9277), .ZN(n6260) );
  NAND2_X1 U8078 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  XNOR2_X1 U8079 ( .A(n6262), .B(n8965), .ZN(n8924) );
  INV_X1 U8080 ( .A(n8924), .ZN(n6265) );
  NAND2_X1 U8081 ( .A1(n9708), .A2(n8961), .ZN(n6264) );
  INV_X1 U8082 ( .A(n9277), .ZN(n9057) );
  OR2_X1 U8083 ( .A1(n9057), .A2(n6047), .ZN(n6263) );
  NAND2_X1 U8084 ( .A1(n6264), .A2(n6263), .ZN(n6291) );
  INV_X1 U8085 ( .A(n6291), .ZN(n8923) );
  NAND2_X1 U8086 ( .A1(n6265), .A2(n8923), .ZN(n6295) );
  NAND2_X1 U8087 ( .A1(n8926), .A2(n6295), .ZN(n9011) );
  NAND2_X1 U8088 ( .A1(n7174), .A2(n8078), .ZN(n6270) );
  NOR2_X1 U8089 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6266) );
  NAND2_X1 U8090 ( .A1(n6267), .A2(n6266), .ZN(n6276) );
  NAND2_X1 U8091 ( .A1(n6278), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6268) );
  XNOR2_X1 U8092 ( .A(n6268), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9225) );
  AOI22_X1 U8093 ( .A1(n9225), .A2(n4427), .B1(n8087), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U8094 ( .A1(n6284), .A2(n9022), .ZN(n6271) );
  NAND2_X1 U8095 ( .A1(n6298), .A2(n6271), .ZN(n9537) );
  AOI22_X1 U8096 ( .A1(n6121), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8069), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U8097 ( .A1(n4282), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6272) );
  OAI211_X1 U8098 ( .C1(n9537), .C2(n8054), .A(n6273), .B(n6272), .ZN(n9282)
         );
  INV_X1 U8099 ( .A(n9282), .ZN(n9033) );
  XNOR2_X1 U8100 ( .A(n6274), .B(n8916), .ZN(n6311) );
  OAI22_X1 U8101 ( .A1(n9540), .A2(n8969), .B1(n9033), .B2(n6047), .ZN(n6312)
         );
  INV_X1 U8102 ( .A(n6312), .ZN(n6275) );
  NAND2_X1 U8103 ( .A1(n7083), .A2(n8078), .ZN(n6281) );
  NAND2_X1 U8104 ( .A1(n6276), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6277) );
  MUX2_X1 U8105 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6277), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6279) );
  AOI22_X1 U8106 ( .A1(n9860), .A2(n4427), .B1(n8087), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n6280) );
  NAND2_X2 U8107 ( .A1(n6281), .A2(n6280), .ZN(n9701) );
  NAND2_X1 U8108 ( .A1(n6282), .A2(n4544), .ZN(n6283) );
  NAND2_X1 U8109 ( .A1(n6284), .A2(n6283), .ZN(n9561) );
  OR2_X1 U8110 ( .A1(n9561), .A2(n8054), .ZN(n6289) );
  NAND2_X1 U8111 ( .A1(n6121), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U8112 ( .A1(n4282), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6285) );
  AND2_X1 U8113 ( .A1(n6286), .A2(n6285), .ZN(n6288) );
  NAND2_X1 U8114 ( .A1(n8069), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6287) );
  NOR2_X1 U8115 ( .A1(n9020), .A2(n6047), .ZN(n6290) );
  AOI21_X1 U8116 ( .B1(n9701), .B2(n8961), .A(n6290), .ZN(n9012) );
  INV_X1 U8117 ( .A(n9012), .ZN(n9114) );
  NAND2_X1 U8118 ( .A1(n9026), .A2(n9114), .ZN(n6318) );
  NAND2_X1 U8119 ( .A1(n9701), .A2(n8967), .ZN(n6293) );
  NAND2_X1 U8120 ( .A1(n9279), .A2(n8961), .ZN(n6292) );
  NAND2_X1 U8121 ( .A1(n6293), .A2(n6292), .ZN(n6294) );
  XNOR2_X1 U8122 ( .A(n6294), .B(n8965), .ZN(n6309) );
  AND2_X1 U8123 ( .A1(n6309), .A2(n6295), .ZN(n9013) );
  NAND3_X1 U8124 ( .A1(n9014), .A2(n9013), .A3(n9026), .ZN(n6317) );
  NAND2_X1 U8125 ( .A1(n7386), .A2(n8078), .ZN(n6297) );
  XNOR2_X1 U8126 ( .A(n6337), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9229) );
  AOI22_X1 U8127 ( .A1(n8087), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4427), .B2(
        n9229), .ZN(n6296) );
  NAND2_X1 U8128 ( .A1(n9530), .A2(n8967), .ZN(n6306) );
  NAND2_X1 U8129 ( .A1(n6298), .A2(n4545), .ZN(n6299) );
  NAND2_X1 U8130 ( .A1(n6342), .A2(n6299), .ZN(n9524) );
  OR2_X1 U8131 ( .A1(n9524), .A2(n8054), .ZN(n6304) );
  INV_X1 U8132 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9228) );
  NAND2_X1 U8133 ( .A1(n4282), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U8134 ( .A1(n8069), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6300) );
  OAI211_X1 U8135 ( .C1(n8085), .C2(n9228), .A(n6301), .B(n6300), .ZN(n6302)
         );
  INV_X1 U8136 ( .A(n6302), .ZN(n6303) );
  NAND2_X1 U8137 ( .A1(n9284), .A2(n8961), .ZN(n6305) );
  NAND2_X1 U8138 ( .A1(n6306), .A2(n6305), .ZN(n6307) );
  XNOR2_X1 U8139 ( .A(n6307), .B(n8965), .ZN(n6319) );
  NOR2_X1 U8140 ( .A1(n9021), .A2(n6047), .ZN(n6308) );
  AOI21_X1 U8141 ( .B1(n9530), .B2(n8961), .A(n6308), .ZN(n6320) );
  XNOR2_X1 U8142 ( .A(n6319), .B(n6320), .ZN(n9027) );
  INV_X1 U8143 ( .A(n6309), .ZN(n6310) );
  AND2_X1 U8144 ( .A1(n6310), .A2(n4366), .ZN(n9010) );
  INV_X1 U8145 ( .A(n6311), .ZN(n6313) );
  NAND2_X1 U8146 ( .A1(n6313), .A2(n6312), .ZN(n9015) );
  OAI21_X1 U8147 ( .B1(n9012), .B2(n9010), .A(n9015), .ZN(n6314) );
  NAND2_X1 U8148 ( .A1(n6314), .A2(n9026), .ZN(n6315) );
  AND2_X1 U8149 ( .A1(n9027), .A2(n6315), .ZN(n6316) );
  OAI211_X1 U8150 ( .C1(n9011), .C2(n6318), .A(n6317), .B(n6316), .ZN(n9030)
         );
  INV_X1 U8151 ( .A(n6319), .ZN(n6321) );
  NAND2_X1 U8152 ( .A1(n6321), .A2(n6320), .ZN(n6322) );
  NAND2_X1 U8153 ( .A1(n7557), .A2(n8078), .ZN(n6324) );
  AOI22_X1 U8154 ( .A1(n8087), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4427), .B2(
        n9444), .ZN(n6323) );
  NAND2_X1 U8155 ( .A1(n9678), .A2(n8967), .ZN(n6332) );
  NAND2_X1 U8156 ( .A1(n6344), .A2(n8954), .ZN(n6325) );
  NAND2_X1 U8157 ( .A1(n6366), .A2(n6325), .ZN(n8953) );
  INV_X1 U8158 ( .A(n8953), .ZN(n9493) );
  NAND2_X1 U8159 ( .A1(n9493), .A2(n7968), .ZN(n6330) );
  INV_X1 U8160 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9247) );
  NAND2_X1 U8161 ( .A1(n4282), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U8162 ( .A1(n8069), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6326) );
  OAI211_X1 U8163 ( .C1(n8085), .C2(n9247), .A(n6327), .B(n6326), .ZN(n6328)
         );
  INV_X1 U8164 ( .A(n6328), .ZN(n6329) );
  NAND2_X1 U8165 ( .A1(n9287), .A2(n8961), .ZN(n6331) );
  NAND2_X1 U8166 ( .A1(n6332), .A2(n6331), .ZN(n6333) );
  XNOR2_X1 U8167 ( .A(n6333), .B(n8965), .ZN(n8946) );
  NAND2_X1 U8168 ( .A1(n9678), .A2(n8961), .ZN(n6335) );
  INV_X1 U8169 ( .A(n6047), .ZN(n8962) );
  NAND2_X1 U8170 ( .A1(n9287), .A2(n8962), .ZN(n6334) );
  NAND2_X1 U8171 ( .A1(n6335), .A2(n6334), .ZN(n6359) );
  NAND2_X1 U8172 ( .A1(n7485), .A2(n8078), .ZN(n6341) );
  INV_X1 U8173 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U8174 ( .A1(n6337), .A2(n6336), .ZN(n6338) );
  NAND2_X1 U8175 ( .A1(n6338), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6339) );
  XNOR2_X1 U8176 ( .A(n6339), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9237) );
  AOI22_X1 U8177 ( .A1(n8087), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9237), .B2(
        n4427), .ZN(n6340) );
  NAND2_X1 U8178 ( .A1(n9510), .A2(n8967), .ZN(n6351) );
  NAND2_X1 U8179 ( .A1(n6342), .A2(n9094), .ZN(n6343) );
  NAND2_X1 U8180 ( .A1(n6344), .A2(n6343), .ZN(n9093) );
  OR2_X1 U8181 ( .A1(n9093), .A2(n8054), .ZN(n6349) );
  INV_X1 U8182 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9245) );
  NAND2_X1 U8183 ( .A1(n4282), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6346) );
  INV_X1 U8184 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10256) );
  OR2_X1 U8185 ( .A1(n6442), .A2(n10256), .ZN(n6345) );
  OAI211_X1 U8186 ( .C1(n8085), .C2(n9245), .A(n6346), .B(n6345), .ZN(n6347)
         );
  INV_X1 U8187 ( .A(n6347), .ZN(n6348) );
  INV_X1 U8188 ( .A(n9285), .ZN(n9128) );
  NAND2_X1 U8189 ( .A1(n9128), .A2(n8961), .ZN(n6350) );
  NAND2_X1 U8190 ( .A1(n6351), .A2(n6350), .ZN(n6352) );
  XNOR2_X1 U8191 ( .A(n6352), .B(n8965), .ZN(n6356) );
  NAND2_X1 U8192 ( .A1(n9510), .A2(n8961), .ZN(n6354) );
  NAND2_X1 U8193 ( .A1(n9128), .A2(n8962), .ZN(n6353) );
  NAND2_X1 U8194 ( .A1(n6354), .A2(n6353), .ZN(n9087) );
  AOI22_X1 U8195 ( .A1(n8946), .A2(n6359), .B1(n6356), .B2(n9087), .ZN(n6355)
         );
  INV_X1 U8196 ( .A(n8946), .ZN(n6362) );
  INV_X1 U8197 ( .A(n6356), .ZN(n8944) );
  INV_X1 U8198 ( .A(n9087), .ZN(n6357) );
  NAND2_X1 U8199 ( .A1(n8944), .A2(n6357), .ZN(n6358) );
  NAND2_X1 U8200 ( .A1(n6358), .A2(n6359), .ZN(n6361) );
  INV_X1 U8201 ( .A(n6358), .ZN(n6360) );
  INV_X1 U8202 ( .A(n6359), .ZN(n8945) );
  AOI22_X1 U8203 ( .A1(n6362), .A2(n6361), .B1(n6360), .B2(n8945), .ZN(n6363)
         );
  NAND2_X1 U8204 ( .A1(n7647), .A2(n8078), .ZN(n6365) );
  NAND2_X1 U8205 ( .A1(n8087), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U8206 ( .A1(n9675), .A2(n8967), .ZN(n6373) );
  NAND2_X1 U8207 ( .A1(n6366), .A2(n4547), .ZN(n6367) );
  AND2_X1 U8208 ( .A1(n6382), .A2(n6367), .ZN(n9483) );
  INV_X1 U8209 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U8210 ( .A1(n4282), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U8211 ( .A1(n8069), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6368) );
  OAI211_X1 U8212 ( .C1(n8085), .C2(n6370), .A(n6369), .B(n6368), .ZN(n6371)
         );
  AOI21_X2 U8213 ( .B1(n9483), .B2(n7968), .A(n6371), .ZN(n9290) );
  OR2_X1 U8214 ( .A1(n9290), .A2(n8969), .ZN(n6372) );
  NAND2_X1 U8215 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  XNOR2_X1 U8216 ( .A(n6374), .B(n8916), .ZN(n6376) );
  NOR2_X1 U8217 ( .A1(n9290), .A2(n6047), .ZN(n6375) );
  AOI21_X1 U8218 ( .B1(n9675), .B2(n8961), .A(n6375), .ZN(n6377) );
  INV_X1 U8219 ( .A(n6376), .ZN(n6379) );
  INV_X1 U8220 ( .A(n6377), .ZN(n6378) );
  NAND2_X1 U8221 ( .A1(n6379), .A2(n6378), .ZN(n9045) );
  NAND2_X1 U8222 ( .A1(n7680), .A2(n8078), .ZN(n6381) );
  NAND2_X1 U8223 ( .A1(n8087), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6380) );
  NAND2_X1 U8224 ( .A1(n9669), .A2(n8967), .ZN(n6391) );
  INV_X1 U8225 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U8226 ( .A1(n6382), .A2(n8994), .ZN(n6383) );
  NAND2_X1 U8227 ( .A1(n6401), .A2(n6383), .ZN(n9473) );
  OR2_X1 U8228 ( .A1(n9473), .A2(n8054), .ZN(n6389) );
  INV_X1 U8229 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U8230 ( .A1(n4282), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U8231 ( .A1(n8069), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6384) );
  OAI211_X1 U8232 ( .C1(n8085), .C2(n6386), .A(n6385), .B(n6384), .ZN(n6387)
         );
  INV_X1 U8233 ( .A(n6387), .ZN(n6388) );
  NAND2_X1 U8234 ( .A1(n9294), .A2(n8961), .ZN(n6390) );
  NAND2_X1 U8235 ( .A1(n6391), .A2(n6390), .ZN(n6392) );
  XNOR2_X1 U8236 ( .A(n6392), .B(n8965), .ZN(n6395) );
  NAND2_X1 U8237 ( .A1(n9669), .A2(n8961), .ZN(n6394) );
  NAND2_X1 U8238 ( .A1(n9294), .A2(n8962), .ZN(n6393) );
  NAND2_X1 U8239 ( .A1(n6394), .A2(n6393), .ZN(n6396) );
  AND2_X1 U8240 ( .A1(n6395), .A2(n6396), .ZN(n8990) );
  INV_X1 U8241 ( .A(n6395), .ZN(n6398) );
  INV_X1 U8242 ( .A(n6396), .ZN(n6397) );
  NAND2_X1 U8243 ( .A1(n6398), .A2(n6397), .ZN(n8989) );
  NAND2_X1 U8244 ( .A1(n7830), .A2(n8078), .ZN(n6400) );
  NAND2_X1 U8245 ( .A1(n8087), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U8246 ( .A1(n6401), .A2(n9071), .ZN(n6402) );
  AND2_X1 U8247 ( .A1(n6403), .A2(n6402), .ZN(n9452) );
  NAND2_X1 U8248 ( .A1(n9452), .A2(n7968), .ZN(n6409) );
  INV_X1 U8249 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U8250 ( .A1(n8069), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U8251 ( .A1(n4282), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6404) );
  OAI211_X1 U8252 ( .C1(n8085), .C2(n6406), .A(n6405), .B(n6404), .ZN(n6407)
         );
  INV_X1 U8253 ( .A(n6407), .ZN(n6408) );
  NOR2_X1 U8254 ( .A1(n9296), .A2(n6047), .ZN(n6410) );
  AOI21_X1 U8255 ( .B1(n9663), .B2(n8961), .A(n6410), .ZN(n6412) );
  INV_X1 U8256 ( .A(n9663), .ZN(n9454) );
  XOR2_X1 U8257 ( .A(n8916), .B(n6411), .Z(n9068) );
  NAND2_X1 U8258 ( .A1(n6413), .A2(n6412), .ZN(n9065) );
  OAI21_X1 U8259 ( .B1(n9067), .B2(n9068), .A(n9065), .ZN(n6449) );
  INV_X1 U8260 ( .A(n6449), .ZN(n6417) );
  NAND2_X1 U8261 ( .A1(n9433), .A2(n8967), .ZN(n6415) );
  NAND2_X1 U8262 ( .A1(n9300), .A2(n8961), .ZN(n6414) );
  NAND2_X1 U8263 ( .A1(n6415), .A2(n6414), .ZN(n6416) );
  XNOR2_X1 U8264 ( .A(n6416), .B(n8916), .ZN(n6447) );
  INV_X1 U8265 ( .A(n6447), .ZN(n6452) );
  NAND2_X1 U8266 ( .A1(n6417), .A2(n6452), .ZN(n8933) );
  NAND2_X1 U8267 ( .A1(n7884), .A2(n8078), .ZN(n6419) );
  NAND2_X1 U8268 ( .A1(n8087), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U8269 ( .A1(n9417), .A2(n8967), .ZN(n6430) );
  INV_X1 U8270 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U8271 ( .A1(n6421), .A2(n6420), .ZN(n6422) );
  AND2_X1 U8272 ( .A1(n6438), .A2(n6422), .ZN(n9426) );
  NAND2_X1 U8273 ( .A1(n9426), .A2(n7968), .ZN(n6428) );
  INV_X1 U8274 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U8275 ( .A1(n8069), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U8276 ( .A1(n4282), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6423) );
  OAI211_X1 U8277 ( .C1(n8085), .C2(n6425), .A(n6424), .B(n6423), .ZN(n6426)
         );
  INV_X1 U8278 ( .A(n6426), .ZN(n6427) );
  NAND2_X1 U8279 ( .A1(n9303), .A2(n8961), .ZN(n6429) );
  NAND2_X1 U8280 ( .A1(n6430), .A2(n6429), .ZN(n6431) );
  XNOR2_X1 U8281 ( .A(n6431), .B(n8916), .ZN(n6434) );
  NOR2_X1 U8282 ( .A1(n9302), .A2(n6047), .ZN(n6432) );
  AOI21_X1 U8283 ( .B1(n9417), .B2(n8961), .A(n6432), .ZN(n6433) );
  INV_X1 U8284 ( .A(n6454), .ZN(n6435) );
  OR2_X1 U8285 ( .A1(n6434), .A2(n6433), .ZN(n6450) );
  NAND2_X1 U8286 ( .A1(n6435), .A2(n6450), .ZN(n9038) );
  NOR2_X1 U8287 ( .A1(n9039), .A2(n9038), .ZN(n9037) );
  NAND2_X1 U8288 ( .A1(n8901), .A2(n8078), .ZN(n6437) );
  NAND2_X1 U8289 ( .A1(n8087), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6436) );
  INV_X1 U8290 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U8291 ( .A1(n6438), .A2(n10218), .ZN(n6439) );
  NAND2_X1 U8292 ( .A1(n9409), .A2(n7968), .ZN(n6445) );
  INV_X1 U8293 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n10160) );
  NAND2_X1 U8294 ( .A1(n6121), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U8295 ( .A1(n4282), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6440) );
  OAI211_X1 U8296 ( .C1(n6442), .C2(n10160), .A(n6441), .B(n6440), .ZN(n6443)
         );
  INV_X1 U8297 ( .A(n6443), .ZN(n6444) );
  OAI22_X1 U8298 ( .A1(n9407), .A2(n8969), .B1(n9306), .B2(n6047), .ZN(n8906)
         );
  XNOR2_X1 U8299 ( .A(n6446), .B(n8916), .ZN(n8908) );
  NAND2_X1 U8300 ( .A1(n6449), .A2(n4984), .ZN(n6457) );
  INV_X1 U8301 ( .A(n6450), .ZN(n6453) );
  INV_X1 U8302 ( .A(n8935), .ZN(n6451) );
  NOR3_X1 U8303 ( .A1(n6453), .A2(n6452), .A3(n6451), .ZN(n6455) );
  NOR2_X1 U8304 ( .A1(n6455), .A2(n6454), .ZN(n6456) );
  INV_X1 U8305 ( .A(n6466), .ZN(n7886) );
  NAND2_X1 U8306 ( .A1(n7886), .A2(P1_B_REG_SCAN_IN), .ZN(n6460) );
  INV_X1 U8307 ( .A(P1_B_REG_SCAN_IN), .ZN(n9257) );
  NAND2_X1 U8308 ( .A1(n6466), .A2(n9257), .ZN(n6459) );
  OAI211_X1 U8309 ( .C1(n9772), .C2(n6460), .A(n6458), .B(n6459), .ZN(n9931)
         );
  OR2_X1 U8310 ( .A1(n9931), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6462) );
  OR2_X1 U8311 ( .A1(n6458), .A2(n9772), .ZN(n6461) );
  NAND2_X1 U8312 ( .A1(n6462), .A2(n6461), .ZN(n6868) );
  NAND2_X1 U8313 ( .A1(n5943), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6464) );
  XNOR2_X1 U8314 ( .A(n6464), .B(n6463), .ZN(n7837) );
  AND2_X1 U8315 ( .A1(n7837), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6465) );
  INV_X1 U8316 ( .A(n9935), .ZN(n8225) );
  OR2_X1 U8317 ( .A1(n9931), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6468) );
  OR2_X1 U8318 ( .A1(n6458), .A2(n6466), .ZN(n6467) );
  NOR4_X1 U8319 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6472) );
  NOR4_X1 U8320 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6471) );
  NOR4_X1 U8321 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n6470) );
  NOR4_X1 U8322 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6469) );
  NAND4_X1 U8323 ( .A1(n6472), .A2(n6471), .A3(n6470), .A4(n6469), .ZN(n6477)
         );
  NOR2_X1 U8324 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .ZN(
        n10149) );
  NOR4_X1 U8325 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6475) );
  NOR4_X1 U8326 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6474) );
  NOR4_X1 U8327 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6473) );
  NAND4_X1 U8328 ( .A1(n10149), .A2(n6475), .A3(n6474), .A4(n6473), .ZN(n6476)
         );
  NOR2_X1 U8329 ( .A1(n6477), .A2(n6476), .ZN(n6478) );
  OR2_X1 U8330 ( .A1(n9931), .A2(n6478), .ZN(n6796) );
  NAND3_X1 U8331 ( .A1(n6799), .A2(n7144), .A3(n6873), .ZN(n6482) );
  INV_X1 U8332 ( .A(n7149), .ZN(n6481) );
  INV_X1 U8333 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8334 ( .A1(n6484), .A2(n6483), .ZN(n6485) );
  NAND2_X1 U8335 ( .A1(n7962), .A2(n6485), .ZN(n9103) );
  INV_X1 U8336 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U8337 ( .A1(n4282), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U8338 ( .A1(n8069), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6486) );
  OAI211_X1 U8339 ( .C1(n8085), .C2(n6488), .A(n6487), .B(n6486), .ZN(n6489)
         );
  INV_X1 U8340 ( .A(n6489), .ZN(n6490) );
  INV_X1 U8341 ( .A(n4426), .ZN(n6906) );
  INV_X1 U8342 ( .A(n6873), .ZN(n8156) );
  NOR2_X1 U8343 ( .A1(n9302), .A2(n9102), .ZN(n6493) );
  AOI21_X1 U8344 ( .B1(n9126), .B2(n9116), .A(n6493), .ZN(n9643) );
  INV_X1 U8345 ( .A(n9643), .ZN(n6502) );
  AND2_X1 U8346 ( .A1(n7144), .A2(n6497), .ZN(n6494) );
  NAND2_X1 U8347 ( .A1(n6494), .A2(n6799), .ZN(n9106) );
  INV_X1 U8348 ( .A(n9409), .ZN(n6500) );
  INV_X1 U8349 ( .A(n6868), .ZN(n6495) );
  NAND2_X1 U8350 ( .A1(n7144), .A2(n6495), .ZN(n6496) );
  NAND2_X1 U8351 ( .A1(n6870), .A2(n6496), .ZN(n6503) );
  AND3_X1 U8352 ( .A1(n7145), .A2(n5969), .A3(n7837), .ZN(n6498) );
  NAND2_X1 U8353 ( .A1(n6503), .A2(n6498), .ZN(n6499) );
  OAI22_X1 U8354 ( .A1(n6500), .A2(n9842), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10218), .ZN(n6501) );
  AOI21_X1 U8355 ( .B1(n6502), .B2(n9832), .A(n6501), .ZN(n6504) );
  INV_X1 U8356 ( .A(n9837), .ZN(n8938) );
  NAND3_X1 U8357 ( .A1(n6505), .A2(n6504), .A3(n4989), .ZN(P1_U3223) );
  INV_X1 U8358 ( .A(SI_28_), .ZN(n6506) );
  NAND2_X1 U8359 ( .A1(n6507), .A2(n6506), .ZN(n6511) );
  AND2_X1 U8360 ( .A1(n6508), .A2(n6511), .ZN(n6509) );
  INV_X1 U8361 ( .A(n6511), .ZN(n6513) );
  INV_X1 U8362 ( .A(SI_29_), .ZN(n6558) );
  NAND2_X1 U8363 ( .A1(n6561), .A2(n6558), .ZN(n6514) );
  MUX2_X1 U8364 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4277), .Z(n6559) );
  NAND2_X1 U8365 ( .A1(n6514), .A2(n6559), .ZN(n6516) );
  MUX2_X1 U8366 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n5061), .Z(n6538) );
  XNOR2_X1 U8367 ( .A(n6538), .B(SI_30_), .ZN(n6517) );
  NAND2_X1 U8368 ( .A1(n8079), .A2(n5787), .ZN(n6519) );
  INV_X1 U8369 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7939) );
  OR2_X1 U8370 ( .A1(n6547), .A2(n7939), .ZN(n6518) );
  INV_X1 U8371 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U8372 ( .A1(n6520), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U8373 ( .A1(n6524), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6521) );
  OAI211_X1 U8374 ( .C1(n6527), .C2(n6523), .A(n6522), .B(n6521), .ZN(n8495)
         );
  INV_X1 U8375 ( .A(n8495), .ZN(n6550) );
  OR2_X1 U8376 ( .A1(n8490), .A2(n6550), .ZN(n6742) );
  INV_X1 U8377 ( .A(n6742), .ZN(n6531) );
  NAND2_X1 U8378 ( .A1(n6524), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6530) );
  INV_X1 U8379 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6525) );
  OR2_X1 U8380 ( .A1(n6526), .A2(n6525), .ZN(n6529) );
  INV_X1 U8381 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7942) );
  OR2_X1 U8382 ( .A1(n6527), .A2(n7942), .ZN(n6528) );
  AND3_X1 U8383 ( .A1(n6530), .A2(n6529), .A3(n6528), .ZN(n6568) );
  INV_X1 U8384 ( .A(n6568), .ZN(n7945) );
  OR2_X1 U8385 ( .A1(n7945), .A2(n7684), .ZN(n6574) );
  NAND3_X1 U8386 ( .A1(n6531), .A2(n8646), .A3(n6574), .ZN(n6580) );
  MUX2_X1 U8387 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n5061), .Z(n6532) );
  XNOR2_X1 U8388 ( .A(n6532), .B(SI_31_), .ZN(n6540) );
  INV_X1 U8389 ( .A(n6540), .ZN(n6534) );
  INV_X1 U8390 ( .A(n6538), .ZN(n6533) );
  AOI21_X1 U8391 ( .B1(n6534), .B2(SI_30_), .A(n6533), .ZN(n6546) );
  INV_X1 U8392 ( .A(SI_30_), .ZN(n6535) );
  AOI21_X1 U8393 ( .B1(n6540), .B2(n6535), .A(n6538), .ZN(n6545) );
  NAND2_X1 U8394 ( .A1(n6538), .A2(SI_30_), .ZN(n6536) );
  NAND2_X1 U8395 ( .A1(n6540), .A2(n6536), .ZN(n6537) );
  NOR2_X1 U8396 ( .A1(n6538), .A2(SI_30_), .ZN(n6539) );
  NOR2_X1 U8397 ( .A1(n6540), .A2(n6539), .ZN(n6541) );
  NAND2_X1 U8398 ( .A1(n6542), .A2(n6541), .ZN(n6543) );
  INV_X1 U8399 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8242) );
  OR2_X1 U8400 ( .A1(n6547), .A2(n8242), .ZN(n6548) );
  OR2_X1 U8401 ( .A1(n8737), .A2(n6568), .ZN(n6744) );
  NAND2_X1 U8402 ( .A1(n8490), .A2(n6550), .ZN(n6743) );
  NAND2_X1 U8403 ( .A1(n6744), .A2(n6743), .ZN(n6611) );
  OR2_X1 U8404 ( .A1(n6733), .A2(n8501), .ZN(n6730) );
  AND3_X1 U8405 ( .A1(n6730), .A2(n6729), .A3(n6551), .ZN(n6554) );
  INV_X1 U8406 ( .A(n6612), .ZN(n6552) );
  NAND2_X1 U8407 ( .A1(n8551), .A2(n6552), .ZN(n6553) );
  NAND2_X1 U8408 ( .A1(n6726), .A2(n8417), .ZN(n6556) );
  INV_X1 U8409 ( .A(n8250), .ZN(n8418) );
  NOR2_X1 U8410 ( .A1(n8417), .A2(n8418), .ZN(n6555) );
  AOI22_X1 U8411 ( .A1(n6556), .A2(n6733), .B1(n6555), .B2(n8762), .ZN(n6557)
         );
  NAND2_X1 U8412 ( .A1(n8755), .A2(n8416), .ZN(n6736) );
  XNOR2_X1 U8413 ( .A(n6559), .B(n6558), .ZN(n6560) );
  NAND2_X1 U8414 ( .A1(n8265), .A2(n5787), .ZN(n6564) );
  NAND2_X1 U8415 ( .A1(n6562), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6563) );
  OR2_X1 U8416 ( .A1(n8746), .A2(n6565), .ZN(n6739) );
  NAND2_X1 U8417 ( .A1(n8746), .A2(n6565), .ZN(n6740) );
  NAND2_X1 U8418 ( .A1(n6566), .A2(n6740), .ZN(n6576) );
  OAI21_X1 U8419 ( .B1(n8743), .B2(n6574), .A(n8646), .ZN(n6567) );
  AND2_X1 U8420 ( .A1(n8737), .A2(n6568), .ZN(n6745) );
  INV_X1 U8421 ( .A(n6745), .ZN(n6586) );
  INV_X1 U8422 ( .A(n8737), .ZN(n7941) );
  NAND4_X1 U8423 ( .A1(n7941), .A2(n6628), .A3(n7558), .A4(n8490), .ZN(n6569)
         );
  OAI21_X1 U8424 ( .B1(n6586), .B2(n7558), .A(n6569), .ZN(n6570) );
  NOR2_X1 U8425 ( .A1(n6745), .A2(n8646), .ZN(n6575) );
  OAI21_X1 U8426 ( .B1(n6576), .B2(n4986), .A(n4987), .ZN(n6573) );
  INV_X1 U8427 ( .A(n6573), .ZN(n6579) );
  INV_X1 U8428 ( .A(n6574), .ZN(n6577) );
  OAI211_X1 U8429 ( .C1(n6577), .C2(n6742), .A(n6576), .B(n6575), .ZN(n6578)
         );
  OAI211_X1 U8430 ( .C1(n6580), .C2(n6611), .A(n6579), .B(n6578), .ZN(n6585)
         );
  INV_X1 U8431 ( .A(n6581), .ZN(n6582) );
  NAND2_X1 U8432 ( .A1(n6585), .A2(n6584), .ZN(n6760) );
  INV_X1 U8433 ( .A(n6611), .ZN(n6605) );
  NAND2_X1 U8434 ( .A1(n6586), .A2(n6742), .ZN(n6610) );
  INV_X1 U8435 ( .A(n6610), .ZN(n6604) );
  INV_X1 U8436 ( .A(n8745), .ZN(n6603) );
  INV_X1 U8437 ( .A(n6587), .ZN(n6600) );
  INV_X1 U8438 ( .A(n6995), .ZN(n6993) );
  CLKBUF_X1 U8439 ( .A(n6590), .Z(n8437) );
  NAND2_X1 U8440 ( .A1(n8437), .A2(n10052), .ZN(n6637) );
  AND2_X1 U8441 ( .A1(n6589), .A2(n6637), .ZN(n7179) );
  NAND4_X1 U8442 ( .A1(n6993), .A2(n7009), .A3(n6607), .A4(n7179), .ZN(n6591)
         );
  NOR4_X1 U8443 ( .A1(n6591), .A2(n7056), .A3(n7235), .A4(n10023), .ZN(n6592)
         );
  NAND4_X1 U8444 ( .A1(n6592), .A2(n7623), .A3(n7360), .A4(n7371), .ZN(n6593)
         );
  NOR4_X1 U8445 ( .A1(n7727), .A2(n5582), .A3(n7702), .A4(n6593), .ZN(n6594)
         );
  NAND4_X1 U8446 ( .A1(n7892), .A2(n7854), .A3(n7812), .A4(n6594), .ZN(n6595)
         );
  NOR4_X1 U8447 ( .A1(n5593), .A2(n8696), .A3(n8721), .A4(n6595), .ZN(n6596)
         );
  NAND3_X1 U8448 ( .A1(n8635), .A2(n4982), .A3(n6596), .ZN(n6597) );
  NOR4_X1 U8449 ( .A1(n6598), .A2(n8610), .A3(n8627), .A4(n6597), .ZN(n6599)
         );
  INV_X1 U8450 ( .A(n8581), .ZN(n6717) );
  NAND4_X1 U8451 ( .A1(n6600), .A2(n8559), .A3(n6599), .A4(n6717), .ZN(n6601)
         );
  NOR4_X1 U8452 ( .A1(n8521), .A2(n8499), .A3(n6601), .A4(n4880), .ZN(n6602)
         );
  NAND4_X1 U8453 ( .A1(n6605), .A2(n6604), .A3(n6603), .A4(n6602), .ZN(n6606)
         );
  XNOR2_X1 U8454 ( .A(n6606), .B(n7558), .ZN(n6608) );
  OAI22_X1 U8455 ( .A1(n6608), .A2(n6628), .B1(n6607), .B2(n6757), .ZN(n6750)
         );
  NAND2_X1 U8456 ( .A1(n6628), .A2(n8646), .ZN(n6609) );
  MUX2_X1 U8457 ( .A(n6611), .B(n6610), .S(n6727), .Z(n6749) );
  MUX2_X1 U8458 ( .A(n6613), .B(n6612), .S(n6727), .Z(n6722) );
  AND2_X1 U8459 ( .A1(n6705), .A2(n6614), .ZN(n6615) );
  MUX2_X1 U8460 ( .A(n6616), .B(n6615), .S(n4633), .Z(n6698) );
  INV_X1 U8461 ( .A(n8696), .ZN(n6694) );
  INV_X1 U8462 ( .A(n6634), .ZN(n6619) );
  NAND2_X1 U8463 ( .A1(n6619), .A2(n6618), .ZN(n6624) );
  NAND2_X1 U8464 ( .A1(n6621), .A2(n6620), .ZN(n6623) );
  INV_X1 U8465 ( .A(n6644), .ZN(n6622) );
  AOI21_X1 U8466 ( .B1(n6624), .B2(n6623), .A(n6622), .ZN(n6647) );
  NAND2_X1 U8467 ( .A1(n6649), .A2(n6625), .ZN(n6626) );
  AOI21_X1 U8468 ( .B1(n6634), .B2(n6627), .A(n6626), .ZN(n6636) );
  AND2_X1 U8469 ( .A1(n6637), .A2(n6628), .ZN(n6631) );
  OAI211_X1 U8470 ( .C1(n6631), .C2(n6629), .A(n6630), .B(n6638), .ZN(n6632)
         );
  NAND3_X1 U8471 ( .A1(n6632), .A2(n6640), .A3(n6727), .ZN(n6633) );
  NAND3_X1 U8472 ( .A1(n6634), .A2(n10019), .A3(n6633), .ZN(n6635) );
  OAI21_X1 U8473 ( .B1(n6636), .B2(n4633), .A(n6635), .ZN(n6645) );
  NAND2_X1 U8474 ( .A1(n6638), .A2(n6637), .ZN(n6641) );
  NAND3_X1 U8475 ( .A1(n6641), .A2(n6640), .A3(n6639), .ZN(n6642) );
  NAND3_X1 U8476 ( .A1(n6642), .A2(n4633), .A3(n6630), .ZN(n6643) );
  NAND3_X1 U8477 ( .A1(n6645), .A2(n6644), .A3(n6643), .ZN(n6646) );
  OAI21_X1 U8478 ( .B1(n6647), .B2(n6727), .A(n6646), .ZN(n6648) );
  OAI211_X1 U8479 ( .C1(n6649), .C2(n6727), .A(n6648), .B(n7360), .ZN(n6653)
         );
  MUX2_X1 U8480 ( .A(n6651), .B(n6650), .S(n6727), .Z(n6652) );
  NAND3_X1 U8481 ( .A1(n6653), .A2(n7623), .A3(n6652), .ZN(n6657) );
  MUX2_X1 U8482 ( .A(n6655), .B(n6654), .S(n6727), .Z(n6656) );
  NAND3_X1 U8483 ( .A1(n6657), .A2(n6658), .A3(n6656), .ZN(n6662) );
  AOI21_X1 U8484 ( .B1(n6667), .B2(n6658), .A(n4633), .ZN(n6660) );
  NAND2_X1 U8485 ( .A1(n6665), .A2(n6663), .ZN(n6659) );
  NOR2_X1 U8486 ( .A1(n6660), .A2(n6659), .ZN(n6661) );
  NAND2_X1 U8487 ( .A1(n6662), .A2(n6661), .ZN(n6672) );
  INV_X1 U8488 ( .A(n6663), .ZN(n6664) );
  NAND2_X1 U8489 ( .A1(n6667), .A2(n6664), .ZN(n6666) );
  NAND3_X1 U8490 ( .A1(n6666), .A2(n6673), .A3(n6665), .ZN(n6669) );
  NAND2_X1 U8491 ( .A1(n6675), .A2(n6667), .ZN(n6668) );
  MUX2_X1 U8492 ( .A(n6669), .B(n6668), .S(n4633), .Z(n6670) );
  INV_X1 U8493 ( .A(n6670), .ZN(n6671) );
  NAND2_X1 U8494 ( .A1(n6672), .A2(n6671), .ZN(n6677) );
  NAND3_X1 U8495 ( .A1(n6677), .A2(n6678), .A3(n6673), .ZN(n6674) );
  NAND3_X1 U8496 ( .A1(n6674), .A2(n4633), .A3(n6676), .ZN(n6681) );
  NAND3_X1 U8497 ( .A1(n6677), .A2(n6676), .A3(n6675), .ZN(n6679) );
  NAND3_X1 U8498 ( .A1(n6679), .A2(n6678), .A3(n6727), .ZN(n6680) );
  NAND3_X1 U8499 ( .A1(n6681), .A2(n6680), .A3(n7854), .ZN(n6684) );
  MUX2_X1 U8500 ( .A(n6682), .B(n7890), .S(n4633), .Z(n6683) );
  NAND3_X1 U8501 ( .A1(n6684), .A2(n7892), .A3(n6683), .ZN(n6688) );
  MUX2_X1 U8502 ( .A(n6686), .B(n6685), .S(n4633), .Z(n6687) );
  NAND3_X1 U8503 ( .A1(n6689), .A2(n6688), .A3(n6687), .ZN(n6693) );
  MUX2_X1 U8504 ( .A(n6691), .B(n6690), .S(n6727), .Z(n6692) );
  MUX2_X1 U8505 ( .A(n6696), .B(n6695), .S(n6727), .Z(n6697) );
  NAND2_X1 U8506 ( .A1(n6706), .A2(n6699), .ZN(n6700) );
  NAND2_X1 U8507 ( .A1(n6700), .A2(n6709), .ZN(n6701) );
  NAND3_X1 U8508 ( .A1(n6701), .A2(n8605), .A3(n6707), .ZN(n6702) );
  NAND3_X1 U8509 ( .A1(n6702), .A2(n6710), .A3(n6714), .ZN(n6703) );
  NAND2_X1 U8510 ( .A1(n6706), .A2(n6705), .ZN(n6708) );
  NAND2_X1 U8511 ( .A1(n6708), .A2(n6707), .ZN(n6711) );
  NAND3_X1 U8512 ( .A1(n6711), .A2(n6710), .A3(n6709), .ZN(n6713) );
  NAND3_X1 U8513 ( .A1(n6713), .A2(n8605), .A3(n6712), .ZN(n6715) );
  NAND2_X1 U8514 ( .A1(n8598), .A2(n4633), .ZN(n6719) );
  NAND2_X1 U8515 ( .A1(n8564), .A2(n6727), .ZN(n6718) );
  MUX2_X1 U8516 ( .A(n6719), .B(n6718), .S(n8781), .Z(n6720) );
  NAND3_X1 U8517 ( .A1(n8551), .A2(n6722), .A3(n6721), .ZN(n6724) );
  OR3_X1 U8518 ( .A1(n8769), .A2(n8352), .A3(n6727), .ZN(n6723) );
  NAND3_X1 U8519 ( .A1(n6724), .A2(n6729), .A3(n6723), .ZN(n6725) );
  OAI21_X1 U8520 ( .B1(n8545), .B2(n8571), .A(n6726), .ZN(n6728) );
  INV_X1 U8521 ( .A(n6730), .ZN(n6731) );
  NAND2_X1 U8522 ( .A1(n6731), .A2(n4633), .ZN(n6732) );
  NAND2_X1 U8523 ( .A1(n6733), .A2(n8501), .ZN(n6734) );
  AOI21_X1 U8524 ( .B1(n6736), .B2(n6734), .A(n4633), .ZN(n6735) );
  NOR2_X1 U8525 ( .A1(n6737), .A2(n4633), .ZN(n6738) );
  MUX2_X1 U8526 ( .A(n6740), .B(n6739), .S(n4633), .Z(n6741) );
  INV_X1 U8527 ( .A(n6744), .ZN(n6746) );
  MUX2_X1 U8528 ( .A(n6746), .B(n6745), .S(n4633), .Z(n6747) );
  INV_X1 U8529 ( .A(n6747), .ZN(n6748) );
  NAND4_X1 U8530 ( .A1(n10044), .A2(n8663), .A3(n6752), .A4(n6751), .ZN(n6753)
         );
  OAI211_X1 U8531 ( .C1(n6755), .C2(n6754), .A(n6753), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6759) );
  INV_X1 U8532 ( .A(n7837), .ZN(n6762) );
  OR2_X1 U8533 ( .A1(n6873), .A2(n6762), .ZN(n6763) );
  NAND2_X1 U8534 ( .A1(n6763), .A2(n6882), .ZN(n6914) );
  OR2_X1 U8535 ( .A1(n6914), .A2(n4427), .ZN(n6765) );
  NAND2_X1 U8536 ( .A1(n6765), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  MUX2_X1 U8537 ( .A(n8389), .B(P2_U3152), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n6776) );
  OAI211_X1 U8538 ( .C1(n6768), .C2(n6766), .A(n7842), .B(n6767), .ZN(n6769)
         );
  INV_X1 U8539 ( .A(n6769), .ZN(n6775) );
  NAND2_X1 U8540 ( .A1(n8433), .A2(n8665), .ZN(n6772) );
  NAND2_X1 U8541 ( .A1(n5657), .A2(n8663), .ZN(n6771) );
  NAND2_X1 U8542 ( .A1(n6772), .A2(n6771), .ZN(n10020) );
  INV_X1 U8543 ( .A(n10020), .ZN(n6773) );
  OAI22_X1 U8544 ( .A1(n8300), .A2(n10035), .B1(n6773), .B2(n8392), .ZN(n6774)
         );
  OR3_X1 U8545 ( .A1(n6776), .A2(n6775), .A3(n6774), .ZN(P2_U3220) );
  INV_X1 U8546 ( .A(n6778), .ZN(n6777) );
  NAND2_X1 U8547 ( .A1(n6778), .A2(n9938), .ZN(n8117) );
  INV_X1 U8548 ( .A(n8169), .ZN(n6780) );
  NAND2_X1 U8549 ( .A1(n9140), .A2(n7454), .ZN(n8116) );
  OAI21_X1 U8550 ( .B1(n6780), .B2(n6779), .A(n7403), .ZN(n6784) );
  NAND2_X1 U8551 ( .A1(n6781), .A2(n9444), .ZN(n6783) );
  NAND2_X1 U8552 ( .A1(n6480), .A2(n8216), .ZN(n6782) );
  NAND2_X1 U8553 ( .A1(n6784), .A2(n9553), .ZN(n6794) );
  NAND2_X1 U8554 ( .A1(n9347), .A2(n9140), .ZN(n6787) );
  OR2_X1 U8555 ( .A1(n9260), .A2(n6785), .ZN(n6786) );
  AND2_X1 U8556 ( .A1(n6787), .A2(n6786), .ZN(n7021) );
  NAND2_X1 U8557 ( .A1(n9140), .A2(n7158), .ZN(n6789) );
  NAND2_X1 U8558 ( .A1(n6788), .A2(n7541), .ZN(n7148) );
  NAND2_X1 U8559 ( .A1(n6874), .A2(n7454), .ZN(n6790) );
  XNOR2_X1 U8560 ( .A(n8169), .B(n7420), .ZN(n9941) );
  NAND3_X1 U8561 ( .A1(n6873), .A2(n6792), .A3(n9471), .ZN(n7796) );
  INV_X1 U8562 ( .A(n7796), .ZN(n9895) );
  NAND2_X1 U8563 ( .A1(n9941), .A2(n9895), .ZN(n6793) );
  NAND3_X1 U8564 ( .A1(n6794), .A2(n7021), .A3(n6793), .ZN(n9939) );
  INV_X1 U8565 ( .A(n6796), .ZN(n6797) );
  NOR2_X1 U8566 ( .A1(n9759), .A2(n6797), .ZN(n6798) );
  MUX2_X1 U8567 ( .A(n9939), .B(P1_REG2_REG_2__SCAN_IN), .S(n9603), .Z(n6806)
         );
  OR2_X1 U8568 ( .A1(n7149), .A2(n8101), .ZN(n6800) );
  OAI22_X1 U8569 ( .A1(n9899), .A2(n4433), .B1(n9814), .B2(n7022), .ZN(n6805)
         );
  INV_X1 U8570 ( .A(n9941), .ZN(n6803) );
  OR2_X1 U8571 ( .A1(n5990), .A2(n9471), .ZN(n7432) );
  OR2_X1 U8572 ( .A1(n9925), .A2(n7432), .ZN(n9566) );
  OR2_X1 U8573 ( .A1(n7149), .A2(n8226), .ZN(n6801) );
  NAND2_X1 U8574 ( .A1(n7151), .A2(n4433), .ZN(n7611) );
  OR2_X1 U8575 ( .A1(n7151), .A2(n4433), .ZN(n6802) );
  NAND2_X1 U8576 ( .A1(n7611), .A2(n6802), .ZN(n9937) );
  OAI22_X1 U8577 ( .A1(n6803), .A2(n9566), .B1(n9527), .B2(n9937), .ZN(n6804)
         );
  OR3_X1 U8578 ( .A1(n6806), .A2(n6805), .A3(n6804), .ZN(P1_U3289) );
  INV_X1 U8579 ( .A(n7186), .ZN(n7193) );
  NAND2_X1 U8580 ( .A1(n4277), .A2(P2_U3152), .ZN(n8904) );
  OAI222_X1 U8581 ( .A1(n7193), .A2(P2_U3152), .B1(n8894), .B2(n6811), .C1(
        n6808), .C2(n8904), .ZN(P2_U3356) );
  INV_X1 U8582 ( .A(n7259), .ZN(n7269) );
  OAI222_X1 U8583 ( .A1(n7269), .A2(P2_U3152), .B1(n8894), .B2(n6816), .C1(
        n6809), .C2(n8904), .ZN(P2_U3357) );
  INV_X1 U8584 ( .A(n9847), .ZN(n6901) );
  NOR2_X1 U8585 ( .A1(n5061), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8257) );
  INV_X2 U8586 ( .A(n8257), .ZN(n9774) );
  AND2_X1 U8587 ( .A1(n5061), .A2(P1_U3084), .ZN(n9771) );
  OAI222_X1 U8588 ( .A1(n6901), .A2(P1_U3084), .B1(n9774), .B2(n6811), .C1(
        n6810), .C2(n7832), .ZN(P1_U3351) );
  INV_X1 U8589 ( .A(n7072), .ZN(n7079) );
  OAI222_X1 U8590 ( .A1(n7832), .A2(n6812), .B1(n9774), .B2(n6814), .C1(
        P1_U3084), .C2(n7079), .ZN(P1_U3350) );
  INV_X1 U8591 ( .A(n8904), .ZN(n8891) );
  AOI22_X1 U8592 ( .A1(n7295), .A2(P2_STATE_REG_SCAN_IN), .B1(n8891), .B2(
        P1_DATAO_REG_3__SCAN_IN), .ZN(n6813) );
  OAI21_X1 U8593 ( .B1(n6814), .B2(n8894), .A(n6813), .ZN(P2_U3355) );
  INV_X1 U8594 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6815) );
  OAI222_X1 U8595 ( .A1(n6942), .A2(P1_U3084), .B1(n9774), .B2(n6816), .C1(
        n6815), .C2(n7832), .ZN(P1_U3352) );
  INV_X1 U8596 ( .A(n6817), .ZN(n6819) );
  AOI22_X1 U8597 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n8891), .B1(n7282), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n6818) );
  OAI21_X1 U8598 ( .B1(n6819), .B2(n8894), .A(n6818), .ZN(P2_U3354) );
  INV_X1 U8599 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6820) );
  INV_X1 U8600 ( .A(n6905), .ZN(n6980) );
  OAI222_X1 U8601 ( .A1(n7832), .A2(n6820), .B1(n9774), .B2(n6819), .C1(
        P1_U3084), .C2(n6980), .ZN(P1_U3349) );
  INV_X1 U8602 ( .A(n6821), .ZN(n6824) );
  AOI22_X1 U8603 ( .A1(n6931), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9771), .ZN(n6822) );
  OAI21_X1 U8604 ( .B1(n6824), .B2(n9774), .A(n6822), .ZN(P1_U3348) );
  AOI22_X1 U8605 ( .A1(n7336), .A2(P2_STATE_REG_SCAN_IN), .B1(n8891), .B2(
        P1_DATAO_REG_5__SCAN_IN), .ZN(n6823) );
  OAI21_X1 U8606 ( .B1(n6824), .B2(n8894), .A(n6823), .ZN(P2_U3353) );
  INV_X1 U8607 ( .A(n6080), .ZN(n6827) );
  AOI22_X1 U8608 ( .A1(n7310), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n8891), .ZN(n6825) );
  OAI21_X1 U8609 ( .B1(n6827), .B2(n8894), .A(n6825), .ZN(P2_U3352) );
  INV_X1 U8610 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6828) );
  INV_X1 U8611 ( .A(n7036), .ZN(n6826) );
  OAI222_X1 U8612 ( .A1(n7832), .A2(n6828), .B1(n9774), .B2(n6827), .C1(
        P1_U3084), .C2(n6826), .ZN(P1_U3347) );
  INV_X1 U8613 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6831) );
  INV_X1 U8614 ( .A(n6829), .ZN(n6832) );
  OAI222_X1 U8615 ( .A1(n8904), .A2(n6831), .B1(n8894), .B2(n6832), .C1(
        P2_U3152), .C2(n6830), .ZN(P2_U3351) );
  INV_X1 U8616 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6833) );
  INV_X1 U8617 ( .A(n9143), .ZN(n7038) );
  OAI222_X1 U8618 ( .A1(n7832), .A2(n6833), .B1(n9774), .B2(n6832), .C1(
        P1_U3084), .C2(n7038), .ZN(P1_U3346) );
  INV_X1 U8619 ( .A(n6834), .ZN(n6838) );
  AOI22_X1 U8620 ( .A1(n7201), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n8891), .ZN(n6835) );
  OAI21_X1 U8621 ( .B1(n6838), .B2(n8894), .A(n6835), .ZN(P2_U3350) );
  INV_X1 U8622 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U8623 ( .A1(n7945), .A2(P2_U3966), .ZN(n6836) );
  OAI21_X1 U8624 ( .B1(n6837), .B2(P2_U3966), .A(n6836), .ZN(P2_U3583) );
  INV_X1 U8625 ( .A(n7040), .ZN(n9160) );
  OAI222_X1 U8626 ( .A1(n7832), .A2(n6839), .B1(n9774), .B2(n6838), .C1(
        P1_U3084), .C2(n9160), .ZN(P1_U3345) );
  INV_X1 U8627 ( .A(n6840), .ZN(n6847) );
  AOI22_X1 U8628 ( .A1(n7495), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n8891), .ZN(n6841) );
  OAI21_X1 U8629 ( .B1(n6847), .B2(n8894), .A(n6841), .ZN(P2_U3348) );
  INV_X1 U8630 ( .A(n6842), .ZN(n6846) );
  OAI222_X1 U8631 ( .A1(n8904), .A2(n6844), .B1(n8894), .B2(n6846), .C1(n6843), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8632 ( .A(n7042), .ZN(n9174) );
  OAI222_X1 U8633 ( .A1(P1_U3084), .A2(n9174), .B1(n9774), .B2(n6846), .C1(
        n6845), .C2(n7832), .ZN(P1_U3344) );
  INV_X1 U8634 ( .A(n7108), .ZN(n7113) );
  OAI222_X1 U8635 ( .A1(n7832), .A2(n6848), .B1(n9774), .B2(n6847), .C1(n7113), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8636 ( .A(n7132), .ZN(n7125) );
  INV_X1 U8637 ( .A(n6849), .ZN(n6851) );
  OAI222_X1 U8638 ( .A1(P1_U3084), .A2(n7125), .B1(n9774), .B2(n6851), .C1(
        n6850), .C2(n7832), .ZN(P1_U3342) );
  OAI222_X1 U8639 ( .A1(n8904), .A2(n6852), .B1(n8894), .B2(n6851), .C1(n7641), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  NOR2_X1 U8640 ( .A1(n10009), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U8641 ( .A1(n8069), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6856) );
  INV_X1 U8642 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9608) );
  OR2_X1 U8643 ( .A1(n8085), .A2(n9608), .ZN(n6855) );
  INV_X1 U8644 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9733) );
  OR2_X1 U8645 ( .A1(n6853), .A2(n9733), .ZN(n6854) );
  AND3_X1 U8646 ( .A1(n6856), .A2(n6855), .A3(n6854), .ZN(n8096) );
  INV_X1 U8647 ( .A(n8096), .ZN(n9261) );
  NAND2_X1 U8648 ( .A1(n9261), .A2(P1_U4006), .ZN(n6857) );
  OAI21_X1 U8649 ( .B1(P1_U4006), .B2(n8242), .A(n6857), .ZN(P1_U3586) );
  INV_X1 U8650 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U8651 ( .A1(n6788), .A2(P1_U4006), .ZN(n6858) );
  OAI21_X1 U8652 ( .B1(P1_U4006), .B2(n6859), .A(n6858), .ZN(P1_U3555) );
  INV_X1 U8653 ( .A(n6860), .ZN(n6867) );
  AOI22_X1 U8654 ( .A1(n7870), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8891), .ZN(n6861) );
  OAI21_X1 U8655 ( .B1(n6867), .B2(n8894), .A(n6861), .ZN(P2_U3345) );
  INV_X1 U8656 ( .A(n6862), .ZN(n6864) );
  OAI222_X1 U8657 ( .A1(n8904), .A2(n10220), .B1(n8894), .B2(n6864), .C1(
        P2_U3152), .C2(n6863), .ZN(P2_U3346) );
  INV_X1 U8658 ( .A(n7133), .ZN(n9188) );
  OAI222_X1 U8659 ( .A1(n7832), .A2(n6865), .B1(n9774), .B2(n6864), .C1(
        P1_U3084), .C2(n9188), .ZN(P1_U3341) );
  INV_X1 U8660 ( .A(n7136), .ZN(n7514) );
  OAI222_X1 U8661 ( .A1(P1_U3084), .A2(n7514), .B1(n9774), .B2(n6867), .C1(
        n6866), .C2(n7832), .ZN(P1_U3340) );
  AND2_X1 U8662 ( .A1(n6868), .A2(n9935), .ZN(n6869) );
  NAND2_X1 U8663 ( .A1(n6788), .A2(n7150), .ZN(n8115) );
  NAND2_X1 U8664 ( .A1(n6872), .A2(n8115), .ZN(n8167) );
  NAND3_X1 U8665 ( .A1(n8167), .A2(n7149), .A3(n6873), .ZN(n6876) );
  OR2_X1 U8666 ( .A1(n9260), .A2(n4446), .ZN(n6875) );
  AND2_X1 U8667 ( .A1(n6876), .A2(n6875), .ZN(n7543) );
  OAI21_X1 U8668 ( .B1(n7149), .B2(n7150), .A(n7543), .ZN(n9731) );
  NAND2_X1 U8669 ( .A1(n9995), .A2(n9731), .ZN(n6877) );
  OAI21_X1 U8670 ( .B1(n9995), .B2(n5996), .A(n6877), .ZN(P1_U3454) );
  INV_X1 U8671 ( .A(n6878), .ZN(n6881) );
  OAI222_X1 U8672 ( .A1(n8904), .A2(n6879), .B1(n8894), .B2(n6881), .C1(n7934), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8673 ( .A(n9210), .ZN(n9200) );
  OAI222_X1 U8674 ( .A1(P1_U3084), .A2(n9200), .B1(n9774), .B2(n6881), .C1(
        n6880), .C2(n7832), .ZN(P1_U3339) );
  INV_X1 U8675 ( .A(n6882), .ZN(n6883) );
  NOR2_X2 U8676 ( .A1(P1_U3083), .A2(n6883), .ZN(n9874) );
  INV_X1 U8677 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6913) );
  INV_X1 U8678 ( .A(n9258), .ZN(n6915) );
  NAND2_X1 U8679 ( .A1(n6915), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9766) );
  NOR2_X1 U8680 ( .A1(n6914), .A2(n9766), .ZN(n6907) );
  INV_X1 U8681 ( .A(n6907), .ZN(n9252) );
  MUX2_X1 U8682 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6884), .S(n9847), .Z(n9854)
         );
  INV_X1 U8683 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7162) );
  MUX2_X1 U8684 ( .A(n7162), .B(P1_REG1_REG_1__SCAN_IN), .S(n6942), .Z(n6938)
         );
  AND2_X1 U8685 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6939) );
  NAND2_X1 U8686 ( .A1(n6938), .A2(n6939), .ZN(n6937) );
  OAI21_X1 U8687 ( .B1(n7162), .B2(n6942), .A(n6937), .ZN(n9855) );
  NAND2_X1 U8688 ( .A1(n9854), .A2(n9855), .ZN(n9853) );
  NAND2_X1 U8689 ( .A1(n9847), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7074) );
  NAND2_X1 U8690 ( .A1(n9853), .A2(n7074), .ZN(n6887) );
  MUX2_X1 U8691 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6885), .S(n7072), .Z(n6886)
         );
  NAND2_X1 U8692 ( .A1(n6887), .A2(n6886), .ZN(n7076) );
  NAND2_X1 U8693 ( .A1(n7072), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6888) );
  NAND2_X1 U8694 ( .A1(n7076), .A2(n6888), .ZN(n6969) );
  INV_X1 U8695 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6890) );
  MUX2_X1 U8696 ( .A(n6890), .B(P1_REG1_REG_4__SCAN_IN), .S(n6905), .Z(n6889)
         );
  NAND2_X1 U8697 ( .A1(n6980), .A2(n6890), .ZN(n6971) );
  MUX2_X1 U8698 ( .A(n6090), .B(P1_REG1_REG_5__SCAN_IN), .S(n6931), .Z(n6927)
         );
  NOR2_X1 U8699 ( .A1(n6928), .A2(n6927), .ZN(n6926) );
  INV_X1 U8700 ( .A(n6892), .ZN(n6895) );
  MUX2_X1 U8701 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6074), .S(n7036), .Z(n6891)
         );
  INV_X1 U8702 ( .A(n6891), .ZN(n6894) );
  NAND2_X1 U8703 ( .A1(n6892), .A2(n6891), .ZN(n9147) );
  INV_X1 U8704 ( .A(n9147), .ZN(n6893) );
  AOI21_X1 U8705 ( .B1(n6895), .B2(n6894), .A(n6893), .ZN(n6898) );
  NOR2_X1 U8706 ( .A1(n4426), .A2(P1_U3084), .ZN(n9763) );
  NAND2_X1 U8707 ( .A1(n9763), .A2(n9258), .ZN(n6896) );
  NAND2_X1 U8708 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3084), .ZN(n6897) );
  OAI21_X1 U8709 ( .B1(n6898), .B2(n9249), .A(n6897), .ZN(n6911) );
  INV_X1 U8710 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6899) );
  MUX2_X1 U8711 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6899), .S(n9847), .Z(n9846)
         );
  INV_X1 U8712 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7453) );
  MUX2_X1 U8713 ( .A(n7453), .B(P1_REG2_REG_1__SCAN_IN), .S(n6942), .Z(n6945)
         );
  AND2_X1 U8714 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6900) );
  NAND2_X1 U8715 ( .A1(n6945), .A2(n6900), .ZN(n6944) );
  OAI21_X1 U8716 ( .B1(n7453), .B2(n6942), .A(n6944), .ZN(n9845) );
  AND2_X1 U8717 ( .A1(n9846), .A2(n9845), .ZN(n9843) );
  NOR2_X1 U8718 ( .A1(n6901), .A2(n6899), .ZN(n7069) );
  MUX2_X1 U8719 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6902), .S(n7072), .Z(n7068)
         );
  OAI21_X1 U8720 ( .B1(n9843), .B2(n7069), .A(n7068), .ZN(n7067) );
  OAI21_X1 U8721 ( .B1(n6902), .B2(n7079), .A(n7067), .ZN(n6967) );
  MUX2_X1 U8722 ( .A(n6903), .B(P1_REG2_REG_4__SCAN_IN), .S(n6905), .Z(n6904)
         );
  NOR2_X1 U8723 ( .A1(n6967), .A2(n6904), .ZN(n6966) );
  NOR2_X1 U8724 ( .A1(n6905), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6968) );
  MUX2_X1 U8725 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6095), .S(n6931), .Z(n6932)
         );
  MUX2_X1 U8726 ( .A(n7444), .B(P1_REG2_REG_6__SCAN_IN), .S(n7036), .Z(n6908)
         );
  NAND2_X1 U8727 ( .A1(n6907), .A2(n6906), .ZN(n9850) );
  AOI211_X1 U8728 ( .C1(n6909), .C2(n6908), .A(n4393), .B(n9850), .ZN(n6910)
         );
  AOI211_X1 U8729 ( .C1(n9861), .C2(n7036), .A(n6911), .B(n6910), .ZN(n6912)
         );
  OAI21_X1 U8730 ( .B1(n9241), .B2(n6913), .A(n6912), .ZN(P1_U3247) );
  INV_X1 U8731 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6925) );
  INV_X1 U8732 ( .A(n6914), .ZN(n6923) );
  INV_X1 U8733 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7547) );
  AOI21_X1 U8734 ( .B1(n6915), .B2(n7547), .A(n4426), .ZN(n6918) );
  INV_X1 U8735 ( .A(n9766), .ZN(n6916) );
  AOI21_X1 U8736 ( .B1(n9763), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6916), .ZN(
        n6917) );
  NOR2_X1 U8737 ( .A1(n6918), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6964) );
  AOI211_X1 U8738 ( .C1(n6918), .C2(P1_IR_REG_0__SCAN_IN), .A(n6917), .B(n6964), .ZN(n6922) );
  NOR2_X1 U8739 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7542), .ZN(n6921) );
  NOR3_X1 U8740 ( .A1(n9249), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6919), .ZN(
        n6920) );
  AOI211_X1 U8741 ( .C1(n6923), .C2(n6922), .A(n6921), .B(n6920), .ZN(n6924)
         );
  OAI21_X1 U8742 ( .B1(n9241), .B2(n6925), .A(n6924), .ZN(P1_U3241) );
  INV_X1 U8743 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6936) );
  AND2_X1 U8744 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n6930) );
  AOI211_X1 U8745 ( .C1(n6928), .C2(n6927), .A(n6926), .B(n9249), .ZN(n6929)
         );
  AOI211_X1 U8746 ( .C1(n9861), .C2(n6931), .A(n6930), .B(n6929), .ZN(n6935)
         );
  NOR3_X1 U8747 ( .A1(n6966), .A2(n6932), .A3(n6968), .ZN(n6933) );
  OAI21_X1 U8748 ( .B1(n4391), .B2(n6933), .A(n9879), .ZN(n6934) );
  OAI211_X1 U8749 ( .C1(n6936), .C2(n9241), .A(n6935), .B(n6934), .ZN(P1_U3246) );
  NAND2_X1 U8750 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n6941) );
  OAI211_X1 U8751 ( .C1(n6939), .C2(n6938), .A(n9878), .B(n6937), .ZN(n6940)
         );
  OAI211_X1 U8752 ( .C1(n9871), .C2(n6942), .A(n6941), .B(n6940), .ZN(n6943)
         );
  INV_X1 U8753 ( .A(n6943), .ZN(n6947) );
  NAND2_X1 U8754 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6962) );
  OAI211_X1 U8755 ( .C1(n6900), .C2(n6945), .A(n9879), .B(n6944), .ZN(n6946)
         );
  OAI211_X1 U8756 ( .C1(n10185), .C2(n9241), .A(n6947), .B(n6946), .ZN(
        P1_U3242) );
  XNOR2_X1 U8757 ( .A(n6949), .B(n6948), .ZN(n6951) );
  XNOR2_X1 U8758 ( .A(n6951), .B(n6950), .ZN(n6956) );
  NAND2_X1 U8759 ( .A1(n9837), .A2(n7145), .ZN(n7028) );
  OAI22_X1 U8760 ( .A1(n9102), .A2(n6953), .B1(n6952), .B2(n9260), .ZN(n7154)
         );
  AOI22_X1 U8761 ( .A1(n7028), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n7154), .B2(
        n9832), .ZN(n6955) );
  NAND2_X1 U8762 ( .A1(n9121), .A2(n7158), .ZN(n6954) );
  OAI211_X1 U8763 ( .C1(n6956), .C2(n9110), .A(n6955), .B(n6954), .ZN(P1_U3220) );
  NAND3_X1 U8764 ( .A1(n9879), .A2(P1_REG2_REG_4__SCAN_IN), .A3(n6967), .ZN(
        n6958) );
  NAND3_X1 U8765 ( .A1(n9878), .A2(P1_REG1_REG_4__SCAN_IN), .A3(n6969), .ZN(
        n6957) );
  AND3_X1 U8766 ( .A1(n6958), .A2(n9871), .A3(n6957), .ZN(n6981) );
  OAI21_X1 U8767 ( .B1(n6961), .B2(n6960), .A(n6959), .ZN(n7027) );
  MUX2_X1 U8768 ( .A(n6962), .B(n7027), .S(n9258), .Z(n6963) );
  NOR2_X1 U8769 ( .A1(n6963), .A2(n4426), .ZN(n6965) );
  NOR3_X1 U8770 ( .A1(n6965), .A2(n6964), .A3(n9129), .ZN(n9851) );
  INV_X1 U8771 ( .A(n9851), .ZN(n6979) );
  AOI21_X1 U8772 ( .B1(n6968), .B2(n6967), .A(n6966), .ZN(n6976) );
  NAND2_X1 U8773 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n6975) );
  INV_X1 U8774 ( .A(n6969), .ZN(n6972) );
  OAI21_X1 U8775 ( .B1(n6972), .B2(n6971), .A(n6970), .ZN(n6973) );
  NAND2_X1 U8776 ( .A1(n9878), .A2(n6973), .ZN(n6974) );
  OAI211_X1 U8777 ( .C1(n9850), .C2(n6976), .A(n6975), .B(n6974), .ZN(n6977)
         );
  AOI21_X1 U8778 ( .B1(n9874), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6977), .ZN(
        n6978) );
  OAI211_X1 U8779 ( .C1(n6981), .C2(n6980), .A(n6979), .B(n6978), .ZN(P1_U3245) );
  XNOR2_X1 U8780 ( .A(n7089), .B(n4416), .ZN(n6984) );
  NOR2_X1 U8781 ( .A1(n6984), .A2(n6983), .ZN(n7087) );
  AOI21_X1 U8782 ( .B1(n6984), .B2(n6983), .A(n7087), .ZN(n6990) );
  INV_X1 U8783 ( .A(n8392), .ZN(n8407) );
  INV_X1 U8784 ( .A(n8437), .ZN(n7101) );
  OAI22_X1 U8785 ( .A1(n7101), .A2(n8563), .B1(n6770), .B2(n8336), .ZN(n6996)
         );
  INV_X1 U8786 ( .A(n6985), .ZN(n6986) );
  NAND2_X1 U8787 ( .A1(n6986), .A2(n10050), .ZN(n7098) );
  AOI22_X1 U8788 ( .A1(n8407), .A2(n6996), .B1(n7098), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6989) );
  INV_X1 U8789 ( .A(n6987), .ZN(n7223) );
  NAND2_X1 U8790 ( .A1(n8411), .A2(n7223), .ZN(n6988) );
  OAI211_X1 U8791 ( .C1(n6990), .C2(n8413), .A(n6989), .B(n6988), .ZN(P2_U3224) );
  INV_X1 U8792 ( .A(n6991), .ZN(n6992) );
  AOI21_X1 U8793 ( .B1(n6994), .B2(n6993), .A(n6992), .ZN(n7222) );
  XNOR2_X1 U8794 ( .A(n6995), .B(n6589), .ZN(n6997) );
  AOI21_X1 U8795 ( .B1(n10021), .B2(n6997), .A(n6996), .ZN(n7227) );
  INV_X1 U8796 ( .A(n7011), .ZN(n6998) );
  AOI211_X1 U8797 ( .C1(n7099), .C2(n7223), .A(n8816), .B(n6998), .ZN(n7219)
         );
  AOI21_X1 U8798 ( .B1(n8840), .B2(n7223), .A(n7219), .ZN(n6999) );
  OAI211_X1 U8799 ( .C1(n7222), .C2(n8849), .A(n7227), .B(n6999), .ZN(n7001)
         );
  NAND2_X1 U8800 ( .A1(n10082), .A2(n7001), .ZN(n7000) );
  OAI21_X1 U8801 ( .B1(n10082), .B2(n5858), .A(n7000), .ZN(P2_U3521) );
  INV_X1 U8802 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7003) );
  NAND2_X1 U8803 ( .A1(n10076), .A2(n7001), .ZN(n7002) );
  OAI21_X1 U8804 ( .B1(n10076), .B2(n7003), .A(n7002), .ZN(P2_U3454) );
  OAI21_X1 U8805 ( .B1(n7006), .B2(n7005), .A(n7004), .ZN(n7475) );
  INV_X1 U8806 ( .A(n7475), .ZN(n7014) );
  OAI21_X1 U8807 ( .B1(n7009), .B2(n7008), .A(n7007), .ZN(n7010) );
  INV_X1 U8808 ( .A(n8434), .ZN(n7248) );
  OAI22_X1 U8809 ( .A1(n7248), .A2(n8336), .B1(n5649), .B2(n8563), .ZN(n7095)
         );
  AOI21_X1 U8810 ( .B1(n7010), .B2(n10021), .A(n7095), .ZN(n7471) );
  OR2_X1 U8811 ( .A1(n10034), .A2(n8816), .ZN(n10036) );
  AOI21_X1 U8812 ( .B1(n7012), .B2(n7011), .A(n10036), .ZN(n7469) );
  AOI21_X1 U8813 ( .B1(n8840), .B2(n7012), .A(n7469), .ZN(n7013) );
  OAI211_X1 U8814 ( .C1(n7014), .C2(n8849), .A(n7471), .B(n7013), .ZN(n7016)
         );
  NAND2_X1 U8815 ( .A1(n10082), .A2(n7016), .ZN(n7015) );
  OAI21_X1 U8816 ( .B1(n10082), .B2(n5857), .A(n7015), .ZN(P2_U3522) );
  INV_X1 U8817 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7018) );
  NAND2_X1 U8818 ( .A1(n10076), .A2(n7016), .ZN(n7017) );
  OAI21_X1 U8819 ( .B1(n10076), .B2(n7018), .A(n7017), .ZN(P2_U3457) );
  XOR2_X1 U8820 ( .A(n7019), .B(n7020), .Z(n7026) );
  INV_X1 U8821 ( .A(n7028), .ZN(n7023) );
  OAI22_X1 U8822 ( .A1(n7023), .A2(n7022), .B1(n7021), .B2(n9106), .ZN(n7024)
         );
  AOI21_X1 U8823 ( .B1(n9121), .B2(n4428), .A(n7024), .ZN(n7025) );
  OAI21_X1 U8824 ( .B1(n7026), .B2(n9110), .A(n7025), .ZN(P1_U3235) );
  INV_X1 U8825 ( .A(n7027), .ZN(n7031) );
  AOI22_X1 U8826 ( .A1(n9121), .A2(n7541), .B1(n7028), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n7030) );
  NAND3_X1 U8827 ( .A1(n9832), .A2(n9116), .A3(n9140), .ZN(n7029) );
  OAI211_X1 U8828 ( .C1(n7031), .C2(n9110), .A(n7030), .B(n7029), .ZN(P1_U3230) );
  MUX2_X1 U8829 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7417), .S(n9143), .Z(n9141)
         );
  NAND2_X1 U8830 ( .A1(n9142), .A2(n9141), .ZN(n9155) );
  NAND2_X1 U8831 ( .A1(n7038), .A2(n7417), .ZN(n9153) );
  MUX2_X1 U8832 ( .A(n7032), .B(P1_REG2_REG_8__SCAN_IN), .S(n7040), .Z(n9154)
         );
  AOI21_X1 U8833 ( .B1(n9155), .B2(n9153), .A(n9154), .ZN(n9157) );
  MUX2_X1 U8834 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n7598), .S(n7042), .Z(n9171)
         );
  NAND2_X1 U8835 ( .A1(n9172), .A2(n9171), .ZN(n9170) );
  NAND2_X1 U8836 ( .A1(n7042), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7034) );
  MUX2_X1 U8837 ( .A(n6181), .B(P1_REG2_REG_10__SCAN_IN), .S(n7108), .Z(n7033)
         );
  AOI21_X1 U8838 ( .B1(n9170), .B2(n7034), .A(n7033), .ZN(n7107) );
  AND3_X1 U8839 ( .A1(n9170), .A2(n7034), .A3(n7033), .ZN(n7035) );
  NOR3_X1 U8840 ( .A1(n7107), .A2(n7035), .A3(n9850), .ZN(n7050) );
  OR2_X1 U8841 ( .A1(n7036), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U8842 ( .A1(n7038), .A2(n7037), .ZN(n7039) );
  OAI21_X1 U8843 ( .B1(n7038), .B2(n7037), .A(n7039), .ZN(n9145) );
  INV_X1 U8844 ( .A(n7039), .ZN(n9162) );
  INV_X1 U8845 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10002) );
  MUX2_X1 U8846 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10002), .S(n7040), .Z(n9163)
         );
  OAI21_X1 U8847 ( .B1(n9164), .B2(n9162), .A(n9163), .ZN(n9178) );
  NAND2_X1 U8848 ( .A1(n9160), .A2(n10002), .ZN(n9176) );
  MUX2_X1 U8849 ( .A(n7041), .B(P1_REG1_REG_9__SCAN_IN), .S(n7042), .Z(n9177)
         );
  AOI21_X1 U8850 ( .B1(n9178), .B2(n9176), .A(n9177), .ZN(n9180) );
  NOR2_X1 U8851 ( .A1(n7042), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7043) );
  MUX2_X1 U8852 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6180), .S(n7108), .Z(n7044)
         );
  OAI21_X1 U8853 ( .B1(n9180), .B2(n7043), .A(n7044), .ZN(n7117) );
  OR3_X1 U8854 ( .A1(n9180), .A2(n7044), .A3(n7043), .ZN(n7045) );
  AOI21_X1 U8855 ( .B1(n7117), .B2(n7045), .A(n9249), .ZN(n7049) );
  NAND2_X1 U8856 ( .A1(n9874), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U8857 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3084), .ZN(n7046) );
  OAI211_X1 U8858 ( .C1(n9871), .C2(n7113), .A(n7047), .B(n7046), .ZN(n7048)
         );
  OR3_X1 U8859 ( .A1(n7050), .A2(n7049), .A3(n7048), .ZN(P1_U3251) );
  INV_X1 U8860 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7064) );
  OAI21_X1 U8861 ( .B1(n7051), .B2(n7056), .A(n7358), .ZN(n7053) );
  INV_X1 U8862 ( .A(n7053), .ZN(n7344) );
  NAND2_X1 U8863 ( .A1(n7055), .A2(n7054), .ZN(n7057) );
  XNOR2_X1 U8864 ( .A(n7057), .B(n7056), .ZN(n7060) );
  NAND2_X1 U8865 ( .A1(n8431), .A2(n8665), .ZN(n7059) );
  NAND2_X1 U8866 ( .A1(n8433), .A2(n8663), .ZN(n7058) );
  NAND2_X1 U8867 ( .A1(n7059), .A2(n7058), .ZN(n7391) );
  AOI21_X1 U8868 ( .B1(n7060), .B2(n10021), .A(n7391), .ZN(n7340) );
  AOI21_X1 U8869 ( .B1(n7238), .B2(n4635), .A(n8816), .ZN(n7061) );
  AND2_X1 U8870 ( .A1(n7376), .A2(n7061), .ZN(n7338) );
  AOI21_X1 U8871 ( .B1(n8840), .B2(n4635), .A(n7338), .ZN(n7062) );
  OAI211_X1 U8872 ( .C1(n7344), .C2(n8849), .A(n7340), .B(n7062), .ZN(n7065)
         );
  NAND2_X1 U8873 ( .A1(n7065), .A2(n10076), .ZN(n7063) );
  OAI21_X1 U8874 ( .B1(n10076), .B2(n7064), .A(n7063), .ZN(P2_U3466) );
  NAND2_X1 U8875 ( .A1(n7065), .A2(n10082), .ZN(n7066) );
  OAI21_X1 U8876 ( .B1(n10082), .B2(n5868), .A(n7066), .ZN(P2_U3525) );
  INV_X1 U8877 ( .A(n7067), .ZN(n7071) );
  NOR3_X1 U8878 ( .A1(n9843), .A2(n7069), .A3(n7068), .ZN(n7070) );
  NOR3_X1 U8879 ( .A1(n9850), .A2(n7071), .A3(n7070), .ZN(n7081) );
  NAND2_X1 U8880 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3084), .ZN(n7078) );
  MUX2_X1 U8881 ( .A(n6885), .B(P1_REG1_REG_3__SCAN_IN), .S(n7072), .Z(n7073)
         );
  NAND3_X1 U8882 ( .A1(n9853), .A2(n7074), .A3(n7073), .ZN(n7075) );
  NAND3_X1 U8883 ( .A1(n9878), .A2(n7076), .A3(n7075), .ZN(n7077) );
  OAI211_X1 U8884 ( .C1(n9871), .C2(n7079), .A(n7078), .B(n7077), .ZN(n7080)
         );
  AOI211_X1 U8885 ( .C1(P1_ADDR_REG_3__SCAN_IN), .C2(n9874), .A(n7081), .B(
        n7080), .ZN(n7082) );
  INV_X1 U8886 ( .A(n7082), .ZN(P1_U3244) );
  INV_X1 U8887 ( .A(n7083), .ZN(n7085) );
  INV_X1 U8888 ( .A(n9860), .ZN(n9204) );
  OAI222_X1 U8889 ( .A1(n7832), .A2(n7084), .B1(n9774), .B2(n7085), .C1(
        P1_U3084), .C2(n9204), .ZN(P1_U3338) );
  OAI222_X1 U8890 ( .A1(n8904), .A2(n7086), .B1(n8894), .B2(n7085), .C1(
        P2_U3152), .C2(n8445), .ZN(P2_U3343) );
  AOI21_X1 U8891 ( .B1(n7089), .B2(n4416), .A(n7087), .ZN(n7093) );
  NAND2_X1 U8892 ( .A1(n7091), .A2(n7090), .ZN(n7092) );
  XNOR2_X1 U8893 ( .A(n7093), .B(n7092), .ZN(n7094) );
  NAND2_X1 U8894 ( .A1(n7094), .A2(n7842), .ZN(n7097) );
  AOI22_X1 U8895 ( .A1(n8407), .A2(n7095), .B1(n7098), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7096) );
  OAI211_X1 U8896 ( .C1(n7472), .C2(n8300), .A(n7097), .B(n7096), .ZN(P2_U3239) );
  INV_X1 U8897 ( .A(n7098), .ZN(n7106) );
  INV_X1 U8898 ( .A(n8381), .ZN(n7771) );
  AOI22_X1 U8899 ( .A1(n7099), .A2(n8411), .B1(n7771), .B2(n8435), .ZN(n7105)
         );
  OAI21_X1 U8900 ( .B1(n7101), .B2(n7100), .A(n10052), .ZN(n7102) );
  NAND3_X1 U8901 ( .A1(n7842), .A2(n7103), .A3(n7102), .ZN(n7104) );
  OAI211_X1 U8902 ( .C1(n7106), .C2(n5009), .A(n7105), .B(n7104), .ZN(P2_U3234) );
  MUX2_X1 U8903 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n6201), .S(n7132), .Z(n7109)
         );
  NOR2_X1 U8904 ( .A1(n7110), .A2(n7109), .ZN(n7111) );
  OAI21_X1 U8905 ( .B1(n7111), .B2(n7124), .A(n9879), .ZN(n7123) );
  NAND2_X1 U8906 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n7112) );
  OAI21_X1 U8907 ( .B1(n9871), .B2(n7125), .A(n7112), .ZN(n7121) );
  NAND2_X1 U8908 ( .A1(n7113), .A2(n6180), .ZN(n7115) );
  MUX2_X1 U8909 ( .A(n7114), .B(P1_REG1_REG_11__SCAN_IN), .S(n7132), .Z(n7116)
         );
  INV_X1 U8910 ( .A(n9193), .ZN(n7119) );
  NAND3_X1 U8911 ( .A1(n7117), .A2(n7116), .A3(n7115), .ZN(n7118) );
  AOI21_X1 U8912 ( .B1(n7119), .B2(n7118), .A(n9249), .ZN(n7120) );
  AOI211_X1 U8913 ( .C1(n9874), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7121), .B(
        n7120), .ZN(n7122) );
  NAND2_X1 U8914 ( .A1(n7123), .A2(n7122), .ZN(P1_U3252) );
  MUX2_X1 U8915 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n7797), .S(n7133), .Z(n9185)
         );
  NAND2_X1 U8916 ( .A1(n7133), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7126) );
  MUX2_X1 U8917 ( .A(n7515), .B(P1_REG2_REG_13__SCAN_IN), .S(n7136), .Z(n7127)
         );
  INV_X1 U8918 ( .A(n9184), .ZN(n7129) );
  NAND2_X1 U8919 ( .A1(n7127), .A2(n7126), .ZN(n7128) );
  OAI21_X1 U8920 ( .B1(n7129), .B2(n7128), .A(n9879), .ZN(n7143) );
  NOR2_X1 U8921 ( .A1(n7130), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9060) );
  NOR2_X1 U8922 ( .A1(n9871), .A2(n7514), .ZN(n7131) );
  AOI211_X1 U8923 ( .C1(n9874), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n9060), .B(
        n7131), .ZN(n7142) );
  NOR2_X1 U8924 ( .A1(n7132), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9192) );
  INV_X1 U8925 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U8926 ( .A1(n9188), .A2(n9723), .ZN(n7139) );
  NAND2_X1 U8927 ( .A1(n7133), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7134) );
  AND2_X1 U8928 ( .A1(n7139), .A2(n7134), .ZN(n9191) );
  OAI21_X1 U8929 ( .B1(n9193), .B2(n9192), .A(n9191), .ZN(n9190) );
  NAND2_X1 U8930 ( .A1(n7514), .A2(n7135), .ZN(n7518) );
  NAND2_X1 U8931 ( .A1(n7136), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U8932 ( .A1(n7518), .A2(n7137), .ZN(n7138) );
  AOI21_X1 U8933 ( .B1(n9190), .B2(n7139), .A(n7138), .ZN(n7520) );
  AND3_X1 U8934 ( .A1(n9190), .A2(n7139), .A3(n7138), .ZN(n7140) );
  OAI21_X1 U8935 ( .B1(n7520), .B2(n7140), .A(n9878), .ZN(n7141) );
  OAI211_X1 U8936 ( .C1(n7513), .C2(n7143), .A(n7142), .B(n7141), .ZN(P1_U3254) );
  XNOR2_X1 U8937 ( .A(n9140), .B(n7454), .ZN(n8170) );
  XNOR2_X1 U8938 ( .A(n8170), .B(n7148), .ZN(n7456) );
  INV_X1 U8939 ( .A(n7456), .ZN(n7160) );
  NOR2_X1 U8940 ( .A1(n7454), .A2(n7150), .ZN(n7152) );
  NOR2_X1 U8941 ( .A1(n7152), .A2(n7151), .ZN(n7153) );
  NAND2_X1 U8942 ( .A1(n9986), .A2(n7153), .ZN(n7449) );
  INV_X1 U8943 ( .A(n7449), .ZN(n7157) );
  XOR2_X1 U8944 ( .A(n6872), .B(n8170), .Z(n7156) );
  INV_X1 U8945 ( .A(n7154), .ZN(n7155) );
  OAI21_X1 U8946 ( .B1(n7156), .B2(n9908), .A(n7155), .ZN(n7451) );
  AOI211_X1 U8947 ( .C1(n9726), .C2(n7158), .A(n7157), .B(n7451), .ZN(n7159)
         );
  OAI21_X1 U8948 ( .B1(n9991), .B2(n7160), .A(n7159), .ZN(n7163) );
  NAND2_X1 U8949 ( .A1(n7163), .A2(n10006), .ZN(n7161) );
  OAI21_X1 U8950 ( .B1(n10006), .B2(n7162), .A(n7161), .ZN(P1_U3524) );
  NAND2_X1 U8951 ( .A1(n7163), .A2(n9995), .ZN(n7164) );
  OAI21_X1 U8952 ( .B1(n9995), .B2(n5978), .A(n7164), .ZN(P1_U3457) );
  XNOR2_X1 U8953 ( .A(n7166), .B(n7165), .ZN(n7172) );
  NAND2_X1 U8954 ( .A1(n9347), .A2(n9138), .ZN(n7168) );
  OR2_X1 U8955 ( .A1(n9260), .A2(n7428), .ZN(n7167) );
  NAND2_X1 U8956 ( .A1(n7168), .A2(n7167), .ZN(n9910) );
  AOI22_X1 U8957 ( .A1(n9910), .A2(n9832), .B1(P1_REG3_REG_4__SCAN_IN), .B2(
        P1_U3084), .ZN(n7170) );
  AND2_X1 U8958 ( .A1(n9726), .A2(n9920), .ZN(n9948) );
  NAND2_X1 U8959 ( .A1(n9837), .A2(n9948), .ZN(n7169) );
  OAI211_X1 U8960 ( .C1(n9842), .C2(n9922), .A(n7170), .B(n7169), .ZN(n7171)
         );
  AOI21_X1 U8961 ( .B1(n7172), .B2(n9838), .A(n7171), .ZN(n7173) );
  INV_X1 U8962 ( .A(n7173), .ZN(P1_U3228) );
  INV_X1 U8963 ( .A(n7174), .ZN(n7177) );
  AOI22_X1 U8964 ( .A1(n9225), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9771), .ZN(n7175) );
  OAI21_X1 U8965 ( .B1(n7177), .B2(n9774), .A(n7175), .ZN(P1_U3337) );
  AOI22_X1 U8966 ( .A1(n8460), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8891), .ZN(n7176) );
  OAI21_X1 U8967 ( .B1(n7177), .B2(n8894), .A(n7176), .ZN(P2_U3342) );
  NOR2_X2 U8968 ( .A1(n8512), .A2(n8816), .ZN(n8670) );
  NOR2_X1 U8969 ( .A1(n8670), .A2(n8727), .ZN(n10038) );
  INV_X1 U8970 ( .A(n7179), .ZN(n10054) );
  AOI22_X1 U8971 ( .A1(n10054), .A2(n10021), .B1(n8665), .B2(n8435), .ZN(
        n10051) );
  OAI21_X1 U8972 ( .B1(n5009), .B2(n10041), .A(n10051), .ZN(n7180) );
  MUX2_X1 U8973 ( .A(P2_REG2_REG_0__SCAN_IN), .B(n7180), .S(n10029), .Z(n7181)
         );
  AOI21_X1 U8974 ( .B1(n8531), .B2(n10054), .A(n7181), .ZN(n7182) );
  OAI21_X1 U8975 ( .B1(n10038), .B2(n10052), .A(n7182), .ZN(P2_U3296) );
  AOI211_X1 U8976 ( .C1(n7185), .C2(n7184), .A(n7183), .B(n8481), .ZN(n7195)
         );
  AOI22_X1 U8977 ( .A1(n10009), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n7192) );
  MUX2_X1 U8978 ( .A(n5857), .B(P2_REG1_REG_2__SCAN_IN), .S(n7186), .Z(n7188)
         );
  NAND3_X1 U8979 ( .A1(n7188), .A2(n7261), .A3(n7187), .ZN(n7189) );
  NAND3_X1 U8980 ( .A1(n10007), .A2(n7190), .A3(n7189), .ZN(n7191) );
  OAI211_X1 U8981 ( .C1(n10010), .C2(n7193), .A(n7192), .B(n7191), .ZN(n7194)
         );
  OR2_X1 U8982 ( .A1(n7195), .A2(n7194), .ZN(P2_U3247) );
  AOI211_X1 U8983 ( .C1(n7198), .C2(n7197), .A(n8481), .B(n7196), .ZN(n7206)
         );
  XNOR2_X1 U8984 ( .A(n7200), .B(n7199), .ZN(n7204) );
  AND2_X1 U8985 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7585) );
  AOI21_X1 U8986 ( .B1(n10009), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n7585), .ZN(
        n7203) );
  NAND2_X1 U8987 ( .A1(n8487), .A2(n7201), .ZN(n7202) );
  OAI211_X1 U8988 ( .C1(n10011), .C2(n7204), .A(n7203), .B(n7202), .ZN(n7205)
         );
  OR2_X1 U8989 ( .A1(n7206), .A2(n7205), .ZN(P2_U3253) );
  AOI211_X1 U8990 ( .C1(n7209), .C2(n7208), .A(n8481), .B(n7207), .ZN(n7218)
         );
  XNOR2_X1 U8991 ( .A(n7211), .B(n7210), .ZN(n7216) );
  NAND2_X1 U8992 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7690) );
  INV_X1 U8993 ( .A(n7690), .ZN(n7212) );
  AOI21_X1 U8994 ( .B1(n10009), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7212), .ZN(
        n7215) );
  NAND2_X1 U8995 ( .A1(n8487), .A2(n7213), .ZN(n7214) );
  OAI211_X1 U8996 ( .C1(n7216), .C2(n10011), .A(n7215), .B(n7214), .ZN(n7217)
         );
  OR2_X1 U8997 ( .A1(n7218), .A2(n7217), .ZN(P2_U3254) );
  INV_X1 U8998 ( .A(n7219), .ZN(n7220) );
  OAI22_X1 U8999 ( .A1(n8512), .A2(n7220), .B1(n7263), .B2(n10041), .ZN(n7221)
         );
  AOI21_X1 U9000 ( .B1(n10031), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7221), .ZN(
        n7226) );
  INV_X1 U9001 ( .A(n7222), .ZN(n7224) );
  AOI22_X1 U9002 ( .A1(n8531), .A2(n7224), .B1(n8727), .B2(n7223), .ZN(n7225)
         );
  OAI211_X1 U9003 ( .C1(n10031), .C2(n7227), .A(n7226), .B(n7225), .ZN(
        P2_U3295) );
  NAND2_X1 U9004 ( .A1(n7004), .A2(n7228), .ZN(n10024) );
  NAND2_X1 U9005 ( .A1(n10024), .A2(n10023), .ZN(n10026) );
  INV_X1 U9006 ( .A(n7235), .ZN(n7230) );
  NAND3_X1 U9007 ( .A1(n10026), .A2(n7230), .A3(n7229), .ZN(n7232) );
  NAND2_X1 U9008 ( .A1(n7232), .A2(n7231), .ZN(n10066) );
  INV_X1 U9009 ( .A(n10066), .ZN(n7244) );
  NAND2_X1 U9010 ( .A1(n7233), .A2(n7234), .ZN(n7236) );
  XNOR2_X1 U9011 ( .A(n7236), .B(n7235), .ZN(n7237) );
  INV_X1 U9012 ( .A(n10021), .ZN(n8673) );
  OAI222_X1 U9013 ( .A1(n8336), .A2(n4636), .B1(n8563), .B2(n7248), .C1(n7237), 
        .C2(n8673), .ZN(n10064) );
  NAND2_X1 U9014 ( .A1(n10064), .A2(n10029), .ZN(n7243) );
  OAI211_X1 U9015 ( .C1(n4392), .C2(n10063), .A(n8861), .B(n7238), .ZN(n10062)
         );
  NOR2_X1 U9016 ( .A1(n8512), .A2(n10062), .ZN(n7241) );
  OAI22_X1 U9017 ( .A1(n10029), .A2(n7239), .B1(n7250), .B2(n10041), .ZN(n7240) );
  AOI211_X1 U9018 ( .C1(n8727), .C2(n4278), .A(n7241), .B(n7240), .ZN(n7242)
         );
  OAI211_X1 U9019 ( .C1(n7244), .C2(n8734), .A(n7243), .B(n7242), .ZN(P2_U3292) );
  OAI21_X1 U9020 ( .B1(n7247), .B2(n7246), .A(n7245), .ZN(n7253) );
  OAI22_X1 U9021 ( .A1(n7248), .A2(n8383), .B1(n8381), .B2(n4636), .ZN(n7252)
         );
  NAND2_X1 U9022 ( .A1(n8411), .A2(n4278), .ZN(n7249) );
  NAND2_X1 U9023 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7273) );
  OAI211_X1 U9024 ( .C1(n8409), .C2(n7250), .A(n7249), .B(n7273), .ZN(n7251)
         );
  AOI211_X1 U9025 ( .C1(n7842), .C2(n7253), .A(n7252), .B(n7251), .ZN(n7254)
         );
  INV_X1 U9026 ( .A(n7254), .ZN(P2_U3232) );
  AOI211_X1 U9027 ( .C1(n7257), .C2(n7256), .A(n7255), .B(n8481), .ZN(n7258)
         );
  INV_X1 U9028 ( .A(n7258), .ZN(n7268) );
  MUX2_X1 U9029 ( .A(n5858), .B(P2_REG1_REG_1__SCAN_IN), .S(n7259), .Z(n7260)
         );
  OAI21_X1 U9030 ( .B1(n5005), .B2(n4692), .A(n7260), .ZN(n7262) );
  AND2_X1 U9031 ( .A1(n7262), .A2(n7261), .ZN(n7266) );
  INV_X1 U9032 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7264) );
  OAI22_X1 U9033 ( .A1(n8480), .A2(n7264), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7263), .ZN(n7265) );
  AOI21_X1 U9034 ( .B1(n10007), .B2(n7266), .A(n7265), .ZN(n7267) );
  OAI211_X1 U9035 ( .C1(n10010), .C2(n7269), .A(n7268), .B(n7267), .ZN(
        P2_U3246) );
  MUX2_X1 U9036 ( .A(n5865), .B(P2_REG1_REG_4__SCAN_IN), .S(n7282), .Z(n7270)
         );
  NAND3_X1 U9037 ( .A1(n7284), .A2(n7271), .A3(n7270), .ZN(n7272) );
  NAND3_X1 U9038 ( .A1(n10007), .A2(n7326), .A3(n7272), .ZN(n7276) );
  INV_X1 U9039 ( .A(n7273), .ZN(n7274) );
  AOI21_X1 U9040 ( .B1(n10009), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n7274), .ZN(
        n7275) );
  NAND2_X1 U9041 ( .A1(n7276), .A2(n7275), .ZN(n7281) );
  AOI211_X1 U9042 ( .C1(n7279), .C2(n7278), .A(n7277), .B(n8481), .ZN(n7280)
         );
  AOI211_X1 U9043 ( .C1(n8487), .C2(n7282), .A(n7281), .B(n7280), .ZN(n7283)
         );
  INV_X1 U9044 ( .A(n7283), .ZN(P2_U3249) );
  OAI211_X1 U9045 ( .C1(n7286), .C2(n7285), .A(n10007), .B(n7284), .ZN(n7289)
         );
  AND2_X1 U9046 ( .A1(P2_U3152), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7287) );
  AOI21_X1 U9047 ( .B1(n10009), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7287), .ZN(
        n7288) );
  NAND2_X1 U9048 ( .A1(n7289), .A2(n7288), .ZN(n7294) );
  AOI211_X1 U9049 ( .C1(n7292), .C2(n7291), .A(n7290), .B(n8481), .ZN(n7293)
         );
  AOI211_X1 U9050 ( .C1(n8487), .C2(n7295), .A(n7294), .B(n7293), .ZN(n7296)
         );
  INV_X1 U9051 ( .A(n7296), .ZN(P2_U3248) );
  INV_X1 U9052 ( .A(n7297), .ZN(n7301) );
  NAND3_X1 U9053 ( .A1(n7328), .A2(n7299), .A3(n7298), .ZN(n7300) );
  NAND3_X1 U9054 ( .A1(n10007), .A2(n7301), .A3(n7300), .ZN(n7304) );
  NAND2_X1 U9055 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7349) );
  INV_X1 U9056 ( .A(n7349), .ZN(n7302) );
  AOI21_X1 U9057 ( .B1(n10009), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7302), .ZN(
        n7303) );
  NAND2_X1 U9058 ( .A1(n7304), .A2(n7303), .ZN(n7309) );
  AOI211_X1 U9059 ( .C1(n7307), .C2(n7306), .A(n8481), .B(n7305), .ZN(n7308)
         );
  AOI211_X1 U9060 ( .C1(n8487), .C2(n7310), .A(n7309), .B(n7308), .ZN(n7311)
         );
  INV_X1 U9061 ( .A(n7311), .ZN(P2_U3251) );
  XNOR2_X1 U9062 ( .A(n7313), .B(n7312), .ZN(n7316) );
  NOR2_X1 U9063 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5149), .ZN(n7314) );
  AOI21_X1 U9064 ( .B1(n10009), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7314), .ZN(
        n7315) );
  OAI21_X1 U9065 ( .B1(n10011), .B2(n7316), .A(n7315), .ZN(n7321) );
  AOI211_X1 U9066 ( .C1(n7319), .C2(n7318), .A(n8481), .B(n7317), .ZN(n7320)
         );
  AOI211_X1 U9067 ( .C1(n8487), .C2(n7322), .A(n7321), .B(n7320), .ZN(n7323)
         );
  INV_X1 U9068 ( .A(n7323), .ZN(P2_U3252) );
  MUX2_X1 U9069 ( .A(n5868), .B(P2_REG1_REG_5__SCAN_IN), .S(n7336), .Z(n7324)
         );
  NAND3_X1 U9070 ( .A1(n7326), .A2(n7325), .A3(n7324), .ZN(n7327) );
  NAND3_X1 U9071 ( .A1(n10007), .A2(n7328), .A3(n7327), .ZN(n7331) );
  AND2_X1 U9072 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7329) );
  AOI21_X1 U9073 ( .B1(n10009), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7329), .ZN(
        n7330) );
  NAND2_X1 U9074 ( .A1(n7331), .A2(n7330), .ZN(n7335) );
  AOI211_X1 U9075 ( .C1(n7333), .C2(n7332), .A(n8481), .B(n4618), .ZN(n7334)
         );
  AOI211_X1 U9076 ( .C1(n8487), .C2(n7336), .A(n7335), .B(n7334), .ZN(n7337)
         );
  INV_X1 U9077 ( .A(n7337), .ZN(P2_U3250) );
  NAND2_X1 U9078 ( .A1(n7338), .A2(n7558), .ZN(n7339) );
  OAI211_X1 U9079 ( .C1(n10041), .C2(n7390), .A(n7340), .B(n7339), .ZN(n7341)
         );
  NAND2_X1 U9080 ( .A1(n7341), .A2(n10029), .ZN(n7343) );
  AOI22_X1 U9081 ( .A1(n8727), .A2(n4635), .B1(n10031), .B2(
        P2_REG2_REG_5__SCAN_IN), .ZN(n7342) );
  OAI211_X1 U9082 ( .C1(n7344), .C2(n8734), .A(n7343), .B(n7342), .ZN(P2_U3291) );
  OAI21_X1 U9083 ( .B1(n4429), .B2(n7346), .A(n7345), .ZN(n7348) );
  NAND2_X1 U9084 ( .A1(n7348), .A2(n7842), .ZN(n7353) );
  OAI21_X1 U9085 ( .B1(n8381), .B2(n7624), .A(n7349), .ZN(n7351) );
  OAI22_X1 U9086 ( .A1(n8409), .A2(n7380), .B1(n8383), .B2(n4636), .ZN(n7350)
         );
  AOI211_X1 U9087 ( .C1(n7382), .C2(n8411), .A(n7351), .B(n7350), .ZN(n7352)
         );
  NAND2_X1 U9088 ( .A1(n7353), .A2(n7352), .ZN(P2_U3241) );
  OAI21_X1 U9089 ( .B1(n7360), .B2(n7355), .A(n7354), .ZN(n7356) );
  AOI222_X1 U9090 ( .A1(n10021), .A2(n7356), .B1(n8429), .B2(n8665), .C1(n8431), .C2(n8663), .ZN(n7550) );
  NAND2_X1 U9091 ( .A1(n7358), .A2(n7357), .ZN(n7375) );
  NAND2_X1 U9092 ( .A1(n7375), .A2(n7374), .ZN(n7373) );
  NAND3_X1 U9093 ( .A1(n7373), .A2(n7360), .A3(n7359), .ZN(n7362) );
  NAND2_X1 U9094 ( .A1(n7362), .A2(n7361), .ZN(n7553) );
  OAI211_X1 U9095 ( .C1(n7377), .C2(n7549), .A(n7363), .B(n8861), .ZN(n7548)
         );
  OAI22_X1 U9096 ( .A1(n10029), .A2(n7364), .B1(n7463), .B2(n10041), .ZN(n7365) );
  AOI21_X1 U9097 ( .B1(n8727), .B2(n7466), .A(n7365), .ZN(n7366) );
  OAI21_X1 U9098 ( .B1(n8512), .B2(n7548), .A(n7366), .ZN(n7367) );
  AOI21_X1 U9099 ( .B1(n7553), .B2(n8531), .A(n7367), .ZN(n7368) );
  OAI21_X1 U9100 ( .B1(n7550), .B2(n10031), .A(n7368), .ZN(P2_U3289) );
  OAI21_X1 U9101 ( .B1(n7371), .B2(n7370), .A(n7369), .ZN(n7372) );
  AOI222_X1 U9102 ( .A1(n10021), .A2(n7372), .B1(n8430), .B2(n8665), .C1(n8432), .C2(n8663), .ZN(n10069) );
  OAI21_X1 U9103 ( .B1(n7375), .B2(n7374), .A(n7373), .ZN(n10073) );
  INV_X1 U9104 ( .A(n7376), .ZN(n7379) );
  INV_X1 U9105 ( .A(n7377), .ZN(n7378) );
  OAI211_X1 U9106 ( .C1(n10071), .C2(n7379), .A(n7378), .B(n8861), .ZN(n10068)
         );
  OAI22_X1 U9107 ( .A1(n10029), .A2(n5132), .B1(n7380), .B2(n10041), .ZN(n7381) );
  AOI21_X1 U9108 ( .B1(n8727), .B2(n7382), .A(n7381), .ZN(n7383) );
  OAI21_X1 U9109 ( .B1(n8512), .B2(n10068), .A(n7383), .ZN(n7384) );
  AOI21_X1 U9110 ( .B1(n10073), .B2(n8531), .A(n7384), .ZN(n7385) );
  OAI21_X1 U9111 ( .B1(n10069), .B2(n10031), .A(n7385), .ZN(P2_U3290) );
  INV_X1 U9112 ( .A(n7386), .ZN(n7389) );
  OAI222_X1 U9113 ( .A1(n8904), .A2(n7387), .B1(n8894), .B2(n7389), .C1(n8473), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U9114 ( .A(n9229), .ZN(n9870) );
  OAI222_X1 U9115 ( .A1(P1_U3084), .A2(n9870), .B1(n9774), .B2(n7389), .C1(
        n7388), .C2(n7832), .ZN(P1_U3336) );
  INV_X1 U9116 ( .A(n7390), .ZN(n7400) );
  AOI22_X1 U9117 ( .A1(n8407), .A2(n7391), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n7392) );
  OAI21_X1 U9118 ( .B1(n7393), .B2(n8300), .A(n7392), .ZN(n7399) );
  INV_X1 U9119 ( .A(n7394), .ZN(n7395) );
  AOI211_X1 U9120 ( .C1(n7397), .C2(n7396), .A(n8413), .B(n7395), .ZN(n7398)
         );
  AOI211_X1 U9121 ( .C1(n8389), .C2(n7400), .A(n7399), .B(n7398), .ZN(n7401)
         );
  INV_X1 U9122 ( .A(n7401), .ZN(P2_U3229) );
  NAND2_X1 U9123 ( .A1(n9138), .A2(n9836), .ZN(n7991) );
  INV_X1 U9124 ( .A(n8168), .ZN(n7604) );
  INV_X1 U9125 ( .A(n8120), .ZN(n7404) );
  OR2_X1 U9126 ( .A1(n9137), .A2(n7405), .ZN(n8124) );
  NAND2_X1 U9127 ( .A1(n9137), .A2(n7405), .ZN(n7992) );
  AND2_X1 U9128 ( .A1(n8124), .A2(n7992), .ZN(n8174) );
  NAND2_X1 U9129 ( .A1(n9907), .A2(n8174), .ZN(n7528) );
  NAND2_X1 U9130 ( .A1(n9136), .A2(n7535), .ZN(n7988) );
  AND2_X1 U9131 ( .A1(n7992), .A2(n7988), .ZN(n7998) );
  NAND2_X1 U9132 ( .A1(n7528), .A2(n7998), .ZN(n7406) );
  OR2_X1 U9133 ( .A1(n9136), .A2(n7535), .ZN(n7995) );
  NAND2_X1 U9134 ( .A1(n7406), .A2(n7995), .ZN(n7439) );
  INV_X1 U9135 ( .A(n7439), .ZN(n7407) );
  INV_X1 U9136 ( .A(n7996), .ZN(n7989) );
  NAND2_X1 U9137 ( .A1(n7407), .A2(n7996), .ZN(n7740) );
  NAND2_X1 U9138 ( .A1(n7740), .A2(n7986), .ZN(n7408) );
  OR2_X1 U9139 ( .A1(n7589), .A2(n7441), .ZN(n7987) );
  NAND2_X1 U9140 ( .A1(n7589), .A2(n7441), .ZN(n8109) );
  NAND2_X1 U9141 ( .A1(n7987), .A2(n8109), .ZN(n8176) );
  XNOR2_X1 U9142 ( .A(n7408), .B(n8176), .ZN(n7411) );
  NAND2_X1 U9143 ( .A1(n9347), .A2(n9135), .ZN(n7410) );
  OR2_X1 U9144 ( .A1(n9260), .A2(n7596), .ZN(n7409) );
  NAND2_X1 U9145 ( .A1(n7410), .A2(n7409), .ZN(n7479) );
  AOI21_X1 U9146 ( .B1(n7411), .B2(n9553), .A(n7479), .ZN(n9972) );
  AOI211_X1 U9147 ( .C1(n7589), .C2(n7415), .A(n9977), .B(n4390), .ZN(n9968)
         );
  NOR2_X1 U9148 ( .A1(n7416), .A2(n9444), .ZN(n9819) );
  NOR2_X1 U9149 ( .A1(n9899), .A2(n7413), .ZN(n7419) );
  OAI22_X1 U9150 ( .A1(n9583), .A2(n7417), .B1(n7481), .B2(n9814), .ZN(n7418)
         );
  AOI211_X1 U9151 ( .C1(n9968), .C2(n9819), .A(n7419), .B(n7418), .ZN(n7435)
         );
  OR2_X1 U9152 ( .A1(n9139), .A2(n4428), .ZN(n7421) );
  NAND2_X1 U9153 ( .A1(n7422), .A2(n7421), .ZN(n7603) );
  NAND2_X1 U9154 ( .A1(n7603), .A2(n8168), .ZN(n7424) );
  OR2_X1 U9155 ( .A1(n9138), .A2(n7612), .ZN(n7423) );
  NAND2_X1 U9156 ( .A1(n7424), .A2(n7423), .ZN(n9912) );
  NAND2_X1 U9157 ( .A1(n9912), .A2(n9913), .ZN(n7426) );
  OR2_X1 U9158 ( .A1(n9137), .A2(n9920), .ZN(n7425) );
  NAND2_X1 U9159 ( .A1(n9136), .A2(n7538), .ZN(n7437) );
  NAND2_X1 U9160 ( .A1(n7436), .A2(n7427), .ZN(n7431) );
  NAND3_X1 U9161 ( .A1(n7440), .A2(n7535), .A3(n7428), .ZN(n7429) );
  NAND2_X1 U9162 ( .A1(n7431), .A2(n7430), .ZN(n7588) );
  XNOR2_X1 U9163 ( .A(n7588), .B(n8176), .ZN(n9970) );
  AND2_X1 U9164 ( .A1(n7796), .A2(n7432), .ZN(n7433) );
  INV_X1 U9165 ( .A(n9585), .ZN(n9914) );
  NAND2_X1 U9166 ( .A1(n9970), .A2(n9914), .ZN(n7434) );
  OAI211_X1 U9167 ( .C1(n9972), .C2(n9925), .A(n7435), .B(n7434), .ZN(P1_U3284) );
  XNOR2_X1 U9168 ( .A(n7538), .B(n9136), .ZN(n8171) );
  OR2_X1 U9169 ( .A1(n7436), .A2(n8171), .ZN(n9955) );
  NAND2_X1 U9170 ( .A1(n9955), .A2(n7437), .ZN(n7438) );
  XNOR2_X1 U9171 ( .A(n7440), .B(n7438), .ZN(n9961) );
  INV_X1 U9172 ( .A(n7440), .ZN(n8172) );
  XNOR2_X1 U9173 ( .A(n7439), .B(n8172), .ZN(n7443) );
  INV_X1 U9174 ( .A(n7441), .ZN(n9134) );
  AOI22_X1 U9175 ( .A1(n9116), .A2(n9134), .B1(n9347), .B2(n9136), .ZN(n7576)
         );
  INV_X1 U9176 ( .A(n7576), .ZN(n7442) );
  AOI21_X1 U9177 ( .B1(n7443), .B2(n9553), .A(n7442), .ZN(n9964) );
  MUX2_X1 U9178 ( .A(n7444), .B(n9964), .S(n9583), .Z(n7448) );
  XNOR2_X1 U9179 ( .A(n7533), .B(n7562), .ZN(n9962) );
  OAI22_X1 U9180 ( .A1(n9899), .A2(n7445), .B1(n9814), .B2(n7574), .ZN(n7446)
         );
  AOI21_X1 U9181 ( .B1(n9919), .B2(n9962), .A(n7446), .ZN(n7447) );
  OAI211_X1 U9182 ( .C1(n9585), .C2(n9961), .A(n7448), .B(n7447), .ZN(P1_U3285) );
  OAI22_X1 U9183 ( .A1(n9814), .A2(n7450), .B1(n9444), .B2(n7449), .ZN(n7452)
         );
  AOI211_X1 U9184 ( .C1(n9895), .C2(n7456), .A(n7452), .B(n7451), .ZN(n7458)
         );
  INV_X1 U9185 ( .A(n9566), .ZN(n9904) );
  OAI22_X1 U9186 ( .A1(n7454), .A2(n9899), .B1(n9583), .B2(n7453), .ZN(n7455)
         );
  AOI21_X1 U9187 ( .B1(n9904), .B2(n7456), .A(n7455), .ZN(n7457) );
  OAI21_X1 U9188 ( .B1(n7458), .B2(n9603), .A(n7457), .ZN(P1_U3290) );
  OAI211_X1 U9189 ( .C1(n7461), .C2(n7460), .A(n7459), .B(n7842), .ZN(n7468)
         );
  OAI22_X1 U9190 ( .A1(n8381), .A2(n7691), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5149), .ZN(n7465) );
  OAI22_X1 U9191 ( .A1(n8409), .A2(n7463), .B1(n8383), .B2(n7462), .ZN(n7464)
         );
  AOI211_X1 U9192 ( .C1(n7466), .C2(n8411), .A(n7465), .B(n7464), .ZN(n7467)
         );
  NAND2_X1 U9193 ( .A1(n7468), .A2(n7467), .ZN(P2_U3215) );
  INV_X1 U9194 ( .A(n8512), .ZN(n8731) );
  AOI22_X1 U9195 ( .A1(n8731), .A2(n7469), .B1(n8678), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7470) );
  OAI21_X1 U9196 ( .B1(n5896), .B2(n10029), .A(n7470), .ZN(n7474) );
  OAI22_X1 U9197 ( .A1(n8681), .A2(n7472), .B1(n7471), .B2(n10031), .ZN(n7473)
         );
  AOI211_X1 U9198 ( .C1(n8531), .C2(n7475), .A(n7474), .B(n7473), .ZN(n7476)
         );
  INV_X1 U9199 ( .A(n7476), .ZN(P2_U3294) );
  XOR2_X1 U9200 ( .A(n7478), .B(n7477), .Z(n7484) );
  NOR2_X1 U9201 ( .A1(n9617), .A2(n7413), .ZN(n9969) );
  AOI22_X1 U9202 ( .A1(n7479), .A2(n9832), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3084), .ZN(n7480) );
  OAI21_X1 U9203 ( .B1(n9842), .B2(n7481), .A(n7480), .ZN(n7482) );
  AOI21_X1 U9204 ( .B1(n9837), .B2(n9969), .A(n7482), .ZN(n7483) );
  OAI21_X1 U9205 ( .B1(n7484), .B2(n9110), .A(n7483), .ZN(P1_U3211) );
  INV_X1 U9206 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7487) );
  INV_X1 U9207 ( .A(n7485), .ZN(n7488) );
  OAI222_X1 U9208 ( .A1(n8904), .A2(n7487), .B1(n8894), .B2(n7488), .C1(
        P2_U3152), .C2(n7486), .ZN(P2_U3340) );
  INV_X1 U9209 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7489) );
  INV_X1 U9210 ( .A(n9237), .ZN(n9246) );
  OAI222_X1 U9211 ( .A1(n7832), .A2(n7489), .B1(n9774), .B2(n7488), .C1(
        P1_U3084), .C2(n9246), .ZN(P1_U3335) );
  AOI211_X1 U9212 ( .C1(n7492), .C2(n7491), .A(n8481), .B(n7490), .ZN(n7500)
         );
  XNOR2_X1 U9213 ( .A(n7494), .B(n7493), .ZN(n7498) );
  AND2_X1 U9214 ( .A1(P2_U3152), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7770) );
  AOI21_X1 U9215 ( .B1(n10009), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7770), .ZN(
        n7497) );
  NAND2_X1 U9216 ( .A1(n8487), .A2(n7495), .ZN(n7496) );
  OAI211_X1 U9217 ( .C1(n7498), .C2(n10011), .A(n7497), .B(n7496), .ZN(n7499)
         );
  OR2_X1 U9218 ( .A1(n7500), .A2(n7499), .ZN(P2_U3255) );
  INV_X1 U9219 ( .A(n7501), .ZN(n7504) );
  XNOR2_X1 U9220 ( .A(n7502), .B(n7563), .ZN(n7503) );
  NOR2_X1 U9221 ( .A1(n7503), .A2(n7504), .ZN(n7566) );
  AOI21_X1 U9222 ( .B1(n7504), .B2(n7503), .A(n7566), .ZN(n7512) );
  INV_X1 U9223 ( .A(n7532), .ZN(n7510) );
  NAND2_X1 U9224 ( .A1(n9726), .A2(n7538), .ZN(n9958) );
  NAND2_X1 U9225 ( .A1(n9347), .A2(n9137), .ZN(n7507) );
  OR2_X1 U9226 ( .A1(n9260), .A2(n7505), .ZN(n7506) );
  NAND2_X1 U9227 ( .A1(n7507), .A2(n7506), .ZN(n7530) );
  AOI22_X1 U9228 ( .A1(n7530), .A2(n9832), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3084), .ZN(n7508) );
  OAI21_X1 U9229 ( .B1(n8938), .B2(n9958), .A(n7508), .ZN(n7509) );
  AOI21_X1 U9230 ( .B1(n7510), .B2(n9104), .A(n7509), .ZN(n7511) );
  OAI21_X1 U9231 ( .B1(n7512), .B2(n9110), .A(n7511), .ZN(P1_U3225) );
  XNOR2_X1 U9232 ( .A(n9209), .B(n9210), .ZN(n7516) );
  AOI21_X1 U9233 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7516), .A(n9211), .ZN(
        n7527) );
  NAND2_X1 U9234 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7517) );
  OAI21_X1 U9235 ( .B1(n9871), .B2(n9200), .A(n7517), .ZN(n7525) );
  INV_X1 U9236 ( .A(n7518), .ZN(n7519) );
  NOR2_X1 U9237 ( .A1(n7520), .A2(n7519), .ZN(n7522) );
  XNOR2_X1 U9238 ( .A(n9210), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7521) );
  AOI21_X1 U9239 ( .B1(n7522), .B2(n7521), .A(n9199), .ZN(n7523) );
  NOR2_X1 U9240 ( .A1(n7523), .A2(n9249), .ZN(n7524) );
  AOI211_X1 U9241 ( .C1(n9874), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7525), .B(
        n7524), .ZN(n7526) );
  OAI21_X1 U9242 ( .B1(n7527), .B2(n9850), .A(n7526), .ZN(P1_U3255) );
  NAND2_X1 U9243 ( .A1(n7528), .A2(n7992), .ZN(n7529) );
  XOR2_X1 U9244 ( .A(n8171), .B(n7529), .Z(n7531) );
  AOI21_X1 U9245 ( .B1(n7531), .B2(n9553), .A(n7530), .ZN(n9959) );
  OAI22_X1 U9246 ( .A1(n9583), .A2(n6095), .B1(n7532), .B2(n9814), .ZN(n7537)
         );
  INV_X1 U9247 ( .A(n9819), .ZN(n7801) );
  INV_X1 U9248 ( .A(n7533), .ZN(n7534) );
  OAI211_X1 U9249 ( .C1(n7535), .C2(n9916), .A(n7534), .B(n9986), .ZN(n9957)
         );
  NOR2_X1 U9250 ( .A1(n7801), .A2(n9957), .ZN(n7536) );
  AOI211_X1 U9251 ( .C1(n9921), .C2(n7538), .A(n7537), .B(n7536), .ZN(n7540)
         );
  NAND2_X1 U9252 ( .A1(n7436), .A2(n8171), .ZN(n9954) );
  NAND3_X1 U9253 ( .A1(n9955), .A2(n9954), .A3(n9914), .ZN(n7539) );
  OAI211_X1 U9254 ( .C1(n9959), .C2(n9925), .A(n7540), .B(n7539), .ZN(P1_U3286) );
  OAI21_X1 U9255 ( .B1(n9919), .B2(n9921), .A(n7541), .ZN(n7546) );
  OAI22_X1 U9256 ( .A1(n9603), .A2(n7543), .B1(n7542), .B2(n9814), .ZN(n7544)
         );
  INV_X1 U9257 ( .A(n7544), .ZN(n7545) );
  OAI211_X1 U9258 ( .C1(n7547), .C2(n9583), .A(n7546), .B(n7545), .ZN(P1_U3291) );
  OAI21_X1 U9259 ( .B1(n7549), .B2(n10070), .A(n7548), .ZN(n7552) );
  INV_X1 U9260 ( .A(n7550), .ZN(n7551) );
  AOI211_X1 U9261 ( .C1(n10074), .C2(n7553), .A(n7552), .B(n7551), .ZN(n7556)
         );
  NAND2_X1 U9262 ( .A1(n10075), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7554) );
  OAI21_X1 U9263 ( .B1(n7556), .B2(n10075), .A(n7554), .ZN(P2_U3472) );
  NAND2_X1 U9264 ( .A1(n10080), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7555) );
  OAI21_X1 U9265 ( .B1(n7556), .B2(n10080), .A(n7555), .ZN(P2_U3527) );
  INV_X1 U9266 ( .A(n7557), .ZN(n7560) );
  OAI222_X1 U9267 ( .A1(n8904), .A2(n7559), .B1(n8894), .B2(n7560), .C1(n7558), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U9268 ( .A1(n7561), .A2(n7832), .B1(P1_U3084), .B2(n9471), .C1(
        n9774), .C2(n7560), .ZN(P1_U3334) );
  NAND2_X1 U9269 ( .A1(n9726), .A2(n7562), .ZN(n9963) );
  AND2_X1 U9270 ( .A1(n7502), .A2(n7563), .ZN(n7567) );
  XNOR2_X1 U9271 ( .A(n7565), .B(n7564), .ZN(n7568) );
  NOR3_X1 U9272 ( .A1(n7566), .A2(n7567), .A3(n7568), .ZN(n7573) );
  INV_X1 U9273 ( .A(n7566), .ZN(n7571) );
  INV_X1 U9274 ( .A(n7567), .ZN(n7570) );
  INV_X1 U9275 ( .A(n7568), .ZN(n7569) );
  AOI21_X1 U9276 ( .B1(n7571), .B2(n7570), .A(n7569), .ZN(n7572) );
  OAI21_X1 U9277 ( .B1(n7573), .B2(n7572), .A(n9838), .ZN(n7580) );
  INV_X1 U9278 ( .A(n7574), .ZN(n7578) );
  OAI22_X1 U9279 ( .A1(n7576), .A2(n9106), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7575), .ZN(n7577) );
  AOI21_X1 U9280 ( .B1(n7578), .B2(n9104), .A(n7577), .ZN(n7579) );
  OAI211_X1 U9281 ( .C1(n8938), .C2(n9963), .A(n7580), .B(n7579), .ZN(P1_U3237) );
  INV_X1 U9282 ( .A(n8860), .ZN(n7631) );
  OAI211_X1 U9283 ( .C1(n7583), .C2(n7582), .A(n7581), .B(n7842), .ZN(n7587)
         );
  OAI22_X1 U9284 ( .A1(n8409), .A2(n7630), .B1(n8383), .B2(n7624), .ZN(n7584)
         );
  AOI211_X1 U9285 ( .C1(n7771), .C2(n8428), .A(n7585), .B(n7584), .ZN(n7586)
         );
  OAI211_X1 U9286 ( .C1(n7631), .C2(n8300), .A(n7587), .B(n7586), .ZN(P2_U3223) );
  NAND2_X1 U9287 ( .A1(n7588), .A2(n8176), .ZN(n7591) );
  OR2_X1 U9288 ( .A1(n7589), .A2(n9134), .ZN(n7590) );
  INV_X1 U9289 ( .A(n7596), .ZN(n9133) );
  NAND2_X1 U9290 ( .A1(n7653), .A2(n9133), .ZN(n7592) );
  OR2_X1 U9291 ( .A1(n7749), .A2(n7778), .ZN(n9805) );
  NAND2_X1 U9292 ( .A1(n7749), .A2(n7778), .ZN(n9806) );
  NAND2_X1 U9293 ( .A1(n9805), .A2(n9806), .ZN(n8177) );
  XNOR2_X1 U9294 ( .A(n7593), .B(n8177), .ZN(n9990) );
  AND2_X1 U9295 ( .A1(n7986), .A2(n7987), .ZN(n7594) );
  AND2_X1 U9296 ( .A1(n7594), .A2(n7978), .ZN(n7738) );
  NAND2_X1 U9297 ( .A1(n7740), .A2(n7738), .ZN(n7595) );
  INV_X1 U9298 ( .A(n7978), .ZN(n8004) );
  AND2_X1 U9299 ( .A1(n7595), .A2(n7735), .ZN(n9808) );
  XNOR2_X1 U9300 ( .A(n9808), .B(n8177), .ZN(n7597) );
  OAI22_X1 U9301 ( .A1(n9102), .A2(n7596), .B1(n7744), .B2(n9260), .ZN(n7719)
         );
  AOI21_X1 U9302 ( .B1(n7597), .B2(n9553), .A(n7719), .ZN(n9989) );
  MUX2_X1 U9303 ( .A(n7598), .B(n9989), .S(n9583), .Z(n7602) );
  AND2_X1 U9304 ( .A1(n9901), .A2(n7749), .ZN(n7599) );
  NOR2_X1 U9305 ( .A1(n9816), .A2(n7599), .ZN(n9987) );
  OAI22_X1 U9306 ( .A1(n9899), .A2(n4652), .B1(n9814), .B2(n7721), .ZN(n7600)
         );
  AOI21_X1 U9307 ( .B1(n9987), .B2(n9919), .A(n7600), .ZN(n7601) );
  OAI211_X1 U9308 ( .C1(n9585), .C2(n9990), .A(n7602), .B(n7601), .ZN(P1_U3282) );
  XNOR2_X1 U9309 ( .A(n7603), .B(n7604), .ZN(n7610) );
  INV_X1 U9310 ( .A(n7610), .ZN(n9947) );
  XNOR2_X1 U9311 ( .A(n7994), .B(n7604), .ZN(n7605) );
  NAND2_X1 U9312 ( .A1(n7605), .A2(n9553), .ZN(n7609) );
  NAND2_X1 U9313 ( .A1(n9347), .A2(n9139), .ZN(n7608) );
  OR2_X1 U9314 ( .A1(n9260), .A2(n7606), .ZN(n7607) );
  AND2_X1 U9315 ( .A1(n7608), .A2(n7607), .ZN(n9831) );
  OAI211_X1 U9316 ( .C1(n7610), .C2(n7796), .A(n7609), .B(n9831), .ZN(n9945)
         );
  MUX2_X1 U9317 ( .A(n9945), .B(P1_REG2_REG_3__SCAN_IN), .S(n9925), .Z(n7615)
         );
  XNOR2_X1 U9318 ( .A(n7611), .B(n7612), .ZN(n9944) );
  INV_X1 U9319 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U9320 ( .A1(n9921), .A2(n7612), .B1(n10198), .B2(n9924), .ZN(n7613)
         );
  OAI21_X1 U9321 ( .B1(n9527), .B2(n9944), .A(n7613), .ZN(n7614) );
  AOI211_X1 U9322 ( .C1(n9904), .C2(n9947), .A(n7615), .B(n7614), .ZN(n7616)
         );
  INV_X1 U9323 ( .A(n7616), .ZN(P1_U3288) );
  OAI21_X1 U9324 ( .B1(n7618), .B2(n5580), .A(n7617), .ZN(n8865) );
  INV_X1 U9325 ( .A(n7619), .ZN(n7620) );
  NAND2_X1 U9326 ( .A1(n10029), .A2(n7620), .ZN(n8702) );
  OAI21_X1 U9327 ( .B1(n7623), .B2(n7622), .A(n7621), .ZN(n7627) );
  OAI22_X1 U9328 ( .A1(n7624), .A2(n8563), .B1(n7767), .B2(n8336), .ZN(n7626)
         );
  NOR2_X1 U9329 ( .A1(n8865), .A2(n8693), .ZN(n7625) );
  AOI211_X1 U9330 ( .C1(n10021), .C2(n7627), .A(n7626), .B(n7625), .ZN(n8864)
         );
  MUX2_X1 U9331 ( .A(n7628), .B(n8864), .S(n10029), .Z(n7634) );
  INV_X1 U9332 ( .A(n7673), .ZN(n7629) );
  AOI21_X1 U9333 ( .B1(n8860), .B2(n7363), .A(n7629), .ZN(n8862) );
  OAI22_X1 U9334 ( .A1(n8681), .A2(n7631), .B1(n7630), .B2(n10041), .ZN(n7632)
         );
  AOI21_X1 U9335 ( .B1(n8862), .B2(n8670), .A(n7632), .ZN(n7633) );
  OAI211_X1 U9336 ( .C1(n8865), .C2(n8702), .A(n7634), .B(n7633), .ZN(P2_U3288) );
  XNOR2_X1 U9337 ( .A(n7636), .B(n7635), .ZN(n7646) );
  OAI21_X1 U9338 ( .B1(n7639), .B2(n7638), .A(n7637), .ZN(n7640) );
  NAND2_X1 U9339 ( .A1(n7640), .A2(n10008), .ZN(n7645) );
  NOR2_X1 U9340 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7846), .ZN(n7643) );
  NOR2_X1 U9341 ( .A1(n10010), .A2(n7641), .ZN(n7642) );
  AOI211_X1 U9342 ( .C1(n10009), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7643), .B(
        n7642), .ZN(n7644) );
  OAI211_X1 U9343 ( .C1(n7646), .C2(n10011), .A(n7645), .B(n7644), .ZN(
        P2_U3256) );
  INV_X1 U9344 ( .A(n7647), .ZN(n7661) );
  OAI222_X1 U9345 ( .A1(n7832), .A2(n7648), .B1(n9774), .B2(n7661), .C1(n8101), 
        .C2(P1_U3084), .ZN(P1_U3333) );
  NAND2_X1 U9346 ( .A1(n7650), .A2(n7649), .ZN(n7651) );
  XOR2_X1 U9347 ( .A(n7652), .B(n7651), .Z(n7660) );
  INV_X1 U9348 ( .A(n7653), .ZN(n9902) );
  NOR2_X1 U9349 ( .A1(n9902), .A2(n9617), .ZN(n9975) );
  NAND2_X1 U9350 ( .A1(n9347), .A2(n9134), .ZN(n7655) );
  OR2_X1 U9351 ( .A1(n9260), .A2(n7778), .ZN(n7654) );
  NAND2_X1 U9352 ( .A1(n7655), .A2(n7654), .ZN(n9894) );
  NOR2_X1 U9353 ( .A1(n7656), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9158) );
  AOI21_X1 U9354 ( .B1(n9894), .B2(n9832), .A(n9158), .ZN(n7657) );
  OAI21_X1 U9355 ( .B1(n9842), .B2(n9896), .A(n7657), .ZN(n7658) );
  AOI21_X1 U9356 ( .B1(n9837), .B2(n9975), .A(n7658), .ZN(n7659) );
  OAI21_X1 U9357 ( .B1(n7660), .B2(n9110), .A(n7659), .ZN(P1_U3219) );
  OAI222_X1 U9358 ( .A1(n8904), .A2(n7663), .B1(P2_U3152), .B2(n7662), .C1(
        n8894), .C2(n7661), .ZN(P2_U3338) );
  OAI21_X1 U9359 ( .B1(n7669), .B2(n7665), .A(n7664), .ZN(n7672) );
  OAI22_X1 U9360 ( .A1(n7691), .A2(n8563), .B1(n7847), .B2(n8336), .ZN(n7671)
         );
  INV_X1 U9361 ( .A(n7666), .ZN(n7667) );
  AOI21_X1 U9362 ( .B1(n7669), .B2(n7668), .A(n7667), .ZN(n8859) );
  NOR2_X1 U9363 ( .A1(n8859), .A2(n8693), .ZN(n7670) );
  AOI211_X1 U9364 ( .C1(n10021), .C2(n7672), .A(n7671), .B(n7670), .ZN(n8858)
         );
  AOI21_X1 U9365 ( .B1(n8855), .B2(n7673), .A(n7709), .ZN(n8856) );
  INV_X1 U9366 ( .A(n8855), .ZN(n7676) );
  INV_X1 U9367 ( .A(n7692), .ZN(n7674) );
  AOI22_X1 U9368 ( .A1(n10031), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7674), .B2(
        n8678), .ZN(n7675) );
  OAI21_X1 U9369 ( .B1(n8681), .B2(n7676), .A(n7675), .ZN(n7678) );
  NOR2_X1 U9370 ( .A1(n8859), .A2(n8702), .ZN(n7677) );
  AOI211_X1 U9371 ( .C1(n8856), .C2(n8670), .A(n7678), .B(n7677), .ZN(n7679)
         );
  OAI21_X1 U9372 ( .B1(n8858), .B2(n10031), .A(n7679), .ZN(P2_U3287) );
  INV_X1 U9373 ( .A(n7680), .ZN(n7683) );
  OAI222_X1 U9374 ( .A1(n7832), .A2(n7682), .B1(n9774), .B2(n7683), .C1(n7681), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  OAI222_X1 U9375 ( .A1(n8904), .A2(n7685), .B1(P2_U3152), .B2(n7684), .C1(
        n8894), .C2(n7683), .ZN(P2_U3337) );
  INV_X1 U9376 ( .A(n7686), .ZN(n7687) );
  AOI21_X1 U9377 ( .B1(n7689), .B2(n7688), .A(n7687), .ZN(n7696) );
  OAI21_X1 U9378 ( .B1(n8381), .B2(n7847), .A(n7690), .ZN(n7694) );
  OAI22_X1 U9379 ( .A1(n8409), .A2(n7692), .B1(n8383), .B2(n7691), .ZN(n7693)
         );
  AOI211_X1 U9380 ( .C1(n8855), .C2(n8411), .A(n7694), .B(n7693), .ZN(n7695)
         );
  OAI21_X1 U9381 ( .B1(n7696), .B2(n8413), .A(n7695), .ZN(P2_U3233) );
  OAI21_X1 U9382 ( .B1(n7699), .B2(n7698), .A(n7697), .ZN(n7706) );
  OAI22_X1 U9383 ( .A1(n7767), .A2(n8563), .B1(n7908), .B2(n8336), .ZN(n7705)
         );
  AND2_X1 U9384 ( .A1(n7666), .A2(n7700), .ZN(n7703) );
  OAI21_X1 U9385 ( .B1(n7703), .B2(n7702), .A(n7701), .ZN(n8854) );
  NOR2_X1 U9386 ( .A1(n8854), .A2(n8693), .ZN(n7704) );
  AOI211_X1 U9387 ( .C1(n10021), .C2(n7706), .A(n7705), .B(n7704), .ZN(n8853)
         );
  OAI22_X1 U9388 ( .A1(n10029), .A2(n7707), .B1(n7768), .B2(n10041), .ZN(n7708) );
  AOI21_X1 U9389 ( .B1(n8727), .B2(n8850), .A(n7708), .ZN(n7712) );
  OR2_X1 U9390 ( .A1(n7709), .A2(n7774), .ZN(n7710) );
  AND2_X1 U9391 ( .A1(n7730), .A2(n7710), .ZN(n8851) );
  NAND2_X1 U9392 ( .A1(n8851), .A2(n8670), .ZN(n7711) );
  OAI211_X1 U9393 ( .C1(n8854), .C2(n8702), .A(n7712), .B(n7711), .ZN(n7713)
         );
  INV_X1 U9394 ( .A(n7713), .ZN(n7714) );
  OAI21_X1 U9395 ( .B1(n8853), .B2(n10031), .A(n7714), .ZN(P2_U3286) );
  INV_X1 U9396 ( .A(n7715), .ZN(n7716) );
  AOI21_X1 U9397 ( .B1(n7718), .B2(n7717), .A(n7716), .ZN(n7724) );
  AND2_X1 U9398 ( .A1(n7749), .A2(n9726), .ZN(n9985) );
  AOI22_X1 U9399 ( .A1(n7719), .A2(n9832), .B1(P1_REG3_REG_9__SCAN_IN), .B2(
        P1_U3084), .ZN(n7720) );
  OAI21_X1 U9400 ( .B1(n7721), .B2(n9842), .A(n7720), .ZN(n7722) );
  AOI21_X1 U9401 ( .B1(n9837), .B2(n9985), .A(n7722), .ZN(n7723) );
  OAI21_X1 U9402 ( .B1(n7724), .B2(n9110), .A(n7723), .ZN(P1_U3229) );
  XNOR2_X1 U9403 ( .A(n7725), .B(n7727), .ZN(n8848) );
  XOR2_X1 U9404 ( .A(n7727), .B(n7726), .Z(n7728) );
  AOI222_X1 U9405 ( .A1(n10021), .A2(n7728), .B1(n8425), .B2(n8665), .C1(n8427), .C2(n8663), .ZN(n8847) );
  MUX2_X1 U9406 ( .A(n7729), .B(n8847), .S(n10029), .Z(n7734) );
  AOI21_X1 U9407 ( .B1(n8844), .B2(n7730), .A(n4700), .ZN(n8845) );
  INV_X1 U9408 ( .A(n8844), .ZN(n7731) );
  OAI22_X1 U9409 ( .A1(n8681), .A2(n7731), .B1(n7848), .B2(n10041), .ZN(n7732)
         );
  AOI21_X1 U9410 ( .B1(n8845), .B2(n8670), .A(n7732), .ZN(n7733) );
  OAI211_X1 U9411 ( .C1(n8848), .C2(n8734), .A(n7734), .B(n7733), .ZN(P2_U3285) );
  INV_X1 U9412 ( .A(n7983), .ZN(n7737) );
  INV_X1 U9413 ( .A(n7735), .ZN(n7736) );
  AND2_X1 U9414 ( .A1(n7738), .A2(n7737), .ZN(n7739) );
  NAND2_X1 U9415 ( .A1(n7740), .A2(n7739), .ZN(n7741) );
  NAND2_X1 U9416 ( .A1(n9818), .A2(n7744), .ZN(n7984) );
  NAND2_X1 U9417 ( .A1(n7984), .A2(n9806), .ZN(n7980) );
  NAND2_X1 U9418 ( .A1(n7980), .A2(n7743), .ZN(n8106) );
  XNOR2_X1 U9419 ( .A(n9725), .B(n9130), .ZN(n8179) );
  XNOR2_X1 U9420 ( .A(n7790), .B(n8179), .ZN(n7754) );
  NAND2_X1 U9421 ( .A1(n9347), .A2(n9131), .ZN(n7746) );
  OR2_X1 U9422 ( .A1(n9260), .A2(n9056), .ZN(n7745) );
  NAND2_X1 U9423 ( .A1(n7746), .A2(n7745), .ZN(n9077) );
  INV_X1 U9424 ( .A(n7778), .ZN(n9132) );
  OR2_X1 U9425 ( .A1(n7749), .A2(n9132), .ZN(n7747) );
  NAND2_X1 U9426 ( .A1(n7749), .A2(n9132), .ZN(n7750) );
  XNOR2_X1 U9427 ( .A(n9818), .B(n9131), .ZN(n9810) );
  OR2_X1 U9428 ( .A1(n9818), .A2(n9131), .ZN(n7752) );
  XNOR2_X1 U9429 ( .A(n7784), .B(n8179), .ZN(n9730) );
  NOR2_X1 U9430 ( .A1(n9730), .A2(n7796), .ZN(n7753) );
  AOI211_X1 U9431 ( .C1(n9553), .C2(n7754), .A(n9077), .B(n7753), .ZN(n9729)
         );
  INV_X1 U9432 ( .A(n9818), .ZN(n7777) );
  INV_X1 U9433 ( .A(n7799), .ZN(n7758) );
  AOI21_X1 U9434 ( .B1(n9725), .B2(n7755), .A(n7758), .ZN(n9727) );
  INV_X1 U9435 ( .A(n9583), .ZN(n9925) );
  INV_X1 U9436 ( .A(n9079), .ZN(n7759) );
  AOI22_X1 U9437 ( .A1(n9925), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9924), .B2(
        n7759), .ZN(n7760) );
  OAI21_X1 U9438 ( .B1(n7756), .B2(n9899), .A(n7760), .ZN(n7762) );
  NOR2_X1 U9439 ( .A1(n9730), .A2(n9566), .ZN(n7761) );
  AOI211_X1 U9440 ( .C1(n9727), .C2(n9919), .A(n7762), .B(n7761), .ZN(n7763)
         );
  OAI21_X1 U9441 ( .B1(n9729), .B2(n9603), .A(n7763), .ZN(P1_U3280) );
  OAI211_X1 U9442 ( .C1(n7766), .C2(n7765), .A(n7764), .B(n7842), .ZN(n7773)
         );
  OAI22_X1 U9443 ( .A1(n8409), .A2(n7768), .B1(n8383), .B2(n7767), .ZN(n7769)
         );
  AOI211_X1 U9444 ( .C1(n7771), .C2(n8426), .A(n7770), .B(n7769), .ZN(n7772)
         );
  OAI211_X1 U9445 ( .C1(n7774), .C2(n8300), .A(n7773), .B(n7772), .ZN(P2_U3219) );
  XOR2_X1 U9446 ( .A(n7776), .B(n7775), .Z(n7782) );
  NOR2_X1 U9447 ( .A1(n7777), .A2(n9617), .ZN(n9824) );
  OAI22_X1 U9448 ( .A1(n9102), .A2(n7778), .B1(n7791), .B2(n9260), .ZN(n9823)
         );
  AOI22_X1 U9449 ( .A1(n9823), .A2(n9832), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3084), .ZN(n7779) );
  OAI21_X1 U9450 ( .B1(n9813), .B2(n9842), .A(n7779), .ZN(n7780) );
  AOI21_X1 U9451 ( .B1(n9824), .B2(n9837), .A(n7780), .ZN(n7781) );
  OAI21_X1 U9452 ( .B1(n7782), .B2(n9110), .A(n7781), .ZN(P1_U3215) );
  NAND2_X1 U9453 ( .A1(n9725), .A2(n9130), .ZN(n7783) );
  OR2_X1 U9454 ( .A1(n9725), .A2(n9130), .ZN(n7785) );
  NAND2_X1 U9455 ( .A1(n9717), .A2(n9056), .ZN(n8015) );
  NAND2_X1 U9456 ( .A1(n8016), .A2(n8015), .ZN(n7792) );
  NAND2_X1 U9457 ( .A1(n7786), .A2(n8181), .ZN(n7787) );
  NAND2_X1 U9458 ( .A1(n9272), .A2(n7787), .ZN(n9720) );
  NAND2_X1 U9459 ( .A1(n9347), .A2(n9130), .ZN(n7789) );
  OR2_X1 U9460 ( .A1(n8008), .A2(n9260), .ZN(n7788) );
  AND2_X1 U9461 ( .A1(n7789), .A2(n7788), .ZN(n9003) );
  NAND2_X1 U9462 ( .A1(n9725), .A2(n7791), .ZN(n8006) );
  NAND2_X1 U9463 ( .A1(n7793), .A2(n7792), .ZN(n7794) );
  NAND3_X1 U9464 ( .A1(n9313), .A2(n9553), .A3(n7794), .ZN(n7795) );
  OAI211_X1 U9465 ( .C1(n9720), .C2(n7796), .A(n9003), .B(n7795), .ZN(n9722)
         );
  NAND2_X1 U9466 ( .A1(n9722), .A2(n9583), .ZN(n7805) );
  OAI22_X1 U9467 ( .A1(n9583), .A2(n7797), .B1(n9006), .B2(n9814), .ZN(n7803)
         );
  NAND2_X1 U9468 ( .A1(n7799), .A2(n9717), .ZN(n7798) );
  NAND2_X1 U9469 ( .A1(n7798), .A2(n9986), .ZN(n7800) );
  NOR2_X2 U9470 ( .A1(n7799), .A2(n9717), .ZN(n9593) );
  OR2_X1 U9471 ( .A1(n7800), .A2(n9593), .ZN(n9718) );
  NOR2_X1 U9472 ( .A1(n9718), .A2(n7801), .ZN(n7802) );
  AOI211_X1 U9473 ( .C1(n9921), .C2(n9717), .A(n7803), .B(n7802), .ZN(n7804)
         );
  OAI211_X1 U9474 ( .C1(n9720), .C2(n9566), .A(n7805), .B(n7804), .ZN(P1_U3279) );
  XOR2_X1 U9475 ( .A(n7806), .B(n7812), .Z(n7807) );
  AOI222_X1 U9476 ( .A1(n10021), .A2(n7807), .B1(n8424), .B2(n8665), .C1(n8426), .C2(n8663), .ZN(n8842) );
  AOI211_X1 U9477 ( .C1(n8839), .C2(n7808), .A(n8816), .B(n7861), .ZN(n8838)
         );
  INV_X1 U9478 ( .A(n8839), .ZN(n7811) );
  INV_X1 U9479 ( .A(n7909), .ZN(n7809) );
  AOI22_X1 U9480 ( .A1(n10031), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7809), .B2(
        n8678), .ZN(n7810) );
  OAI21_X1 U9481 ( .B1(n7811), .B2(n8681), .A(n7810), .ZN(n7815) );
  XOR2_X1 U9482 ( .A(n7813), .B(n7812), .Z(n8843) );
  NOR2_X1 U9483 ( .A1(n8843), .A2(n8734), .ZN(n7814) );
  AOI211_X1 U9484 ( .C1(n8838), .C2(n8731), .A(n7815), .B(n7814), .ZN(n7816)
         );
  OAI21_X1 U9485 ( .B1(n10031), .B2(n8842), .A(n7816), .ZN(P2_U3284) );
  AOI21_X1 U9486 ( .B1(n7819), .B2(n7818), .A(n7817), .ZN(n7829) );
  AOI211_X1 U9487 ( .C1(n7822), .C2(n7821), .A(n7820), .B(n8481), .ZN(n7823)
         );
  INV_X1 U9488 ( .A(n7823), .ZN(n7828) );
  INV_X1 U9489 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U9490 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7907) );
  OAI21_X1 U9491 ( .B1(n8480), .B2(n7824), .A(n7907), .ZN(n7825) );
  AOI21_X1 U9492 ( .B1(n8487), .B2(n7826), .A(n7825), .ZN(n7827) );
  OAI211_X1 U9493 ( .C1(n7829), .C2(n10011), .A(n7828), .B(n7827), .ZN(
        P2_U3257) );
  INV_X1 U9494 ( .A(n7830), .ZN(n7834) );
  OAI222_X1 U9495 ( .A1(n7832), .A2(n7831), .B1(n9774), .B2(n7834), .C1(
        P1_U3084), .C2(n6479), .ZN(P1_U3331) );
  OAI222_X1 U9496 ( .A1(n8904), .A2(n7835), .B1(n8894), .B2(n7834), .C1(n7833), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9497 ( .A(n7836), .ZN(n7841) );
  OR2_X1 U9498 ( .A1(n7837), .A2(P1_U3084), .ZN(n8217) );
  INV_X1 U9499 ( .A(n8217), .ZN(n8231) );
  AOI21_X1 U9500 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9771), .A(n8231), .ZN(
        n7838) );
  OAI21_X1 U9501 ( .B1(n7841), .B2(n9774), .A(n7838), .ZN(P1_U3330) );
  AOI21_X1 U9502 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8891), .A(n7839), .ZN(
        n7840) );
  OAI21_X1 U9503 ( .B1(n7841), .B2(n8894), .A(n7840), .ZN(P2_U3335) );
  OAI211_X1 U9504 ( .C1(n7845), .C2(n7844), .A(n7843), .B(n7842), .ZN(n7852)
         );
  OAI22_X1 U9505 ( .A1(n8381), .A2(n7919), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7846), .ZN(n7850) );
  OAI22_X1 U9506 ( .A1(n8409), .A2(n7848), .B1(n8383), .B2(n7847), .ZN(n7849)
         );
  AOI211_X1 U9507 ( .C1(n8844), .C2(n8411), .A(n7850), .B(n7849), .ZN(n7851)
         );
  NAND2_X1 U9508 ( .A1(n7852), .A2(n7851), .ZN(P2_U3238) );
  OAI21_X1 U9509 ( .B1(n7854), .B2(n7853), .A(n7891), .ZN(n7860) );
  OAI22_X1 U9510 ( .A1(n7919), .A2(n8563), .B1(n8404), .B2(n8336), .ZN(n7859)
         );
  NAND2_X1 U9511 ( .A1(n7855), .A2(n7854), .ZN(n7856) );
  NAND2_X1 U9512 ( .A1(n7857), .A2(n7856), .ZN(n8837) );
  NOR2_X1 U9513 ( .A1(n8837), .A2(n8693), .ZN(n7858) );
  AOI211_X1 U9514 ( .C1(n10021), .C2(n7860), .A(n7859), .B(n7858), .ZN(n8836)
         );
  INV_X1 U9515 ( .A(n7861), .ZN(n7863) );
  AOI21_X1 U9516 ( .B1(n8833), .B2(n7863), .A(n7862), .ZN(n8834) );
  INV_X1 U9517 ( .A(n7920), .ZN(n7864) );
  AOI22_X1 U9518 ( .A1(n10031), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7864), .B2(
        n8678), .ZN(n7865) );
  OAI21_X1 U9519 ( .B1(n7866), .B2(n8681), .A(n7865), .ZN(n7868) );
  NOR2_X1 U9520 ( .A1(n8837), .A2(n8702), .ZN(n7867) );
  AOI211_X1 U9521 ( .C1(n8834), .C2(n8670), .A(n7868), .B(n7867), .ZN(n7869)
         );
  OAI21_X1 U9522 ( .B1(n8836), .B2(n10031), .A(n7869), .ZN(P2_U3283) );
  INV_X1 U9523 ( .A(n7870), .ZN(n7883) );
  OAI21_X1 U9524 ( .B1(n7873), .B2(n7872), .A(n7871), .ZN(n7874) );
  NAND2_X1 U9525 ( .A1(n10008), .A2(n7874), .ZN(n7882) );
  OAI21_X1 U9526 ( .B1(n7877), .B2(n7876), .A(n7875), .ZN(n7880) );
  INV_X1 U9527 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7878) );
  NAND2_X1 U9528 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7918) );
  OAI21_X1 U9529 ( .B1(n8480), .B2(n7878), .A(n7918), .ZN(n7879) );
  AOI21_X1 U9530 ( .B1(n10007), .B2(n7880), .A(n7879), .ZN(n7881) );
  OAI211_X1 U9531 ( .C1(n10010), .C2(n7883), .A(n7882), .B(n7881), .ZN(
        P2_U3258) );
  INV_X1 U9532 ( .A(n7884), .ZN(n7888) );
  OAI222_X1 U9533 ( .A1(P1_U3084), .A2(n7886), .B1(n9774), .B2(n7888), .C1(
        n7885), .C2(n7832), .ZN(P1_U3329) );
  OAI222_X1 U9534 ( .A1(P2_U3152), .A2(n7889), .B1(n8894), .B2(n7888), .C1(
        n7887), .C2(n8904), .ZN(P2_U3334) );
  NAND2_X1 U9535 ( .A1(n7891), .A2(n7890), .ZN(n7893) );
  XNOR2_X1 U9536 ( .A(n7893), .B(n7892), .ZN(n7894) );
  AOI222_X1 U9537 ( .A1(n10021), .A2(n7894), .B1(n8422), .B2(n8665), .C1(n8424), .C2(n8663), .ZN(n8831) );
  INV_X1 U9538 ( .A(n7862), .ZN(n7896) );
  INV_X1 U9539 ( .A(n8728), .ZN(n7895) );
  AOI21_X1 U9540 ( .B1(n8828), .B2(n7896), .A(n7895), .ZN(n8829) );
  INV_X1 U9541 ( .A(n8274), .ZN(n7897) );
  AOI22_X1 U9542 ( .A1(n10031), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7897), .B2(
        n8678), .ZN(n7898) );
  OAI21_X1 U9543 ( .B1(n7899), .B2(n8681), .A(n7898), .ZN(n7902) );
  XNOR2_X1 U9544 ( .A(n7900), .B(n5587), .ZN(n8832) );
  NOR2_X1 U9545 ( .A1(n8832), .A2(n8734), .ZN(n7901) );
  AOI211_X1 U9546 ( .C1(n8829), .C2(n8670), .A(n7902), .B(n7901), .ZN(n7903)
         );
  OAI21_X1 U9547 ( .B1(n10031), .B2(n8831), .A(n7903), .ZN(P2_U3282) );
  NAND2_X1 U9548 ( .A1(n7904), .A2(n7914), .ZN(n7906) );
  XOR2_X1 U9549 ( .A(n7906), .B(n7905), .Z(n7913) );
  OAI21_X1 U9550 ( .B1(n8383), .B2(n7908), .A(n7907), .ZN(n7911) );
  OAI22_X1 U9551 ( .A1(n8409), .A2(n7909), .B1(n8381), .B2(n8273), .ZN(n7910)
         );
  AOI211_X1 U9552 ( .C1(n8839), .C2(n8411), .A(n7911), .B(n7910), .ZN(n7912)
         );
  OAI21_X1 U9553 ( .B1(n7913), .B2(n8413), .A(n7912), .ZN(P2_U3226) );
  NAND2_X1 U9554 ( .A1(n7915), .A2(n7914), .ZN(n7917) );
  XNOR2_X1 U9555 ( .A(n7917), .B(n7916), .ZN(n7924) );
  OAI21_X1 U9556 ( .B1(n8381), .B2(n8404), .A(n7918), .ZN(n7922) );
  OAI22_X1 U9557 ( .A1(n8409), .A2(n7920), .B1(n8383), .B2(n7919), .ZN(n7921)
         );
  AOI211_X1 U9558 ( .C1(n8833), .C2(n8411), .A(n7922), .B(n7921), .ZN(n7923)
         );
  OAI21_X1 U9559 ( .B1(n7924), .B2(n8413), .A(n7923), .ZN(P2_U3236) );
  OAI21_X1 U9560 ( .B1(n7927), .B2(n7926), .A(n7925), .ZN(n7937) );
  INV_X1 U9561 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7933) );
  NOR2_X1 U9562 ( .A1(n7929), .A2(n7928), .ZN(n7930) );
  OAI21_X1 U9563 ( .B1(n7931), .B2(n7930), .A(n10007), .ZN(n7932) );
  NAND2_X1 U9564 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8272) );
  OAI211_X1 U9565 ( .C1(n7933), .C2(n8480), .A(n7932), .B(n8272), .ZN(n7936)
         );
  NOR2_X1 U9566 ( .A1(n10010), .A2(n7934), .ZN(n7935) );
  AOI211_X1 U9567 ( .C1(n10008), .C2(n7937), .A(n7936), .B(n7935), .ZN(n7938)
         );
  INV_X1 U9568 ( .A(n7938), .ZN(P2_U3259) );
  INV_X1 U9569 ( .A(n8079), .ZN(n8263) );
  OAI222_X1 U9570 ( .A1(n8904), .A2(n7939), .B1(n8894), .B2(n8263), .C1(n5008), 
        .C2(P2_U3152), .ZN(P2_U3328) );
  INV_X1 U9571 ( .A(n8746), .ZN(n7940) );
  NOR2_X2 U9572 ( .A1(n8510), .A2(n8490), .ZN(n8489) );
  INV_X1 U9573 ( .A(n8670), .ZN(n8711) );
  NOR2_X1 U9574 ( .A1(n10029), .A2(n7942), .ZN(n7946) );
  NOR2_X1 U9575 ( .A1(n8897), .A2(n7943), .ZN(n7944) );
  NOR2_X1 U9576 ( .A1(n8336), .A2(n7944), .ZN(n8496) );
  NAND2_X1 U9577 ( .A1(n7945), .A2(n8496), .ZN(n8741) );
  NOR2_X1 U9578 ( .A1(n10031), .A2(n8741), .ZN(n8491) );
  AOI211_X1 U9579 ( .C1(n8737), .C2(n8727), .A(n7946), .B(n8491), .ZN(n7947)
         );
  OAI21_X1 U9580 ( .B1(n8739), .B2(n8711), .A(n7947), .ZN(P2_U3265) );
  INV_X1 U9581 ( .A(n8066), .ZN(n8097) );
  NAND2_X1 U9582 ( .A1(n8898), .A2(n8078), .ZN(n7949) );
  NAND2_X1 U9583 ( .A1(n8087), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n7948) );
  NOR2_X1 U9584 ( .A1(n9336), .A2(n9126), .ZN(n7950) );
  OR2_X1 U9585 ( .A1(n9339), .A2(n7950), .ZN(n7951) );
  AND2_X1 U9586 ( .A1(n9337), .A2(n9126), .ZN(n7958) );
  NOR2_X1 U9587 ( .A1(n7952), .A2(n9336), .ZN(n7957) );
  MUX2_X1 U9588 ( .A(n7958), .B(n7957), .S(n8097), .Z(n8045) );
  NAND2_X1 U9589 ( .A1(n8895), .A2(n8078), .ZN(n7960) );
  NAND2_X1 U9590 ( .A1(n8087), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7959) );
  INV_X1 U9591 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7961) );
  NAND2_X1 U9592 ( .A1(n7962), .A2(n7961), .ZN(n7963) );
  INV_X1 U9593 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n7966) );
  NAND2_X1 U9594 ( .A1(n8069), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n7965) );
  NAND2_X1 U9595 ( .A1(n4282), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n7964) );
  OAI211_X1 U9596 ( .C1(n7966), .C2(n8085), .A(n7965), .B(n7964), .ZN(n7967)
         );
  NAND2_X1 U9597 ( .A1(n9631), .A2(n4281), .ZN(n8103) );
  NAND2_X1 U9598 ( .A1(n9417), .A2(n9302), .ZN(n9333) );
  NAND2_X1 U9599 ( .A1(n9433), .A2(n9298), .ZN(n8160) );
  AND2_X1 U9600 ( .A1(n9333), .A2(n8160), .ZN(n7974) );
  OR2_X1 U9601 ( .A1(n7974), .A2(n9335), .ZN(n7969) );
  NAND2_X1 U9602 ( .A1(n7969), .A2(n9337), .ZN(n8204) );
  INV_X1 U9603 ( .A(n8204), .ZN(n7973) );
  INV_X1 U9604 ( .A(n9420), .ZN(n7970) );
  NAND2_X1 U9605 ( .A1(n9333), .A2(n7970), .ZN(n9334) );
  NAND2_X1 U9606 ( .A1(n4918), .A2(n9334), .ZN(n7971) );
  NOR2_X1 U9607 ( .A1(n9336), .A2(n7971), .ZN(n7972) );
  MUX2_X1 U9608 ( .A(n7973), .B(n7972), .S(n8066), .Z(n8043) );
  INV_X1 U9609 ( .A(n7974), .ZN(n8146) );
  OR2_X2 U9610 ( .A1(n9669), .A2(n9070), .ZN(n8161) );
  AND2_X1 U9611 ( .A1(n9675), .A2(n9290), .ZN(n9327) );
  NAND2_X1 U9612 ( .A1(n8161), .A2(n9327), .ZN(n7975) );
  NAND2_X1 U9613 ( .A1(n9669), .A2(n9070), .ZN(n9329) );
  AND2_X1 U9614 ( .A1(n7975), .A2(n9329), .ZN(n7976) );
  NAND2_X1 U9615 ( .A1(n9663), .A2(n9296), .ZN(n9331) );
  NAND2_X1 U9616 ( .A1(n7976), .A2(n9331), .ZN(n8198) );
  NAND2_X1 U9617 ( .A1(n9712), .A2(n8008), .ZN(n9316) );
  INV_X1 U9618 ( .A(n9316), .ZN(n8011) );
  NAND2_X1 U9619 ( .A1(n7439), .A2(n7986), .ZN(n7977) );
  NAND3_X1 U9620 ( .A1(n7977), .A2(n8109), .A3(n7996), .ZN(n7979) );
  NAND3_X1 U9621 ( .A1(n7979), .A2(n7978), .A3(n7987), .ZN(n7982) );
  INV_X1 U9622 ( .A(n7980), .ZN(n7981) );
  NAND2_X1 U9623 ( .A1(n7983), .A2(n7984), .ZN(n7985) );
  NAND2_X1 U9624 ( .A1(n7987), .A2(n7986), .ZN(n7999) );
  NOR2_X1 U9625 ( .A1(n7989), .A2(n7988), .ZN(n7990) );
  AND2_X1 U9626 ( .A1(n7992), .A2(n7991), .ZN(n7993) );
  NAND2_X1 U9627 ( .A1(n8125), .A2(n7993), .ZN(n8114) );
  INV_X1 U9628 ( .A(n7994), .ZN(n8003) );
  NAND2_X1 U9629 ( .A1(n7996), .A2(n7995), .ZN(n8126) );
  NAND2_X1 U9630 ( .A1(n8120), .A2(n8124), .ZN(n7997) );
  AND2_X1 U9631 ( .A1(n7998), .A2(n7997), .ZN(n8001) );
  INV_X1 U9632 ( .A(n7999), .ZN(n8000) );
  OAI21_X1 U9633 ( .B1(n8126), .B2(n8001), .A(n8000), .ZN(n8002) );
  OAI21_X1 U9634 ( .B1(n8114), .B2(n8003), .A(n8002), .ZN(n8192) );
  INV_X1 U9635 ( .A(n8192), .ZN(n9888) );
  NAND2_X1 U9636 ( .A1(n9887), .A2(n8110), .ZN(n8005) );
  NOR2_X1 U9637 ( .A1(n7983), .A2(n8004), .ZN(n8131) );
  NAND2_X1 U9638 ( .A1(n8015), .A2(n8006), .ZN(n8108) );
  INV_X1 U9639 ( .A(n8108), .ZN(n8007) );
  NAND3_X1 U9640 ( .A1(n8019), .A2(n8007), .A3(n9316), .ZN(n8010) );
  OR2_X1 U9641 ( .A1(n9712), .A2(n8008), .ZN(n8166) );
  NAND2_X1 U9642 ( .A1(n9541), .A2(n8166), .ZN(n8135) );
  INV_X1 U9643 ( .A(n8135), .ZN(n8009) );
  OAI211_X1 U9644 ( .C1(n8011), .C2(n8016), .A(n8010), .B(n8009), .ZN(n8012)
         );
  NAND2_X1 U9645 ( .A1(n9708), .A2(n9057), .ZN(n8165) );
  INV_X1 U9646 ( .A(n8015), .ZN(n8018) );
  INV_X1 U9647 ( .A(n8013), .ZN(n8014) );
  NAND2_X1 U9648 ( .A1(n8015), .A2(n8014), .ZN(n8017) );
  OAI211_X1 U9649 ( .C1(n8019), .C2(n8018), .A(n9312), .B(n8166), .ZN(n8021)
         );
  NAND2_X1 U9650 ( .A1(n8165), .A2(n9316), .ZN(n8112) );
  INV_X1 U9651 ( .A(n8112), .ZN(n8020) );
  NAND2_X1 U9652 ( .A1(n8021), .A2(n8020), .ZN(n8022) );
  INV_X1 U9653 ( .A(n9543), .ZN(n8023) );
  NAND2_X1 U9654 ( .A1(n9540), .A2(n9282), .ZN(n9318) );
  NAND2_X1 U9655 ( .A1(n9697), .A2(n9033), .ZN(n9319) );
  NAND2_X1 U9656 ( .A1(n9318), .A2(n9319), .ZN(n9544) );
  INV_X1 U9657 ( .A(n9544), .ZN(n8026) );
  INV_X1 U9658 ( .A(n9317), .ZN(n8024) );
  MUX2_X1 U9659 ( .A(n9543), .B(n8024), .S(n8097), .Z(n8025) );
  OR2_X1 U9660 ( .A1(n9530), .A2(n9021), .ZN(n9503) );
  NAND2_X1 U9661 ( .A1(n9530), .A2(n9021), .ZN(n9321) );
  NAND2_X1 U9662 ( .A1(n9503), .A2(n9321), .ZN(n9519) );
  INV_X1 U9663 ( .A(n9519), .ZN(n9523) );
  MUX2_X1 U9664 ( .A(n9318), .B(n9319), .S(n8066), .Z(n8027) );
  NAND3_X1 U9665 ( .A1(n8028), .A2(n9523), .A3(n8027), .ZN(n8030) );
  OR2_X1 U9666 ( .A1(n9510), .A2(n9285), .ZN(n8164) );
  AND2_X1 U9667 ( .A1(n8164), .A2(n9503), .ZN(n9322) );
  NAND2_X1 U9668 ( .A1(n9510), .A2(n9285), .ZN(n9323) );
  NAND2_X1 U9669 ( .A1(n9323), .A2(n9321), .ZN(n8140) );
  MUX2_X1 U9670 ( .A(n9322), .B(n4292), .S(n8097), .Z(n8029) );
  NAND2_X1 U9671 ( .A1(n8030), .A2(n8029), .ZN(n8034) );
  NAND2_X1 U9672 ( .A1(n9678), .A2(n9286), .ZN(n9324) );
  NAND2_X1 U9673 ( .A1(n9324), .A2(n9323), .ZN(n8105) );
  INV_X1 U9674 ( .A(n8105), .ZN(n8031) );
  OR2_X1 U9675 ( .A1(n9675), .A2(n9290), .ZN(n9326) );
  OR2_X1 U9676 ( .A1(n9678), .A2(n9286), .ZN(n8162) );
  AND2_X1 U9677 ( .A1(n9326), .A2(n8162), .ZN(n8104) );
  NAND2_X1 U9678 ( .A1(n8032), .A2(n8066), .ZN(n8033) );
  OR4_X1 U9679 ( .A1(n8146), .A2(n9296), .A3(n8097), .A4(n9663), .ZN(n8041) );
  NAND4_X1 U9680 ( .A1(n9420), .A2(n8097), .A3(n9296), .A4(n9663), .ZN(n8040)
         );
  NAND3_X1 U9681 ( .A1(n8034), .A2(n8164), .A3(n8162), .ZN(n8035) );
  INV_X1 U9682 ( .A(n9327), .ZN(n8163) );
  NAND3_X1 U9683 ( .A1(n8035), .A2(n8163), .A3(n9324), .ZN(n8036) );
  AOI21_X1 U9684 ( .B1(n8036), .B2(n9326), .A(n4907), .ZN(n8038) );
  OR2_X1 U9685 ( .A1(n9663), .A2(n9296), .ZN(n9330) );
  NAND3_X1 U9686 ( .A1(n9330), .A2(n8097), .A3(n8161), .ZN(n8037) );
  NOR2_X1 U9687 ( .A1(n8038), .A2(n8037), .ZN(n8039) );
  OR2_X1 U9688 ( .A1(n9636), .A2(n9126), .ZN(n9308) );
  NAND3_X1 U9689 ( .A1(n8046), .A2(n9380), .A3(n9308), .ZN(n8048) );
  MUX2_X1 U9690 ( .A(n8103), .B(n9340), .S(n8066), .Z(n8047) );
  NAND2_X1 U9691 ( .A1(n8890), .A2(n8078), .ZN(n8050) );
  NAND2_X1 U9692 ( .A1(n8087), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U9693 ( .A1(n4538), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9354) );
  INV_X1 U9694 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8051) );
  NAND2_X1 U9695 ( .A1(n8052), .A2(n8051), .ZN(n8053) );
  NAND2_X1 U9696 ( .A1(n9354), .A2(n8053), .ZN(n8979) );
  INV_X1 U9697 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U9698 ( .A1(n4282), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8056) );
  NAND2_X1 U9699 ( .A1(n8069), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8055) );
  OAI211_X1 U9700 ( .C1(n8085), .C2(n8057), .A(n8056), .B(n8055), .ZN(n8058)
         );
  INV_X1 U9701 ( .A(n8058), .ZN(n8059) );
  NAND2_X1 U9702 ( .A1(n9625), .A2(n8970), .ZN(n9341) );
  INV_X1 U9703 ( .A(n9362), .ZN(n8061) );
  MUX2_X1 U9704 ( .A(n8151), .B(n9341), .S(n8097), .Z(n8063) );
  NAND2_X1 U9705 ( .A1(n8265), .A2(n8078), .ZN(n8065) );
  NAND2_X1 U9706 ( .A1(n8087), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8064) );
  NAND2_X1 U9707 ( .A1(n9614), .A2(n8066), .ZN(n8077) );
  OR2_X1 U9708 ( .A1(n9354), .A2(n8067), .ZN(n8075) );
  INV_X1 U9709 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8072) );
  NAND2_X1 U9710 ( .A1(n4282), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8071) );
  NAND2_X1 U9711 ( .A1(n8069), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8070) );
  OAI211_X1 U9712 ( .C1(n8085), .C2(n8072), .A(n8071), .B(n8070), .ZN(n8073)
         );
  INV_X1 U9713 ( .A(n8073), .ZN(n8074) );
  INV_X1 U9714 ( .A(n8978), .ZN(n9124) );
  MUX2_X1 U9715 ( .A(n9124), .B(n9614), .S(n8097), .Z(n8076) );
  NAND2_X1 U9716 ( .A1(n8079), .A2(n8078), .ZN(n8081) );
  NAND2_X1 U9717 ( .A1(n8087), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8080) );
  INV_X1 U9718 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8084) );
  NAND2_X1 U9719 ( .A1(n4282), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8083) );
  NAND2_X1 U9720 ( .A1(n8069), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8082) );
  OAI211_X1 U9721 ( .C1(n8085), .C2(n8084), .A(n8083), .B(n8082), .ZN(n9343)
         );
  NAND2_X1 U9722 ( .A1(n9261), .A2(n9343), .ZN(n8086) );
  NAND2_X1 U9723 ( .A1(n9610), .A2(n8086), .ZN(n8208) );
  NAND2_X1 U9724 ( .A1(n8087), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U9725 ( .A1(n9604), .A2(n8096), .ZN(n8091) );
  OR2_X1 U9726 ( .A1(n9610), .A2(n9344), .ZN(n8090) );
  INV_X1 U9727 ( .A(n8189), .ZN(n8092) );
  NAND2_X1 U9728 ( .A1(n8092), .A2(n9604), .ZN(n8215) );
  NAND4_X1 U9729 ( .A1(n8095), .A2(n8978), .A3(n9616), .A4(n8208), .ZN(n8093)
         );
  NAND3_X1 U9730 ( .A1(n8094), .A2(n8215), .A3(n8093), .ZN(n8100) );
  OR2_X1 U9731 ( .A1(n9604), .A2(n8096), .ZN(n8232) );
  AOI21_X1 U9732 ( .B1(n8098), .B2(n8097), .A(n8187), .ZN(n8099) );
  INV_X1 U9733 ( .A(n8234), .ZN(n8239) );
  NAND2_X1 U9734 ( .A1(n8101), .A2(n9444), .ZN(n8155) );
  NAND2_X1 U9735 ( .A1(n9340), .A2(n9339), .ZN(n8102) );
  NAND3_X1 U9736 ( .A1(n9341), .A2(n8103), .A3(n8102), .ZN(n8206) );
  NAND2_X1 U9737 ( .A1(n9420), .A2(n9330), .ZN(n8200) );
  OAI211_X1 U9738 ( .C1(n9322), .C2(n8105), .A(n8161), .B(n8104), .ZN(n8196)
         );
  INV_X1 U9739 ( .A(n9319), .ZN(n8139) );
  INV_X1 U9740 ( .A(n8106), .ZN(n8107) );
  NOR2_X1 U9741 ( .A1(n8108), .A2(n8107), .ZN(n8130) );
  NAND3_X1 U9742 ( .A1(n8130), .A2(n8110), .A3(n8109), .ZN(n8111) );
  OR3_X1 U9743 ( .A1(n9317), .A2(n8112), .A3(n8111), .ZN(n8113) );
  OR3_X1 U9744 ( .A1(n8140), .A2(n8139), .A3(n8113), .ZN(n8193) );
  INV_X1 U9745 ( .A(n8114), .ZN(n8123) );
  AND2_X1 U9746 ( .A1(n8115), .A2(n6480), .ZN(n8119) );
  OAI211_X1 U9747 ( .C1(n8119), .C2(n8118), .A(n8117), .B(n8116), .ZN(n8121)
         );
  NAND3_X1 U9748 ( .A1(n8121), .A2(n8120), .A3(n7402), .ZN(n8122) );
  NAND2_X1 U9749 ( .A1(n8123), .A2(n8122), .ZN(n8129) );
  INV_X1 U9750 ( .A(n8124), .ZN(n8127) );
  OAI21_X1 U9751 ( .B1(n8127), .B2(n8126), .A(n8125), .ZN(n8128) );
  NAND2_X1 U9752 ( .A1(n8129), .A2(n8128), .ZN(n8141) );
  INV_X1 U9753 ( .A(n8130), .ZN(n8132) );
  OAI21_X1 U9754 ( .B1(n8132), .B2(n8131), .A(n9312), .ZN(n8133) );
  AND2_X1 U9755 ( .A1(n8133), .A2(n9316), .ZN(n8134) );
  OAI21_X1 U9756 ( .B1(n8135), .B2(n8134), .A(n8165), .ZN(n8136) );
  OAI211_X1 U9757 ( .C1(n9317), .C2(n8136), .A(n9318), .B(n9543), .ZN(n8137)
         );
  INV_X1 U9758 ( .A(n8137), .ZN(n8138) );
  OAI21_X1 U9759 ( .B1(n8193), .B2(n8141), .A(n8191), .ZN(n8142) );
  AND2_X1 U9760 ( .A1(n8142), .A2(n9324), .ZN(n8143) );
  NOR2_X1 U9761 ( .A1(n8196), .A2(n8143), .ZN(n8144) );
  NOR2_X1 U9762 ( .A1(n8198), .A2(n8144), .ZN(n8145) );
  NOR2_X1 U9763 ( .A1(n8200), .A2(n8145), .ZN(n8147) );
  NOR2_X1 U9764 ( .A1(n8147), .A2(n8146), .ZN(n8148) );
  NAND2_X1 U9765 ( .A1(n8149), .A2(n9337), .ZN(n8150) );
  NAND2_X1 U9766 ( .A1(n8158), .A2(n8151), .ZN(n8210) );
  NAND2_X1 U9767 ( .A1(n9610), .A2(n9344), .ZN(n8188) );
  NAND2_X1 U9768 ( .A1(n9614), .A2(n8978), .ZN(n8209) );
  OAI211_X1 U9769 ( .C1(n8152), .C2(n8210), .A(n8188), .B(n8209), .ZN(n8153)
         );
  AOI21_X1 U9770 ( .B1(n8189), .B2(n8153), .A(n8187), .ZN(n8154) );
  MUX2_X1 U9771 ( .A(n8155), .B(n8226), .S(n8154), .Z(n8230) );
  NAND4_X1 U9772 ( .A1(n8230), .A2(n8156), .A3(n8231), .A4(n9444), .ZN(n8238)
         );
  AND2_X1 U9773 ( .A1(n8216), .A2(n9471), .ZN(n8212) );
  INV_X1 U9774 ( .A(n8212), .ZN(n8157) );
  NOR2_X1 U9775 ( .A1(n6480), .A2(n8157), .ZN(n8224) );
  NAND2_X1 U9776 ( .A1(n9420), .A2(n8160), .ZN(n9437) );
  NAND2_X1 U9777 ( .A1(n9330), .A2(n9331), .ZN(n9455) );
  NAND2_X1 U9778 ( .A1(n8161), .A2(n9329), .ZN(n9328) );
  INV_X1 U9779 ( .A(n9328), .ZN(n9466) );
  NAND2_X1 U9780 ( .A1(n8164), .A2(n9323), .ZN(n9513) );
  INV_X1 U9781 ( .A(n9572), .ZN(n9571) );
  NAND2_X1 U9782 ( .A1(n8166), .A2(n9316), .ZN(n9587) );
  NOR4_X1 U9783 ( .A1(n8170), .A2(n8169), .A3(n8168), .A4(n8167), .ZN(n8173)
         );
  NAND4_X1 U9784 ( .A1(n8174), .A2(n8173), .A3(n8172), .A4(n8171), .ZN(n8178)
         );
  INV_X1 U9785 ( .A(n8175), .ZN(n9891) );
  NOR4_X1 U9786 ( .A1(n9513), .A2(n9544), .A3(n9519), .A4(n8182), .ZN(n8183)
         );
  NAND4_X1 U9787 ( .A1(n9466), .A2(n9496), .A3(n9479), .A4(n8183), .ZN(n8184)
         );
  NOR4_X1 U9788 ( .A1(n9403), .A2(n9437), .A3(n9455), .A4(n8184), .ZN(n8185)
         );
  XNOR2_X1 U9789 ( .A(n9417), .B(n9303), .ZN(n9424) );
  NAND4_X1 U9790 ( .A1(n9380), .A2(n9393), .A3(n8185), .A4(n9424), .ZN(n8186)
         );
  NAND3_X1 U9791 ( .A1(n8190), .A2(n8189), .A3(n8188), .ZN(n8223) );
  OAI21_X1 U9792 ( .B1(n8193), .B2(n8192), .A(n8191), .ZN(n8194) );
  AND2_X1 U9793 ( .A1(n8194), .A2(n9324), .ZN(n8195) );
  NOR2_X1 U9794 ( .A1(n8196), .A2(n8195), .ZN(n8197) );
  NOR2_X1 U9795 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  OR2_X1 U9796 ( .A1(n8200), .A2(n8199), .ZN(n8201) );
  NOR2_X1 U9797 ( .A1(n9335), .A2(n8201), .ZN(n8203) );
  OAI211_X1 U9798 ( .C1(n8204), .C2(n8203), .A(n8202), .B(n9338), .ZN(n8205)
         );
  INV_X1 U9799 ( .A(n8205), .ZN(n8207) );
  AOI21_X1 U9800 ( .B1(n8207), .B2(n9340), .A(n8206), .ZN(n8211) );
  OAI211_X1 U9801 ( .C1(n8211), .C2(n8210), .A(n8209), .B(n8208), .ZN(n8214)
         );
  NAND3_X1 U9802 ( .A1(n8232), .A2(n6480), .A3(n8212), .ZN(n8213) );
  AOI21_X1 U9803 ( .B1(n8215), .B2(n8214), .A(n8213), .ZN(n8222) );
  AND2_X1 U9804 ( .A1(n8216), .A2(n9444), .ZN(n8218) );
  INV_X1 U9805 ( .A(n8218), .ZN(n8220) );
  AOI21_X1 U9806 ( .B1(n6480), .B2(n8218), .A(n8217), .ZN(n8219) );
  OAI21_X1 U9807 ( .B1(n8223), .B2(n8220), .A(n8219), .ZN(n8221) );
  AOI211_X1 U9808 ( .C1(n8224), .C2(n8223), .A(n8222), .B(n8221), .ZN(n8229)
         );
  NOR4_X1 U9809 ( .A1(n9102), .A2(n9258), .A3(n8226), .A4(n8225), .ZN(n8227)
         );
  AOI211_X1 U9810 ( .C1(n8231), .C2(n6479), .A(n9257), .B(n8227), .ZN(n8228)
         );
  AOI21_X1 U9811 ( .B1(n8229), .B2(n8230), .A(n8228), .ZN(n8237) );
  INV_X1 U9812 ( .A(n8230), .ZN(n8235) );
  NAND4_X1 U9813 ( .A1(n8232), .A2(n6480), .A3(n8231), .A4(n6479), .ZN(n8233)
         );
  OAI211_X1 U9814 ( .C1(n8239), .C2(n8238), .A(n8237), .B(n8236), .ZN(P1_U3240) );
  NAND3_X1 U9815 ( .A1(n8241), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8243) );
  OAI22_X1 U9816 ( .A1(n8240), .A2(n8243), .B1(n8242), .B2(n8904), .ZN(n8244)
         );
  INV_X1 U9817 ( .A(n8244), .ZN(n8245) );
  OAI21_X1 U9818 ( .B1(n8256), .B2(n8894), .A(n8245), .ZN(P2_U3327) );
  OAI22_X1 U9819 ( .A1(n8250), .A2(n8383), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8249), .ZN(n8252) );
  NOR2_X1 U9820 ( .A1(n8416), .A2(n8381), .ZN(n8251) );
  AOI211_X1 U9821 ( .C1(n8389), .C2(n8533), .A(n8252), .B(n8251), .ZN(n8253)
         );
  INV_X1 U9822 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8255) );
  NAND3_X1 U9823 ( .A1(n8255), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n8261) );
  INV_X1 U9824 ( .A(n8256), .ZN(n8258) );
  NAND2_X1 U9825 ( .A1(n8258), .A2(n8257), .ZN(n8260) );
  NAND2_X1 U9826 ( .A1(n9771), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8259) );
  OAI211_X1 U9827 ( .C1(n8254), .C2(n8261), .A(n8260), .B(n8259), .ZN(P1_U3322) );
  INV_X1 U9828 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8264) );
  OAI222_X1 U9829 ( .A1(n7832), .A2(n8264), .B1(n9774), .B2(n8263), .C1(
        P1_U3084), .C2(n8262), .ZN(P1_U3323) );
  INV_X1 U9830 ( .A(n8265), .ZN(n9761) );
  INV_X1 U9831 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8266) );
  OAI222_X1 U9832 ( .A1(n8894), .A2(n9761), .B1(P2_U3152), .B2(n8267), .C1(
        n8266), .C2(n8904), .ZN(P2_U3329) );
  INV_X1 U9833 ( .A(n8316), .ZN(n8269) );
  AOI21_X1 U9834 ( .B1(n8271), .B2(n8270), .A(n8269), .ZN(n8278) );
  OAI21_X1 U9835 ( .B1(n8381), .B2(n8324), .A(n8272), .ZN(n8276) );
  OAI22_X1 U9836 ( .A1(n8409), .A2(n8274), .B1(n8383), .B2(n8273), .ZN(n8275)
         );
  AOI211_X1 U9837 ( .C1(n8828), .C2(n8411), .A(n8276), .B(n8275), .ZN(n8277)
         );
  OAI21_X1 U9838 ( .B1(n8278), .B2(n8413), .A(n8277), .ZN(P2_U3217) );
  NAND2_X1 U9839 ( .A1(n8279), .A2(n8343), .ZN(n8280) );
  XNOR2_X1 U9840 ( .A(n8280), .B(n8344), .ZN(n8286) );
  OAI22_X1 U9841 ( .A1(n8309), .A2(n8336), .B1(n8281), .B2(n8563), .ZN(n8583)
         );
  OAI22_X1 U9842 ( .A1(n8409), .A2(n8585), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8282), .ZN(n8284) );
  NOR2_X1 U9843 ( .A1(n8579), .A2(n8300), .ZN(n8283) );
  AOI211_X1 U9844 ( .C1(n8407), .C2(n8583), .A(n8284), .B(n8283), .ZN(n8285)
         );
  OAI21_X1 U9845 ( .B1(n8286), .B2(n8413), .A(n8285), .ZN(P2_U3218) );
  INV_X1 U9846 ( .A(n4447), .ZN(n8288) );
  AOI21_X1 U9847 ( .B1(n8290), .B2(n8289), .A(n8288), .ZN(n8296) );
  OAI22_X1 U9848 ( .A1(n8291), .A2(n8336), .B1(n8337), .B2(n8563), .ZN(n8639)
         );
  NAND2_X1 U9849 ( .A1(n8407), .A2(n8639), .ZN(n8292) );
  OAI211_X1 U9850 ( .C1(n8409), .C2(n8648), .A(n8293), .B(n8292), .ZN(n8294)
         );
  AOI21_X1 U9851 ( .B1(n8802), .B2(n8411), .A(n8294), .ZN(n8295) );
  OAI21_X1 U9852 ( .B1(n8296), .B2(n8413), .A(n8295), .ZN(P2_U3221) );
  XNOR2_X1 U9853 ( .A(n8298), .B(n8297), .ZN(n8304) );
  AOI22_X1 U9854 ( .A1(n5600), .A2(n8665), .B1(n8663), .B2(n8419), .ZN(n8611)
         );
  OAI22_X1 U9855 ( .A1(n8611), .A2(n8392), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8299), .ZN(n8302) );
  NOR2_X1 U9856 ( .A1(n8617), .A2(n8300), .ZN(n8301) );
  AOI211_X1 U9857 ( .C1(n8389), .C2(n8614), .A(n8302), .B(n8301), .ZN(n8303)
         );
  OAI21_X1 U9858 ( .B1(n8304), .B2(n8413), .A(n8303), .ZN(P2_U3225) );
  XOR2_X1 U9859 ( .A(n8306), .B(n8305), .Z(n8307) );
  XNOR2_X1 U9860 ( .A(n8308), .B(n8307), .ZN(n8314) );
  AOI22_X1 U9861 ( .A1(n8418), .A2(n8665), .B1(n8663), .B2(n5602), .ZN(n8553)
         );
  NOR2_X1 U9862 ( .A1(n8553), .A2(n8392), .ZN(n8312) );
  OAI22_X1 U9863 ( .A1(n8547), .A2(n8409), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8310), .ZN(n8311) );
  AOI211_X1 U9864 ( .C1(n8769), .C2(n8411), .A(n8312), .B(n8311), .ZN(n8313)
         );
  OAI21_X1 U9865 ( .B1(n8314), .B2(n8413), .A(n8313), .ZN(P2_U3227) );
  NAND2_X1 U9866 ( .A1(n8316), .A2(n8315), .ZN(n8318) );
  NAND2_X1 U9867 ( .A1(n8318), .A2(n8317), .ZN(n8400) );
  NOR2_X1 U9868 ( .A1(n8318), .A2(n8317), .ZN(n8399) );
  AOI21_X1 U9869 ( .B1(n8319), .B2(n8400), .A(n8399), .ZN(n8323) );
  XNOR2_X1 U9870 ( .A(n8321), .B(n8320), .ZN(n8322) );
  XNOR2_X1 U9871 ( .A(n8323), .B(n8322), .ZN(n8328) );
  OAI22_X1 U9872 ( .A1(n8382), .A2(n8336), .B1(n8324), .B2(n8563), .ZN(n8694)
         );
  AOI22_X1 U9873 ( .A1(n8407), .A2(n8694), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n8325) );
  OAI21_X1 U9874 ( .B1(n8409), .B2(n8706), .A(n8325), .ZN(n8326) );
  AOI21_X1 U9875 ( .B1(n8709), .B2(n8411), .A(n8326), .ZN(n8327) );
  OAI21_X1 U9876 ( .B1(n8328), .B2(n8413), .A(n8327), .ZN(P2_U3228) );
  NAND2_X1 U9877 ( .A1(n8330), .A2(n8329), .ZN(n8332) );
  NAND2_X1 U9878 ( .A1(n8332), .A2(n8331), .ZN(n8334) );
  XNOR2_X1 U9879 ( .A(n8334), .B(n8333), .ZN(n8342) );
  INV_X1 U9880 ( .A(n8679), .ZN(n8339) );
  OAI22_X1 U9881 ( .A1(n8337), .A2(n8336), .B1(n8335), .B2(n8563), .ZN(n8674)
         );
  AOI22_X1 U9882 ( .A1(n8407), .A2(n8674), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8338) );
  OAI21_X1 U9883 ( .B1(n8409), .B2(n8339), .A(n8338), .ZN(n8340) );
  AOI21_X1 U9884 ( .B1(n8811), .B2(n8411), .A(n8340), .ZN(n8341) );
  OAI21_X1 U9885 ( .B1(n8342), .B2(n8413), .A(n8341), .ZN(P2_U3230) );
  INV_X1 U9886 ( .A(n8279), .ZN(n8345) );
  OAI21_X1 U9887 ( .B1(n8345), .B2(n8344), .A(n8343), .ZN(n8349) );
  XOR2_X1 U9888 ( .A(n8347), .B(n8346), .Z(n8348) );
  XNOR2_X1 U9889 ( .A(n8349), .B(n8348), .ZN(n8356) );
  OAI22_X1 U9890 ( .A1(n8564), .A2(n8383), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8350), .ZN(n8354) );
  INV_X1 U9891 ( .A(n8560), .ZN(n8351) );
  OAI22_X1 U9892 ( .A1(n8352), .A2(n8381), .B1(n8409), .B2(n8351), .ZN(n8353)
         );
  AOI211_X1 U9893 ( .C1(n8776), .C2(n8411), .A(n8354), .B(n8353), .ZN(n8355)
         );
  OAI21_X1 U9894 ( .B1(n8356), .B2(n8413), .A(n8355), .ZN(P2_U3231) );
  XNOR2_X1 U9895 ( .A(n8358), .B(n8357), .ZN(n8362) );
  OAI22_X1 U9896 ( .A1(n8381), .A2(n8371), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10232), .ZN(n8360) );
  OAI22_X1 U9897 ( .A1(n8409), .A2(n8622), .B1(n8383), .B2(n8380), .ZN(n8359)
         );
  AOI211_X1 U9898 ( .C1(n8796), .C2(n8411), .A(n8360), .B(n8359), .ZN(n8361)
         );
  OAI21_X1 U9899 ( .B1(n8362), .B2(n8413), .A(n8361), .ZN(P2_U3235) );
  INV_X1 U9900 ( .A(n8363), .ZN(n8364) );
  NOR2_X1 U9901 ( .A1(n8365), .A2(n8364), .ZN(n8369) );
  XNOR2_X1 U9902 ( .A(n8367), .B(n8366), .ZN(n8368) );
  XNOR2_X1 U9903 ( .A(n8369), .B(n8368), .ZN(n8375) );
  OAI22_X1 U9904 ( .A1(n8564), .A2(n8381), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8370), .ZN(n8373) );
  OAI22_X1 U9905 ( .A1(n8409), .A2(n8591), .B1(n8383), .B2(n8371), .ZN(n8372)
         );
  AOI211_X1 U9906 ( .C1(n8786), .C2(n8411), .A(n8373), .B(n8372), .ZN(n8374)
         );
  OAI21_X1 U9907 ( .B1(n8375), .B2(n8413), .A(n8374), .ZN(P2_U3237) );
  NAND2_X1 U9908 ( .A1(n8377), .A2(n8376), .ZN(n8379) );
  XNOR2_X1 U9909 ( .A(n8379), .B(n8378), .ZN(n8387) );
  NAND2_X1 U9910 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8478) );
  OAI21_X1 U9911 ( .B1(n8381), .B2(n8380), .A(n8478), .ZN(n8385) );
  OAI22_X1 U9912 ( .A1(n8409), .A2(n8657), .B1(n8383), .B2(n8382), .ZN(n8384)
         );
  AOI211_X1 U9913 ( .C1(n8805), .C2(n8411), .A(n8385), .B(n8384), .ZN(n8386)
         );
  OAI21_X1 U9914 ( .B1(n8387), .B2(n8413), .A(n8386), .ZN(P2_U3240) );
  INV_X1 U9915 ( .A(n8388), .ZN(n8393) );
  AOI22_X1 U9916 ( .A1(n8390), .A2(n8389), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8391) );
  OAI21_X1 U9917 ( .B1(n8393), .B2(n8392), .A(n8391), .ZN(n8397) );
  INV_X1 U9918 ( .A(n8398), .ZN(P2_U3242) );
  INV_X1 U9919 ( .A(n8399), .ZN(n8401) );
  NAND2_X1 U9920 ( .A1(n8401), .A2(n8400), .ZN(n8403) );
  XNOR2_X1 U9921 ( .A(n8403), .B(n8402), .ZN(n8414) );
  OR2_X1 U9922 ( .A1(n8404), .A2(n8563), .ZN(n8406) );
  NAND2_X1 U9923 ( .A1(n8421), .A2(n8665), .ZN(n8405) );
  NAND2_X1 U9924 ( .A1(n8406), .A2(n8405), .ZN(n8716) );
  AOI22_X1 U9925 ( .A1(n8407), .A2(n8716), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n8408) );
  OAI21_X1 U9926 ( .B1(n8409), .B2(n8724), .A(n8408), .ZN(n8410) );
  AOI21_X1 U9927 ( .B1(n8824), .B2(n8411), .A(n8410), .ZN(n8412) );
  OAI21_X1 U9928 ( .B1(n8414), .B2(n8413), .A(n8412), .ZN(P2_U3243) );
  MUX2_X1 U9929 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8495), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9930 ( .A(n8415), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8436), .Z(
        P2_U3581) );
  INV_X1 U9931 ( .A(n8416), .ZN(n8503) );
  MUX2_X1 U9932 ( .A(n8503), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8436), .Z(
        P2_U3580) );
  MUX2_X1 U9933 ( .A(n8417), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8436), .Z(
        P2_U3579) );
  MUX2_X1 U9934 ( .A(n8418), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8436), .Z(
        P2_U3578) );
  MUX2_X1 U9935 ( .A(n8571), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8436), .Z(
        P2_U3577) );
  MUX2_X1 U9936 ( .A(n5602), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8436), .Z(
        P2_U3576) );
  MUX2_X1 U9937 ( .A(n8598), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8436), .Z(
        P2_U3575) );
  MUX2_X1 U9938 ( .A(n5600), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8436), .Z(
        P2_U3574) );
  MUX2_X1 U9939 ( .A(n8628), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8436), .Z(
        P2_U3573) );
  MUX2_X1 U9940 ( .A(n8419), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8436), .Z(
        P2_U3572) );
  MUX2_X1 U9941 ( .A(n8666), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8436), .Z(
        P2_U3571) );
  MUX2_X1 U9942 ( .A(n8420), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8436), .Z(
        P2_U3570) );
  MUX2_X1 U9943 ( .A(n8664), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8436), .Z(
        P2_U3569) );
  MUX2_X1 U9944 ( .A(n8421), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8436), .Z(
        P2_U3568) );
  MUX2_X1 U9945 ( .A(n8422), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8436), .Z(
        P2_U3567) );
  MUX2_X1 U9946 ( .A(n8423), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8436), .Z(
        P2_U3566) );
  MUX2_X1 U9947 ( .A(n8424), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8436), .Z(
        P2_U3565) );
  MUX2_X1 U9948 ( .A(n8425), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8436), .Z(
        P2_U3564) );
  MUX2_X1 U9949 ( .A(n8426), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8436), .Z(
        P2_U3563) );
  MUX2_X1 U9950 ( .A(n8427), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8436), .Z(
        P2_U3562) );
  MUX2_X1 U9951 ( .A(n8428), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8436), .Z(
        P2_U3561) );
  MUX2_X1 U9952 ( .A(n8429), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8436), .Z(
        P2_U3560) );
  MUX2_X1 U9953 ( .A(n8430), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8436), .Z(
        P2_U3559) );
  MUX2_X1 U9954 ( .A(n8431), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8436), .Z(
        P2_U3558) );
  MUX2_X1 U9955 ( .A(n8432), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8436), .Z(
        P2_U3557) );
  MUX2_X1 U9956 ( .A(n8433), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8436), .Z(
        P2_U3556) );
  MUX2_X1 U9957 ( .A(n8434), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8436), .Z(
        P2_U3555) );
  MUX2_X1 U9958 ( .A(n5657), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8436), .Z(
        P2_U3554) );
  MUX2_X1 U9959 ( .A(n8435), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8436), .Z(
        P2_U3553) );
  MUX2_X1 U9960 ( .A(n8437), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8436), .Z(
        P2_U3552) );
  OAI21_X1 U9961 ( .B1(n8439), .B2(n8725), .A(n8438), .ZN(n8447) );
  AND2_X1 U9962 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8440) );
  AOI21_X1 U9963 ( .B1(n10009), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8440), .ZN(
        n8444) );
  OAI211_X1 U9964 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n8442), .A(n10007), .B(
        n8441), .ZN(n8443) );
  OAI211_X1 U9965 ( .C1(n10010), .C2(n8445), .A(n8444), .B(n8443), .ZN(n8446)
         );
  AOI21_X1 U9966 ( .B1(n10008), .B2(n8447), .A(n8446), .ZN(n8448) );
  INV_X1 U9967 ( .A(n8448), .ZN(P2_U3260) );
  AOI21_X1 U9968 ( .B1(n8451), .B2(n8450), .A(n8449), .ZN(n8462) );
  INV_X1 U9969 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8454) );
  OR2_X1 U9970 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8452), .ZN(n8453) );
  OAI21_X1 U9971 ( .B1(n8480), .B2(n8454), .A(n8453), .ZN(n8459) );
  AOI211_X1 U9972 ( .C1(n8457), .C2(n8456), .A(n8455), .B(n8481), .ZN(n8458)
         );
  AOI211_X1 U9973 ( .C1(n8487), .C2(n8460), .A(n8459), .B(n8458), .ZN(n8461)
         );
  OAI21_X1 U9974 ( .B1(n8462), .B2(n10011), .A(n8461), .ZN(P2_U3261) );
  AND2_X1 U9975 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8469) );
  INV_X1 U9976 ( .A(n8463), .ZN(n8467) );
  INV_X1 U9977 ( .A(n8464), .ZN(n8466) );
  AOI211_X1 U9978 ( .C1(n8467), .C2(n8466), .A(n8465), .B(n10011), .ZN(n8468)
         );
  AOI211_X1 U9979 ( .C1(n10009), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n8469), .B(
        n8468), .ZN(n8472) );
  OAI211_X1 U9980 ( .C1(n4394), .C2(n4622), .A(n10008), .B(n8470), .ZN(n8471)
         );
  OAI211_X1 U9981 ( .C1(n10010), .C2(n8473), .A(n8472), .B(n8471), .ZN(
        P2_U3262) );
  INV_X1 U9982 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10120) );
  AND2_X1 U9983 ( .A1(n8475), .A2(n8474), .ZN(n8476) );
  OAI21_X1 U9984 ( .B1(n8477), .B2(n8476), .A(n10007), .ZN(n8479) );
  OAI211_X1 U9985 ( .C1(n10120), .C2(n8480), .A(n8479), .B(n8478), .ZN(n8485)
         );
  AOI211_X1 U9986 ( .C1(n8483), .C2(n5378), .A(n8482), .B(n8481), .ZN(n8484)
         );
  AOI211_X1 U9987 ( .C1(n8487), .C2(n8486), .A(n8485), .B(n8484), .ZN(n8488)
         );
  INV_X1 U9988 ( .A(n8488), .ZN(P2_U3263) );
  AOI21_X1 U9989 ( .B1(n8490), .B2(n8510), .A(n8489), .ZN(n8740) );
  NAND2_X1 U9990 ( .A1(n8740), .A2(n8670), .ZN(n8493) );
  AOI21_X1 U9991 ( .B1(n10031), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8491), .ZN(
        n8492) );
  OAI211_X1 U9992 ( .C1(n8743), .C2(n8681), .A(n8493), .B(n8492), .ZN(P2_U3266) );
  AOI22_X1 U9993 ( .A1(n8503), .A2(n8663), .B1(n8496), .B2(n8495), .ZN(n8497)
         );
  NAND2_X1 U9994 ( .A1(n8535), .A2(n8501), .ZN(n8502) );
  NOR2_X1 U9995 ( .A1(n8755), .A2(n8503), .ZN(n8744) );
  INV_X1 U9996 ( .A(n8744), .ZN(n8504) );
  NAND2_X1 U9997 ( .A1(n8751), .A2(n8504), .ZN(n8505) );
  XNOR2_X1 U9998 ( .A(n8505), .B(n8745), .ZN(n8506) );
  NAND2_X1 U9999 ( .A1(n8506), .A2(n8531), .ZN(n8516) );
  OAI22_X1 U10000 ( .A1(n8508), .A2(n10041), .B1(n8507), .B2(n10029), .ZN(
        n8514) );
  AOI21_X1 U10001 ( .B1(n8746), .B2(n8509), .A(n8816), .ZN(n8511) );
  NOR2_X1 U10002 ( .A1(n8748), .A2(n8512), .ZN(n8513) );
  AOI211_X1 U10003 ( .C1(n8727), .C2(n8746), .A(n8514), .B(n8513), .ZN(n8515)
         );
  OAI211_X1 U10004 ( .C1(n8517), .C2(n10031), .A(n8516), .B(n8515), .ZN(
        P2_U3267) );
  XNOR2_X1 U10005 ( .A(n8518), .B(n8521), .ZN(n8520) );
  OAI21_X1 U10006 ( .B1(n8520), .B2(n8673), .A(n8519), .ZN(n8752) );
  INV_X1 U10007 ( .A(n8752), .ZN(n8530) );
  XNOR2_X1 U10008 ( .A(n8522), .B(n8521), .ZN(n8753) );
  NAND2_X1 U10009 ( .A1(n8753), .A2(n8531), .ZN(n8529) );
  AOI211_X1 U10010 ( .C1(n8755), .C2(n8524), .A(n8816), .B(n8523), .ZN(n8754)
         );
  AOI22_X1 U10011 ( .A1(n8525), .A2(n8678), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10031), .ZN(n8526) );
  OAI21_X1 U10012 ( .B1(n4680), .B2(n8681), .A(n8526), .ZN(n8527) );
  AOI21_X1 U10013 ( .B1(n8754), .B2(n8731), .A(n8527), .ZN(n8528) );
  OAI211_X1 U10014 ( .C1(n8530), .C2(n10031), .A(n8529), .B(n8528), .ZN(
        P2_U3268) );
  NAND2_X1 U10015 ( .A1(n8532), .A2(n8531), .ZN(n8539) );
  AOI22_X1 U10016 ( .A1(n8533), .A2(n8678), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n10031), .ZN(n8534) );
  OAI21_X1 U10017 ( .B1(n8535), .B2(n8681), .A(n8534), .ZN(n8536) );
  AOI21_X1 U10018 ( .B1(n8537), .B2(n8670), .A(n8536), .ZN(n8538) );
  OAI211_X1 U10019 ( .C1(n8540), .C2(n10031), .A(n8539), .B(n8538), .ZN(
        P2_U3269) );
  XNOR2_X1 U10020 ( .A(n4316), .B(n4880), .ZN(n8767) );
  INV_X1 U10021 ( .A(n8541), .ZN(n8544) );
  INV_X1 U10022 ( .A(n8542), .ZN(n8543) );
  AOI211_X1 U10023 ( .C1(n8769), .C2(n8544), .A(n8816), .B(n8543), .ZN(n8768)
         );
  NOR2_X1 U10024 ( .A1(n8545), .A2(n8681), .ZN(n8549) );
  OAI22_X1 U10025 ( .A1(n8547), .A2(n10041), .B1(n8546), .B2(n10029), .ZN(
        n8548) );
  AOI211_X1 U10026 ( .C1(n8768), .C2(n8689), .A(n8549), .B(n8548), .ZN(n8556)
         );
  OAI211_X1 U10027 ( .C1(n8552), .C2(n8551), .A(n8550), .B(n10021), .ZN(n8554)
         );
  NAND2_X1 U10028 ( .A1(n8554), .A2(n8553), .ZN(n8766) );
  NAND2_X1 U10029 ( .A1(n8766), .A2(n10029), .ZN(n8555) );
  OAI211_X1 U10030 ( .C1(n8767), .C2(n8734), .A(n8556), .B(n8555), .ZN(
        P2_U3271) );
  AOI21_X1 U10031 ( .B1(n8559), .B2(n8558), .A(n8557), .ZN(n8780) );
  XNOR2_X1 U10032 ( .A(n8562), .B(n8577), .ZN(n8777) );
  AOI22_X1 U10033 ( .A1(n8560), .A2(n8678), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10031), .ZN(n8561) );
  OAI21_X1 U10034 ( .B1(n8562), .B2(n8681), .A(n8561), .ZN(n8573) );
  NOR2_X1 U10035 ( .A1(n8564), .A2(n8563), .ZN(n8570) );
  INV_X1 U10036 ( .A(n8565), .ZN(n8566) );
  AOI211_X1 U10037 ( .C1(n8568), .C2(n8567), .A(n8673), .B(n8566), .ZN(n8569)
         );
  AOI211_X2 U10038 ( .C1(n8665), .C2(n8571), .A(n8570), .B(n8569), .ZN(n8779)
         );
  NOR2_X1 U10039 ( .A1(n8779), .A2(n10031), .ZN(n8572) );
  OAI21_X1 U10040 ( .B1(n8780), .B2(n8734), .A(n8574), .ZN(P2_U3272) );
  OAI21_X1 U10041 ( .B1(n8576), .B2(n8581), .A(n8575), .ZN(n8785) );
  AOI21_X1 U10042 ( .B1(n8781), .B2(n8590), .A(n5606), .ZN(n8782) );
  OAI22_X1 U10043 ( .A1(n8579), .A2(n8681), .B1(n8578), .B2(n10029), .ZN(n8580) );
  AOI21_X1 U10044 ( .B1(n8782), .B2(n8670), .A(n8580), .ZN(n8588) );
  XNOR2_X1 U10045 ( .A(n8582), .B(n8581), .ZN(n8584) );
  AOI21_X1 U10046 ( .B1(n8584), .B2(n10021), .A(n8583), .ZN(n8784) );
  OAI21_X1 U10047 ( .B1(n8585), .B2(n10041), .A(n8784), .ZN(n8586) );
  NAND2_X1 U10048 ( .A1(n8586), .A2(n10029), .ZN(n8587) );
  OAI211_X1 U10049 ( .C1(n8785), .C2(n8734), .A(n8588), .B(n8587), .ZN(
        P2_U3273) );
  XNOR2_X1 U10050 ( .A(n8589), .B(n8596), .ZN(n8790) );
  AOI21_X1 U10051 ( .B1(n8786), .B2(n4297), .A(n4685), .ZN(n8787) );
  INV_X1 U10052 ( .A(n8591), .ZN(n8592) );
  AOI22_X1 U10053 ( .A1(n10031), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8592), 
        .B2(n8678), .ZN(n8593) );
  OAI21_X1 U10054 ( .B1(n8594), .B2(n8681), .A(n8593), .ZN(n8602) );
  OAI211_X1 U10055 ( .C1(n8597), .C2(n8596), .A(n8595), .B(n10021), .ZN(n8600)
         );
  AOI22_X1 U10056 ( .A1(n8598), .A2(n8665), .B1(n8663), .B2(n8628), .ZN(n8599)
         );
  NOR2_X1 U10057 ( .A1(n8789), .A2(n10031), .ZN(n8601) );
  AOI211_X1 U10058 ( .C1(n8787), .C2(n8670), .A(n8602), .B(n8601), .ZN(n8603)
         );
  OAI21_X1 U10059 ( .B1(n8790), .B2(n8734), .A(n8603), .ZN(P2_U3274) );
  XOR2_X1 U10060 ( .A(n8604), .B(n8610), .Z(n8795) );
  NAND2_X1 U10061 ( .A1(n8606), .A2(n8605), .ZN(n8609) );
  INV_X1 U10062 ( .A(n8607), .ZN(n8608) );
  AOI21_X1 U10063 ( .B1(n8610), .B2(n8609), .A(n8608), .ZN(n8612) );
  OAI21_X1 U10064 ( .B1(n8612), .B2(n8673), .A(n8611), .ZN(n8791) );
  XNOR2_X1 U10065 ( .A(n8621), .B(n8617), .ZN(n8613) );
  NOR2_X1 U10066 ( .A1(n8613), .A2(n8816), .ZN(n8792) );
  NAND2_X1 U10067 ( .A1(n8792), .A2(n8731), .ZN(n8616) );
  AOI22_X1 U10068 ( .A1(n10031), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8614), 
        .B2(n8678), .ZN(n8615) );
  OAI211_X1 U10069 ( .C1(n8617), .C2(n8681), .A(n8616), .B(n8615), .ZN(n8618)
         );
  AOI21_X1 U10070 ( .B1(n8791), .B2(n10029), .A(n8618), .ZN(n8619) );
  OAI21_X1 U10071 ( .B1(n8795), .B2(n8734), .A(n8619), .ZN(P2_U3275) );
  XNOR2_X1 U10072 ( .A(n8620), .B(n8627), .ZN(n8800) );
  AOI21_X1 U10073 ( .B1(n8796), .B2(n4983), .A(n8621), .ZN(n8797) );
  INV_X1 U10074 ( .A(n8796), .ZN(n8625) );
  INV_X1 U10075 ( .A(n8622), .ZN(n8623) );
  AOI22_X1 U10076 ( .A1(n10031), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8623), 
        .B2(n8678), .ZN(n8624) );
  OAI21_X1 U10077 ( .B1(n8625), .B2(n8681), .A(n8624), .ZN(n8631) );
  XOR2_X1 U10078 ( .A(n8626), .B(n8627), .Z(n8629) );
  AOI222_X1 U10079 ( .A1(n10021), .A2(n8629), .B1(n8628), .B2(n8665), .C1(
        n8666), .C2(n8663), .ZN(n8799) );
  NOR2_X1 U10080 ( .A1(n8799), .A2(n10031), .ZN(n8630) );
  AOI211_X1 U10081 ( .C1(n8797), .C2(n8670), .A(n8631), .B(n8630), .ZN(n8632)
         );
  OAI21_X1 U10082 ( .B1(n8734), .B2(n8800), .A(n8632), .ZN(P2_U3276) );
  INV_X1 U10083 ( .A(n8635), .ZN(n8634) );
  XNOR2_X1 U10084 ( .A(n8633), .B(n8634), .ZN(n8804) );
  XNOR2_X1 U10085 ( .A(n8636), .B(n8635), .ZN(n8637) );
  NAND2_X1 U10086 ( .A1(n8637), .A2(n10021), .ZN(n8645) );
  INV_X1 U10087 ( .A(n8804), .ZN(n8643) );
  XNOR2_X1 U10088 ( .A(n8638), .B(n8654), .ZN(n8640) );
  AOI21_X1 U10089 ( .B1(n8640), .B2(n8861), .A(n8639), .ZN(n8641) );
  NAND2_X1 U10090 ( .A1(n8645), .A2(n8641), .ZN(n8801) );
  AOI21_X1 U10091 ( .B1(n8643), .B2(n8642), .A(n8801), .ZN(n8644) );
  AOI211_X1 U10092 ( .C1(n8646), .C2(n8645), .A(n10031), .B(n8644), .ZN(n8647)
         );
  INV_X1 U10093 ( .A(n8647), .ZN(n8652) );
  INV_X1 U10094 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8649) );
  OAI22_X1 U10095 ( .A1(n10029), .A2(n8649), .B1(n8648), .B2(n10041), .ZN(
        n8650) );
  AOI21_X1 U10096 ( .B1(n8802), .B2(n8727), .A(n8650), .ZN(n8651) );
  OAI211_X1 U10097 ( .C1(n8804), .C2(n8702), .A(n8652), .B(n8651), .ZN(
        P2_U3277) );
  XNOR2_X1 U10098 ( .A(n8653), .B(n4982), .ZN(n8809) );
  INV_X1 U10099 ( .A(n8677), .ZN(n8656) );
  INV_X1 U10100 ( .A(n8654), .ZN(n8655) );
  AOI21_X1 U10101 ( .B1(n8805), .B2(n8656), .A(n8655), .ZN(n8806) );
  INV_X1 U10102 ( .A(n8657), .ZN(n8658) );
  AOI22_X1 U10103 ( .A1(n10031), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8658), 
        .B2(n8678), .ZN(n8659) );
  OAI21_X1 U10104 ( .B1(n8660), .B2(n8681), .A(n8659), .ZN(n8669) );
  OAI21_X1 U10105 ( .B1(n8662), .B2(n4982), .A(n8661), .ZN(n8667) );
  AOI222_X1 U10106 ( .A1(n10021), .A2(n8667), .B1(n8666), .B2(n8665), .C1(
        n8664), .C2(n8663), .ZN(n8808) );
  NOR2_X1 U10107 ( .A1(n8808), .A2(n10031), .ZN(n8668) );
  AOI211_X1 U10108 ( .C1(n8806), .C2(n8670), .A(n8669), .B(n8668), .ZN(n8671)
         );
  OAI21_X1 U10109 ( .B1(n8809), .B2(n8734), .A(n8671), .ZN(P2_U3278) );
  AOI21_X1 U10110 ( .B1(n8672), .B2(n5593), .A(n8673), .ZN(n8676) );
  AOI21_X1 U10111 ( .B1(n8676), .B2(n8675), .A(n8674), .ZN(n8813) );
  AOI211_X1 U10112 ( .C1(n8811), .C2(n8705), .A(n8816), .B(n8677), .ZN(n8810)
         );
  INV_X1 U10113 ( .A(n8811), .ZN(n8682) );
  AOI22_X1 U10114 ( .A1(n10031), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8679), 
        .B2(n8678), .ZN(n8680) );
  OAI21_X1 U10115 ( .B1(n8682), .B2(n8681), .A(n8680), .ZN(n8688) );
  INV_X1 U10116 ( .A(n8684), .ZN(n8685) );
  AOI21_X1 U10117 ( .B1(n8686), .B2(n8683), .A(n8685), .ZN(n8814) );
  NOR2_X1 U10118 ( .A1(n8814), .A2(n8734), .ZN(n8687) );
  AOI211_X1 U10119 ( .C1(n8810), .C2(n8689), .A(n8688), .B(n8687), .ZN(n8690)
         );
  OAI21_X1 U10120 ( .B1(n10031), .B2(n8813), .A(n8690), .ZN(P2_U3279) );
  OAI21_X1 U10121 ( .B1(n8691), .B2(n8696), .A(n4403), .ZN(n8701) );
  OR2_X1 U10122 ( .A1(n8701), .A2(n8693), .ZN(n8700) );
  INV_X1 U10123 ( .A(n8694), .ZN(n8699) );
  XNOR2_X1 U10124 ( .A(n8695), .B(n8696), .ZN(n8697) );
  NAND2_X1 U10125 ( .A1(n8697), .A2(n10021), .ZN(n8698) );
  INV_X1 U10126 ( .A(n8701), .ZN(n8820) );
  INV_X1 U10127 ( .A(n8702), .ZN(n8713) );
  INV_X1 U10128 ( .A(n8703), .ZN(n8729) );
  NAND2_X1 U10129 ( .A1(n8729), .A2(n8709), .ZN(n8704) );
  NAND2_X1 U10130 ( .A1(n8705), .A2(n8704), .ZN(n8817) );
  INV_X1 U10131 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8707) );
  OAI22_X1 U10132 ( .A1(n10029), .A2(n8707), .B1(n8706), .B2(n10041), .ZN(
        n8708) );
  AOI21_X1 U10133 ( .B1(n8709), .B2(n8727), .A(n8708), .ZN(n8710) );
  OAI21_X1 U10134 ( .B1(n8817), .B2(n8711), .A(n8710), .ZN(n8712) );
  AOI21_X1 U10135 ( .B1(n8820), .B2(n8713), .A(n8712), .ZN(n8714) );
  OAI21_X1 U10136 ( .B1(n8822), .B2(n10031), .A(n8714), .ZN(P2_U3280) );
  XNOR2_X1 U10137 ( .A(n8715), .B(n8721), .ZN(n8717) );
  AOI21_X1 U10138 ( .B1(n8717), .B2(n10021), .A(n8716), .ZN(n8826) );
  NAND2_X1 U10139 ( .A1(n8719), .A2(n8718), .ZN(n8722) );
  NAND2_X1 U10140 ( .A1(n8722), .A2(n8721), .ZN(n8720) );
  OAI21_X1 U10141 ( .B1(n8722), .B2(n8721), .A(n8720), .ZN(n8723) );
  INV_X1 U10142 ( .A(n8723), .ZN(n8827) );
  OAI22_X1 U10143 ( .A1(n10029), .A2(n8725), .B1(n8724), .B2(n10041), .ZN(
        n8726) );
  AOI21_X1 U10144 ( .B1(n8824), .B2(n8727), .A(n8726), .ZN(n8733) );
  AOI21_X1 U10145 ( .B1(n8728), .B2(n8824), .A(n8816), .ZN(n8730) );
  AND2_X1 U10146 ( .A1(n8730), .A2(n8729), .ZN(n8823) );
  NAND2_X1 U10147 ( .A1(n8823), .A2(n8731), .ZN(n8732) );
  OAI211_X1 U10148 ( .C1(n8827), .C2(n8734), .A(n8733), .B(n8732), .ZN(n8735)
         );
  INV_X1 U10149 ( .A(n8735), .ZN(n8736) );
  OAI21_X1 U10150 ( .B1(n10031), .B2(n8826), .A(n8736), .ZN(P2_U3281) );
  NAND2_X1 U10151 ( .A1(n8737), .A2(n10032), .ZN(n8738) );
  OAI211_X1 U10152 ( .C1(n8739), .C2(n8816), .A(n8741), .B(n8738), .ZN(n8867)
         );
  MUX2_X1 U10153 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8867), .S(n10082), .Z(
        P2_U3551) );
  NAND2_X1 U10154 ( .A1(n8740), .A2(n8861), .ZN(n8742) );
  OAI211_X1 U10155 ( .C1(n8743), .C2(n10070), .A(n8742), .B(n8741), .ZN(n8868)
         );
  MUX2_X1 U10156 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8868), .S(n10082), .Z(
        P2_U3550) );
  NOR3_X1 U10157 ( .A1(n8745), .A2(n8849), .A3(n8744), .ZN(n8750) );
  NAND3_X1 U10158 ( .A1(n8745), .A2(n8744), .A3(n10074), .ZN(n8749) );
  NAND2_X1 U10159 ( .A1(n8746), .A2(n10032), .ZN(n8747) );
  MUX2_X1 U10160 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8869), .S(n10082), .Z(
        P2_U3549) );
  NAND2_X1 U10161 ( .A1(n8753), .A2(n10074), .ZN(n8759) );
  INV_X1 U10162 ( .A(n8754), .ZN(n8757) );
  NAND3_X1 U10163 ( .A1(n8530), .A2(n8759), .A3(n8758), .ZN(n8870) );
  MUX2_X1 U10164 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8870), .S(n10082), .Z(
        P2_U3548) );
  AOI21_X1 U10165 ( .B1(n8840), .B2(n8762), .A(n8761), .ZN(n8763) );
  MUX2_X1 U10166 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8871), .S(n10082), .Z(
        P2_U3546) );
  MUX2_X1 U10167 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8872), .S(n10082), .Z(
        P2_U3545) );
  AOI22_X1 U10168 ( .A1(n8777), .A2(n8861), .B1(n8840), .B2(n8776), .ZN(n8778)
         );
  OAI211_X1 U10169 ( .C1(n8849), .C2(n8780), .A(n8779), .B(n8778), .ZN(n8873)
         );
  MUX2_X1 U10170 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8873), .S(n10082), .Z(
        P2_U3544) );
  AOI22_X1 U10171 ( .A1(n8782), .A2(n8861), .B1(n10032), .B2(n8781), .ZN(n8783) );
  OAI211_X1 U10172 ( .C1(n8785), .C2(n8849), .A(n8784), .B(n8783), .ZN(n8874)
         );
  MUX2_X1 U10173 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8874), .S(n10082), .Z(
        P2_U3543) );
  AOI22_X1 U10174 ( .A1(n8787), .A2(n8861), .B1(n8840), .B2(n8786), .ZN(n8788)
         );
  OAI211_X1 U10175 ( .C1(n8790), .C2(n8849), .A(n8789), .B(n8788), .ZN(n8875)
         );
  MUX2_X1 U10176 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8875), .S(n10082), .Z(
        P2_U3542) );
  AOI211_X1 U10177 ( .C1(n8840), .C2(n8793), .A(n8792), .B(n8791), .ZN(n8794)
         );
  OAI21_X1 U10178 ( .B1(n8849), .B2(n8795), .A(n8794), .ZN(n8876) );
  MUX2_X1 U10179 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8876), .S(n10082), .Z(
        P2_U3541) );
  AOI22_X1 U10180 ( .A1(n8797), .A2(n8861), .B1(n8840), .B2(n8796), .ZN(n8798)
         );
  OAI211_X1 U10181 ( .C1(n8849), .C2(n8800), .A(n8799), .B(n8798), .ZN(n8877)
         );
  MUX2_X1 U10182 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8877), .S(n10082), .Z(
        P2_U3540) );
  AOI21_X1 U10183 ( .B1(n8840), .B2(n8802), .A(n8801), .ZN(n8803) );
  OAI21_X1 U10184 ( .B1(n8804), .B2(n8849), .A(n8803), .ZN(n8878) );
  MUX2_X1 U10185 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8878), .S(n10082), .Z(
        P2_U3539) );
  AOI22_X1 U10186 ( .A1(n8806), .A2(n8861), .B1(n10032), .B2(n8805), .ZN(n8807) );
  OAI211_X1 U10187 ( .C1(n8849), .C2(n8809), .A(n8808), .B(n8807), .ZN(n8879)
         );
  MUX2_X1 U10188 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8879), .S(n10082), .Z(
        P2_U3538) );
  AOI21_X1 U10189 ( .B1(n8840), .B2(n8811), .A(n8810), .ZN(n8812) );
  OAI211_X1 U10190 ( .C1(n8814), .C2(n8849), .A(n8813), .B(n8812), .ZN(n8880)
         );
  MUX2_X1 U10191 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8880), .S(n10082), .Z(
        P2_U3537) );
  INV_X1 U10192 ( .A(n8866), .ZN(n8819) );
  OAI22_X1 U10193 ( .A1(n8817), .A2(n8816), .B1(n8815), .B2(n10070), .ZN(n8818) );
  AOI21_X1 U10194 ( .B1(n8820), .B2(n8819), .A(n8818), .ZN(n8821) );
  NAND2_X1 U10195 ( .A1(n8822), .A2(n8821), .ZN(n8881) );
  MUX2_X1 U10196 ( .A(n8881), .B(P2_REG1_REG_16__SCAN_IN), .S(n10080), .Z(
        P2_U3536) );
  AOI21_X1 U10197 ( .B1(n8840), .B2(n8824), .A(n8823), .ZN(n8825) );
  OAI211_X1 U10198 ( .C1(n8827), .C2(n8849), .A(n8826), .B(n8825), .ZN(n8882)
         );
  MUX2_X1 U10199 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8882), .S(n10082), .Z(
        P2_U3535) );
  AOI22_X1 U10200 ( .A1(n8829), .A2(n8861), .B1(n8840), .B2(n8828), .ZN(n8830)
         );
  OAI211_X1 U10201 ( .C1(n8849), .C2(n8832), .A(n8831), .B(n8830), .ZN(n8883)
         );
  MUX2_X1 U10202 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8883), .S(n10082), .Z(
        P2_U3534) );
  AOI22_X1 U10203 ( .A1(n8834), .A2(n8861), .B1(n10032), .B2(n8833), .ZN(n8835) );
  OAI211_X1 U10204 ( .C1(n8866), .C2(n8837), .A(n8836), .B(n8835), .ZN(n8884)
         );
  MUX2_X1 U10205 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8884), .S(n10082), .Z(
        P2_U3533) );
  AOI21_X1 U10206 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(n8841) );
  OAI211_X1 U10207 ( .C1(n8849), .C2(n8843), .A(n8842), .B(n8841), .ZN(n8885)
         );
  MUX2_X1 U10208 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8885), .S(n10082), .Z(
        P2_U3532) );
  AOI22_X1 U10209 ( .A1(n8845), .A2(n8861), .B1(n10032), .B2(n8844), .ZN(n8846) );
  OAI211_X1 U10210 ( .C1(n8849), .C2(n8848), .A(n8847), .B(n8846), .ZN(n8886)
         );
  MUX2_X1 U10211 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8886), .S(n10082), .Z(
        P2_U3531) );
  AOI22_X1 U10212 ( .A1(n8851), .A2(n8861), .B1(n10032), .B2(n8850), .ZN(n8852) );
  OAI211_X1 U10213 ( .C1(n8866), .C2(n8854), .A(n8853), .B(n8852), .ZN(n8887)
         );
  MUX2_X1 U10214 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n8887), .S(n10082), .Z(
        P2_U3530) );
  AOI22_X1 U10215 ( .A1(n8856), .A2(n8861), .B1(n10032), .B2(n8855), .ZN(n8857) );
  OAI211_X1 U10216 ( .C1(n8859), .C2(n8866), .A(n8858), .B(n8857), .ZN(n8888)
         );
  MUX2_X1 U10217 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8888), .S(n10082), .Z(
        P2_U3529) );
  AOI22_X1 U10218 ( .A1(n8862), .A2(n8861), .B1(n10032), .B2(n8860), .ZN(n8863) );
  OAI211_X1 U10219 ( .C1(n8866), .C2(n8865), .A(n8864), .B(n8863), .ZN(n8889)
         );
  MUX2_X1 U10220 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n8889), .S(n10082), .Z(
        P2_U3528) );
  MUX2_X1 U10221 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8867), .S(n10076), .Z(
        P2_U3519) );
  MUX2_X1 U10222 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8868), .S(n10076), .Z(
        P2_U3518) );
  MUX2_X1 U10223 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8869), .S(n10076), .Z(
        P2_U3517) );
  MUX2_X1 U10224 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8870), .S(n10076), .Z(
        P2_U3516) );
  MUX2_X1 U10225 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8871), .S(n10076), .Z(
        P2_U3514) );
  MUX2_X1 U10226 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8872), .S(n10076), .Z(
        P2_U3513) );
  MUX2_X1 U10227 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8873), .S(n10076), .Z(
        P2_U3512) );
  MUX2_X1 U10228 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8874), .S(n10076), .Z(
        P2_U3511) );
  MUX2_X1 U10229 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8875), .S(n10076), .Z(
        P2_U3510) );
  MUX2_X1 U10230 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8876), .S(n10076), .Z(
        P2_U3509) );
  MUX2_X1 U10231 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8877), .S(n10076), .Z(
        P2_U3508) );
  MUX2_X1 U10232 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8878), .S(n10076), .Z(
        P2_U3507) );
  MUX2_X1 U10233 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8879), .S(n10076), .Z(
        P2_U3505) );
  MUX2_X1 U10234 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8880), .S(n10076), .Z(
        P2_U3502) );
  MUX2_X1 U10235 ( .A(n8881), .B(P2_REG0_REG_16__SCAN_IN), .S(n10075), .Z(
        P2_U3499) );
  MUX2_X1 U10236 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8882), .S(n10076), .Z(
        P2_U3496) );
  MUX2_X1 U10237 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8883), .S(n10076), .Z(
        P2_U3493) );
  MUX2_X1 U10238 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8884), .S(n10076), .Z(
        P2_U3490) );
  MUX2_X1 U10239 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n8885), .S(n10076), .Z(
        P2_U3487) );
  MUX2_X1 U10240 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8886), .S(n10076), .Z(
        P2_U3484) );
  MUX2_X1 U10241 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n8887), .S(n10076), .Z(
        P2_U3481) );
  MUX2_X1 U10242 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n8888), .S(n10076), .Z(
        P2_U3478) );
  MUX2_X1 U10243 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n8889), .S(n10076), .Z(
        P2_U3475) );
  INV_X1 U10244 ( .A(n8890), .ZN(n9765) );
  NAND2_X1 U10245 ( .A1(n8891), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8892) );
  OAI211_X1 U10246 ( .C1(n9765), .C2(n8894), .A(n8893), .B(n8892), .ZN(
        P2_U3330) );
  INV_X1 U10247 ( .A(n8895), .ZN(n9768) );
  OAI222_X1 U10248 ( .A1(n8897), .A2(P2_U3152), .B1(n8894), .B2(n9768), .C1(
        n8896), .C2(n8904), .ZN(P2_U3331) );
  INV_X1 U10249 ( .A(n8898), .ZN(n9770) );
  OAI222_X1 U10250 ( .A1(P2_U3152), .A2(n8900), .B1(n8894), .B2(n9770), .C1(
        n8899), .C2(n8904), .ZN(P2_U3332) );
  INV_X1 U10251 ( .A(n8901), .ZN(n9775) );
  OAI222_X1 U10252 ( .A1(n8904), .A2(n8903), .B1(n8894), .B2(n9775), .C1(
        P2_U3152), .C2(n8902), .ZN(P2_U3333) );
  MUX2_X1 U10253 ( .A(n8905), .B(n4407), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10254 ( .A(n8906), .ZN(n8909) );
  NAND2_X1 U10255 ( .A1(n9636), .A2(n8967), .ZN(n8911) );
  NAND2_X1 U10256 ( .A1(n9126), .A2(n8961), .ZN(n8910) );
  NAND2_X1 U10257 ( .A1(n8911), .A2(n8910), .ZN(n8912) );
  XNOR2_X1 U10258 ( .A(n8912), .B(n8916), .ZN(n8915) );
  NOR2_X1 U10259 ( .A1(n9307), .A2(n6047), .ZN(n8913) );
  AOI21_X1 U10260 ( .B1(n9636), .B2(n8961), .A(n8913), .ZN(n8914) );
  NOR2_X1 U10261 ( .A1(n8915), .A2(n8914), .ZN(n9099) );
  INV_X1 U10262 ( .A(n9631), .ZN(n9378) );
  OAI22_X1 U10263 ( .A1(n9378), .A2(n8969), .B1(n4281), .B2(n6047), .ZN(n8974)
         );
  XNOR2_X1 U10264 ( .A(n8917), .B(n8916), .ZN(n8973) );
  XOR2_X1 U10265 ( .A(n8974), .B(n8973), .Z(n8918) );
  XNOR2_X1 U10266 ( .A(n8960), .B(n8918), .ZN(n8922) );
  AOI22_X1 U10267 ( .A1(n9348), .A2(n9116), .B1(n9347), .B2(n9126), .ZN(n9382)
         );
  AOI22_X1 U10268 ( .A1(n9376), .A2(n9104), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8919) );
  OAI21_X1 U10269 ( .B1(n9382), .B2(n9106), .A(n8919), .ZN(n8920) );
  AOI21_X1 U10270 ( .B1(n9631), .B2(n9121), .A(n8920), .ZN(n8921) );
  OAI21_X1 U10271 ( .B1(n8922), .B2(n9110), .A(n8921), .ZN(P1_U3212) );
  XNOR2_X1 U10272 ( .A(n8924), .B(n8923), .ZN(n8925) );
  XNOR2_X1 U10273 ( .A(n8926), .B(n8925), .ZN(n8931) );
  AOI22_X1 U10274 ( .A1(n9279), .A2(n9116), .B1(n9347), .B2(n9274), .ZN(n9574)
         );
  OAI22_X1 U10275 ( .A1(n9574), .A2(n9106), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8927), .ZN(n8929) );
  INV_X1 U10276 ( .A(n9708), .ZN(n9581) );
  NOR2_X1 U10277 ( .A1(n9581), .A2(n9098), .ZN(n8928) );
  AOI211_X1 U10278 ( .C1(n9104), .C2(n9578), .A(n8929), .B(n8928), .ZN(n8930)
         );
  OAI21_X1 U10279 ( .B1(n8931), .B2(n9110), .A(n8930), .ZN(P1_U3213) );
  INV_X1 U10280 ( .A(n8932), .ZN(n8934) );
  NAND2_X1 U10281 ( .A1(n8934), .A2(n8933), .ZN(n8936) );
  XNOR2_X1 U10282 ( .A(n8936), .B(n8935), .ZN(n8942) );
  OAI22_X1 U10283 ( .A1(n9302), .A2(n9260), .B1(n9296), .B2(n9102), .ZN(n9655)
         );
  OAI22_X1 U10284 ( .A1(n9441), .A2(n9842), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8937), .ZN(n8940) );
  NAND2_X1 U10285 ( .A1(n9433), .A2(n9726), .ZN(n9656) );
  NOR2_X1 U10286 ( .A1(n9656), .A2(n8938), .ZN(n8939) );
  AOI211_X1 U10287 ( .C1(n9832), .C2(n9655), .A(n8940), .B(n8939), .ZN(n8941)
         );
  OAI21_X1 U10288 ( .B1(n8942), .B2(n9110), .A(n8941), .ZN(P1_U3214) );
  INV_X1 U10289 ( .A(n9678), .ZN(n9495) );
  NOR2_X1 U10290 ( .A1(n8943), .A2(n8944), .ZN(n9088) );
  NOR2_X1 U10291 ( .A1(n9088), .A2(n9087), .ZN(n8947) );
  XNOR2_X1 U10292 ( .A(n8946), .B(n8945), .ZN(n8948) );
  NOR3_X1 U10293 ( .A1(n8947), .A2(n9090), .A3(n8948), .ZN(n8952) );
  INV_X1 U10294 ( .A(n8947), .ZN(n9091) );
  INV_X1 U10295 ( .A(n9090), .ZN(n8950) );
  INV_X1 U10296 ( .A(n8948), .ZN(n8949) );
  AOI21_X1 U10297 ( .B1(n9091), .B2(n8950), .A(n8949), .ZN(n8951) );
  OAI21_X1 U10298 ( .B1(n8952), .B2(n8951), .A(n9838), .ZN(n8957) );
  OAI22_X1 U10299 ( .A1(n9290), .A2(n9260), .B1(n9285), .B2(n9102), .ZN(n9498)
         );
  NOR2_X1 U10300 ( .A1(n9842), .A2(n8953), .ZN(n8955) );
  NOR2_X1 U10301 ( .A1(n8954), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9254) );
  AOI211_X1 U10302 ( .C1(n9498), .C2(n9832), .A(n8955), .B(n9254), .ZN(n8956)
         );
  OAI211_X1 U10303 ( .C1(n9495), .C2(n9098), .A(n8957), .B(n8956), .ZN(
        P1_U3217) );
  INV_X1 U10304 ( .A(n8974), .ZN(n8958) );
  NAND2_X1 U10305 ( .A1(n9625), .A2(n8961), .ZN(n8964) );
  NAND2_X1 U10306 ( .A1(n9348), .A2(n8962), .ZN(n8963) );
  NAND2_X1 U10307 ( .A1(n8964), .A2(n8963), .ZN(n8966) );
  XNOR2_X1 U10308 ( .A(n8966), .B(n8965), .ZN(n8972) );
  NAND2_X1 U10309 ( .A1(n9625), .A2(n8967), .ZN(n8968) );
  OAI21_X1 U10310 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(n8971) );
  XNOR2_X1 U10311 ( .A(n8972), .B(n8971), .ZN(n8976) );
  INV_X1 U10312 ( .A(n8976), .ZN(n8982) );
  INV_X1 U10313 ( .A(n8973), .ZN(n8975) );
  NAND2_X1 U10314 ( .A1(n8975), .A2(n8974), .ZN(n8981) );
  NAND3_X1 U10315 ( .A1(n8982), .A2(n8981), .A3(n9838), .ZN(n8987) );
  NAND3_X1 U10316 ( .A1(n8988), .A2(n9838), .A3(n8976), .ZN(n8986) );
  OR2_X1 U10317 ( .A1(n4281), .A2(n9102), .ZN(n8977) );
  OAI21_X1 U10318 ( .B1(n8978), .B2(n9260), .A(n8977), .ZN(n9364) );
  INV_X1 U10319 ( .A(n8979), .ZN(n9369) );
  AOI22_X1 U10320 ( .A1(n9369), .A2(n9104), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8980) );
  OAI21_X1 U10321 ( .B1(n4496), .B2(n9106), .A(n8980), .ZN(n8984) );
  NOR3_X1 U10322 ( .A1(n8982), .A2(n8981), .A3(n9110), .ZN(n8983) );
  AOI211_X1 U10323 ( .C1(n9121), .C2(n9625), .A(n8984), .B(n8983), .ZN(n8985)
         );
  OAI211_X1 U10324 ( .C1(n8988), .C2(n8987), .A(n8986), .B(n8985), .ZN(
        P1_U3218) );
  INV_X1 U10325 ( .A(n8989), .ZN(n8991) );
  NOR2_X1 U10326 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  XNOR2_X1 U10327 ( .A(n8993), .B(n8992), .ZN(n8998) );
  OAI22_X1 U10328 ( .A1(n9296), .A2(n9260), .B1(n9290), .B2(n9102), .ZN(n9467)
         );
  OAI22_X1 U10329 ( .A1(n9473), .A2(n9842), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8994), .ZN(n8995) );
  AOI21_X1 U10330 ( .B1(n9467), .B2(n9832), .A(n8995), .ZN(n8997) );
  NAND2_X1 U10331 ( .A1(n9669), .A2(n9121), .ZN(n8996) );
  OAI211_X1 U10332 ( .C1(n8998), .C2(n9110), .A(n8997), .B(n8996), .ZN(
        P1_U3221) );
  INV_X1 U10333 ( .A(n8999), .ZN(n9000) );
  AOI21_X1 U10334 ( .B1(n9002), .B2(n9001), .A(n9000), .ZN(n9009) );
  INV_X1 U10335 ( .A(n9003), .ZN(n9004) );
  AOI22_X1 U10336 ( .A1(n9004), .A2(n9832), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n9005) );
  OAI21_X1 U10337 ( .B1(n9006), .B2(n9842), .A(n9005), .ZN(n9007) );
  AOI21_X1 U10338 ( .B1(n9717), .B2(n9121), .A(n9007), .ZN(n9008) );
  OAI21_X1 U10339 ( .B1(n9009), .B2(n9110), .A(n9008), .ZN(P1_U3222) );
  AND2_X1 U10340 ( .A1(n9011), .A2(n9010), .ZN(n9112) );
  NOR2_X1 U10341 ( .A1(n9112), .A2(n9012), .ZN(n9017) );
  NAND2_X1 U10342 ( .A1(n9026), .A2(n9015), .ZN(n9016) );
  NOR3_X1 U10343 ( .A1(n9017), .A2(n9113), .A3(n9016), .ZN(n9029) );
  OAI21_X1 U10344 ( .B1(n9017), .B2(n9113), .A(n9016), .ZN(n9018) );
  INV_X1 U10345 ( .A(n9018), .ZN(n9019) );
  OAI21_X1 U10346 ( .B1(n9029), .B2(n9019), .A(n9838), .ZN(n9025) );
  OAI22_X1 U10347 ( .A1(n9021), .A2(n9260), .B1(n9102), .B2(n9020), .ZN(n9546)
         );
  NOR2_X1 U10348 ( .A1(n9022), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9218) );
  NOR2_X1 U10349 ( .A1(n9842), .A2(n9537), .ZN(n9023) );
  AOI211_X1 U10350 ( .C1(n9832), .C2(n9546), .A(n9218), .B(n9023), .ZN(n9024)
         );
  OAI211_X1 U10351 ( .C1(n9540), .C2(n9098), .A(n9025), .B(n9024), .ZN(
        P1_U3224) );
  INV_X1 U10352 ( .A(n9026), .ZN(n9028) );
  NOR3_X1 U10353 ( .A1(n9029), .A2(n9028), .A3(n9027), .ZN(n9032) );
  INV_X1 U10354 ( .A(n9030), .ZN(n9031) );
  OAI21_X1 U10355 ( .B1(n9032), .B2(n9031), .A(n9838), .ZN(n9036) );
  OAI22_X1 U10356 ( .A1(n9285), .A2(n9260), .B1(n9033), .B2(n9102), .ZN(n9521)
         );
  AND2_X1 U10357 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9873) );
  NOR2_X1 U10358 ( .A1(n9842), .A2(n9524), .ZN(n9034) );
  AOI211_X1 U10359 ( .C1(n9832), .C2(n9521), .A(n9873), .B(n9034), .ZN(n9035)
         );
  OAI211_X1 U10360 ( .C1(n9690), .C2(n9098), .A(n9036), .B(n9035), .ZN(
        P1_U3226) );
  AOI21_X1 U10361 ( .B1(n9039), .B2(n9038), .A(n9037), .ZN(n9044) );
  AND2_X1 U10362 ( .A1(n9417), .A2(n9726), .ZN(n9650) );
  NOR2_X1 U10363 ( .A1(n9298), .A2(n9102), .ZN(n9040) );
  AOI21_X1 U10364 ( .B1(n9127), .B2(n9116), .A(n9040), .ZN(n9425) );
  AOI22_X1 U10365 ( .A1(n9426), .A2(n9104), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9041) );
  OAI21_X1 U10366 ( .B1(n9425), .B2(n9106), .A(n9041), .ZN(n9042) );
  AOI21_X1 U10367 ( .B1(n9650), .B2(n9837), .A(n9042), .ZN(n9043) );
  OAI21_X1 U10368 ( .B1(n9044), .B2(n9110), .A(n9043), .ZN(P1_U3227) );
  NAND2_X1 U10369 ( .A1(n4308), .A2(n9045), .ZN(n9046) );
  XNOR2_X1 U10370 ( .A(n9047), .B(n9046), .ZN(n9051) );
  AOI22_X1 U10371 ( .A1(n9294), .A2(n9116), .B1(n9347), .B2(n9287), .ZN(n9480)
         );
  OAI22_X1 U10372 ( .A1(n9480), .A2(n9106), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n4547), .ZN(n9049) );
  INV_X1 U10373 ( .A(n9675), .ZN(n9486) );
  NOR2_X1 U10374 ( .A1(n9486), .A2(n9098), .ZN(n9048) );
  AOI211_X1 U10375 ( .C1(n9104), .C2(n9483), .A(n9049), .B(n9048), .ZN(n9050)
         );
  OAI21_X1 U10376 ( .B1(n9051), .B2(n9110), .A(n9050), .ZN(P1_U3231) );
  XNOR2_X1 U10377 ( .A(n9053), .B(n9052), .ZN(n9054) );
  XNOR2_X1 U10378 ( .A(n9055), .B(n9054), .ZN(n9064) );
  INV_X1 U10379 ( .A(n9056), .ZN(n9270) );
  NAND2_X1 U10380 ( .A1(n9347), .A2(n9270), .ZN(n9059) );
  OR2_X1 U10381 ( .A1(n9260), .A2(n9057), .ZN(n9058) );
  NAND2_X1 U10382 ( .A1(n9059), .A2(n9058), .ZN(n9592) );
  AOI21_X1 U10383 ( .B1(n9592), .B2(n9832), .A(n9060), .ZN(n9061) );
  OAI21_X1 U10384 ( .B1(n9842), .B2(n9596), .A(n9061), .ZN(n9062) );
  AOI21_X1 U10385 ( .B1(n9712), .B2(n9121), .A(n9062), .ZN(n9063) );
  OAI21_X1 U10386 ( .B1(n9064), .B2(n9110), .A(n9063), .ZN(P1_U3232) );
  INV_X1 U10387 ( .A(n9065), .ZN(n9066) );
  NOR2_X1 U10388 ( .A1(n9067), .A2(n9066), .ZN(n9069) );
  XNOR2_X1 U10389 ( .A(n9069), .B(n9068), .ZN(n9076) );
  OAI22_X1 U10390 ( .A1(n9298), .A2(n9260), .B1(n9070), .B2(n9102), .ZN(n9457)
         );
  INV_X1 U10391 ( .A(n9452), .ZN(n9072) );
  OAI22_X1 U10392 ( .A1(n9072), .A2(n9842), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9071), .ZN(n9073) );
  AOI21_X1 U10393 ( .B1(n9457), .B2(n9832), .A(n9073), .ZN(n9075) );
  NAND2_X1 U10394 ( .A1(n9663), .A2(n9121), .ZN(n9074) );
  OAI211_X1 U10395 ( .C1(n9076), .C2(n9110), .A(n9075), .B(n9074), .ZN(
        P1_U3233) );
  AOI22_X1 U10396 ( .A1(n9077), .A2(n9832), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3084), .ZN(n9078) );
  OAI21_X1 U10397 ( .B1(n9842), .B2(n9079), .A(n9078), .ZN(n9085) );
  INV_X1 U10398 ( .A(n9080), .ZN(n9081) );
  AOI211_X1 U10399 ( .C1(n9083), .C2(n9082), .A(n9110), .B(n9081), .ZN(n9084)
         );
  AOI211_X1 U10400 ( .C1(n9121), .C2(n9725), .A(n9085), .B(n9084), .ZN(n9086)
         );
  INV_X1 U10401 ( .A(n9086), .ZN(P1_U3234) );
  OAI21_X1 U10402 ( .B1(n9088), .B2(n9090), .A(n9087), .ZN(n9089) );
  OAI21_X1 U10403 ( .B1(n9091), .B2(n9090), .A(n9089), .ZN(n9092) );
  NAND2_X1 U10404 ( .A1(n9092), .A2(n9838), .ZN(n9097) );
  INV_X1 U10405 ( .A(n9093), .ZN(n9509) );
  AOI22_X1 U10406 ( .A1(n9287), .A2(n9116), .B1(n9347), .B2(n9284), .ZN(n9506)
         );
  OAI22_X1 U10407 ( .A1(n9506), .A2(n9106), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9094), .ZN(n9095) );
  AOI21_X1 U10408 ( .B1(n9509), .B2(n9104), .A(n9095), .ZN(n9096) );
  OAI211_X1 U10409 ( .C1(n9685), .C2(n9098), .A(n9097), .B(n9096), .ZN(
        P1_U3236) );
  NOR2_X1 U10410 ( .A1(n9099), .A2(n4383), .ZN(n9100) );
  XNOR2_X1 U10411 ( .A(n9101), .B(n9100), .ZN(n9111) );
  OAI22_X1 U10412 ( .A1(n4281), .A2(n9260), .B1(n9306), .B2(n9102), .ZN(n9395)
         );
  INV_X1 U10413 ( .A(n9395), .ZN(n9107) );
  INV_X1 U10414 ( .A(n9103), .ZN(n9391) );
  AOI22_X1 U10415 ( .A1(n9391), .A2(n9104), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9105) );
  OAI21_X1 U10416 ( .B1(n9107), .B2(n9106), .A(n9105), .ZN(n9108) );
  AOI21_X1 U10417 ( .B1(n9636), .B2(n9121), .A(n9108), .ZN(n9109) );
  OAI21_X1 U10418 ( .B1(n9111), .B2(n9110), .A(n9109), .ZN(P1_U3238) );
  NOR2_X1 U10419 ( .A1(n9113), .A2(n9112), .ZN(n9115) );
  XNOR2_X1 U10420 ( .A(n9115), .B(n9114), .ZN(n9123) );
  NAND2_X1 U10421 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U10422 ( .A1(n9282), .A2(n9116), .ZN(n9118) );
  NAND2_X1 U10423 ( .A1(n9347), .A2(n9277), .ZN(n9117) );
  NAND2_X1 U10424 ( .A1(n9118), .A2(n9117), .ZN(n9558) );
  NAND2_X1 U10425 ( .A1(n9558), .A2(n9832), .ZN(n9119) );
  OAI211_X1 U10426 ( .C1(n9842), .C2(n9561), .A(n9858), .B(n9119), .ZN(n9120)
         );
  AOI21_X1 U10427 ( .B1(n9701), .B2(n9121), .A(n9120), .ZN(n9122) );
  OAI21_X1 U10428 ( .B1(n9123), .B2(n9110), .A(n9122), .ZN(P1_U3239) );
  MUX2_X1 U10429 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9343), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10430 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9124), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10431 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9348), .S(P1_U4006), .Z(
        P1_U3583) );
  INV_X1 U10432 ( .A(n4281), .ZN(n9310) );
  MUX2_X1 U10433 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9310), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10434 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9126), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10435 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9127), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10436 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9303), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9300), .S(P1_U4006), .Z(
        P1_U3578) );
  INV_X1 U10438 ( .A(n9296), .ZN(n9295) );
  MUX2_X1 U10439 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9295), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10440 ( .A(n9294), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9129), .Z(
        P1_U3576) );
  INV_X1 U10441 ( .A(n9290), .ZN(n9291) );
  MUX2_X1 U10442 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9291), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10443 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9287), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10444 ( .A(n9128), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9129), .Z(
        P1_U3573) );
  MUX2_X1 U10445 ( .A(n9284), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9129), .Z(
        P1_U3572) );
  MUX2_X1 U10446 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9282), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10447 ( .A(n9279), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9129), .Z(
        P1_U3570) );
  MUX2_X1 U10448 ( .A(n9277), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9129), .Z(
        P1_U3569) );
  MUX2_X1 U10449 ( .A(n9274), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9129), .Z(
        P1_U3568) );
  MUX2_X1 U10450 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9270), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10451 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9130), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10452 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9131), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10453 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9132), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10454 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9133), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10455 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9134), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10456 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9135), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10457 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9136), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10458 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9137), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10459 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9138), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10460 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9139), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10461 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9140), .S(P1_U4006), .Z(
        P1_U3556) );
  OAI21_X1 U10462 ( .B1(n9142), .B2(n9141), .A(n9155), .ZN(n9144) );
  AOI22_X1 U10463 ( .A1(n9144), .A2(n9879), .B1(n9143), .B2(n9861), .ZN(n9152)
         );
  NAND2_X1 U10464 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n9151) );
  NAND2_X1 U10465 ( .A1(n9874), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n9150) );
  AND3_X1 U10466 ( .A1(n9147), .A2(n9146), .A3(n9145), .ZN(n9148) );
  OAI21_X1 U10467 ( .B1(n9164), .B2(n9148), .A(n9878), .ZN(n9149) );
  NAND4_X1 U10468 ( .A1(n9152), .A2(n9151), .A3(n9150), .A4(n9149), .ZN(
        P1_U3248) );
  AND3_X1 U10469 ( .A1(n9155), .A2(n9154), .A3(n9153), .ZN(n9156) );
  OAI21_X1 U10470 ( .B1(n9157), .B2(n9156), .A(n9879), .ZN(n9169) );
  INV_X1 U10471 ( .A(n9158), .ZN(n9159) );
  OAI21_X1 U10472 ( .B1(n9871), .B2(n9160), .A(n9159), .ZN(n9161) );
  AOI21_X1 U10473 ( .B1(n9874), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n9161), .ZN(
        n9168) );
  INV_X1 U10474 ( .A(n9178), .ZN(n9166) );
  NOR3_X1 U10475 ( .A1(n9164), .A2(n9163), .A3(n9162), .ZN(n9165) );
  OAI21_X1 U10476 ( .B1(n9166), .B2(n9165), .A(n9878), .ZN(n9167) );
  NAND3_X1 U10477 ( .A1(n9169), .A2(n9168), .A3(n9167), .ZN(P1_U3249) );
  OAI211_X1 U10478 ( .C1(n9172), .C2(n9171), .A(n9170), .B(n9879), .ZN(n9183)
         );
  NAND2_X1 U10479 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n9173) );
  OAI21_X1 U10480 ( .B1(n9871), .B2(n9174), .A(n9173), .ZN(n9175) );
  AOI21_X1 U10481 ( .B1(n9874), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9175), .ZN(
        n9182) );
  AND3_X1 U10482 ( .A1(n9178), .A2(n9177), .A3(n9176), .ZN(n9179) );
  OAI21_X1 U10483 ( .B1(n9180), .B2(n9179), .A(n9878), .ZN(n9181) );
  NAND3_X1 U10484 ( .A1(n9183), .A2(n9182), .A3(n9181), .ZN(P1_U3250) );
  OAI211_X1 U10485 ( .C1(n9186), .C2(n9185), .A(n9184), .B(n9879), .ZN(n9198)
         );
  NAND2_X1 U10486 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n9187) );
  OAI21_X1 U10487 ( .B1(n9871), .B2(n9188), .A(n9187), .ZN(n9189) );
  AOI21_X1 U10488 ( .B1(n9874), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9189), .ZN(
        n9197) );
  INV_X1 U10489 ( .A(n9190), .ZN(n9195) );
  NOR3_X1 U10490 ( .A1(n9193), .A2(n9192), .A3(n9191), .ZN(n9194) );
  OAI21_X1 U10491 ( .B1(n9195), .B2(n9194), .A(n9878), .ZN(n9196) );
  NAND3_X1 U10492 ( .A1(n9198), .A2(n9197), .A3(n9196), .ZN(P1_U3253) );
  XOR2_X1 U10493 ( .A(n9225), .B(P1_REG1_REG_16__SCAN_IN), .Z(n9206) );
  AOI21_X1 U10494 ( .B1(n9200), .B2(n10135), .A(n9199), .ZN(n9201) );
  INV_X1 U10495 ( .A(n9201), .ZN(n9203) );
  INV_X1 U10496 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9202) );
  XNOR2_X1 U10497 ( .A(n9201), .B(n9860), .ZN(n9862) );
  OAI22_X1 U10498 ( .A1(n9204), .A2(n9203), .B1(n9202), .B2(n9862), .ZN(n9205)
         );
  NAND2_X1 U10499 ( .A1(n9206), .A2(n9205), .ZN(n9226) );
  OAI211_X1 U10500 ( .C1(n9206), .C2(n9205), .A(n9226), .B(n9878), .ZN(n9216)
         );
  INV_X1 U10501 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9207) );
  MUX2_X1 U10502 ( .A(n9207), .B(P1_REG2_REG_16__SCAN_IN), .S(n9225), .Z(n9208) );
  INV_X1 U10503 ( .A(n9208), .ZN(n9214) );
  INV_X1 U10504 ( .A(n9212), .ZN(n9213) );
  NAND2_X1 U10505 ( .A1(n9214), .A2(n9213), .ZN(n9220) );
  OAI211_X1 U10506 ( .C1(n9214), .C2(n9213), .A(n9879), .B(n9220), .ZN(n9215)
         );
  NAND2_X1 U10507 ( .A1(n9216), .A2(n9215), .ZN(n9217) );
  AOI211_X1 U10508 ( .C1(n9861), .C2(n9225), .A(n9218), .B(n9217), .ZN(n9219)
         );
  OAI21_X1 U10509 ( .B1(n9241), .B2(n4455), .A(n9219), .ZN(P1_U3257) );
  INV_X1 U10510 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9240) );
  INV_X1 U10511 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U10512 ( .A1(n9225), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U10513 ( .A1(n9221), .A2(n9220), .ZN(n9882) );
  MUX2_X1 U10514 ( .A(n9525), .B(P1_REG2_REG_17__SCAN_IN), .S(n9229), .Z(n9222) );
  INV_X1 U10515 ( .A(n9222), .ZN(n9881) );
  NAND2_X1 U10516 ( .A1(n9882), .A2(n9881), .ZN(n9880) );
  OAI21_X1 U10517 ( .B1(n9525), .B2(n9870), .A(n9880), .ZN(n9224) );
  XNOR2_X1 U10518 ( .A(n9246), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n9223) );
  NAND2_X1 U10519 ( .A1(n9223), .A2(n9224), .ZN(n9242) );
  OAI211_X1 U10520 ( .C1(n9224), .C2(n9223), .A(n9879), .B(n9242), .ZN(n9239)
         );
  NAND2_X1 U10521 ( .A1(n9225), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9227) );
  NAND2_X1 U10522 ( .A1(n9227), .A2(n9226), .ZN(n9875) );
  XNOR2_X1 U10523 ( .A(n9229), .B(n9228), .ZN(n9876) );
  NAND2_X1 U10524 ( .A1(n9875), .A2(n9876), .ZN(n9231) );
  NAND2_X1 U10525 ( .A1(n9229), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U10526 ( .A1(n9231), .A2(n9230), .ZN(n9233) );
  AOI22_X1 U10527 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n9246), .B1(n9237), .B2(
        n9245), .ZN(n9232) );
  NOR2_X1 U10528 ( .A1(n9232), .A2(n9233), .ZN(n9244) );
  AOI21_X1 U10529 ( .B1(n9233), .B2(n9232), .A(n9244), .ZN(n9235) );
  NAND2_X1 U10530 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3084), .ZN(n9234) );
  OAI21_X1 U10531 ( .B1(n9235), .B2(n9249), .A(n9234), .ZN(n9236) );
  AOI21_X1 U10532 ( .B1(n9237), .B2(n9861), .A(n9236), .ZN(n9238) );
  OAI211_X1 U10533 ( .C1(n9241), .C2(n9240), .A(n9239), .B(n9238), .ZN(
        P1_U3259) );
  OAI21_X1 U10534 ( .B1(n9246), .B2(n10256), .A(n9242), .ZN(n9243) );
  AOI21_X1 U10535 ( .B1(n9246), .B2(n9245), .A(n9244), .ZN(n9248) );
  XOR2_X1 U10536 ( .A(n9248), .B(n9247), .Z(n9250) );
  AOI21_X1 U10537 ( .B1(n9250), .B2(n9878), .A(n9861), .ZN(n9251) );
  INV_X1 U10538 ( .A(n9604), .ZN(n9264) );
  INV_X1 U10539 ( .A(n9712), .ZN(n9600) );
  AND2_X2 U10540 ( .A1(n9593), .A2(n9600), .ZN(n9594) );
  NAND2_X1 U10541 ( .A1(n9508), .A2(n9685), .ZN(n9490) );
  OR2_X2 U10542 ( .A1(n9490), .A2(n9678), .ZN(n9491) );
  INV_X1 U10543 ( .A(n9669), .ZN(n9255) );
  NAND2_X1 U10544 ( .A1(n9482), .A2(n9255), .ZN(n9450) );
  NOR2_X2 U10545 ( .A1(n9418), .A2(n9402), .ZN(n9388) );
  NAND2_X1 U10546 ( .A1(n9607), .A2(n9919), .ZN(n9263) );
  NOR2_X1 U10547 ( .A1(n9258), .A2(n9257), .ZN(n9259) );
  NOR2_X1 U10548 ( .A1(n9260), .A2(n9259), .ZN(n9342) );
  NAND2_X1 U10549 ( .A1(n9342), .A2(n9261), .ZN(n9612) );
  NOR2_X1 U10550 ( .A1(n9925), .A2(n9612), .ZN(n9268) );
  AOI21_X1 U10551 ( .B1(n9603), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9268), .ZN(
        n9262) );
  OAI211_X1 U10552 ( .C1(n9264), .C2(n9899), .A(n9263), .B(n9262), .ZN(
        P1_U3261) );
  INV_X1 U10553 ( .A(n9610), .ZN(n9266) );
  INV_X1 U10554 ( .A(n9352), .ZN(n9265) );
  NOR2_X1 U10555 ( .A1(n9266), .A2(n9899), .ZN(n9267) );
  AOI211_X1 U10556 ( .C1(n9603), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9268), .B(
        n9267), .ZN(n9269) );
  OAI21_X1 U10557 ( .B1(n9527), .B2(n9613), .A(n9269), .ZN(P1_U3262) );
  NAND2_X1 U10558 ( .A1(n9717), .A2(n9270), .ZN(n9271) );
  NAND2_X1 U10559 ( .A1(n9272), .A2(n9271), .ZN(n9586) );
  OR2_X1 U10560 ( .A1(n9712), .A2(n9274), .ZN(n9273) );
  NAND2_X1 U10561 ( .A1(n9712), .A2(n9274), .ZN(n9275) );
  AND2_X1 U10562 ( .A1(n9708), .A2(n9277), .ZN(n9278) );
  NAND2_X1 U10563 ( .A1(n9701), .A2(n9279), .ZN(n9280) );
  AND2_X1 U10564 ( .A1(n9697), .A2(n9282), .ZN(n9283) );
  NAND2_X1 U10565 ( .A1(n9495), .A2(n9286), .ZN(n9289) );
  NOR2_X1 U10566 ( .A1(n9663), .A2(n9295), .ZN(n9297) );
  INV_X1 U10567 ( .A(n9433), .ZN(n9299) );
  NAND2_X1 U10568 ( .A1(n9299), .A2(n9298), .ZN(n9301) );
  NAND2_X1 U10569 ( .A1(n9416), .A2(n4976), .ZN(n9305) );
  NAND2_X1 U10570 ( .A1(n9305), .A2(n9304), .ZN(n9400) );
  NOR2_X1 U10571 ( .A1(n7952), .A2(n9307), .ZN(n9309) );
  INV_X1 U10572 ( .A(n9380), .ZN(n9311) );
  NAND2_X1 U10573 ( .A1(n9625), .A2(n9348), .ZN(n9619) );
  XNOR2_X1 U10574 ( .A(n4969), .B(n9620), .ZN(n9359) );
  NAND2_X1 U10575 ( .A1(n9313), .A2(n9312), .ZN(n9588) );
  INV_X1 U10576 ( .A(n9588), .ZN(n9315) );
  NAND2_X1 U10577 ( .A1(n9318), .A2(n9317), .ZN(n9320) );
  NAND2_X1 U10578 ( .A1(n9497), .A2(n9496), .ZN(n9325) );
  NAND2_X1 U10579 ( .A1(n9332), .A2(n9331), .ZN(n9438) );
  NAND2_X1 U10580 ( .A1(n9381), .A2(n9380), .ZN(n9379) );
  NAND2_X1 U10581 ( .A1(n9379), .A2(n9340), .ZN(n9363) );
  INV_X1 U10582 ( .A(n9342), .ZN(n9345) );
  NOR2_X1 U10583 ( .A1(n9345), .A2(n9344), .ZN(n9346) );
  INV_X1 U10584 ( .A(n9367), .ZN(n9350) );
  NAND2_X1 U10585 ( .A1(n9614), .A2(n9350), .ZN(n9351) );
  INV_X1 U10586 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9353) );
  OAI22_X1 U10587 ( .A1(n9354), .A2(n9814), .B1(n9353), .B2(n9583), .ZN(n9355)
         );
  AOI21_X1 U10588 ( .B1(n9614), .B2(n9921), .A(n9355), .ZN(n9356) );
  OAI21_X1 U10589 ( .B1(n9615), .B2(n9527), .A(n9356), .ZN(n9357) );
  AOI21_X1 U10590 ( .B1(n9618), .B2(n9583), .A(n9357), .ZN(n9358) );
  OAI21_X1 U10591 ( .B1(n9359), .B2(n9585), .A(n9358), .ZN(P1_U3355) );
  NAND2_X1 U10592 ( .A1(n9361), .A2(n9622), .ZN(n9630) );
  XNOR2_X1 U10593 ( .A(n9363), .B(n9362), .ZN(n9365) );
  INV_X1 U10594 ( .A(n9627), .ZN(n9373) );
  INV_X1 U10595 ( .A(n9366), .ZN(n9368) );
  AOI211_X1 U10596 ( .C1(n9625), .C2(n9368), .A(n9977), .B(n9367), .ZN(n9626)
         );
  NAND2_X1 U10597 ( .A1(n9626), .A2(n9819), .ZN(n9371) );
  AOI22_X1 U10598 ( .A1(n9369), .A2(n9924), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9603), .ZN(n9370) );
  OAI211_X1 U10599 ( .C1(n9629), .C2(n9899), .A(n9371), .B(n9370), .ZN(n9372)
         );
  AOI21_X1 U10600 ( .B1(n9373), .B2(n9583), .A(n9372), .ZN(n9374) );
  OAI21_X1 U10601 ( .B1(n9630), .B2(n9585), .A(n9374), .ZN(P1_U3263) );
  XNOR2_X1 U10602 ( .A(n9375), .B(n9380), .ZN(n9635) );
  AOI21_X1 U10603 ( .B1(n9631), .B2(n9389), .A(n9366), .ZN(n9632) );
  AOI22_X1 U10604 ( .A1(n9376), .A2(n9924), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9603), .ZN(n9377) );
  OAI21_X1 U10605 ( .B1(n9378), .B2(n9899), .A(n9377), .ZN(n9385) );
  OAI211_X1 U10606 ( .C1(n9381), .C2(n9380), .A(n9379), .B(n9553), .ZN(n9383)
         );
  NOR2_X1 U10607 ( .A1(n9634), .A2(n9925), .ZN(n9384) );
  AOI211_X1 U10608 ( .C1(n9919), .C2(n9632), .A(n9385), .B(n9384), .ZN(n9386)
         );
  OAI21_X1 U10609 ( .B1(n9635), .B2(n9585), .A(n9386), .ZN(P1_U3264) );
  XOR2_X1 U10610 ( .A(n9393), .B(n9387), .Z(n9640) );
  INV_X1 U10611 ( .A(n9389), .ZN(n9390) );
  AOI21_X1 U10612 ( .B1(n9636), .B2(n9406), .A(n9390), .ZN(n9637) );
  AOI22_X1 U10613 ( .A1(n9391), .A2(n9924), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9603), .ZN(n9392) );
  OAI21_X1 U10614 ( .B1(n7952), .B2(n9899), .A(n9392), .ZN(n9398) );
  XNOR2_X1 U10615 ( .A(n9394), .B(n9393), .ZN(n9396) );
  AOI21_X1 U10616 ( .B1(n9396), .B2(n9553), .A(n9395), .ZN(n9639) );
  NOR2_X1 U10617 ( .A1(n9639), .A2(n9603), .ZN(n9397) );
  AOI211_X1 U10618 ( .C1(n9637), .C2(n9919), .A(n9398), .B(n9397), .ZN(n9399)
         );
  OAI21_X1 U10619 ( .B1(n9640), .B2(n9585), .A(n9399), .ZN(P1_U3265) );
  XNOR2_X1 U10620 ( .A(n9401), .B(n9403), .ZN(n9646) );
  INV_X1 U10621 ( .A(n9646), .ZN(n9415) );
  AOI22_X1 U10622 ( .A1(n9402), .A2(n9921), .B1(n9925), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n9414) );
  XNOR2_X1 U10623 ( .A(n9404), .B(n9403), .ZN(n9405) );
  NAND2_X1 U10624 ( .A1(n9405), .A2(n9553), .ZN(n9644) );
  INV_X1 U10625 ( .A(n9644), .ZN(n9412) );
  INV_X1 U10626 ( .A(n9418), .ZN(n9408) );
  OAI211_X1 U10627 ( .C1(n9408), .C2(n9407), .A(n9986), .B(n9406), .ZN(n9642)
         );
  NAND2_X1 U10628 ( .A1(n9409), .A2(n9924), .ZN(n9410) );
  OAI211_X1 U10629 ( .C1(n9642), .C2(n9444), .A(n9643), .B(n9410), .ZN(n9411)
         );
  OAI21_X1 U10630 ( .B1(n9412), .B2(n9411), .A(n9583), .ZN(n9413) );
  OAI211_X1 U10631 ( .C1(n9415), .C2(n9585), .A(n9414), .B(n9413), .ZN(
        P1_U3266) );
  XOR2_X1 U10632 ( .A(n9424), .B(n9416), .Z(n9648) );
  INV_X1 U10633 ( .A(n9648), .ZN(n9431) );
  AOI22_X1 U10634 ( .A1(n9417), .A2(n9921), .B1(n9603), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9430) );
  OAI211_X1 U10635 ( .C1(n9419), .C2(n9436), .A(n9986), .B(n9418), .ZN(n9651)
         );
  NAND2_X1 U10636 ( .A1(n9439), .A2(n9420), .ZN(n9423) );
  NAND2_X1 U10637 ( .A1(n9421), .A2(n4918), .ZN(n9422) );
  OAI211_X1 U10638 ( .C1(n9424), .C2(n9423), .A(n9422), .B(n9553), .ZN(n9652)
         );
  INV_X1 U10639 ( .A(n9425), .ZN(n9649) );
  AOI21_X1 U10640 ( .B1(n9426), .B2(n9924), .A(n9649), .ZN(n9427) );
  OAI211_X1 U10641 ( .C1(n9444), .C2(n9651), .A(n9652), .B(n9427), .ZN(n9428)
         );
  NAND2_X1 U10642 ( .A1(n9428), .A2(n9583), .ZN(n9429) );
  OAI211_X1 U10643 ( .C1(n9431), .C2(n9585), .A(n9430), .B(n9429), .ZN(
        P1_U3267) );
  XOR2_X1 U10644 ( .A(n9432), .B(n9437), .Z(n9661) );
  INV_X1 U10645 ( .A(n9661), .ZN(n9448) );
  AOI22_X1 U10646 ( .A1(n9433), .A2(n9921), .B1(n9603), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9447) );
  NAND2_X1 U10647 ( .A1(n9433), .A2(n9451), .ZN(n9434) );
  NAND2_X1 U10648 ( .A1(n9434), .A2(n9986), .ZN(n9435) );
  OR2_X1 U10649 ( .A1(n9436), .A2(n9435), .ZN(n9657) );
  AOI21_X1 U10650 ( .B1(n9438), .B2(n9437), .A(n9908), .ZN(n9440) );
  NAND2_X1 U10651 ( .A1(n9440), .A2(n9439), .ZN(n9659) );
  INV_X1 U10652 ( .A(n9441), .ZN(n9442) );
  AOI21_X1 U10653 ( .B1(n9442), .B2(n9924), .A(n9655), .ZN(n9443) );
  OAI211_X1 U10654 ( .C1(n9444), .C2(n9657), .A(n9659), .B(n9443), .ZN(n9445)
         );
  NAND2_X1 U10655 ( .A1(n9445), .A2(n9583), .ZN(n9446) );
  OAI211_X1 U10656 ( .C1(n9448), .C2(n9585), .A(n9447), .B(n9446), .ZN(
        P1_U3268) );
  XOR2_X1 U10657 ( .A(n9455), .B(n9449), .Z(n9667) );
  AOI21_X1 U10658 ( .B1(n9663), .B2(n9450), .A(n9256), .ZN(n9664) );
  AOI22_X1 U10659 ( .A1(n9452), .A2(n9924), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9603), .ZN(n9453) );
  OAI21_X1 U10660 ( .B1(n9454), .B2(n9899), .A(n9453), .ZN(n9460) );
  XOR2_X1 U10661 ( .A(n9456), .B(n9455), .Z(n9458) );
  AOI21_X1 U10662 ( .B1(n9458), .B2(n9553), .A(n9457), .ZN(n9666) );
  NOR2_X1 U10663 ( .A1(n9666), .A2(n9925), .ZN(n9459) );
  AOI211_X1 U10664 ( .C1(n9664), .C2(n9919), .A(n9460), .B(n9459), .ZN(n9461)
         );
  OAI21_X1 U10665 ( .B1(n9667), .B2(n9585), .A(n9461), .ZN(P1_U3269) );
  AOI21_X1 U10666 ( .B1(n9466), .B2(n9463), .A(n9462), .ZN(n9464) );
  INV_X1 U10667 ( .A(n9464), .ZN(n9672) );
  AOI22_X1 U10668 ( .A1(n9669), .A2(n9921), .B1(n9603), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9476) );
  OAI21_X1 U10669 ( .B1(n4328), .B2(n9466), .A(n9465), .ZN(n9468) );
  AOI21_X1 U10670 ( .B1(n9468), .B2(n9553), .A(n9467), .ZN(n9671) );
  INV_X1 U10671 ( .A(n9482), .ZN(n9470) );
  INV_X1 U10672 ( .A(n9450), .ZN(n9469) );
  AOI211_X1 U10673 ( .C1(n9669), .C2(n9470), .A(n9977), .B(n9469), .ZN(n9668)
         );
  NAND2_X1 U10674 ( .A1(n9668), .A2(n9471), .ZN(n9472) );
  OAI211_X1 U10675 ( .C1(n9814), .C2(n9473), .A(n9671), .B(n9472), .ZN(n9474)
         );
  NAND2_X1 U10676 ( .A1(n9474), .A2(n9583), .ZN(n9475) );
  OAI211_X1 U10677 ( .C1(n9672), .C2(n9585), .A(n9476), .B(n9475), .ZN(
        P1_U3270) );
  XNOR2_X1 U10678 ( .A(n9478), .B(n9479), .ZN(n9677) );
  OAI21_X1 U10679 ( .B1(n9481), .B2(n9908), .A(n9480), .ZN(n9673) );
  AOI211_X1 U10680 ( .C1(n9675), .C2(n9491), .A(n9977), .B(n9482), .ZN(n9674)
         );
  NAND2_X1 U10681 ( .A1(n9674), .A2(n9819), .ZN(n9485) );
  AOI22_X1 U10682 ( .A1(n9483), .A2(n9924), .B1(n9925), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9484) );
  OAI211_X1 U10683 ( .C1(n9486), .C2(n9899), .A(n9485), .B(n9484), .ZN(n9487)
         );
  AOI21_X1 U10684 ( .B1(n9673), .B2(n9583), .A(n9487), .ZN(n9488) );
  OAI21_X1 U10685 ( .B1(n9677), .B2(n9585), .A(n9488), .ZN(P1_U3271) );
  XOR2_X1 U10686 ( .A(n9489), .B(n9496), .Z(n9682) );
  INV_X1 U10687 ( .A(n9491), .ZN(n9492) );
  AOI21_X1 U10688 ( .B1(n9678), .B2(n9490), .A(n9492), .ZN(n9679) );
  AOI22_X1 U10689 ( .A1(n9925), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9924), .B2(
        n9493), .ZN(n9494) );
  OAI21_X1 U10690 ( .B1(n9495), .B2(n9899), .A(n9494), .ZN(n9501) );
  XNOR2_X1 U10691 ( .A(n9497), .B(n9496), .ZN(n9499) );
  AOI21_X1 U10692 ( .B1(n9499), .B2(n9553), .A(n9498), .ZN(n9681) );
  NOR2_X1 U10693 ( .A1(n9681), .A2(n9925), .ZN(n9500) );
  AOI211_X1 U10694 ( .C1(n9679), .C2(n9919), .A(n9501), .B(n9500), .ZN(n9502)
         );
  OAI21_X1 U10695 ( .B1(n9585), .B2(n9682), .A(n9502), .ZN(P1_U3272) );
  NAND2_X1 U10696 ( .A1(n9504), .A2(n9503), .ZN(n9505) );
  XOR2_X1 U10697 ( .A(n9513), .B(n9505), .Z(n9507) );
  OAI21_X1 U10698 ( .B1(n9507), .B2(n9908), .A(n9506), .ZN(n9688) );
  OAI21_X1 U10699 ( .B1(n9508), .B2(n9685), .A(n9490), .ZN(n9686) );
  AOI22_X1 U10700 ( .A1(n9925), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9924), .B2(
        n9509), .ZN(n9512) );
  NAND2_X1 U10701 ( .A1(n9510), .A2(n9921), .ZN(n9511) );
  OAI211_X1 U10702 ( .C1(n9686), .C2(n9527), .A(n9512), .B(n9511), .ZN(n9517)
         );
  NOR2_X1 U10703 ( .A1(n9514), .A2(n9513), .ZN(n9684) );
  INV_X1 U10704 ( .A(n9515), .ZN(n9683) );
  NOR3_X1 U10705 ( .A1(n9684), .A2(n9683), .A3(n9585), .ZN(n9516) );
  AOI211_X1 U10706 ( .C1(n9583), .C2(n9688), .A(n9517), .B(n9516), .ZN(n9518)
         );
  INV_X1 U10707 ( .A(n9518), .ZN(P1_U3273) );
  XNOR2_X1 U10708 ( .A(n9520), .B(n9519), .ZN(n9522) );
  AOI21_X1 U10709 ( .B1(n9522), .B2(n9553), .A(n9521), .ZN(n9694) );
  XNOR2_X1 U10710 ( .A(n4365), .B(n9523), .ZN(n9695) );
  OR2_X1 U10711 ( .A1(n9695), .A2(n9585), .ZN(n9532) );
  OAI22_X1 U10712 ( .A1(n9583), .A2(n9525), .B1(n9524), .B2(n9814), .ZN(n9529)
         );
  NOR2_X1 U10713 ( .A1(n9536), .A2(n9690), .ZN(n9526) );
  OR2_X1 U10714 ( .A1(n9508), .A2(n9526), .ZN(n9691) );
  NOR2_X1 U10715 ( .A1(n9691), .A2(n9527), .ZN(n9528) );
  AOI211_X1 U10716 ( .C1(n9921), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9531)
         );
  OAI211_X1 U10717 ( .C1(n9694), .C2(n9603), .A(n9532), .B(n9531), .ZN(
        P1_U3274) );
  XNOR2_X1 U10718 ( .A(n9533), .B(n9544), .ZN(n9700) );
  NAND2_X1 U10719 ( .A1(n9559), .A2(n9697), .ZN(n9534) );
  NAND2_X1 U10720 ( .A1(n9534), .A2(n9986), .ZN(n9535) );
  NOR2_X1 U10721 ( .A1(n9536), .A2(n9535), .ZN(n9696) );
  INV_X1 U10722 ( .A(n9537), .ZN(n9538) );
  AOI22_X1 U10723 ( .A1(n9925), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9924), .B2(
        n9538), .ZN(n9539) );
  OAI21_X1 U10724 ( .B1(n9540), .B2(n9899), .A(n9539), .ZN(n9549) );
  NAND2_X1 U10725 ( .A1(n9542), .A2(n9541), .ZN(n9555) );
  NAND2_X1 U10726 ( .A1(n9555), .A2(n4419), .ZN(n9554) );
  NAND2_X1 U10727 ( .A1(n9554), .A2(n9543), .ZN(n9545) );
  XNOR2_X1 U10728 ( .A(n9545), .B(n9544), .ZN(n9547) );
  AOI21_X1 U10729 ( .B1(n9547), .B2(n9553), .A(n9546), .ZN(n9699) );
  NOR2_X1 U10730 ( .A1(n9699), .A2(n9925), .ZN(n9548) );
  AOI211_X1 U10731 ( .C1(n9696), .C2(n9819), .A(n9549), .B(n9548), .ZN(n9550)
         );
  OAI21_X1 U10732 ( .B1(n9585), .B2(n9700), .A(n9550), .ZN(P1_U3275) );
  XNOR2_X1 U10733 ( .A(n9552), .B(n9551), .ZN(n9565) );
  OAI211_X1 U10734 ( .C1(n9555), .C2(n4419), .A(n9554), .B(n9553), .ZN(n9556)
         );
  INV_X1 U10735 ( .A(n9556), .ZN(n9557) );
  AOI211_X1 U10736 ( .C1(n9895), .C2(n9565), .A(n9558), .B(n9557), .ZN(n9704)
         );
  INV_X1 U10737 ( .A(n9559), .ZN(n9560) );
  AOI21_X1 U10738 ( .B1(n9701), .B2(n9577), .A(n9560), .ZN(n9702) );
  INV_X1 U10739 ( .A(n9701), .ZN(n9564) );
  INV_X1 U10740 ( .A(n9561), .ZN(n9562) );
  AOI22_X1 U10741 ( .A1(n9925), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9924), .B2(
        n9562), .ZN(n9563) );
  OAI21_X1 U10742 ( .B1(n9564), .B2(n9899), .A(n9563), .ZN(n9568) );
  INV_X1 U10743 ( .A(n9565), .ZN(n9705) );
  NOR2_X1 U10744 ( .A1(n9705), .A2(n9566), .ZN(n9567) );
  AOI211_X1 U10745 ( .C1(n9702), .C2(n9919), .A(n9568), .B(n9567), .ZN(n9569)
         );
  OAI21_X1 U10746 ( .B1(n9704), .B2(n9603), .A(n9569), .ZN(P1_U3276) );
  XNOR2_X1 U10747 ( .A(n9570), .B(n9571), .ZN(n9710) );
  XNOR2_X1 U10748 ( .A(n9573), .B(n9572), .ZN(n9575) );
  OAI21_X1 U10749 ( .B1(n9575), .B2(n9908), .A(n9574), .ZN(n9706) );
  OR2_X1 U10750 ( .A1(n9594), .A2(n9581), .ZN(n9576) );
  AND3_X1 U10751 ( .A1(n9577), .A2(n9576), .A3(n9986), .ZN(n9707) );
  NAND2_X1 U10752 ( .A1(n9707), .A2(n9819), .ZN(n9580) );
  AOI22_X1 U10753 ( .A1(n9925), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9924), .B2(
        n9578), .ZN(n9579) );
  OAI211_X1 U10754 ( .C1(n9581), .C2(n9899), .A(n9580), .B(n9579), .ZN(n9582)
         );
  AOI21_X1 U10755 ( .B1(n9706), .B2(n9583), .A(n9582), .ZN(n9584) );
  OAI21_X1 U10756 ( .B1(n9585), .B2(n9710), .A(n9584), .ZN(P1_U3277) );
  XOR2_X1 U10757 ( .A(n9586), .B(n9587), .Z(n9711) );
  NAND2_X1 U10758 ( .A1(n9588), .A2(n9587), .ZN(n9589) );
  AOI21_X1 U10759 ( .B1(n9590), .B2(n9589), .A(n9908), .ZN(n9591) );
  AOI211_X1 U10760 ( .C1(n9895), .C2(n9711), .A(n9592), .B(n9591), .ZN(n9715)
         );
  INV_X1 U10761 ( .A(n9593), .ZN(n9595) );
  AOI21_X1 U10762 ( .B1(n9712), .B2(n9595), .A(n9594), .ZN(n9713) );
  NAND2_X1 U10763 ( .A1(n9713), .A2(n9919), .ZN(n9599) );
  INV_X1 U10764 ( .A(n9596), .ZN(n9597) );
  AOI22_X1 U10765 ( .A1(n9925), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9924), .B2(
        n9597), .ZN(n9598) );
  OAI211_X1 U10766 ( .C1(n9600), .C2(n9899), .A(n9599), .B(n9598), .ZN(n9601)
         );
  AOI21_X1 U10767 ( .B1(n9711), .B2(n9904), .A(n9601), .ZN(n9602) );
  OAI21_X1 U10768 ( .B1(n9715), .B2(n9603), .A(n9602), .ZN(P1_U3278) );
  NAND2_X1 U10769 ( .A1(n9604), .A2(n9726), .ZN(n9605) );
  NAND2_X1 U10770 ( .A1(n9605), .A2(n9612), .ZN(n9606) );
  AOI21_X1 U10771 ( .B1(n9607), .B2(n9986), .A(n9606), .ZN(n9732) );
  INV_X1 U10772 ( .A(n9609), .ZN(P1_U3554) );
  NAND2_X1 U10773 ( .A1(n9610), .A2(n9726), .ZN(n9611) );
  OAI211_X1 U10774 ( .C1(n9613), .C2(n9977), .A(n9612), .B(n9611), .ZN(n9735)
         );
  MUX2_X1 U10775 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9735), .S(n10006), .Z(
        P1_U3553) );
  INV_X1 U10776 ( .A(n9726), .ZN(n9617) );
  INV_X1 U10777 ( .A(n9614), .ZN(n9616) );
  AND2_X1 U10778 ( .A1(n9620), .A2(n4968), .ZN(n9621) );
  NAND2_X1 U10779 ( .A1(n9622), .A2(n9621), .ZN(n9623) );
  MUX2_X1 U10780 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9736), .S(n10006), .Z(
        P1_U3552) );
  INV_X1 U10781 ( .A(n9625), .ZN(n9629) );
  INV_X1 U10782 ( .A(n9626), .ZN(n9628) );
  MUX2_X1 U10783 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9737), .S(n10006), .Z(
        P1_U3551) );
  AOI22_X1 U10784 ( .A1(n9632), .A2(n9986), .B1(n9726), .B2(n9631), .ZN(n9633)
         );
  OAI211_X1 U10785 ( .C1(n9635), .C2(n9991), .A(n9634), .B(n9633), .ZN(n9738)
         );
  MUX2_X1 U10786 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9738), .S(n10006), .Z(
        P1_U3550) );
  AOI22_X1 U10787 ( .A1(n9637), .A2(n9986), .B1(n9726), .B2(n9636), .ZN(n9638)
         );
  OAI211_X1 U10788 ( .C1(n9640), .C2(n9991), .A(n9639), .B(n9638), .ZN(n9739)
         );
  MUX2_X1 U10789 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9739), .S(n10006), .Z(
        P1_U3549) );
  NAND4_X1 U10790 ( .A1(n9644), .A2(n9643), .A3(n9642), .A4(n9641), .ZN(n9645)
         );
  AOI21_X1 U10791 ( .B1(n9646), .B2(n9971), .A(n9645), .ZN(n9647) );
  INV_X1 U10792 ( .A(n9647), .ZN(n9740) );
  MUX2_X1 U10793 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9740), .S(n10006), .Z(
        P1_U3548) );
  NAND2_X1 U10794 ( .A1(n9648), .A2(n9971), .ZN(n9654) );
  NOR2_X1 U10795 ( .A1(n9650), .A2(n9649), .ZN(n9653) );
  NAND4_X1 U10796 ( .A1(n9654), .A2(n9653), .A3(n9652), .A4(n9651), .ZN(n9741)
         );
  MUX2_X1 U10797 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9741), .S(n10006), .Z(
        P1_U3547) );
  INV_X1 U10798 ( .A(n9655), .ZN(n9658) );
  NAND4_X1 U10799 ( .A1(n9659), .A2(n9658), .A3(n9657), .A4(n9656), .ZN(n9660)
         );
  AOI21_X1 U10800 ( .B1(n9661), .B2(n9971), .A(n9660), .ZN(n9662) );
  INV_X1 U10801 ( .A(n9662), .ZN(n9742) );
  MUX2_X1 U10802 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9742), .S(n10006), .Z(
        P1_U3546) );
  AOI22_X1 U10803 ( .A1(n9664), .A2(n9986), .B1(n9726), .B2(n9663), .ZN(n9665)
         );
  OAI211_X1 U10804 ( .C1(n9667), .C2(n9991), .A(n9666), .B(n9665), .ZN(n9743)
         );
  MUX2_X1 U10805 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9743), .S(n10006), .Z(
        P1_U3545) );
  AOI21_X1 U10806 ( .B1(n9726), .B2(n9669), .A(n9668), .ZN(n9670) );
  OAI211_X1 U10807 ( .C1(n9672), .C2(n9991), .A(n9671), .B(n9670), .ZN(n9744)
         );
  MUX2_X1 U10808 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9744), .S(n10006), .Z(
        P1_U3544) );
  AOI211_X1 U10809 ( .C1(n9726), .C2(n9675), .A(n9674), .B(n9673), .ZN(n9676)
         );
  OAI21_X1 U10810 ( .B1(n9991), .B2(n9677), .A(n9676), .ZN(n9745) );
  MUX2_X1 U10811 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9745), .S(n10006), .Z(
        P1_U3543) );
  AOI22_X1 U10812 ( .A1(n9679), .A2(n9986), .B1(n9726), .B2(n9678), .ZN(n9680)
         );
  OAI211_X1 U10813 ( .C1(n9682), .C2(n9991), .A(n9681), .B(n9680), .ZN(n9746)
         );
  MUX2_X1 U10814 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9746), .S(n10006), .Z(
        P1_U3542) );
  NOR3_X1 U10815 ( .A1(n9684), .A2(n9683), .A3(n9991), .ZN(n9689) );
  OAI22_X1 U10816 ( .A1(n9686), .A2(n9977), .B1(n9685), .B2(n9617), .ZN(n9687)
         );
  MUX2_X1 U10817 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9747), .S(n10006), .Z(
        P1_U3541) );
  OAI22_X1 U10818 ( .A1(n9691), .A2(n9977), .B1(n9690), .B2(n9617), .ZN(n9692)
         );
  INV_X1 U10819 ( .A(n9692), .ZN(n9693) );
  OAI211_X1 U10820 ( .C1(n9695), .C2(n9991), .A(n9694), .B(n9693), .ZN(n9748)
         );
  MUX2_X1 U10821 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9748), .S(n10006), .Z(
        P1_U3540) );
  AOI21_X1 U10822 ( .B1(n9726), .B2(n9697), .A(n9696), .ZN(n9698) );
  OAI211_X1 U10823 ( .C1(n9991), .C2(n9700), .A(n9699), .B(n9698), .ZN(n9749)
         );
  MUX2_X1 U10824 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9749), .S(n10006), .Z(
        P1_U3539) );
  AOI22_X1 U10825 ( .A1(n9702), .A2(n9986), .B1(n9726), .B2(n9701), .ZN(n9703)
         );
  OAI211_X1 U10826 ( .C1(n9705), .C2(n9936), .A(n9704), .B(n9703), .ZN(n9750)
         );
  MUX2_X1 U10827 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9750), .S(n10006), .Z(
        P1_U3538) );
  AOI211_X1 U10828 ( .C1(n9726), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9709)
         );
  OAI21_X1 U10829 ( .B1(n9991), .B2(n9710), .A(n9709), .ZN(n9751) );
  MUX2_X1 U10830 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9751), .S(n10006), .Z(
        P1_U3537) );
  INV_X1 U10831 ( .A(n9711), .ZN(n9716) );
  AOI22_X1 U10832 ( .A1(n9713), .A2(n9986), .B1(n9726), .B2(n9712), .ZN(n9714)
         );
  OAI211_X1 U10833 ( .C1(n9936), .C2(n9716), .A(n9715), .B(n9714), .ZN(n9752)
         );
  MUX2_X1 U10834 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9752), .S(n10006), .Z(
        P1_U3536) );
  NAND2_X1 U10835 ( .A1(n9717), .A2(n9726), .ZN(n9719) );
  OAI211_X1 U10836 ( .C1(n9720), .C2(n9936), .A(n9719), .B(n9718), .ZN(n9721)
         );
  NOR2_X1 U10837 ( .A1(n9722), .A2(n9721), .ZN(n9753) );
  MUX2_X1 U10838 ( .A(n9723), .B(n9753), .S(n10006), .Z(n9724) );
  INV_X1 U10839 ( .A(n9724), .ZN(P1_U3535) );
  AOI22_X1 U10840 ( .A1(n9727), .A2(n9986), .B1(n9726), .B2(n9725), .ZN(n9728)
         );
  OAI211_X1 U10841 ( .C1(n9936), .C2(n9730), .A(n9729), .B(n9728), .ZN(n9756)
         );
  MUX2_X1 U10842 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9756), .S(n10006), .Z(
        P1_U3534) );
  MUX2_X1 U10843 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9731), .S(n10006), .Z(
        P1_U3523) );
  INV_X1 U10844 ( .A(n9734), .ZN(P1_U3522) );
  MUX2_X1 U10845 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9735), .S(n9995), .Z(
        P1_U3521) );
  MUX2_X1 U10846 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9736), .S(n9995), .Z(
        P1_U3520) );
  MUX2_X1 U10847 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9737), .S(n9995), .Z(
        P1_U3519) );
  MUX2_X1 U10848 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9738), .S(n9995), .Z(
        P1_U3518) );
  MUX2_X1 U10849 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9739), .S(n9995), .Z(
        P1_U3517) );
  MUX2_X1 U10850 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9740), .S(n9995), .Z(
        P1_U3516) );
  MUX2_X1 U10851 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9741), .S(n9995), .Z(
        P1_U3515) );
  MUX2_X1 U10852 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9742), .S(n9995), .Z(
        P1_U3514) );
  MUX2_X1 U10853 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9743), .S(n9995), .Z(
        P1_U3513) );
  MUX2_X1 U10854 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9744), .S(n9995), .Z(
        P1_U3512) );
  MUX2_X1 U10855 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9745), .S(n9995), .Z(
        P1_U3511) );
  MUX2_X1 U10856 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9746), .S(n9995), .Z(
        P1_U3510) );
  MUX2_X1 U10857 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9747), .S(n9995), .Z(
        P1_U3508) );
  MUX2_X1 U10858 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9748), .S(n9995), .Z(
        P1_U3505) );
  MUX2_X1 U10859 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9749), .S(n9995), .Z(
        P1_U3502) );
  MUX2_X1 U10860 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9750), .S(n9995), .Z(
        P1_U3499) );
  MUX2_X1 U10861 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9751), .S(n9995), .Z(
        P1_U3496) );
  MUX2_X1 U10862 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9752), .S(n9995), .Z(
        P1_U3493) );
  MUX2_X1 U10863 ( .A(n9754), .B(n9753), .S(n9995), .Z(n9755) );
  INV_X1 U10864 ( .A(n9755), .ZN(P1_U3490) );
  INV_X1 U10865 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U10866 ( .A1(n9756), .A2(n9995), .ZN(n9757) );
  OAI21_X1 U10867 ( .B1(n9995), .B2(n9758), .A(n9757), .ZN(P1_U3487) );
  MUX2_X1 U10868 ( .A(P1_D_REG_0__SCAN_IN), .B(n9759), .S(n9935), .Z(P1_U3440)
         );
  INV_X1 U10869 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9760) );
  OAI222_X1 U10870 ( .A1(P1_U3084), .A2(n9762), .B1(n9774), .B2(n9761), .C1(
        n9760), .C2(n7832), .ZN(P1_U3324) );
  AOI21_X1 U10871 ( .B1(n9771), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9763), .ZN(
        n9764) );
  OAI21_X1 U10872 ( .B1(n9765), .B2(n9774), .A(n9764), .ZN(P1_U3325) );
  NAND2_X1 U10873 ( .A1(n9771), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9767) );
  OAI211_X1 U10874 ( .C1(n9768), .C2(n9774), .A(n9767), .B(n9766), .ZN(
        P1_U3326) );
  AOI22_X1 U10875 ( .A1(n6458), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9771), .ZN(n9769) );
  OAI21_X1 U10876 ( .B1(n9770), .B2(n9774), .A(n9769), .ZN(P1_U3327) );
  AOI22_X1 U10877 ( .A1(n9772), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n9771), .ZN(n9773) );
  OAI21_X1 U10878 ( .B1(n9775), .B2(n9774), .A(n9773), .ZN(P1_U3328) );
  INV_X1 U10879 ( .A(n9776), .ZN(n9777) );
  MUX2_X1 U10880 ( .A(n9777), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NOR2_X1 U10881 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9778) );
  AOI21_X1 U10882 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9778), .ZN(n10089) );
  NOR2_X1 U10883 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9779) );
  AOI21_X1 U10884 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9779), .ZN(n10092) );
  NOR2_X1 U10885 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9780) );
  AOI21_X1 U10886 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9780), .ZN(n10095) );
  NOR2_X1 U10887 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9781) );
  AOI21_X1 U10888 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9781), .ZN(n10098) );
  NOR2_X1 U10889 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9782) );
  AOI21_X1 U10890 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9782), .ZN(n10101) );
  NOR2_X1 U10891 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n9783) );
  AOI21_X1 U10892 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n9783), .ZN(n10134) );
  NAND2_X1 U10893 ( .A1(n10185), .A2(n10085), .ZN(n9784) );
  NOR2_X1 U10894 ( .A1(n10185), .A2(n10085), .ZN(n10083) );
  AOI21_X1 U10895 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(n9784), .A(n10083), .ZN(
        n10128) );
  NAND2_X1 U10896 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9785) );
  OAI21_X1 U10897 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n9785), .ZN(n10127) );
  NOR2_X1 U10898 ( .A1(n10128), .A2(n10127), .ZN(n10126) );
  NAND2_X1 U10899 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9786) );
  OAI21_X1 U10900 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n9786), .ZN(n10130) );
  NOR2_X1 U10901 ( .A1(n10131), .A2(n10130), .ZN(n10129) );
  NAND2_X1 U10902 ( .A1(n10134), .A2(n10133), .ZN(n10132) );
  OAI21_X1 U10903 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10132), .ZN(n9787) );
  INV_X1 U10904 ( .A(n9787), .ZN(n9788) );
  NAND2_X1 U10905 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9788), .ZN(n10117) );
  NAND2_X1 U10906 ( .A1(n6936), .A2(n10117), .ZN(n10114) );
  NOR2_X1 U10907 ( .A1(n9789), .A2(n6913), .ZN(n9790) );
  XNOR2_X1 U10908 ( .A(n9789), .B(n6913), .ZN(n10113) );
  INV_X1 U10909 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10112) );
  NOR2_X1 U10910 ( .A1(n9791), .A2(n10184), .ZN(n9792) );
  INV_X1 U10911 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10241) );
  XNOR2_X1 U10912 ( .A(n10184), .B(n9791), .ZN(n10125) );
  INV_X1 U10913 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9793) );
  NAND2_X1 U10914 ( .A1(n9794), .A2(n9793), .ZN(n10275) );
  INV_X1 U10915 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9796) );
  NOR2_X1 U10916 ( .A1(n9795), .A2(n9796), .ZN(n9797) );
  INV_X1 U10917 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10201) );
  XNOR2_X1 U10918 ( .A(n9796), .B(n9795), .ZN(n10123) );
  NAND2_X1 U10919 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9798) );
  OAI21_X1 U10920 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9798), .ZN(n10109) );
  NAND2_X1 U10921 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9799) );
  OAI21_X1 U10922 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9799), .ZN(n10106) );
  NOR2_X1 U10923 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9800) );
  AOI21_X1 U10924 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9800), .ZN(n10103) );
  NAND2_X1 U10925 ( .A1(n10098), .A2(n10097), .ZN(n10096) );
  NAND2_X1 U10926 ( .A1(n10095), .A2(n10094), .ZN(n10093) );
  NAND2_X1 U10927 ( .A1(n10089), .A2(n10088), .ZN(n10087) );
  NOR2_X1 U10928 ( .A1(n10120), .A2(n10119), .ZN(n9801) );
  NAND2_X1 U10929 ( .A1(n10120), .A2(n10119), .ZN(n10118) );
  XNOR2_X1 U10930 ( .A(n4774), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n9802) );
  XNOR2_X1 U10931 ( .A(n9803), .B(n9802), .ZN(ADD_1071_U4) );
  OAI21_X1 U10932 ( .B1(n4385), .B2(n7751), .A(n9804), .ZN(n9828) );
  INV_X1 U10933 ( .A(n9805), .ZN(n9807) );
  OAI21_X1 U10934 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(n9809) );
  XOR2_X1 U10935 ( .A(n9810), .B(n9809), .Z(n9811) );
  NOR2_X1 U10936 ( .A1(n9811), .A2(n9908), .ZN(n9826) );
  AOI211_X1 U10937 ( .C1(n9895), .C2(n9828), .A(n9823), .B(n9826), .ZN(n9822)
         );
  NAND2_X1 U10938 ( .A1(n9925), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9812) );
  OAI21_X1 U10939 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n9815) );
  AOI21_X1 U10940 ( .B1(n9921), .B2(n9818), .A(n9815), .ZN(n9821) );
  INV_X1 U10941 ( .A(n9816), .ZN(n9817) );
  AOI211_X1 U10942 ( .C1(n9818), .C2(n9817), .A(n9977), .B(n7757), .ZN(n9825)
         );
  AOI22_X1 U10943 ( .A1(n9904), .A2(n9828), .B1(n9825), .B2(n9819), .ZN(n9820)
         );
  OAI211_X1 U10944 ( .C1(n9925), .C2(n9822), .A(n9821), .B(n9820), .ZN(
        P1_U3281) );
  OR3_X1 U10945 ( .A1(n9825), .A2(n9824), .A3(n9823), .ZN(n9827) );
  AOI211_X1 U10946 ( .C1(n9971), .C2(n9828), .A(n9827), .B(n9826), .ZN(n9830)
         );
  INV_X1 U10947 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9829) );
  AOI22_X1 U10948 ( .A1(n9995), .A2(n9830), .B1(n9829), .B2(n9993), .ZN(
        P1_U3484) );
  AOI22_X1 U10949 ( .A1(n10006), .A2(n9830), .B1(n6180), .B2(n10004), .ZN(
        P1_U3533) );
  XNOR2_X1 U10950 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10951 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10952 ( .A(n9831), .ZN(n9833) );
  AOI22_X1 U10953 ( .A1(n9833), .A2(n9832), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3084), .ZN(n9841) );
  XNOR2_X1 U10954 ( .A(n9835), .B(n9834), .ZN(n9839) );
  NOR2_X1 U10955 ( .A1(n9617), .A2(n9836), .ZN(n9942) );
  AOI22_X1 U10956 ( .A1(n9839), .A2(n9838), .B1(n9837), .B2(n9942), .ZN(n9840)
         );
  OAI211_X1 U10957 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9842), .A(n9841), .B(
        n9840), .ZN(P1_U3216) );
  INV_X1 U10958 ( .A(n9843), .ZN(n9844) );
  OAI21_X1 U10959 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(n9849) );
  NAND2_X1 U10960 ( .A1(n9861), .A2(n9847), .ZN(n9848) );
  OAI21_X1 U10961 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9852) );
  AOI211_X1 U10962 ( .C1(n9874), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n9852), .B(
        n9851), .ZN(n9857) );
  OAI211_X1 U10963 ( .C1(n9855), .C2(n9854), .A(n9878), .B(n9853), .ZN(n9856)
         );
  OAI211_X1 U10964 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n7022), .A(n9857), .B(
        n9856), .ZN(P1_U3243) );
  INV_X1 U10965 ( .A(n9858), .ZN(n9859) );
  AOI21_X1 U10966 ( .B1(n9861), .B2(n9860), .A(n9859), .ZN(n9869) );
  NAND2_X1 U10967 ( .A1(n9874), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n9868) );
  XNOR2_X1 U10968 ( .A(n9862), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n9863) );
  NAND2_X1 U10969 ( .A1(n9863), .A2(n9878), .ZN(n9867) );
  XOR2_X1 U10970 ( .A(P1_REG2_REG_15__SCAN_IN), .B(n9864), .Z(n9865) );
  NAND2_X1 U10971 ( .A1(n9865), .A2(n9879), .ZN(n9866) );
  NAND4_X1 U10972 ( .A1(n9869), .A2(n9868), .A3(n9867), .A4(n9866), .ZN(
        P1_U3256) );
  NOR2_X1 U10973 ( .A1(n9871), .A2(n9870), .ZN(n9872) );
  AOI211_X1 U10974 ( .C1(n9874), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9873), .B(
        n9872), .ZN(n9885) );
  XOR2_X1 U10975 ( .A(n9876), .B(n9875), .Z(n9877) );
  NAND2_X1 U10976 ( .A1(n9878), .A2(n9877), .ZN(n9884) );
  OAI211_X1 U10977 ( .C1(n9882), .C2(n9881), .A(n9880), .B(n9879), .ZN(n9883)
         );
  NAND3_X1 U10978 ( .A1(n9885), .A2(n9884), .A3(n9883), .ZN(P1_U3258) );
  XNOR2_X1 U10979 ( .A(n9886), .B(n9891), .ZN(n9982) );
  INV_X1 U10980 ( .A(n9887), .ZN(n9892) );
  AND2_X1 U10981 ( .A1(n9889), .A2(n9888), .ZN(n9890) );
  AOI211_X1 U10982 ( .C1(n9892), .C2(n9891), .A(n9908), .B(n9890), .ZN(n9893)
         );
  AOI211_X1 U10983 ( .C1(n9895), .C2(n9982), .A(n9894), .B(n9893), .ZN(n9979)
         );
  INV_X1 U10984 ( .A(n9896), .ZN(n9897) );
  AOI22_X1 U10985 ( .A1(n9925), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9924), .B2(
        n9897), .ZN(n9898) );
  OAI21_X1 U10986 ( .B1(n9899), .B2(n9902), .A(n9898), .ZN(n9900) );
  INV_X1 U10987 ( .A(n9900), .ZN(n9906) );
  OAI21_X1 U10988 ( .B1(n4390), .B2(n9902), .A(n9901), .ZN(n9978) );
  INV_X1 U10989 ( .A(n9978), .ZN(n9903) );
  AOI22_X1 U10990 ( .A1(n9982), .A2(n9904), .B1(n9919), .B2(n9903), .ZN(n9905)
         );
  OAI211_X1 U10991 ( .C1(n9925), .C2(n9979), .A(n9906), .B(n9905), .ZN(
        P1_U3283) );
  INV_X1 U10992 ( .A(n9907), .ZN(n9909) );
  AOI21_X1 U10993 ( .B1(n9909), .B2(n9913), .A(n9908), .ZN(n9911) );
  AOI21_X1 U10994 ( .B1(n9911), .B2(n7528), .A(n9910), .ZN(n9950) );
  XNOR2_X1 U10995 ( .A(n9913), .B(n9912), .ZN(n9953) );
  NAND2_X1 U10996 ( .A1(n9914), .A2(n9953), .ZN(n9929) );
  AND2_X1 U10997 ( .A1(n9915), .A2(n9920), .ZN(n9917) );
  OR2_X1 U10998 ( .A1(n9917), .A2(n9916), .ZN(n9951) );
  INV_X1 U10999 ( .A(n9951), .ZN(n9918) );
  NAND2_X1 U11000 ( .A1(n9919), .A2(n9918), .ZN(n9928) );
  NAND2_X1 U11001 ( .A1(n9921), .A2(n9920), .ZN(n9927) );
  INV_X1 U11002 ( .A(n9922), .ZN(n9923) );
  AOI22_X1 U11003 ( .A1(n9925), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9924), .B2(
        n9923), .ZN(n9926) );
  AND4_X1 U11004 ( .A1(n9929), .A2(n9928), .A3(n9927), .A4(n9926), .ZN(n9930)
         );
  OAI21_X1 U11005 ( .B1(n9925), .B2(n9950), .A(n9930), .ZN(P1_U3287) );
  AND2_X1 U11006 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9933), .ZN(P1_U3292) );
  AND2_X1 U11007 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9933), .ZN(P1_U3293) );
  AND2_X1 U11008 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9933), .ZN(P1_U3294) );
  AND2_X1 U11009 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9933), .ZN(P1_U3295) );
  AND2_X1 U11010 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9933), .ZN(P1_U3296) );
  AND2_X1 U11011 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9933), .ZN(P1_U3297) );
  AND2_X1 U11012 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9933), .ZN(P1_U3298) );
  AND2_X1 U11013 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9933), .ZN(P1_U3299) );
  AND2_X1 U11014 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9933), .ZN(P1_U3300) );
  AND2_X1 U11015 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9933), .ZN(P1_U3301) );
  AND2_X1 U11016 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9933), .ZN(P1_U3302) );
  AND2_X1 U11017 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9933), .ZN(P1_U3303) );
  AND2_X1 U11018 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9933), .ZN(P1_U3304) );
  AND2_X1 U11019 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9933), .ZN(P1_U3305) );
  AND2_X1 U11020 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9933), .ZN(P1_U3306) );
  AND2_X1 U11021 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9933), .ZN(P1_U3307) );
  AND2_X1 U11022 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9933), .ZN(P1_U3308) );
  AND2_X1 U11023 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9933), .ZN(P1_U3309) );
  AND2_X1 U11024 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9933), .ZN(P1_U3310) );
  AND2_X1 U11025 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9933), .ZN(P1_U3311) );
  INV_X1 U11026 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U11027 ( .A1(n9932), .A2(n10221), .ZN(P1_U3312) );
  INV_X1 U11028 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U11029 ( .A1(n9932), .A2(n10215), .ZN(P1_U3313) );
  AND2_X1 U11030 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9933), .ZN(P1_U3314) );
  AND2_X1 U11031 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9933), .ZN(P1_U3315) );
  INV_X1 U11032 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10229) );
  NOR2_X1 U11033 ( .A1(n9932), .A2(n10229), .ZN(P1_U3316) );
  AND2_X1 U11034 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9933), .ZN(P1_U3317) );
  AND2_X1 U11035 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9933), .ZN(P1_U3318) );
  INV_X1 U11036 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10175) );
  NOR2_X1 U11037 ( .A1(n9932), .A2(n10175), .ZN(P1_U3319) );
  AND2_X1 U11038 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9933), .ZN(P1_U3320) );
  AND2_X1 U11039 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9933), .ZN(P1_U3321) );
  INV_X1 U11040 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10173) );
  OAI21_X1 U11041 ( .B1(n9935), .B2(n10173), .A(n9934), .ZN(P1_U3441) );
  INV_X1 U11042 ( .A(n9936), .ZN(n9983) );
  OAI22_X1 U11043 ( .A1(n9617), .A2(n4433), .B1(n9977), .B2(n9937), .ZN(n9940)
         );
  AOI211_X1 U11044 ( .C1(n9983), .C2(n9941), .A(n9940), .B(n9939), .ZN(n9996)
         );
  AOI22_X1 U11045 ( .A1(n9995), .A2(n9996), .B1(n6015), .B2(n9993), .ZN(
        P1_U3460) );
  INV_X1 U11046 ( .A(n9942), .ZN(n9943) );
  OAI21_X1 U11047 ( .B1(n9977), .B2(n9944), .A(n9943), .ZN(n9946) );
  AOI211_X1 U11048 ( .C1(n9983), .C2(n9947), .A(n9946), .B(n9945), .ZN(n9997)
         );
  AOI22_X1 U11049 ( .A1(n9995), .A2(n9997), .B1(n4558), .B2(n9993), .ZN(
        P1_U3463) );
  INV_X1 U11050 ( .A(n9948), .ZN(n9949) );
  OAI211_X1 U11051 ( .C1(n9977), .C2(n9951), .A(n9950), .B(n9949), .ZN(n9952)
         );
  AOI21_X1 U11052 ( .B1(n9971), .B2(n9953), .A(n9952), .ZN(n9998) );
  AOI22_X1 U11053 ( .A1(n9995), .A2(n9998), .B1(n6056), .B2(n9993), .ZN(
        P1_U3466) );
  NAND3_X1 U11054 ( .A1(n9955), .A2(n9954), .A3(n9971), .ZN(n9956) );
  AND4_X1 U11055 ( .A1(n9959), .A2(n9958), .A3(n9957), .A4(n9956), .ZN(n9999)
         );
  INV_X1 U11056 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U11057 ( .A1(n9995), .A2(n9999), .B1(n9960), .B2(n9993), .ZN(
        P1_U3469) );
  INV_X1 U11058 ( .A(n9961), .ZN(n9967) );
  INV_X1 U11059 ( .A(n9962), .ZN(n9965) );
  OAI211_X1 U11060 ( .C1(n9977), .C2(n9965), .A(n9964), .B(n9963), .ZN(n9966)
         );
  AOI21_X1 U11061 ( .B1(n9967), .B2(n9971), .A(n9966), .ZN(n10000) );
  AOI22_X1 U11062 ( .A1(n9995), .A2(n10000), .B1(n4559), .B2(n9993), .ZN(
        P1_U3472) );
  AOI211_X1 U11063 ( .C1(n9971), .C2(n9970), .A(n9969), .B(n9968), .ZN(n9973)
         );
  AND2_X1 U11064 ( .A1(n9973), .A2(n9972), .ZN(n10001) );
  INV_X1 U11065 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11066 ( .A1(n9995), .A2(n10001), .B1(n9974), .B2(n9993), .ZN(
        P1_U3475) );
  INV_X1 U11067 ( .A(n9975), .ZN(n9976) );
  OAI21_X1 U11068 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(n9981) );
  INV_X1 U11069 ( .A(n9979), .ZN(n9980) );
  AOI211_X1 U11070 ( .C1(n9983), .C2(n9982), .A(n9981), .B(n9980), .ZN(n10003)
         );
  INV_X1 U11071 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U11072 ( .A1(n9995), .A2(n10003), .B1(n9984), .B2(n9993), .ZN(
        P1_U3478) );
  AOI21_X1 U11073 ( .B1(n9987), .B2(n9986), .A(n9985), .ZN(n9988) );
  OAI211_X1 U11074 ( .C1(n9991), .C2(n9990), .A(n9989), .B(n9988), .ZN(n9992)
         );
  INV_X1 U11075 ( .A(n9992), .ZN(n10005) );
  INV_X1 U11076 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U11077 ( .A1(n9995), .A2(n10005), .B1(n9994), .B2(n9993), .ZN(
        P1_U3481) );
  AOI22_X1 U11078 ( .A1(n10006), .A2(n9996), .B1(n6884), .B2(n10004), .ZN(
        P1_U3525) );
  AOI22_X1 U11079 ( .A1(n10006), .A2(n9997), .B1(n6885), .B2(n10004), .ZN(
        P1_U3526) );
  AOI22_X1 U11080 ( .A1(n10006), .A2(n9998), .B1(n6890), .B2(n10004), .ZN(
        P1_U3527) );
  AOI22_X1 U11081 ( .A1(n10006), .A2(n9999), .B1(n6090), .B2(n10004), .ZN(
        P1_U3528) );
  AOI22_X1 U11082 ( .A1(n10006), .A2(n10000), .B1(n6074), .B2(n10004), .ZN(
        P1_U3529) );
  AOI22_X1 U11083 ( .A1(n10006), .A2(n10001), .B1(n7037), .B2(n10004), .ZN(
        P1_U3530) );
  AOI22_X1 U11084 ( .A1(n10006), .A2(n10003), .B1(n10002), .B2(n10004), .ZN(
        P1_U3531) );
  AOI22_X1 U11085 ( .A1(n10006), .A2(n10005), .B1(n7041), .B2(n10004), .ZN(
        P1_U3532) );
  AOI22_X1 U11086 ( .A1(n10008), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10007), .ZN(n10017) );
  AOI22_X1 U11087 ( .A1(n10009), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10016) );
  OAI21_X1 U11088 ( .B1(n10011), .B2(P2_REG1_REG_0__SCAN_IN), .A(n10010), .ZN(
        n10014) );
  NOR2_X1 U11089 ( .A1(n10012), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10013) );
  OAI21_X1 U11090 ( .B1(n10014), .B2(n10013), .A(n4407), .ZN(n10015) );
  OAI211_X1 U11091 ( .C1(n4407), .C2(n10017), .A(n10016), .B(n10015), .ZN(
        P2_U3245) );
  OAI21_X1 U11092 ( .B1(n10019), .B2(n10018), .A(n7233), .ZN(n10022) );
  AOI21_X1 U11093 ( .B1(n10022), .B2(n10021), .A(n10020), .ZN(n10059) );
  OR2_X1 U11094 ( .A1(n10024), .A2(n10023), .ZN(n10025) );
  NAND2_X1 U11095 ( .A1(n10026), .A2(n10025), .ZN(n10056) );
  NAND2_X1 U11096 ( .A1(n10056), .A2(n10027), .ZN(n10028) );
  NAND2_X1 U11097 ( .A1(n10059), .A2(n10028), .ZN(n10030) );
  AOI22_X1 U11098 ( .A1(n10031), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n10030), 
        .B2(n10029), .ZN(n10040) );
  AOI21_X1 U11099 ( .B1(n10034), .B2(n10033), .A(n10032), .ZN(n10037) );
  MUX2_X1 U11100 ( .A(n10037), .B(n10036), .S(n10035), .Z(n10058) );
  OR2_X1 U11101 ( .A1(n10038), .A2(n10058), .ZN(n10039) );
  OAI211_X1 U11102 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n10041), .A(n10040), .B(
        n10039), .ZN(P2_U3293) );
  INV_X1 U11103 ( .A(n10042), .ZN(n10043) );
  AND2_X1 U11104 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10047), .ZN(P2_U3297) );
  AND2_X1 U11105 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10047), .ZN(P2_U3298) );
  INV_X1 U11106 ( .A(n10047), .ZN(n10045) );
  INV_X1 U11107 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10240) );
  NOR2_X1 U11108 ( .A1(n10045), .A2(n10240), .ZN(P2_U3299) );
  AND2_X1 U11109 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10047), .ZN(P2_U3300) );
  AND2_X1 U11110 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10047), .ZN(P2_U3301) );
  AND2_X1 U11111 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10047), .ZN(P2_U3302) );
  AND2_X1 U11112 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10047), .ZN(P2_U3303) );
  AND2_X1 U11113 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10047), .ZN(P2_U3304) );
  INV_X1 U11114 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10227) );
  NOR2_X1 U11115 ( .A1(n10045), .A2(n10227), .ZN(P2_U3305) );
  AND2_X1 U11116 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10047), .ZN(P2_U3306) );
  AND2_X1 U11117 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10047), .ZN(P2_U3307) );
  AND2_X1 U11118 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10047), .ZN(P2_U3308) );
  AND2_X1 U11119 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10047), .ZN(P2_U3309) );
  AND2_X1 U11120 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10047), .ZN(P2_U3310) );
  AND2_X1 U11121 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10047), .ZN(P2_U3311) );
  AND2_X1 U11122 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10047), .ZN(P2_U3312) );
  AND2_X1 U11123 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10047), .ZN(P2_U3313) );
  INV_X1 U11124 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10200) );
  NOR2_X1 U11125 ( .A1(n10045), .A2(n10200), .ZN(P2_U3314) );
  AND2_X1 U11126 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10047), .ZN(P2_U3315) );
  AND2_X1 U11127 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10047), .ZN(P2_U3316) );
  AND2_X1 U11128 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10047), .ZN(P2_U3317) );
  INV_X1 U11129 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10195) );
  NOR2_X1 U11130 ( .A1(n10045), .A2(n10195), .ZN(P2_U3318) );
  AND2_X1 U11131 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10047), .ZN(P2_U3319) );
  AND2_X1 U11132 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10047), .ZN(P2_U3320) );
  AND2_X1 U11133 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10047), .ZN(P2_U3321) );
  AND2_X1 U11134 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10047), .ZN(P2_U3322) );
  AND2_X1 U11135 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10047), .ZN(P2_U3323) );
  AND2_X1 U11136 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10047), .ZN(P2_U3324) );
  AND2_X1 U11137 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10047), .ZN(P2_U3325) );
  AND2_X1 U11138 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10047), .ZN(P2_U3326) );
  AOI22_X1 U11139 ( .A1(n10050), .A2(n10046), .B1(n10140), .B2(n10047), .ZN(
        P2_U3437) );
  AOI22_X1 U11140 ( .A1(n10050), .A2(n10049), .B1(n10048), .B2(n10047), .ZN(
        P2_U3438) );
  OAI21_X1 U11141 ( .B1(n10052), .B2(n6756), .A(n10051), .ZN(n10053) );
  AOI21_X1 U11142 ( .B1(n10074), .B2(n10054), .A(n10053), .ZN(n10077) );
  INV_X1 U11143 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U11144 ( .A1(n10076), .A2(n10077), .B1(n10055), .B2(n10075), .ZN(
        P2_U3451) );
  NAND2_X1 U11145 ( .A1(n10056), .A2(n10074), .ZN(n10057) );
  AND3_X1 U11146 ( .A1(n10059), .A2(n10058), .A3(n10057), .ZN(n10078) );
  INV_X1 U11147 ( .A(n10078), .ZN(n10060) );
  OAI22_X1 U11148 ( .A1(n10075), .A2(n10060), .B1(P2_REG0_REG_3__SCAN_IN), 
        .B2(n10076), .ZN(n10061) );
  INV_X1 U11149 ( .A(n10061), .ZN(P2_U3460) );
  OAI21_X1 U11150 ( .B1(n10063), .B2(n10070), .A(n10062), .ZN(n10065) );
  AOI211_X1 U11151 ( .C1(n10074), .C2(n10066), .A(n10065), .B(n10064), .ZN(
        n10079) );
  INV_X1 U11152 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U11153 ( .A1(n10076), .A2(n10079), .B1(n10067), .B2(n10075), .ZN(
        P2_U3463) );
  OAI211_X1 U11154 ( .C1(n10071), .C2(n10070), .A(n10069), .B(n10068), .ZN(
        n10072) );
  AOI21_X1 U11155 ( .B1(n10074), .B2(n10073), .A(n10072), .ZN(n10081) );
  INV_X1 U11156 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U11157 ( .A1(n10076), .A2(n10081), .B1(n10163), .B2(n10075), .ZN(
        P2_U3469) );
  AOI22_X1 U11158 ( .A1(n10082), .A2(n10077), .B1(n5005), .B2(n10080), .ZN(
        P2_U3520) );
  AOI22_X1 U11159 ( .A1(n10082), .A2(n10078), .B1(n5864), .B2(n10080), .ZN(
        P2_U3523) );
  AOI22_X1 U11160 ( .A1(n10082), .A2(n10079), .B1(n5865), .B2(n10080), .ZN(
        P2_U3524) );
  AOI22_X1 U11161 ( .A1(n10082), .A2(n10081), .B1(n5127), .B2(n10080), .ZN(
        P2_U3526) );
  AOI21_X1 U11162 ( .B1(n10085), .B2(n10185), .A(n10083), .ZN(n10084) );
  XNOR2_X1 U11163 ( .A(n10084), .B(n7264), .ZN(ADD_1071_U5) );
  OAI21_X1 U11164 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(n10085), .ZN(n10086) );
  INV_X1 U11165 ( .A(n10086), .ZN(ADD_1071_U46) );
  OAI21_X1 U11166 ( .B1(n10089), .B2(n10088), .A(n10087), .ZN(ADD_1071_U56) );
  OAI21_X1 U11167 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(ADD_1071_U57) );
  OAI21_X1 U11168 ( .B1(n10095), .B2(n10094), .A(n10093), .ZN(ADD_1071_U58) );
  OAI21_X1 U11169 ( .B1(n10098), .B2(n10097), .A(n10096), .ZN(ADD_1071_U59) );
  OAI21_X1 U11170 ( .B1(n10101), .B2(n10100), .A(n10099), .ZN(ADD_1071_U60) );
  OAI21_X1 U11171 ( .B1(n10104), .B2(n10103), .A(n10102), .ZN(ADD_1071_U61) );
  AOI21_X1 U11172 ( .B1(n10107), .B2(n10106), .A(n10105), .ZN(ADD_1071_U62) );
  AOI21_X1 U11173 ( .B1(n10110), .B2(n10109), .A(n10108), .ZN(ADD_1071_U63) );
  AOI21_X1 U11174 ( .B1(n10113), .B2(n10112), .A(n10111), .ZN(ADD_1071_U50) );
  OAI222_X1 U11175 ( .A1(n6936), .A2(n10117), .B1(n6936), .B2(n10116), .C1(
        n10115), .C2(n10114), .ZN(ADD_1071_U51) );
  OAI21_X1 U11176 ( .B1(n10120), .B2(n10119), .A(n10118), .ZN(n10121) );
  XNOR2_X1 U11177 ( .A(n10121), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11178 ( .B1(n10201), .B2(n10123), .A(n10122), .ZN(ADD_1071_U47) );
  AOI21_X1 U11179 ( .B1(n10241), .B2(n10125), .A(n10124), .ZN(ADD_1071_U49) );
  AOI21_X1 U11180 ( .B1(n10128), .B2(n10127), .A(n10126), .ZN(ADD_1071_U54) );
  AOI21_X1 U11181 ( .B1(n10131), .B2(n10130), .A(n10129), .ZN(ADD_1071_U53) );
  OAI21_X1 U11182 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(ADD_1071_U52) );
  NAND4_X1 U11183 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_DATAO_REG_11__SCAN_IN), 
        .A3(P2_D_REG_14__SCAN_IN), .A4(P1_ADDR_REG_9__SCAN_IN), .ZN(n10146) );
  NOR4_X1 U11184 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(n10232), .A3(n10135), 
        .A4(n10231), .ZN(n10138) );
  NOR4_X1 U11185 ( .A1(SI_13_), .A2(P1_IR_REG_28__SCAN_IN), .A3(
        P1_REG2_REG_5__SCAN_IN), .A4(n10215), .ZN(n10137) );
  NOR4_X1 U11186 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(n10218), .A3(n10220), 
        .A4(n10213), .ZN(n10136) );
  NAND3_X1 U11187 ( .A1(n10138), .A2(n10137), .A3(n10136), .ZN(n10145) );
  INV_X1 U11188 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10246) );
  NAND4_X1 U11189 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(SI_30_), .A3(n10248), 
        .A4(n10246), .ZN(n10144) );
  NOR3_X1 U11190 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_REG2_REG_20__SCAN_IN), .ZN(n10142) );
  NOR4_X1 U11191 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_REG2_REG_18__SCAN_IN), 
        .A3(P2_IR_REG_15__SCAN_IN), .A4(P2_REG2_REG_4__SCAN_IN), .ZN(n10139)
         );
  AND4_X1 U11192 ( .A1(P1_REG1_REG_30__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), 
        .A3(n10139), .A4(P1_REG2_REG_3__SCAN_IN), .ZN(n10141) );
  NAND4_X1 U11193 ( .A1(n10142), .A2(P1_REG2_REG_27__SCAN_IN), .A3(n10141), 
        .A4(n10140), .ZN(n10143) );
  NOR4_X1 U11194 ( .A1(n10146), .A2(n10145), .A3(n10144), .A4(n10143), .ZN(
        n10271) );
  NAND4_X1 U11195 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_1__SCAN_IN), 
        .A3(P1_ADDR_REG_7__SCAN_IN), .A4(n10185), .ZN(n10157) );
  NAND4_X1 U11196 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .A3(n6056), .A4(n5029), .ZN(n10156) );
  NOR4_X1 U11197 ( .A1(P2_REG1_REG_27__SCAN_IN), .A2(n10160), .A3(n10163), 
        .A4(n10241), .ZN(n10147) );
  NAND3_X1 U11198 ( .A1(n10149), .A2(n10148), .A3(n10147), .ZN(n10155) );
  NOR4_X1 U11199 ( .A1(P1_D_REG_1__SCAN_IN), .A2(SI_9_), .A3(
        P1_REG1_REG_17__SCAN_IN), .A4(P2_REG1_REG_11__SCAN_IN), .ZN(n10153) );
  NOR4_X1 U11200 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n5628), .A3(n10175), .A4(
        n10176), .ZN(n10152) );
  NOR4_X1 U11201 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(SI_2_), .A3(
        P2_REG3_REG_6__SCAN_IN), .A4(n4746), .ZN(n10151) );
  NOR4_X1 U11202 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .A3(P1_ADDR_REG_11__SCAN_IN), .A4(P2_U3152), .ZN(n10150) );
  NAND4_X1 U11203 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10154) );
  NOR4_X1 U11204 ( .A1(n10157), .A2(n10156), .A3(n10155), .A4(n10154), .ZN(
        n10270) );
  AOI22_X1 U11205 ( .A1(n6056), .A2(keyinput13), .B1(keyinput57), .B2(n7878), 
        .ZN(n10158) );
  OAI221_X1 U11206 ( .B1(n6056), .B2(keyinput13), .C1(n7878), .C2(keyinput57), 
        .A(n10158), .ZN(n10170) );
  AOI22_X1 U11207 ( .A1(n10160), .A2(keyinput45), .B1(keyinput25), .B2(n5029), 
        .ZN(n10159) );
  OAI221_X1 U11208 ( .B1(n10160), .B2(keyinput45), .C1(n5029), .C2(keyinput25), 
        .A(n10159), .ZN(n10169) );
  AOI22_X1 U11209 ( .A1(n10163), .A2(keyinput42), .B1(n10162), .B2(keyinput35), 
        .ZN(n10161) );
  OAI221_X1 U11210 ( .B1(n10163), .B2(keyinput42), .C1(n10162), .C2(keyinput35), .A(n10161), .ZN(n10168) );
  XNOR2_X1 U11211 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput33), .ZN(n10166) );
  XNOR2_X1 U11212 ( .A(P1_REG1_REG_17__SCAN_IN), .B(keyinput18), .ZN(n10165)
         );
  NAND2_X1 U11213 ( .A1(n10166), .A2(n10165), .ZN(n10167) );
  NOR4_X1 U11214 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10211) );
  AOI22_X1 U11215 ( .A1(n5628), .A2(keyinput11), .B1(keyinput28), .B2(n5892), 
        .ZN(n10171) );
  OAI221_X1 U11216 ( .B1(n5628), .B2(keyinput11), .C1(n5892), .C2(keyinput28), 
        .A(n10171), .ZN(n10182) );
  AOI22_X1 U11217 ( .A1(n10173), .A2(keyinput60), .B1(keyinput14), .B2(n7264), 
        .ZN(n10172) );
  OAI221_X1 U11218 ( .B1(n10173), .B2(keyinput60), .C1(n7264), .C2(keyinput14), 
        .A(n10172), .ZN(n10181) );
  AOI22_X1 U11219 ( .A1(n10176), .A2(keyinput12), .B1(n10175), .B2(keyinput15), 
        .ZN(n10174) );
  OAI221_X1 U11220 ( .B1(n10176), .B2(keyinput12), .C1(n10175), .C2(keyinput15), .A(n10174), .ZN(n10180) );
  XNOR2_X1 U11221 ( .A(P2_REG1_REG_11__SCAN_IN), .B(keyinput51), .ZN(n10178)
         );
  XNOR2_X1 U11222 ( .A(SI_9_), .B(keyinput48), .ZN(n10177) );
  NAND2_X1 U11223 ( .A1(n10178), .A2(n10177), .ZN(n10179) );
  NOR4_X1 U11224 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10210) );
  AOI22_X1 U11225 ( .A1(n10184), .A2(keyinput26), .B1(n7037), .B2(keyinput63), 
        .ZN(n10183) );
  OAI221_X1 U11226 ( .B1(n10184), .B2(keyinput26), .C1(n7037), .C2(keyinput63), 
        .A(n10183), .ZN(n10193) );
  XNOR2_X1 U11227 ( .A(keyinput31), .B(n4746), .ZN(n10192) );
  XNOR2_X1 U11228 ( .A(keyinput55), .B(n10185), .ZN(n10191) );
  XNOR2_X1 U11229 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput58), .ZN(n10189) );
  XNOR2_X1 U11230 ( .A(SI_2_), .B(keyinput46), .ZN(n10188) );
  XNOR2_X1 U11231 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput7), .ZN(n10187) );
  XNOR2_X1 U11232 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput43), .ZN(n10186) );
  NAND4_X1 U11233 ( .A1(n10189), .A2(n10188), .A3(n10187), .A4(n10186), .ZN(
        n10190) );
  NOR4_X1 U11234 ( .A1(n10193), .A2(n10192), .A3(n10191), .A4(n10190), .ZN(
        n10209) );
  AOI22_X1 U11235 ( .A1(n6061), .A2(keyinput50), .B1(keyinput4), .B2(n10195), 
        .ZN(n10194) );
  OAI221_X1 U11236 ( .B1(n6061), .B2(keyinput50), .C1(n10195), .C2(keyinput4), 
        .A(n10194), .ZN(n10207) );
  INV_X1 U11237 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U11238 ( .A1(n10198), .A2(keyinput5), .B1(keyinput44), .B2(n10197), 
        .ZN(n10196) );
  OAI221_X1 U11239 ( .B1(n10198), .B2(keyinput5), .C1(n10197), .C2(keyinput44), 
        .A(n10196), .ZN(n10206) );
  AOI22_X1 U11240 ( .A1(n10201), .A2(keyinput62), .B1(n10200), .B2(keyinput40), 
        .ZN(n10199) );
  OAI221_X1 U11241 ( .B1(n10201), .B2(keyinput62), .C1(n10200), .C2(keyinput40), .A(n10199), .ZN(n10205) );
  XNOR2_X1 U11242 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(keyinput3), .ZN(n10203)
         );
  XNOR2_X1 U11243 ( .A(P1_REG1_REG_14__SCAN_IN), .B(keyinput59), .ZN(n10202)
         );
  NAND2_X1 U11244 ( .A1(n10203), .A2(n10202), .ZN(n10204) );
  NOR4_X1 U11245 ( .A1(n10207), .A2(n10206), .A3(n10205), .A4(n10204), .ZN(
        n10208) );
  NAND4_X1 U11246 ( .A1(n10211), .A2(n10210), .A3(n10209), .A4(n10208), .ZN(
        n10269) );
  AOI22_X1 U11247 ( .A1(n10213), .A2(keyinput52), .B1(n5396), .B2(keyinput0), 
        .ZN(n10212) );
  OAI221_X1 U11248 ( .B1(n10213), .B2(keyinput52), .C1(n5396), .C2(keyinput0), 
        .A(n10212), .ZN(n10225) );
  AOI22_X1 U11249 ( .A1(n10216), .A2(keyinput34), .B1(n10215), .B2(keyinput23), 
        .ZN(n10214) );
  OAI221_X1 U11250 ( .B1(n10216), .B2(keyinput34), .C1(n10215), .C2(keyinput23), .A(n10214), .ZN(n10224) );
  AOI22_X1 U11251 ( .A1(n10218), .A2(keyinput9), .B1(n5973), .B2(keyinput8), 
        .ZN(n10217) );
  OAI221_X1 U11252 ( .B1(n10218), .B2(keyinput9), .C1(n5973), .C2(keyinput8), 
        .A(n10217), .ZN(n10223) );
  AOI22_X1 U11253 ( .A1(n10221), .A2(keyinput20), .B1(keyinput30), .B2(n10220), 
        .ZN(n10219) );
  OAI221_X1 U11254 ( .B1(n10221), .B2(keyinput20), .C1(n10220), .C2(keyinput30), .A(n10219), .ZN(n10222) );
  NOR4_X1 U11255 ( .A1(n10225), .A2(n10224), .A3(n10223), .A4(n10222), .ZN(
        n10267) );
  AOI22_X1 U11256 ( .A1(n10227), .A2(keyinput1), .B1(n6095), .B2(keyinput61), 
        .ZN(n10226) );
  OAI221_X1 U11257 ( .B1(n10227), .B2(keyinput1), .C1(n6095), .C2(keyinput61), 
        .A(n10226), .ZN(n10238) );
  AOI22_X1 U11258 ( .A1(n10229), .A2(keyinput36), .B1(keyinput37), .B2(n6925), 
        .ZN(n10228) );
  OAI221_X1 U11259 ( .B1(n10229), .B2(keyinput36), .C1(n6925), .C2(keyinput37), 
        .A(n10228), .ZN(n10237) );
  AOI22_X1 U11260 ( .A1(n10232), .A2(keyinput21), .B1(keyinput29), .B2(n10231), 
        .ZN(n10230) );
  OAI221_X1 U11261 ( .B1(n10232), .B2(keyinput21), .C1(n10231), .C2(keyinput29), .A(n10230), .ZN(n10236) );
  XOR2_X1 U11262 ( .A(n8546), .B(keyinput16), .Z(n10234) );
  XNOR2_X1 U11263 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput53), .ZN(n10233) );
  NAND2_X1 U11264 ( .A1(n10234), .A2(n10233), .ZN(n10235) );
  NOR4_X1 U11265 ( .A1(n10238), .A2(n10237), .A3(n10236), .A4(n10235), .ZN(
        n10266) );
  AOI22_X1 U11266 ( .A1(n10241), .A2(keyinput39), .B1(n10240), .B2(keyinput27), 
        .ZN(n10239) );
  OAI221_X1 U11267 ( .B1(n10241), .B2(keyinput39), .C1(n10240), .C2(keyinput27), .A(n10239), .ZN(n10252) );
  INV_X1 U11268 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U11269 ( .A1(n10243), .A2(keyinput38), .B1(keyinput10), .B2(n5417), 
        .ZN(n10242) );
  OAI221_X1 U11270 ( .B1(n10243), .B2(keyinput38), .C1(n5417), .C2(keyinput10), 
        .A(n10242), .ZN(n10251) );
  AOI22_X1 U11271 ( .A1(n10246), .A2(keyinput54), .B1(n10245), .B2(keyinput47), 
        .ZN(n10244) );
  OAI221_X1 U11272 ( .B1(n10246), .B2(keyinput54), .C1(n10245), .C2(keyinput47), .A(n10244), .ZN(n10250) );
  AOI22_X1 U11273 ( .A1(n6535), .A2(keyinput41), .B1(n10248), .B2(keyinput32), 
        .ZN(n10247) );
  OAI221_X1 U11274 ( .B1(n6535), .B2(keyinput41), .C1(n10248), .C2(keyinput32), 
        .A(n10247), .ZN(n10249) );
  NOR4_X1 U11275 ( .A1(n10252), .A2(n10251), .A3(n10250), .A4(n10249), .ZN(
        n10265) );
  INV_X1 U11276 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U11277 ( .A1(n10254), .A2(keyinput19), .B1(n6902), .B2(keyinput2), 
        .ZN(n10253) );
  OAI221_X1 U11278 ( .B1(n10254), .B2(keyinput19), .C1(n6902), .C2(keyinput2), 
        .A(n10253), .ZN(n10263) );
  AOI22_X1 U11279 ( .A1(n7239), .A2(keyinput17), .B1(n10256), .B2(keyinput6), 
        .ZN(n10255) );
  OAI221_X1 U11280 ( .B1(n7239), .B2(keyinput17), .C1(n10256), .C2(keyinput6), 
        .A(n10255), .ZN(n10262) );
  XNOR2_X1 U11281 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput56), .ZN(n10260) );
  XNOR2_X1 U11282 ( .A(P2_D_REG_0__SCAN_IN), .B(keyinput49), .ZN(n10259) );
  XNOR2_X1 U11283 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput22), .ZN(n10258) );
  XNOR2_X1 U11284 ( .A(P1_REG1_REG_30__SCAN_IN), .B(keyinput24), .ZN(n10257)
         );
  NAND4_X1 U11285 ( .A1(n10260), .A2(n10259), .A3(n10258), .A4(n10257), .ZN(
        n10261) );
  NOR3_X1 U11286 ( .A1(n10263), .A2(n10262), .A3(n10261), .ZN(n10264) );
  NAND4_X1 U11287 ( .A1(n10267), .A2(n10266), .A3(n10265), .A4(n10264), .ZN(
        n10268) );
  AOI211_X1 U11288 ( .C1(n10271), .C2(n10270), .A(n10269), .B(n10268), .ZN(
        n10272) );
  XOR2_X1 U11289 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10272), .Z(n10277) );
  INV_X1 U11290 ( .A(n10273), .ZN(n10274) );
  NAND2_X1 U11291 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  XNOR2_X1 U11292 ( .A(n10277), .B(n10276), .ZN(ADD_1071_U48) );
  CLKBUF_X1 U4786 ( .A(n6807), .Z(n4276) );
  CLKBUF_X1 U4791 ( .A(n5771), .Z(n4404) );
  AND2_X1 U4827 ( .A1(n7662), .A2(n7558), .ZN(n6752) );
  CLKBUF_X1 U5060 ( .A(n5651), .Z(n7100) );
  CLKBUF_X1 U5484 ( .A(n5126), .Z(n6524) );
  CLKBUF_X1 U5795 ( .A(n5075), .Z(n5336) );
  BUF_X2 U6036 ( .A(n8068), .Z(n4282) );
endmodule

