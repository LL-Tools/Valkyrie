

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4282, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165;

  AND2_X1 U4788 ( .A1(n6221), .A2(n6220), .ZN(n8423) );
  INV_X1 U4789 ( .A(n9274), .ZN(n9276) );
  INV_X1 U4790 ( .A(n8106), .ZN(n9686) );
  INV_X1 U4791 ( .A(n5517), .ZN(n5634) );
  OR2_X1 U4792 ( .A1(n6086), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6097) );
  CLKBUF_X2 U4793 ( .A(n5078), .Z(n5616) );
  INV_X1 U4794 ( .A(n6561), .ZN(n5060) );
  NOR2_X1 U4796 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6003) );
  INV_X2 U4797 ( .A(n5065), .ZN(n5105) );
  CLKBUF_X1 U4798 ( .A(n9126), .Z(n4282) );
  OAI21_X1 U4799 ( .B1(n5717), .B2(n7064), .A(n9531), .ZN(n9126) );
  OR2_X2 U4800 ( .A1(n6146), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6161) );
  OAI21_X2 U4802 ( .B1(n4659), .B2(n4658), .A(n4656), .ZN(n9280) );
  NAND2_X1 U4803 ( .A1(n5078), .A2(n5113), .ZN(n5104) );
  INV_X1 U4804 ( .A(n5517), .ZN(n5659) );
  NAND2_X1 U4805 ( .A1(n7193), .A2(n7284), .ZN(n6448) );
  NOR2_X1 U4806 ( .A1(n5860), .A2(n8459), .ZN(n8487) );
  INV_X1 U4807 ( .A(n5991), .ZN(n6132) );
  INV_X1 U4808 ( .A(n7942), .ZN(n7963) );
  OR2_X1 U4809 ( .A1(n6014), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6020) );
  OR2_X1 U4810 ( .A1(n5959), .A2(n5846), .ZN(n5960) );
  CLKBUF_X3 U4811 ( .A(n5125), .Z(n5671) );
  INV_X1 U4812 ( .A(n5128), .ZN(n6364) );
  NAND2_X2 U4813 ( .A1(n6469), .A2(n4285), .ZN(n5128) );
  XNOR2_X1 U4814 ( .A(n8823), .B(n8607), .ZN(n8588) );
  AND2_X2 U4816 ( .A1(n9547), .A2(n9958), .ZN(n4313) );
  XNOR2_X2 U4817 ( .A(n5960), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5961) );
  AND4_X2 U4818 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n6926)
         );
  NOR2_X2 U4819 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5825) );
  BUF_X4 U4820 ( .A(n5723), .Z(n4285) );
  XNOR2_X2 U4821 ( .A(n5763), .B(n5762), .ZN(n7667) );
  NAND2_X2 U4822 ( .A1(n5754), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5763) );
  AND2_X2 U4823 ( .A1(n9119), .A2(n5271), .ZN(n5290) );
  OAI211_X2 U4824 ( .C1(n6873), .C2(n4300), .A(n5267), .B(n9120), .ZN(n9119)
         );
  BUF_X8 U4825 ( .A(n4902), .Z(n6362) );
  NOR4_X2 U4826 ( .A1(n7969), .A2(n7792), .A3(n7791), .A4(n7950), .ZN(n7793)
         );
  XNOR2_X2 U4827 ( .A(n5011), .B(n5010), .ZN(n8049) );
  XNOR2_X1 U4828 ( .A(n5827), .B(n5826), .ZN(n5833) );
  NAND2_X1 U4829 ( .A1(n8336), .A2(n4415), .ZN(n8394) );
  NOR2_X1 U4830 ( .A1(n8536), .A2(n8537), .ZN(n8535) );
  AOI21_X1 U4831 ( .B1(n4291), .B2(n4672), .A(n4671), .ZN(n4670) );
  OR2_X1 U4832 ( .A1(n5867), .A2(n4421), .ZN(n8536) );
  AND2_X1 U4833 ( .A1(n4422), .A2(n6965), .ZN(n5867) );
  NOR2_X1 U4834 ( .A1(n4422), .A2(n6965), .ZN(n4421) );
  NAND2_X1 U4835 ( .A1(n4424), .A2(n4423), .ZN(n4422) );
  OAI21_X1 U4836 ( .B1(n8495), .B2(n4740), .A(n4739), .ZN(n8524) );
  OAI21_X1 U4837 ( .B1(n9666), .B2(n9290), .A(n9289), .ZN(n9456) );
  NOR2_X1 U4838 ( .A1(n8487), .A2(n8486), .ZN(n8485) );
  NOR2_X1 U4839 ( .A1(n9491), .A2(n9474), .ZN(n9473) );
  INV_X1 U4840 ( .A(n7592), .ZN(n4659) );
  AND3_X1 U4841 ( .A1(n4733), .A2(n4363), .A3(n4734), .ZN(n5859) );
  NAND2_X1 U4842 ( .A1(n5409), .A2(n5408), .ZN(n9529) );
  XNOR2_X1 U4843 ( .A(n5855), .B(n7349), .ZN(n7351) );
  NAND2_X1 U4844 ( .A1(n5048), .A2(n4973), .ZN(n5432) );
  OR2_X1 U4845 ( .A1(n6740), .A2(n6739), .ZN(n4306) );
  AND3_X1 U4846 ( .A1(n4418), .A2(n6012), .A3(n4417), .ZN(n10039) );
  NAND2_X1 U4847 ( .A1(n5209), .A2(n5208), .ZN(n7263) );
  NAND2_X1 U4848 ( .A1(n5193), .A2(n5192), .ZN(n7012) );
  INV_X1 U4849 ( .A(n7303), .ZN(n9943) );
  INV_X1 U4850 ( .A(n8452), .ZN(n6987) );
  OR2_X1 U4851 ( .A1(n6576), .A2(n6869), .ZN(n6574) );
  NAND4_X1 U4852 ( .A1(n5998), .A2(n5997), .A3(n5996), .A4(n5995), .ZN(n8452)
         );
  NAND2_X1 U4853 ( .A1(n8453), .A2(n10020), .ZN(n7841) );
  INV_X1 U4854 ( .A(n8051), .ZN(n4629) );
  INV_X1 U4855 ( .A(n5104), .ZN(n5517) );
  INV_X2 U4856 ( .A(n9940), .ZN(n9941) );
  INV_X1 U4857 ( .A(n6925), .ZN(n8453) );
  AND4_X1 U4858 ( .A1(n5989), .A2(n5988), .A3(n5987), .A4(n5986), .ZN(n6925)
         );
  XNOR2_X1 U4860 ( .A(n5785), .B(n5784), .ZN(n7193) );
  NAND4_X1 U4861 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n9184)
         );
  INV_X1 U4862 ( .A(n6666), .ZN(n7025) );
  INV_X2 U4863 ( .A(n5992), .ZN(n7758) );
  XNOR2_X1 U4864 ( .A(n5757), .B(n5756), .ZN(n7731) );
  OR2_X2 U4865 ( .A1(n7541), .A2(n5009), .ZN(n5708) );
  NAND2_X1 U4866 ( .A1(n5790), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U4867 ( .A1(n5755), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5757) );
  INV_X1 U4868 ( .A(n8232), .ZN(n7254) );
  AND2_X1 U4869 ( .A1(n5017), .A2(n5016), .ZN(n8232) );
  XNOR2_X1 U4870 ( .A(n5008), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7568) );
  MUX2_X1 U4871 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5777), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5779) );
  XNOR2_X1 U4872 ( .A(n5029), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U4873 ( .A1(n5007), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5008) );
  XNOR2_X1 U4874 ( .A(n4914), .B(SI_5_), .ZN(n5188) );
  AND2_X1 U4875 ( .A1(n5012), .A2(n4998), .ZN(n5015) );
  OAI21_X1 U4876 ( .B1(n9687), .B2(n9689), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5029) );
  NAND2_X1 U4877 ( .A1(n4460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5006) );
  AND2_X1 U4878 ( .A1(n4997), .A2(n4996), .ZN(n5012) );
  INV_X1 U4879 ( .A(n4892), .ZN(n4902) );
  AND2_X1 U4880 ( .A1(n5752), .A2(n8945), .ZN(n4401) );
  NOR2_X1 U4881 ( .A1(n5320), .A2(n4991), .ZN(n4997) );
  AND4_X1 U4882 ( .A1(n4980), .A2(n5096), .A3(n4307), .A4(n4979), .ZN(n4777)
         );
  NOR2_X1 U4883 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  AND3_X1 U4884 ( .A1(n4998), .A2(n5041), .A3(n5010), .ZN(n4985) );
  AND4_X1 U4885 ( .A1(n4977), .A2(n4976), .A3(n5297), .A4(n4975), .ZN(n4980)
         );
  INV_X1 U4886 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5803) );
  INV_X1 U4887 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5798) );
  INV_X1 U4888 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5796) );
  INV_X1 U4889 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5808) );
  INV_X1 U4890 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5816) );
  INV_X1 U4891 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5826) );
  INV_X1 U4892 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4975) );
  INV_X4 U4893 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U4894 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4977) );
  NOR2_X1 U4895 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n4748) );
  NOR2_X1 U4896 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4623) );
  INV_X4 U4897 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4898 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5372) );
  INV_X1 U4899 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5368) );
  NOR2_X1 U4900 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4624) );
  INV_X1 U4901 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5748) );
  AND2_X4 U4902 ( .A1(n5962), .A2(n7736), .ZN(n6125) );
  OAI22_X2 U4903 ( .A1(n7591), .A2(n7590), .B1(n9176), .B2(n9779), .ZN(n7592)
         );
  OAI21_X2 U4904 ( .B1(n9915), .B2(n4636), .A(n4635), .ZN(n7591) );
  NOR2_X2 U4905 ( .A1(n9093), .A2(n9092), .ZN(n9101) );
  BUF_X4 U4906 ( .A(n5091), .Z(n4287) );
  INV_X1 U4907 ( .A(n5078), .ZN(n5091) );
  INV_X1 U4908 ( .A(n7060), .ZN(n5061) );
  OR2_X1 U4909 ( .A1(n8835), .A2(n8349), .ZN(n7939) );
  XNOR2_X1 U4910 ( .A(n5264), .B(n5616), .ZN(n5268) );
  INV_X1 U4911 ( .A(n7739), .ZN(n5030) );
  OAI21_X1 U4912 ( .B1(n4288), .B2(n4650), .A(n4655), .ZN(n4649) );
  OR2_X1 U4913 ( .A1(n9474), .A2(n9288), .ZN(n4655) );
  NAND2_X1 U4914 ( .A1(n4391), .A2(n5599), .ZN(n5625) );
  NAND2_X1 U4915 ( .A1(n5598), .A2(n5597), .ZN(n4391) );
  NAND2_X1 U4916 ( .A1(n4387), .A2(n4953), .ZN(n5366) );
  NAND2_X1 U4917 ( .A1(n4912), .A2(n4911), .ZN(n5187) );
  AND2_X1 U4918 ( .A1(n5962), .A2(n5961), .ZN(n5993) );
  NAND2_X1 U4919 ( .A1(n5820), .A2(n5835), .ZN(n5837) );
  OAI21_X1 U4920 ( .B1(n8220), .B2(n8219), .A(n8218), .ZN(n8229) );
  NAND2_X1 U4921 ( .A1(n8818), .A2(n7766), .ZN(n7964) );
  NAND2_X1 U4922 ( .A1(n8583), .A2(n8441), .ZN(n7747) );
  INV_X1 U4923 ( .A(n4810), .ZN(n4806) );
  OAI21_X1 U4924 ( .B1(n4711), .B2(n4709), .A(n4968), .ZN(n4708) );
  NAND2_X1 U4925 ( .A1(n4924), .A2(n4923), .ZN(n4927) );
  XNOR2_X1 U4926 ( .A(n6714), .B(n6459), .ZN(n6451) );
  NAND2_X1 U4927 ( .A1(n7964), .A2(n7747), .ZN(n7948) );
  OR2_X1 U4928 ( .A1(n8583), .A2(n8441), .ZN(n7790) );
  INV_X1 U4929 ( .A(n4853), .ZN(n4852) );
  OAI21_X1 U4930 ( .B1(n6693), .B2(n4854), .A(n6398), .ZN(n4853) );
  INV_X1 U4931 ( .A(n5882), .ZN(n4854) );
  AOI21_X1 U4932 ( .B1(n4818), .B2(n4816), .A(n4333), .ZN(n4815) );
  INV_X1 U4933 ( .A(n4820), .ZN(n4816) );
  INV_X1 U4934 ( .A(n4818), .ZN(n4817) );
  INV_X1 U4935 ( .A(n6521), .ZN(n6515) );
  NAND2_X1 U4936 ( .A1(n8454), .A2(n6515), .ZN(n7833) );
  INV_X1 U4937 ( .A(n5992), .ZN(n5985) );
  AND2_X1 U4938 ( .A1(n8829), .A2(n8617), .ZN(n6298) );
  INV_X1 U4939 ( .A(n4827), .ZN(n4826) );
  OAI21_X1 U4940 ( .B1(n8664), .B2(n4828), .A(n6292), .ZN(n4827) );
  OR2_X1 U4941 ( .A1(n8996), .A2(n8270), .ZN(n7921) );
  NAND2_X1 U4942 ( .A1(n6280), .A2(n4310), .ZN(n4840) );
  OR2_X1 U4943 ( .A1(n8253), .A2(n9733), .ZN(n7899) );
  NOR2_X1 U4944 ( .A1(n5865), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n5782) );
  OR2_X1 U4945 ( .A1(n4802), .A2(n4801), .ZN(n4800) );
  INV_X1 U4946 ( .A(n9145), .ZN(n4492) );
  CLKBUF_X1 U4947 ( .A(n5697), .Z(n8225) );
  NAND2_X1 U4948 ( .A1(n5553), .A2(n5552), .ZN(n5576) );
  OAI21_X1 U4949 ( .B1(n5432), .B2(n4699), .A(n4381), .ZN(n5527) );
  AOI21_X1 U4950 ( .B1(n4698), .B2(n4382), .A(n4358), .ZN(n4381) );
  INV_X1 U4951 ( .A(n4702), .ZN(n4382) );
  AOI21_X1 U4952 ( .B1(n4702), .B2(n5431), .A(n4360), .ZN(n4701) );
  NAND2_X1 U4953 ( .A1(n4384), .A2(n4949), .ZN(n5345) );
  NAND2_X1 U4954 ( .A1(n4945), .A2(n4385), .ZN(n4384) );
  XNOR2_X1 U4955 ( .A(n4917), .B(SI_6_), .ZN(n5165) );
  NAND2_X1 U4956 ( .A1(n8406), .A2(n4354), .ZN(n8323) );
  INV_X1 U4957 ( .A(n8321), .ZN(n8263) );
  NAND2_X1 U4958 ( .A1(n4408), .A2(n6915), .ZN(n4407) );
  OR2_X1 U4959 ( .A1(n8818), .A2(n7766), .ZN(n7794) );
  INV_X1 U4960 ( .A(n6013), .ZN(n6243) );
  AND2_X1 U4961 ( .A1(n7737), .A2(n7736), .ZN(n6002) );
  XNOR2_X1 U4962 ( .A(n5918), .B(n5916), .ZN(n4400) );
  OR2_X1 U4963 ( .A1(n6578), .A2(n5881), .ZN(n6692) );
  NOR2_X1 U4964 ( .A1(n6835), .A2(n7132), .ZN(n6945) );
  NAND2_X1 U4965 ( .A1(n7159), .A2(n7160), .ZN(n7158) );
  NAND2_X1 U4966 ( .A1(n4724), .A2(n4722), .ZN(n4729) );
  AND2_X1 U4967 ( .A1(n4725), .A2(n4301), .ZN(n4722) );
  OR2_X1 U4968 ( .A1(n7311), .A2(n5884), .ZN(n5886) );
  NAND2_X1 U4969 ( .A1(n4480), .A2(n4479), .ZN(n4478) );
  INV_X1 U4970 ( .A(n7410), .ZN(n4479) );
  NOR2_X1 U4971 ( .A1(n8497), .A2(n8498), .ZN(n8496) );
  OAI21_X1 U4972 ( .B1(n8533), .B2(n4866), .A(n4865), .ZN(n8555) );
  NAND2_X1 U4973 ( .A1(n4867), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4866) );
  NAND2_X1 U4974 ( .A1(n5896), .A2(n4867), .ZN(n4865) );
  INV_X1 U4975 ( .A(n8556), .ZN(n4867) );
  NAND2_X1 U4976 ( .A1(n6212), .A2(n7939), .ZN(n8602) );
  OR2_X1 U4977 ( .A1(n8799), .A2(n8386), .ZN(n7812) );
  OR2_X1 U4978 ( .A1(n8809), .A2(n8432), .ZN(n7901) );
  INV_X1 U4979 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4403) );
  INV_X1 U4980 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5835) );
  OAI21_X1 U4981 ( .B1(P2_IR_REG_1__SCAN_IN), .B2(n5846), .A(n4486), .ZN(n5830) );
  NAND2_X1 U4982 ( .A1(n4487), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n4486) );
  NAND2_X1 U4983 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4487) );
  XNOR2_X1 U4984 ( .A(n4488), .B(n4287), .ZN(n4776) );
  NAND2_X1 U4985 ( .A1(n5104), .A2(n6666), .ZN(n4372) );
  XNOR2_X1 U4986 ( .A(n5112), .B(n5616), .ZN(n5114) );
  AOI21_X1 U4987 ( .B1(n8229), .B2(n8237), .A(n8049), .ZN(n4556) );
  AND4_X1 U4989 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n9312)
         );
  AND4_X1 U4990 ( .A1(n5380), .A2(n5379), .A3(n5378), .A4(n5377), .ZN(n8111)
         );
  INV_X1 U4991 ( .A(n4649), .ZN(n4648) );
  NAND2_X1 U4992 ( .A1(n6818), .A2(n4633), .ZN(n7299) );
  NAND2_X1 U4993 ( .A1(n7029), .A2(n4634), .ZN(n4633) );
  NAND2_X1 U4994 ( .A1(n8041), .A2(n8040), .ZN(n9253) );
  XNOR2_X1 U4995 ( .A(n5651), .B(n5650), .ZN(n7634) );
  NAND2_X1 U4996 ( .A1(n4494), .A2(n4493), .ZN(n5042) );
  AOI21_X1 U4997 ( .B1(n4496), .B2(n9688), .A(n9688), .ZN(n4493) );
  NAND2_X1 U4998 ( .A1(n4713), .A2(n4958), .ZN(n5384) );
  NAND2_X1 U4999 ( .A1(n4512), .A2(n4907), .ZN(n5144) );
  NAND2_X1 U5000 ( .A1(n4373), .A2(n5126), .ZN(n4512) );
  NAND2_X1 U5001 ( .A1(n9998), .A2(n9997), .ZN(n9996) );
  OAI21_X1 U5002 ( .B1(n6624), .B2(n10083), .A(n5875), .ZN(n9997) );
  NAND2_X1 U5003 ( .A1(n6604), .A2(n6603), .ZN(n6602) );
  OAI21_X1 U5004 ( .B1(n6945), .B2(n6944), .A(n6943), .ZN(n6947) );
  NOR2_X1 U5005 ( .A1(n7345), .A2(n10103), .ZN(n7344) );
  NOR2_X1 U5006 ( .A1(n8458), .A2(n9752), .ZN(n8457) );
  OR2_X1 U5007 ( .A1(n8477), .A2(n8476), .ZN(n4485) );
  OR2_X1 U5008 ( .A1(n8515), .A2(n8514), .ZN(n4482) );
  NOR2_X1 U5009 ( .A1(n8564), .A2(n8563), .ZN(n8562) );
  OAI211_X1 U5010 ( .C1(n8587), .C2(n7610), .A(n6311), .B(n6310), .ZN(n8579)
         );
  NAND2_X1 U5011 ( .A1(n6223), .A2(n6222), .ZN(n8823) );
  NAND2_X1 U5012 ( .A1(n4442), .A2(n4439), .ZN(n7830) );
  INV_X1 U5013 ( .A(n4440), .ZN(n4439) );
  NAND2_X1 U5014 ( .A1(n7822), .A2(n7821), .ZN(n4442) );
  AOI21_X1 U5015 ( .B1(n7826), .B2(n7820), .A(n7821), .ZN(n4440) );
  NAND2_X1 U5016 ( .A1(n7855), .A2(n7963), .ZN(n4438) );
  NAND2_X1 U5017 ( .A1(n4434), .A2(n7942), .ZN(n4433) );
  NAND2_X1 U5018 ( .A1(n4437), .A2(n4435), .ZN(n4434) );
  INV_X1 U5019 ( .A(n4436), .ZN(n4435) );
  OAI21_X1 U5020 ( .B1(n7851), .B2(n7845), .A(n4327), .ZN(n4437) );
  NOR2_X1 U5021 ( .A1(n8161), .A2(n4570), .ZN(n4569) );
  NOR2_X1 U5022 ( .A1(n8153), .A2(n8154), .ZN(n4570) );
  OAI21_X1 U5023 ( .B1(n4453), .B2(n4452), .A(n4451), .ZN(n7898) );
  NAND2_X1 U5024 ( .A1(n7892), .A2(n7891), .ZN(n4452) );
  NAND2_X1 U5025 ( .A1(n8660), .A2(n7923), .ZN(n4447) );
  INV_X1 U5026 ( .A(n7930), .ZN(n4450) );
  NAND2_X1 U5027 ( .A1(n4557), .A2(n8179), .ZN(n8184) );
  INV_X1 U5028 ( .A(n7456), .ZN(n8060) );
  NAND2_X1 U5029 ( .A1(n4710), .A2(n4962), .ZN(n4709) );
  INV_X1 U5030 ( .A(n5405), .ZN(n4710) );
  AND2_X1 U5031 ( .A1(n8847), .A2(n8282), .ZN(n7769) );
  AND2_X1 U5032 ( .A1(n4810), .A2(n9063), .ZN(n4801) );
  INV_X1 U5033 ( .A(n7400), .ZN(n4785) );
  NAND2_X1 U5034 ( .A1(n8202), .A2(n4314), .ZN(n4577) );
  NAND2_X1 U5035 ( .A1(n4580), .A2(n4579), .ZN(n4578) );
  INV_X1 U5036 ( .A(n8202), .ZN(n4579) );
  NAND2_X1 U5037 ( .A1(n4581), .A2(n4319), .ZN(n4580) );
  INV_X1 U5038 ( .A(n6233), .ZN(n4693) );
  INV_X1 U5039 ( .A(n4709), .ZN(n4705) );
  NOR2_X1 U5040 ( .A1(n4950), .A2(n4386), .ZN(n4385) );
  INV_X1 U5041 ( .A(n4944), .ZN(n4386) );
  NAND2_X1 U5042 ( .A1(n8394), .A2(n4355), .ZN(n8280) );
  AOI21_X1 U5043 ( .B1(n7767), .B2(n7284), .A(n6449), .ZN(n6450) );
  NAND2_X1 U5044 ( .A1(n6446), .A2(n4775), .ZN(n4774) );
  INV_X1 U5045 ( .A(n6447), .ZN(n4775) );
  INV_X1 U5046 ( .A(n8418), .ZN(n4759) );
  NOR2_X1 U5047 ( .A1(n7966), .A2(n7792), .ZN(n4679) );
  INV_X1 U5048 ( .A(n6693), .ZN(n4850) );
  AND2_X1 U5049 ( .A1(n5882), .A2(n6842), .ZN(n4855) );
  OR2_X1 U5050 ( .A1(n7321), .A2(n4361), .ZN(n5855) );
  INV_X1 U5051 ( .A(n7943), .ZN(n4616) );
  INV_X1 U5052 ( .A(n4615), .ZN(n4614) );
  OAI21_X1 U5053 ( .B1(n8601), .B2(n4616), .A(n8588), .ZN(n4615) );
  INV_X1 U5054 ( .A(n4847), .ZN(n4846) );
  OAI21_X1 U5055 ( .B1(n8603), .B2(n6298), .A(n4325), .ZN(n4847) );
  OR2_X1 U5056 ( .A1(n10071), .A2(n7559), .ZN(n7885) );
  NAND2_X1 U5057 ( .A1(n6273), .A2(n4311), .ZN(n4842) );
  NAND2_X1 U5058 ( .A1(n4819), .A2(n4822), .ZN(n4818) );
  NAND2_X1 U5059 ( .A1(n4831), .A2(n4830), .ZN(n7126) );
  NAND2_X1 U5060 ( .A1(n4343), .A2(n6268), .ZN(n4830) );
  NAND2_X1 U5061 ( .A1(n7848), .A2(n4605), .ZN(n4609) );
  INV_X1 U5062 ( .A(n7844), .ZN(n4605) );
  INV_X1 U5063 ( .A(n7936), .ZN(n4585) );
  NOR2_X1 U5064 ( .A1(n7769), .A2(n7809), .ZN(n4590) );
  OR2_X1 U5065 ( .A1(n8841), .A2(n8287), .ZN(n7935) );
  OR2_X1 U5066 ( .A1(n8847), .A2(n8282), .ZN(n7933) );
  AND2_X1 U5067 ( .A1(n8320), .A2(n8665), .ZN(n7925) );
  NAND2_X1 U5068 ( .A1(n4838), .A2(n6285), .ZN(n4837) );
  NAND2_X1 U5069 ( .A1(n4318), .A2(n4839), .ZN(n4835) );
  INV_X1 U5070 ( .A(n6285), .ZN(n4839) );
  NAND2_X1 U5071 ( .A1(n5760), .A2(n4457), .ZN(n5776) );
  AND2_X1 U5072 ( .A1(n5759), .A2(n4458), .ZN(n4457) );
  INV_X1 U5073 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4458) );
  AND2_X1 U5074 ( .A1(n4515), .A2(n4514), .ZN(n4892) );
  INV_X1 U5075 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4519) );
  XNOR2_X1 U5076 ( .A(n5492), .B(n5616), .ZN(n5494) );
  OAI22_X1 U5077 ( .A1(n9295), .A2(n5593), .B1(n9293), .B2(n5676), .ZN(n5493)
         );
  XNOR2_X1 U5078 ( .A(n5156), .B(n4287), .ZN(n5159) );
  INV_X1 U5079 ( .A(n5250), .ZN(n4779) );
  NAND2_X1 U5080 ( .A1(n4799), .A2(n4801), .ZN(n4798) );
  INV_X1 U5081 ( .A(n4807), .ZN(n4799) );
  AOI21_X1 U5082 ( .B1(n4804), .B2(n4806), .A(n4803), .ZN(n4802) );
  INV_X1 U5083 ( .A(n9062), .ZN(n4803) );
  INV_X1 U5084 ( .A(n9773), .ZN(n4794) );
  AND2_X1 U5085 ( .A1(n4787), .A2(n4793), .ZN(n4786) );
  AND2_X1 U5086 ( .A1(n4787), .A2(n4794), .ZN(n4791) );
  INV_X1 U5087 ( .A(n9756), .ZN(n4793) );
  OAI21_X1 U5088 ( .B1(n8214), .B2(n8213), .A(n8212), .ZN(n8217) );
  NOR2_X1 U5089 ( .A1(n8211), .A2(n8210), .ZN(n8212) );
  OR2_X1 U5090 ( .A1(n9556), .A2(n9162), .ZN(n8045) );
  NOR2_X1 U5091 ( .A1(n9556), .A2(n9563), .ZN(n4464) );
  OR2_X1 U5092 ( .A1(n9563), .A2(n9312), .ZN(n8198) );
  NAND2_X1 U5093 ( .A1(n4534), .A2(n4532), .ZN(n9434) );
  AOI21_X1 U5094 ( .B1(n4535), .B2(n4536), .A(n4533), .ZN(n4532) );
  INV_X1 U5095 ( .A(n9259), .ZN(n4533) );
  NOR2_X1 U5096 ( .A1(n5410), .A2(n9094), .ZN(n5052) );
  NOR2_X1 U5097 ( .A1(n8110), .A2(n9779), .ZN(n4465) );
  NOR2_X1 U5098 ( .A1(n4644), .A2(n7450), .ZN(n4637) );
  OAI21_X1 U5099 ( .B1(n8064), .B2(n4290), .A(n7523), .ZN(n4642) );
  INV_X1 U5100 ( .A(n4550), .ZN(n4549) );
  OAI21_X1 U5101 ( .B1(n9260), .B2(n9263), .A(n9262), .ZN(n4550) );
  NAND2_X1 U5102 ( .A1(n7662), .A2(n7661), .ZN(n4389) );
  OR2_X1 U5103 ( .A1(n7660), .A2(n7659), .ZN(n7661) );
  INV_X1 U5104 ( .A(n5650), .ZN(n4697) );
  AOI21_X1 U5105 ( .B1(n5650), .B2(n4696), .A(n4695), .ZN(n4694) );
  INV_X1 U5106 ( .A(n5626), .ZN(n4696) );
  INV_X1 U5107 ( .A(n5652), .ZN(n4695) );
  NAND2_X1 U5108 ( .A1(n5625), .A2(n5624), .ZN(n5627) );
  NAND2_X1 U5109 ( .A1(n4677), .A2(n5577), .ZN(n5598) );
  NOR2_X1 U5110 ( .A1(n4963), .A2(n4712), .ZN(n4711) );
  INV_X1 U5111 ( .A(n4958), .ZN(n4712) );
  OR2_X1 U5112 ( .A1(n5366), .A2(n5365), .ZN(n4713) );
  XNOR2_X1 U5113 ( .A(n4947), .B(SI_12_), .ZN(n5319) );
  AND2_X1 U5114 ( .A1(n4942), .A2(n5293), .ZN(n4943) );
  XNOR2_X1 U5115 ( .A(n4940), .B(SI_10_), .ZN(n5272) );
  INV_X1 U5116 ( .A(n4525), .ZN(n4522) );
  OAI21_X1 U5117 ( .B1(n4913), .B2(n4526), .A(n4916), .ZN(n4525) );
  INV_X1 U5118 ( .A(n5165), .ZN(n4916) );
  NAND2_X1 U5119 ( .A1(n4927), .A2(n4926), .ZN(n5227) );
  AOI21_X1 U5120 ( .B1(n4919), .B2(n4690), .A(n4336), .ZN(n4689) );
  INV_X1 U5121 ( .A(n4918), .ZN(n4690) );
  OR2_X1 U5122 ( .A1(n8272), .A2(n8332), .ZN(n8335) );
  INV_X1 U5123 ( .A(n6723), .ZN(n6720) );
  OAI21_X1 U5124 ( .B1(n6915), .B2(n4410), .A(n4408), .ZN(n7274) );
  AND2_X1 U5125 ( .A1(n7434), .A2(n7436), .ZN(n4771) );
  NAND2_X1 U5126 ( .A1(n7544), .A2(n4414), .ZN(n4413) );
  INV_X1 U5127 ( .A(n7439), .ZN(n4414) );
  XNOR2_X1 U5128 ( .A(n6714), .B(n10039), .ZN(n6909) );
  INV_X1 U5129 ( .A(n8451), .ZN(n6766) );
  OAI21_X1 U5130 ( .B1(n7749), .B2(n7748), .A(n7768), .ZN(n7765) );
  INV_X1 U5131 ( .A(n7948), .ZN(n7768) );
  AND3_X1 U5132 ( .A1(n6143), .A2(n6142), .A3(n6141), .ZN(n8386) );
  AND4_X1 U5133 ( .A1(n6037), .A2(n6036), .A3(n6035), .A4(n6034), .ZN(n7271)
         );
  OAI21_X1 U5134 ( .B1(n6832), .B2(n4474), .A(n4472), .ZN(n4477) );
  INV_X1 U5135 ( .A(n4473), .ZN(n4472) );
  OAI21_X1 U5136 ( .B1(n6948), .B2(n4474), .A(n4359), .ZN(n4473) );
  NAND2_X1 U5137 ( .A1(n7158), .A2(n5935), .ZN(n7314) );
  XNOR2_X1 U5138 ( .A(n4477), .B(n4476), .ZN(n7165) );
  NAND2_X1 U5139 ( .A1(n7314), .A2(n7315), .ZN(n7313) );
  NAND2_X1 U5140 ( .A1(n7413), .A2(n7414), .ZN(n7412) );
  NAND2_X1 U5141 ( .A1(n8468), .A2(n5939), .ZN(n8479) );
  NAND2_X1 U5142 ( .A1(n8503), .A2(n5941), .ZN(n8517) );
  NAND2_X1 U5143 ( .A1(n8517), .A2(n8518), .ZN(n8516) );
  AOI21_X1 U5144 ( .B1(n4620), .B2(n8702), .A(n4619), .ZN(n4618) );
  INV_X1 U5145 ( .A(n7917), .ZN(n4619) );
  AND2_X1 U5146 ( .A1(n6152), .A2(n6151), .ZN(n8706) );
  INV_X1 U5147 ( .A(n6118), .ZN(n6117) );
  NAND2_X1 U5148 ( .A1(n6085), .A2(n6084), .ZN(n8248) );
  NAND2_X1 U5149 ( .A1(n4305), .A2(n6083), .ZN(n7563) );
  NAND2_X1 U5150 ( .A1(n6058), .A2(n6057), .ZN(n7526) );
  NAND2_X1 U5151 ( .A1(n7073), .A2(n7864), .ZN(n4617) );
  AND4_X1 U5152 ( .A1(n6025), .A2(n6024), .A3(n6023), .A4(n6022), .ZN(n7072)
         );
  OAI211_X1 U5153 ( .C1(n5991), .C2(n6379), .A(n4308), .B(n4823), .ZN(n6991)
         );
  OR2_X1 U5154 ( .A1(n5990), .A2(n6380), .ZN(n4823) );
  AOI21_X1 U5155 ( .B1(n6927), .B2(n6261), .A(n6260), .ZN(n6984) );
  OAI21_X1 U5156 ( .B1(n4594), .B2(n7822), .A(n7824), .ZN(n4593) );
  AND2_X1 U5157 ( .A1(n7833), .A2(n7832), .ZN(n7772) );
  NAND2_X1 U5158 ( .A1(n7823), .A2(n7824), .ZN(n7828) );
  NAND2_X1 U5159 ( .A1(n4441), .A2(n6849), .ZN(n7826) );
  INV_X1 U5160 ( .A(n10007), .ZN(n4441) );
  NAND2_X1 U5161 ( .A1(n6460), .A2(n10007), .ZN(n7822) );
  AOI21_X1 U5162 ( .B1(n4590), .B2(n4588), .A(n4587), .ZN(n4586) );
  INV_X1 U5163 ( .A(n4592), .ZN(n4588) );
  INV_X1 U5164 ( .A(n7933), .ZN(n4587) );
  INV_X1 U5165 ( .A(n4590), .ZN(n4589) );
  AND2_X1 U5166 ( .A1(n7935), .A2(n7936), .ZN(n8625) );
  NAND2_X1 U5167 ( .A1(n4825), .A2(n4824), .ZN(n8637) );
  AOI21_X1 U5168 ( .B1(n4826), .B2(n4828), .A(n4335), .ZN(n4824) );
  NOR2_X1 U5169 ( .A1(n7925), .A2(n7808), .ZN(n4592) );
  AND2_X1 U5170 ( .A1(n7932), .A2(n7933), .ZN(n8638) );
  NAND2_X1 U5171 ( .A1(n8663), .A2(n8664), .ZN(n8662) );
  OR2_X1 U5172 ( .A1(n7925), .A2(n7809), .ZN(n8651) );
  AND2_X1 U5173 ( .A1(n6288), .A2(n8673), .ZN(n8690) );
  NAND2_X1 U5174 ( .A1(n8708), .A2(n8707), .ZN(n8709) );
  NAND2_X1 U5175 ( .A1(n8747), .A2(n4356), .ZN(n8728) );
  AND2_X1 U5176 ( .A1(n6438), .A2(n7963), .ZN(n8739) );
  NAND2_X1 U5177 ( .A1(n6300), .A2(n6340), .ZN(n8752) );
  AND2_X1 U5178 ( .A1(n7899), .A2(n6103), .ZN(n7896) );
  INV_X1 U5179 ( .A(n5776), .ZN(n5775) );
  NAND2_X1 U5180 ( .A1(n5782), .A2(n5764), .ZN(n6249) );
  OAI21_X1 U5181 ( .B1(n5157), .B2(n4500), .A(n5198), .ZN(n4499) );
  INV_X1 U5182 ( .A(n5364), .ZN(n4504) );
  NAND2_X1 U5183 ( .A1(n5019), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5393) );
  INV_X1 U5184 ( .A(n7401), .ZN(n5292) );
  OR2_X1 U5185 ( .A1(n5211), .A2(n5210), .ZN(n5236) );
  NOR2_X1 U5186 ( .A1(n9099), .A2(n9100), .ZN(n4807) );
  AND2_X1 U5187 ( .A1(n5540), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5560) );
  AND2_X1 U5188 ( .A1(n5560), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5584) );
  XNOR2_X1 U5189 ( .A(n5268), .B(n5269), .ZN(n9120) );
  AND2_X1 U5190 ( .A1(n9134), .A2(n9135), .ZN(n5472) );
  INV_X1 U5191 ( .A(n5574), .ZN(n4783) );
  AND2_X1 U5192 ( .A1(n5592), .A2(n5591), .ZN(n9307) );
  AND4_X1 U5193 ( .A1(n5174), .A2(n5173), .A3(n5172), .A4(n5171), .ZN(n7013)
         );
  OR2_X1 U5194 ( .A1(n9726), .A2(n9725), .ZN(n4376) );
  NOR2_X1 U5195 ( .A1(n9812), .A2(n4383), .ZN(n7217) );
  AND2_X1 U5196 ( .A1(n7215), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4383) );
  NAND2_X1 U5197 ( .A1(n7217), .A2(n7216), .ZN(n7697) );
  AND2_X1 U5198 ( .A1(n9380), .A2(n4296), .ZN(n9320) );
  NAND2_X1 U5199 ( .A1(n9380), .A2(n4462), .ZN(n9335) );
  NAND2_X1 U5200 ( .A1(n9556), .A2(n9162), .ZN(n9328) );
  NAND2_X1 U5201 ( .A1(n4676), .A2(n4294), .ZN(n4674) );
  NAND2_X1 U5202 ( .A1(n4304), .A2(n9314), .ZN(n4675) );
  NAND2_X1 U5203 ( .A1(n4546), .A2(n9264), .ZN(n4545) );
  INV_X1 U5204 ( .A(n4547), .ZN(n4546) );
  AOI21_X1 U5205 ( .B1(n4549), .B2(n9263), .A(n4548), .ZN(n4547) );
  INV_X1 U5206 ( .A(n9409), .ZN(n4548) );
  NAND2_X1 U5207 ( .A1(n9438), .A2(n4309), .ZN(n4540) );
  OAI21_X1 U5208 ( .B1(n9438), .B2(n4544), .A(n4541), .ZN(n9389) );
  AOI21_X1 U5209 ( .B1(n4545), .B2(n4543), .A(n4542), .ZN(n4541) );
  INV_X1 U5210 ( .A(n4545), .ZN(n4544) );
  INV_X1 U5211 ( .A(n4309), .ZN(n4543) );
  AND2_X1 U5212 ( .A1(n8185), .A2(n9264), .ZN(n9409) );
  INV_X1 U5213 ( .A(n4875), .ZN(n4652) );
  AND2_X1 U5214 ( .A1(n8099), .A2(n8173), .ZN(n9471) );
  AND2_X1 U5215 ( .A1(n8046), .A2(n8172), .ZN(n9486) );
  NAND2_X1 U5216 ( .A1(n9506), .A2(n4539), .ZN(n9484) );
  NOR2_X1 U5217 ( .A1(n4323), .A2(n4665), .ZN(n4664) );
  AND2_X1 U5218 ( .A1(n8110), .A2(n9175), .ZN(n4665) );
  NAND2_X1 U5219 ( .A1(n4659), .A2(n4660), .ZN(n4663) );
  OAI21_X1 U5220 ( .B1(n9915), .B2(n4644), .A(n4639), .ZN(n4645) );
  NOR2_X1 U5221 ( .A1(n4640), .A2(n8064), .ZN(n4639) );
  NOR2_X1 U5222 ( .A1(n9914), .A2(n4644), .ZN(n4640) );
  AND2_X1 U5223 ( .A1(n7581), .A2(n8157), .ZN(n8064) );
  NAND2_X1 U5224 ( .A1(n6806), .A2(n6776), .ZN(n6777) );
  XNOR2_X1 U5225 ( .A(n4389), .B(n7751), .ZN(n7743) );
  NAND2_X1 U5226 ( .A1(n4777), .A2(n4778), .ZN(n4460) );
  XNOR2_X1 U5227 ( .A(n5625), .B(n5624), .ZN(n7619) );
  NAND2_X1 U5228 ( .A1(n4700), .A2(n4701), .ZN(n5496) );
  NAND2_X1 U5229 ( .A1(n5432), .A2(n4702), .ZN(n4700) );
  XNOR2_X1 U5230 ( .A(n5457), .B(n5456), .ZN(n7252) );
  NAND2_X1 U5231 ( .A1(n5452), .A2(n5476), .ZN(n5457) );
  XNOR2_X1 U5232 ( .A(n5318), .B(n5319), .ZN(n6527) );
  NAND2_X1 U5233 ( .A1(n4945), .A2(n4944), .ZN(n5318) );
  NAND2_X1 U5234 ( .A1(n4524), .A2(n4915), .ZN(n5164) );
  NAND2_X1 U5235 ( .A1(n5187), .A2(n4913), .ZN(n4524) );
  AND2_X1 U5236 ( .A1(n6169), .A2(n6168), .ZN(n8316) );
  NAND2_X1 U5237 ( .A1(n8428), .A2(n8256), .ZN(n8356) );
  NAND2_X1 U5238 ( .A1(n6125), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U5239 ( .A1(n5993), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5964) );
  AND4_X1 U5240 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n8432)
         );
  INV_X1 U5241 ( .A(n7802), .ZN(n4599) );
  INV_X1 U5242 ( .A(n7973), .ZN(n7971) );
  INV_X1 U5243 ( .A(n7983), .ZN(n4459) );
  NAND2_X1 U5244 ( .A1(n4861), .A2(n4858), .ZN(n6608) );
  OAI21_X1 U5245 ( .B1(n4431), .B2(n9996), .A(n4860), .ZN(n4859) );
  NAND2_X1 U5246 ( .A1(n6602), .A2(n4396), .ZN(n6573) );
  OR2_X1 U5247 ( .A1(n5926), .A2(n5927), .ZN(n4396) );
  AND2_X1 U5248 ( .A1(n5823), .A2(n5822), .ZN(n6703) );
  NAND2_X1 U5249 ( .A1(n6947), .A2(n4726), .ZN(n4725) );
  AND2_X1 U5250 ( .A1(n4724), .A2(n4727), .ZN(n4723) );
  OR2_X1 U5251 ( .A1(n7344), .A2(n5887), .ZN(n4480) );
  INV_X1 U5252 ( .A(n4478), .ZN(n7409) );
  INV_X1 U5253 ( .A(n4864), .ZN(n5889) );
  INV_X1 U5254 ( .A(n5863), .ZN(n4741) );
  NOR2_X1 U5255 ( .A1(n5893), .A2(n8496), .ZN(n8515) );
  INV_X1 U5256 ( .A(n4483), .ZN(n5892) );
  NOR2_X1 U5257 ( .A1(n4747), .A2(n4746), .ZN(n4745) );
  INV_X1 U5258 ( .A(n8563), .ZN(n4746) );
  XNOR2_X1 U5259 ( .A(n4430), .B(n4429), .ZN(n4428) );
  INV_X1 U5260 ( .A(n5947), .ZN(n4429) );
  OR2_X1 U5261 ( .A1(n8562), .A2(n5869), .ZN(n4430) );
  NAND2_X1 U5262 ( .A1(n5905), .A2(n8325), .ZN(n4426) );
  AOI21_X1 U5263 ( .B1(n5904), .B2(n10000), .A(n5903), .ZN(n5905) );
  NAND2_X1 U5264 ( .A1(n6160), .A2(n6159), .ZN(n8788) );
  NAND2_X1 U5265 ( .A1(n6134), .A2(n6133), .ZN(n8799) );
  NAND2_X1 U5266 ( .A1(n6105), .A2(n6104), .ZN(n8809) );
  OAI211_X1 U5267 ( .C1(n6308), .C2(n6623), .A(n6000), .B(n5999), .ZN(n6891)
         );
  NAND2_X1 U5268 ( .A1(n7757), .A2(n7756), .ZN(n8814) );
  NAND2_X1 U5269 ( .A1(n6239), .A2(n7755), .ZN(n6241) );
  NOR2_X1 U5270 ( .A1(n4878), .A2(n8579), .ZN(n6354) );
  NAND2_X1 U5271 ( .A1(n4613), .A2(n7943), .ZN(n8589) );
  NAND2_X1 U5272 ( .A1(n8602), .A2(n8601), .ZN(n4613) );
  NAND2_X2 U5273 ( .A1(n6214), .A2(n6213), .ZN(n8829) );
  XNOR2_X1 U5274 ( .A(n5774), .B(n5773), .ZN(n7657) );
  NAND2_X1 U5275 ( .A1(n5778), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U5276 ( .A1(n5829), .A2(n5830), .ZN(n4718) );
  NAND2_X1 U5277 ( .A1(n9047), .A2(n4510), .ZN(n4509) );
  AND2_X1 U5278 ( .A1(n9112), .A2(n9113), .ZN(n4510) );
  NAND2_X1 U5279 ( .A1(n5256), .A2(n5255), .ZN(n5265) );
  NAND2_X1 U5280 ( .A1(n5391), .A2(n5390), .ZN(n9274) );
  NOR2_X1 U5281 ( .A1(n8233), .A2(n7254), .ZN(n4576) );
  OAI21_X1 U5282 ( .B1(n4556), .B2(n4555), .A(n4554), .ZN(n8231) );
  OAI22_X1 U5283 ( .A1(n8234), .A2(n8232), .B1(n8236), .B2(n8235), .ZN(n4575)
         );
  INV_X1 U5284 ( .A(n8111), .ZN(n9174) );
  INV_X1 U5285 ( .A(n7588), .ZN(n9176) );
  INV_X1 U5286 ( .A(n7234), .ZN(n9760) );
  NOR2_X1 U5287 ( .A1(n9824), .A2(n9825), .ZN(n9823) );
  XNOR2_X1 U5288 ( .A(n4380), .B(n4379), .ZN(n7713) );
  NAND2_X1 U5289 ( .A1(n9893), .A2(n7711), .ZN(n4380) );
  NAND2_X1 U5290 ( .A1(n4553), .A2(n9910), .ZN(n4552) );
  XNOR2_X1 U5291 ( .A(n9270), .B(n8204), .ZN(n4553) );
  AOI211_X1 U5292 ( .C1(n9556), .C2(n9358), .A(n9527), .B(n4316), .ZN(n9558)
         );
  NAND2_X1 U5293 ( .A1(n5559), .A2(n5558), .ZN(n9574) );
  NAND2_X1 U5294 ( .A1(n5128), .A2(n4470), .ZN(n4469) );
  OAI22_X1 U5295 ( .A1(n6376), .A2(n4471), .B1(n4891), .B2(n6362), .ZN(n4470)
         );
  OR2_X1 U5296 ( .A1(n5127), .A2(n6378), .ZN(n5102) );
  OR2_X1 U5297 ( .A1(n6380), .A2(n5101), .ZN(n5131) );
  OR2_X1 U5298 ( .A1(n7840), .A2(n7839), .ZN(n7851) );
  OAI21_X1 U5299 ( .B1(n7846), .B2(n7848), .A(n7852), .ZN(n4436) );
  NAND2_X1 U5300 ( .A1(n4438), .A2(n4433), .ZN(n7874) );
  AOI21_X1 U5301 ( .B1(n4569), .B2(n4571), .A(n4572), .ZN(n4568) );
  NAND2_X1 U5302 ( .A1(n8152), .A2(n8151), .ZN(n4571) );
  NOR2_X1 U5303 ( .A1(n8159), .A2(n8160), .ZN(n4572) );
  AOI21_X1 U5304 ( .B1(n4456), .B2(n4455), .A(n4454), .ZN(n4453) );
  NAND2_X1 U5305 ( .A1(n6083), .A2(n7887), .ZN(n4454) );
  NAND2_X1 U5306 ( .A1(n7883), .A2(n7963), .ZN(n4455) );
  AOI21_X1 U5307 ( .B1(n7884), .B2(n7942), .A(n7888), .ZN(n4456) );
  AND2_X1 U5308 ( .A1(n7896), .A2(n7895), .ZN(n4451) );
  OAI21_X1 U5309 ( .B1(n8175), .B2(n8171), .A(n4351), .ZN(n4566) );
  OAI21_X1 U5310 ( .B1(n8175), .B2(n8174), .A(n4561), .ZN(n4560) );
  NOR2_X1 U5311 ( .A1(n4563), .A2(n4562), .ZN(n4561) );
  NAND2_X1 U5312 ( .A1(n8172), .A2(n8209), .ZN(n4562) );
  NAND2_X1 U5313 ( .A1(n4564), .A2(n4558), .ZN(n4557) );
  AND2_X1 U5314 ( .A1(n4560), .A2(n4559), .ZN(n4558) );
  NAND2_X1 U5315 ( .A1(n4565), .A2(n8223), .ZN(n4564) );
  INV_X1 U5316 ( .A(n8180), .ZN(n4559) );
  OAI211_X1 U5317 ( .C1(n4448), .C2(n7938), .A(n4315), .B(n4444), .ZN(n4445)
         );
  INV_X1 U5318 ( .A(n7931), .ZN(n4448) );
  INV_X1 U5319 ( .A(n4449), .ZN(n4444) );
  NOR2_X1 U5320 ( .A1(n4449), .A2(n4447), .ZN(n4446) );
  AND2_X1 U5321 ( .A1(n8191), .A2(n8190), .ZN(n8194) );
  AOI21_X1 U5322 ( .B1(n7956), .B2(n7955), .A(n7947), .ZN(n7952) );
  INV_X1 U5323 ( .A(n6265), .ZN(n4832) );
  AND2_X1 U5324 ( .A1(n6268), .A2(n6263), .ZN(n4829) );
  OR2_X1 U5325 ( .A1(n9334), .A2(n7996), .ZN(n8201) );
  OR2_X1 U5326 ( .A1(n9529), .A2(n9103), .ZN(n8164) );
  AND2_X1 U5327 ( .A1(n4530), .A2(n8151), .ZN(n7456) );
  INV_X1 U5328 ( .A(n5227), .ZN(n4688) );
  XNOR2_X1 U5329 ( .A(n6714), .B(n6891), .ZN(n6731) );
  OAI21_X1 U5330 ( .B1(n6910), .B2(n4410), .A(n6999), .ZN(n4409) );
  INV_X1 U5331 ( .A(n4409), .ZN(n4408) );
  OAI21_X1 U5332 ( .B1(n6692), .B2(n4854), .A(n4852), .ZN(n6948) );
  INV_X1 U5333 ( .A(n6950), .ZN(n4474) );
  NOR2_X1 U5334 ( .A1(n7416), .A2(n4738), .ZN(n4737) );
  NAND2_X1 U5335 ( .A1(n4736), .A2(n4735), .ZN(n4734) );
  INV_X1 U5336 ( .A(n7416), .ZN(n4735) );
  INV_X1 U5337 ( .A(n5856), .ZN(n4736) );
  NAND2_X1 U5338 ( .A1(n6885), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4423) );
  INV_X1 U5339 ( .A(n8524), .ZN(n4424) );
  NAND2_X1 U5340 ( .A1(n7790), .A2(n7747), .ZN(n7947) );
  NOR2_X1 U5341 ( .A1(n6272), .A2(n4821), .ZN(n4820) );
  INV_X1 U5342 ( .A(n6270), .ZN(n4821) );
  INV_X1 U5343 ( .A(n6291), .ZN(n4828) );
  INV_X1 U5344 ( .A(n5760), .ZN(n5758) );
  INV_X1 U5345 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4622) );
  INV_X1 U5346 ( .A(n5163), .ZN(n4500) );
  OR2_X1 U5347 ( .A1(n5494), .A2(n5493), .ZN(n5495) );
  AND2_X1 U5348 ( .A1(n5018), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U5349 ( .A1(n5424), .A2(n5425), .ZN(n4810) );
  NAND2_X1 U5350 ( .A1(n4578), .A2(n4324), .ZN(n8208) );
  AND2_X1 U5351 ( .A1(n7685), .A2(n9860), .ZN(n7686) );
  NOR2_X1 U5352 ( .A1(n9334), .A2(n4463), .ZN(n4462) );
  INV_X1 U5353 ( .A(n4464), .ZN(n4463) );
  OR2_X1 U5354 ( .A1(n9321), .A2(n7988), .ZN(n8206) );
  NAND2_X1 U5355 ( .A1(n8173), .A2(n8172), .ZN(n4536) );
  NAND2_X1 U5356 ( .A1(n4537), .A2(n8173), .ZN(n4535) );
  AND2_X1 U5357 ( .A1(n4661), .A2(n4657), .ZN(n4656) );
  NAND2_X1 U5358 ( .A1(n8065), .A2(n4664), .ZN(n4657) );
  AND2_X1 U5359 ( .A1(n9277), .A2(n4322), .ZN(n4661) );
  NAND2_X1 U5360 ( .A1(n4529), .A2(n8002), .ZN(n4528) );
  AND2_X1 U5361 ( .A1(n7456), .A2(n8120), .ZN(n8019) );
  NOR2_X1 U5362 ( .A1(n9403), .A2(n9574), .ZN(n7724) );
  NAND2_X1 U5363 ( .A1(n9526), .A2(n9674), .ZN(n9509) );
  INV_X1 U5364 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U5365 ( .A1(n6236), .A2(n6235), .ZN(n7660) );
  AOI21_X1 U5366 ( .B1(n4694), .B2(n4697), .A(n4693), .ZN(n4692) );
  INV_X1 U5367 ( .A(n5430), .ZN(n4703) );
  INV_X1 U5368 ( .A(n4497), .ZN(n4496) );
  OAI21_X1 U5369 ( .B1(n4995), .B2(n9688), .A(n5039), .ZN(n4497) );
  OAI21_X1 U5370 ( .B1(n5366), .B2(n4704), .A(n4707), .ZN(n5046) );
  NAND2_X1 U5371 ( .A1(n4705), .A2(n4714), .ZN(n4704) );
  INV_X1 U5372 ( .A(n4708), .ZN(n4707) );
  AND2_X1 U5373 ( .A1(n4973), .A2(n4972), .ZN(n5045) );
  AND2_X1 U5374 ( .A1(n5252), .A2(n4978), .ZN(n4979) );
  INV_X1 U5375 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U5376 ( .A1(n4937), .A2(n4936), .ZN(n4944) );
  INV_X1 U5377 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U5378 ( .A1(n4395), .A2(n4681), .ZN(n5294) );
  NOR2_X1 U5379 ( .A1(n4683), .A2(n4682), .ZN(n4681) );
  INV_X1 U5380 ( .A(n4934), .ZN(n4682) );
  NAND2_X1 U5381 ( .A1(n5251), .A2(n4302), .ZN(n4395) );
  NAND2_X1 U5382 ( .A1(n4687), .A2(n4685), .ZN(n5251) );
  NAND2_X1 U5383 ( .A1(n4684), .A2(n4390), .ZN(n4687) );
  AND2_X1 U5384 ( .A1(n4686), .A2(n4927), .ZN(n4685) );
  AND2_X1 U5385 ( .A1(n4689), .A2(n4688), .ZN(n4684) );
  OAI21_X1 U5386 ( .B1(n5187), .B2(n4526), .A(n4522), .ZN(n4390) );
  INV_X1 U5387 ( .A(n5188), .ZN(n4913) );
  NAND2_X1 U5388 ( .A1(n4904), .A2(n4903), .ZN(n4905) );
  OAI21_X1 U5389 ( .B1(n4892), .B2(n4891), .A(n4890), .ZN(n4896) );
  NAND2_X1 U5390 ( .A1(n5776), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U5391 ( .A1(n4754), .A2(n4353), .ZN(n4752) );
  AND2_X1 U5392 ( .A1(n6516), .A2(n6453), .ZN(n6455) );
  AND2_X1 U5393 ( .A1(n8417), .A2(n8290), .ZN(n8344) );
  INV_X1 U5394 ( .A(n8629), .ZN(n8349) );
  NOR2_X1 U5395 ( .A1(n8365), .A2(n4767), .ZN(n4766) );
  INV_X1 U5396 ( .A(n4769), .ZN(n4767) );
  NAND2_X1 U5397 ( .A1(n8354), .A2(n8740), .ZN(n4769) );
  NAND2_X1 U5398 ( .A1(n8356), .A2(n4770), .ZN(n4768) );
  OR2_X1 U5399 ( .A1(n8354), .A2(n8740), .ZN(n4770) );
  NAND2_X1 U5400 ( .A1(n8313), .A2(n8397), .ZN(n8373) );
  CLKBUF_X1 U5401 ( .A(n8280), .Z(n8281) );
  NAND2_X1 U5402 ( .A1(n4771), .A2(n7435), .ZN(n7533) );
  NAND2_X1 U5403 ( .A1(n6455), .A2(n6454), .ZN(n6517) );
  NAND2_X1 U5404 ( .A1(n4759), .A2(n4755), .ZN(n4754) );
  INV_X1 U5405 ( .A(n4757), .ZN(n4755) );
  AOI21_X1 U5406 ( .B1(n8344), .B2(n8345), .A(n4758), .ZN(n4757) );
  INV_X1 U5407 ( .A(n8417), .ZN(n4758) );
  OAI211_X1 U5408 ( .C1(n7967), .C2(n4680), .A(n7970), .B(n4678), .ZN(n7973)
         );
  NAND2_X1 U5409 ( .A1(n7968), .A2(n7963), .ZN(n4680) );
  OR4_X1 U5410 ( .A1(n7948), .A2(n8590), .A3(n8603), .A4(n7789), .ZN(n7791) );
  AND2_X1 U5411 ( .A1(n7764), .A2(n7763), .ZN(n7795) );
  AND2_X1 U5412 ( .A1(n7764), .A2(n6247), .ZN(n8441) );
  INV_X1 U5413 ( .A(n5876), .ZN(n4856) );
  NAND2_X1 U5414 ( .A1(n4731), .A2(n4730), .ZN(n6592) );
  OAI21_X1 U5415 ( .B1(n5844), .B2(n6384), .A(n4715), .ZN(n6576) );
  OAI211_X1 U5416 ( .C1(n6692), .C2(n4851), .A(n4849), .B(n4848), .ZN(n6833)
         );
  INV_X1 U5417 ( .A(n4855), .ZN(n4851) );
  AOI22_X1 U5418 ( .A1(n4852), .A2(n4854), .B1(n4855), .B2(n4850), .ZN(n4849)
         );
  AOI21_X1 U5419 ( .B1(n6832), .B2(n6948), .A(n4474), .ZN(n6953) );
  AND2_X1 U5420 ( .A1(n4728), .A2(n4729), .ZN(n7323) );
  INV_X1 U5421 ( .A(n5854), .ZN(n4728) );
  NOR2_X1 U5422 ( .A1(n7323), .A2(n7322), .ZN(n7321) );
  NAND2_X1 U5423 ( .A1(n7351), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7350) );
  NAND2_X1 U5424 ( .A1(n5886), .A2(n6445), .ZN(n5885) );
  AND2_X1 U5425 ( .A1(n7350), .A2(n5856), .ZN(n7417) );
  NAND2_X1 U5426 ( .A1(n7412), .A2(n5938), .ZN(n8469) );
  NAND2_X1 U5427 ( .A1(n8469), .A2(n8470), .ZN(n8468) );
  NAND2_X1 U5428 ( .A1(n4478), .A2(n4368), .ZN(n4864) );
  XNOR2_X1 U5429 ( .A(n4483), .B(n6711), .ZN(n8497) );
  NAND2_X1 U5430 ( .A1(n8504), .A2(n8505), .ZN(n8503) );
  OR2_X1 U5431 ( .A1(n8495), .A2(n8917), .ZN(n4742) );
  NAND2_X1 U5432 ( .A1(n4485), .A2(n4484), .ZN(n4483) );
  NAND2_X1 U5433 ( .A1(n6654), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4484) );
  NAND2_X1 U5434 ( .A1(n4773), .A2(n4772), .ZN(n5865) );
  INV_X1 U5435 ( .A(n5792), .ZN(n4773) );
  NAND2_X1 U5436 ( .A1(n4482), .A2(n4370), .ZN(n4481) );
  NAND2_X1 U5437 ( .A1(n4481), .A2(n6965), .ZN(n5895) );
  NAND2_X1 U5438 ( .A1(n8516), .A2(n5942), .ZN(n8545) );
  NAND2_X1 U5439 ( .A1(n4402), .A2(n8552), .ZN(n8557) );
  INV_X1 U5440 ( .A(n8551), .ZN(n4402) );
  NOR2_X1 U5441 ( .A1(n5945), .A2(n5944), .ZN(n8551) );
  NOR2_X1 U5442 ( .A1(n8555), .A2(n5898), .ZN(n5899) );
  NAND2_X1 U5443 ( .A1(n4612), .A2(n4611), .ZN(n7749) );
  AOI21_X1 U5444 ( .B1(n4614), .B2(n4616), .A(n4334), .ZN(n4611) );
  NAND2_X1 U5445 ( .A1(n8602), .A2(n4614), .ZN(n4612) );
  AOI21_X1 U5446 ( .B1(n4846), .B2(n6298), .A(n4341), .ZN(n4845) );
  NAND2_X1 U5447 ( .A1(n6191), .A2(n6190), .ZN(n6205) );
  INV_X1 U5448 ( .A(n6192), .ZN(n6191) );
  OR2_X1 U5449 ( .A1(n6181), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6192) );
  OR2_X1 U5450 ( .A1(n6172), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U5451 ( .A1(n6096), .A2(n6095), .ZN(n6106) );
  NOR2_X1 U5452 ( .A1(n6068), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6077) );
  OR2_X1 U5453 ( .A1(n6050), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6059) );
  OR2_X1 U5454 ( .A1(n6059), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6068) );
  AND2_X1 U5455 ( .A1(n4887), .A2(n6274), .ZN(n4841) );
  NAND2_X1 U5456 ( .A1(n4842), .A2(n6274), .ZN(n7389) );
  AOI21_X1 U5457 ( .B1(n4815), .B2(n4817), .A(n4320), .ZN(n4813) );
  NAND2_X1 U5458 ( .A1(n4814), .A2(n4818), .ZN(n7289) );
  NAND2_X1 U5459 ( .A1(n6271), .A2(n4820), .ZN(n4814) );
  AOI21_X1 U5460 ( .B1(n4607), .B2(n4604), .A(n4606), .ZN(n4603) );
  AND2_X1 U5461 ( .A1(n7074), .A2(n7865), .ZN(n7778) );
  INV_X1 U5462 ( .A(n4608), .ZN(n4607) );
  NAND2_X1 U5463 ( .A1(n4833), .A2(n6265), .ZN(n7044) );
  NAND2_X1 U5464 ( .A1(n6887), .A2(n6263), .ZN(n4833) );
  AND4_X2 U5465 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n6986)
         );
  NAND2_X1 U5466 ( .A1(n6923), .A2(n7832), .ZN(n6989) );
  NAND2_X1 U5467 ( .A1(n7828), .A2(n6848), .ZN(n6929) );
  NOR2_X1 U5468 ( .A1(n8605), .A2(n6298), .ZN(n8591) );
  OR2_X1 U5469 ( .A1(n8829), .A2(n8423), .ZN(n7943) );
  AOI21_X1 U5470 ( .B1(n4586), .B2(n4589), .A(n4585), .ZN(n4584) );
  AND2_X1 U5471 ( .A1(n7939), .A2(n7940), .ZN(n8615) );
  OR2_X1 U5472 ( .A1(n8624), .A2(n8625), .ZN(n8626) );
  NAND2_X1 U5473 ( .A1(n4836), .A2(n4834), .ZN(n8689) );
  AND2_X1 U5474 ( .A1(n4835), .A2(n6287), .ZN(n4834) );
  NAND2_X1 U5475 ( .A1(n8736), .A2(n6285), .ZN(n8719) );
  NAND2_X1 U5476 ( .A1(n8728), .A2(n4625), .ZN(n8717) );
  NOR2_X1 U5477 ( .A1(n7770), .A2(n4626), .ZN(n4625) );
  INV_X1 U5478 ( .A(n7814), .ZN(n4626) );
  NAND2_X1 U5479 ( .A1(n6284), .A2(n8731), .ZN(n8736) );
  NAND2_X1 U5480 ( .A1(n4840), .A2(n6281), .ZN(n7627) );
  NAND2_X1 U5481 ( .A1(n4840), .A2(n4329), .ZN(n8750) );
  AOI21_X1 U5482 ( .B1(n7571), .B2(n7892), .A(n6092), .ZN(n7626) );
  INV_X1 U5483 ( .A(n6991), .ZN(n10020) );
  AND2_X1 U5484 ( .A1(n5772), .A2(n5773), .ZN(n4627) );
  NAND2_X1 U5485 ( .A1(n5760), .A2(n4420), .ZN(n5778) );
  AND2_X1 U5486 ( .A1(n4457), .A2(n5772), .ZN(n4420) );
  INV_X1 U5487 ( .A(n6249), .ZN(n6248) );
  INV_X1 U5488 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5787) );
  XNOR2_X1 U5489 ( .A(n5133), .B(n4287), .ZN(n5138) );
  AND2_X1 U5490 ( .A1(n5644), .A2(n5643), .ZN(n5703) );
  INV_X1 U5491 ( .A(n6645), .ZN(n5157) );
  XNOR2_X1 U5492 ( .A(n5159), .B(n5160), .ZN(n6645) );
  OR2_X1 U5493 ( .A1(n5236), .A2(n5235), .ZN(n5257) );
  OR2_X1 U5494 ( .A1(n6876), .A2(n4779), .ZN(n4300) );
  AOI21_X1 U5495 ( .B1(n4802), .B2(n4805), .A(n4797), .ZN(n4796) );
  NAND2_X1 U5496 ( .A1(n9059), .A2(n4798), .ZN(n4797) );
  NAND2_X1 U5497 ( .A1(n4791), .A2(n4795), .ZN(n4788) );
  NAND2_X1 U5498 ( .A1(n7401), .A2(n4791), .ZN(n4789) );
  NOR2_X1 U5499 ( .A1(n5508), .A2(n5506), .ZN(n5540) );
  NAND2_X1 U5500 ( .A1(n5522), .A2(n5521), .ZN(n5524) );
  AND2_X1 U5501 ( .A1(n5291), .A2(n4793), .ZN(n4792) );
  INV_X1 U5502 ( .A(n4502), .ZN(n4501) );
  NAND2_X1 U5503 ( .A1(n8222), .A2(n9350), .ZN(n4554) );
  OR2_X1 U5504 ( .A1(n8221), .A2(n9350), .ZN(n4555) );
  AND4_X1 U5505 ( .A1(n5638), .A2(n5637), .A3(n5636), .A4(n5635), .ZN(n9162)
         );
  AND2_X1 U5506 ( .A1(n5516), .A2(n5515), .ZN(n9299) );
  AND4_X1 U5507 ( .A1(n5356), .A2(n5355), .A3(n5354), .A4(n5353), .ZN(n7580)
         );
  AND4_X1 U5508 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n7588)
         );
  AND4_X1 U5509 ( .A1(n5261), .A2(n5260), .A3(n5259), .A4(n5258), .ZN(n7234)
         );
  AND4_X1 U5510 ( .A1(n5241), .A2(n5240), .A3(n5239), .A4(n5238), .ZN(n7238)
         );
  AND4_X1 U5511 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n7093)
         );
  NAND2_X1 U5512 ( .A1(n6492), .A2(n6493), .ZN(n7209) );
  AND2_X1 U5513 ( .A1(n7209), .A2(n4388), .ZN(n9213) );
  NAND2_X1 U5514 ( .A1(n7210), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4388) );
  NOR2_X1 U5515 ( .A1(n9213), .A2(n9212), .ZN(n9211) );
  AND2_X1 U5516 ( .A1(n4376), .A2(n4375), .ZN(n9245) );
  NAND2_X1 U5517 ( .A1(n9729), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4375) );
  NAND2_X1 U5518 ( .A1(n9245), .A2(n9246), .ZN(n9244) );
  NAND2_X1 U5519 ( .A1(n9244), .A2(n4374), .ZN(n9699) );
  OR2_X1 U5520 ( .A1(n9248), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4374) );
  NOR2_X1 U5521 ( .A1(n9823), .A2(n7701), .ZN(n9841) );
  NOR2_X1 U5522 ( .A1(n7706), .A2(n7707), .ZN(n9850) );
  AND2_X1 U5523 ( .A1(n7705), .A2(n9860), .ZN(n7707) );
  NOR2_X1 U5524 ( .A1(n4673), .A2(n4668), .ZN(n4667) );
  INV_X1 U5525 ( .A(n9310), .ZN(n4668) );
  NAND2_X1 U5526 ( .A1(n4291), .A2(n9316), .ZN(n4673) );
  NOR2_X1 U5527 ( .A1(n9332), .A2(n4304), .ZN(n4672) );
  NOR2_X1 U5528 ( .A1(n9334), .A2(n9317), .ZN(n4671) );
  NAND2_X1 U5529 ( .A1(n9380), .A2(n9363), .ZN(n9358) );
  AND2_X1 U5530 ( .A1(n8193), .A2(n9265), .ZN(n9379) );
  AND2_X1 U5531 ( .A1(n7723), .A2(n9655), .ZN(n9423) );
  NAND2_X1 U5532 ( .A1(n9423), .A2(n9407), .ZN(n9403) );
  OR2_X1 U5533 ( .A1(n5441), .A2(n5440), .ZN(n5460) );
  OR2_X1 U5534 ( .A1(n5460), .A2(n9138), .ZN(n5508) );
  NAND2_X1 U5535 ( .A1(n4531), .A2(n4535), .ZN(n9451) );
  OR2_X1 U5536 ( .A1(n9506), .A2(n4536), .ZN(n4531) );
  OR2_X1 U5537 ( .A1(n9509), .A2(n9493), .ZN(n9491) );
  OAI21_X1 U5538 ( .B1(n8081), .B2(n8080), .A(n8079), .ZN(n9521) );
  NAND2_X1 U5539 ( .A1(n9521), .A2(n9524), .ZN(n9520) );
  OR2_X1 U5540 ( .A1(n5393), .A2(n5020), .ZN(n5410) );
  NAND3_X1 U5541 ( .A1(n9276), .A2(n4292), .A3(n7480), .ZN(n9528) );
  NOR2_X1 U5542 ( .A1(n9528), .A2(n9529), .ZN(n9526) );
  NAND2_X1 U5543 ( .A1(n7637), .A2(n8149), .ZN(n8081) );
  OR2_X1 U5544 ( .A1(n7599), .A2(n8067), .ZN(n7637) );
  NAND2_X1 U5545 ( .A1(n7480), .A2(n4465), .ZN(n7604) );
  NOR2_X1 U5546 ( .A1(n4641), .A2(n4637), .ZN(n4636) );
  AOI21_X1 U5547 ( .B1(n4339), .B2(n4641), .A(n4295), .ZN(n4635) );
  INV_X1 U5548 ( .A(n4642), .ZN(n4641) );
  NAND2_X1 U5549 ( .A1(n9906), .A2(n7458), .ZN(n7582) );
  AND2_X1 U5550 ( .A1(n9916), .A2(n7519), .ZN(n7480) );
  AND2_X1 U5551 ( .A1(n9919), .A2(n9956), .ZN(n9916) );
  AND3_X1 U5552 ( .A1(n7020), .A2(n4293), .A3(n4467), .ZN(n9919) );
  NOR2_X1 U5553 ( .A1(n9790), .A2(n5265), .ZN(n4467) );
  NAND2_X1 U5554 ( .A1(n7097), .A2(n4879), .ZN(n7099) );
  INV_X1 U5555 ( .A(n8125), .ZN(n7098) );
  NAND2_X1 U5556 ( .A1(n7099), .A2(n7098), .ZN(n7173) );
  NAND2_X1 U5557 ( .A1(n7011), .A2(n4632), .ZN(n7014) );
  NAND2_X1 U5558 ( .A1(n6976), .A2(n7110), .ZN(n4632) );
  NAND2_X1 U5559 ( .A1(n7014), .A2(n7017), .ZN(n7097) );
  NAND2_X1 U5560 ( .A1(n7020), .A2(n7034), .ZN(n7100) );
  NOR2_X1 U5561 ( .A1(n5180), .A2(n6900), .ZN(n5182) );
  NOR2_X1 U5562 ( .A1(n7300), .A2(n7012), .ZN(n7020) );
  NAND2_X1 U5563 ( .A1(n7299), .A2(n8052), .ZN(n7298) );
  NAND2_X1 U5564 ( .A1(n6788), .A2(n6787), .ZN(n6790) );
  NAND2_X1 U5565 ( .A1(n6790), .A2(n6789), .ZN(n6818) );
  NOR2_X1 U5566 ( .A1(n6814), .A2(n7038), .ZN(n6796) );
  NAND2_X1 U5567 ( .A1(n8051), .A2(n4628), .ZN(n6806) );
  NAND2_X1 U5568 ( .A1(n7721), .A2(n7720), .ZN(n8213) );
  NAND2_X1 U5569 ( .A1(n5583), .A2(n5582), .ZN(n9381) );
  NAND2_X1 U5570 ( .A1(n5539), .A2(n5538), .ZN(n9579) );
  OAI21_X1 U5571 ( .B1(n9438), .B2(n9263), .A(n4549), .ZN(n9408) );
  NAND2_X1 U5572 ( .A1(n5483), .A2(n5482), .ZN(n9444) );
  NAND2_X1 U5573 ( .A1(n5459), .A2(n5458), .ZN(n9460) );
  NAND2_X1 U5574 ( .A1(n5051), .A2(n5050), .ZN(n9512) );
  XNOR2_X1 U5575 ( .A(n7754), .B(n7753), .ZN(n9029) );
  XNOR2_X1 U5576 ( .A(n7660), .B(n7658), .ZN(n6237) );
  NAND2_X1 U5577 ( .A1(n6237), .A2(SI_29_), .ZN(n7662) );
  NAND2_X1 U5578 ( .A1(n9687), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5025) );
  INV_X1 U5579 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5028) );
  XNOR2_X1 U5580 ( .A(n6234), .B(n6233), .ZN(n7655) );
  INV_X1 U5581 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5000) );
  OAI21_X1 U5582 ( .B1(n5527), .B2(n5526), .A(n5525), .ZN(n5535) );
  NAND2_X1 U5583 ( .A1(n5049), .A2(n4995), .ZN(n4495) );
  NAND2_X1 U5584 ( .A1(n4706), .A2(n4962), .ZN(n5406) );
  NAND2_X1 U5585 ( .A1(n4713), .A2(n4711), .ZN(n4706) );
  OAI211_X1 U5586 ( .C1(n4523), .C2(n4521), .A(n4689), .B(n4520), .ZN(n5228)
         );
  INV_X1 U5587 ( .A(n5187), .ZN(n4523) );
  NAND2_X1 U5588 ( .A1(n4522), .A2(n4919), .ZN(n4521) );
  OR2_X1 U5589 ( .A1(n5189), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U5590 ( .A1(n4753), .A2(n4750), .ZN(n8304) );
  NOR2_X1 U5591 ( .A1(n4752), .A2(n4751), .ZN(n4750) );
  INV_X1 U5592 ( .A(n8305), .ZN(n4751) );
  NOR2_X1 U5593 ( .A1(n4749), .A2(n4752), .ZN(n8306) );
  INV_X1 U5594 ( .A(n4753), .ZN(n4749) );
  AND4_X1 U5595 ( .A1(n6102), .A2(n6101), .A3(n6100), .A4(n6099), .ZN(n9733)
         );
  CLKBUF_X1 U5596 ( .A(n8323), .Z(n8383) );
  NAND2_X1 U5597 ( .A1(n8406), .A2(n8262), .ZN(n8322) );
  NAND2_X1 U5598 ( .A1(n7533), .A2(n7439), .ZN(n7545) );
  AND3_X1 U5599 ( .A1(n6122), .A2(n6121), .A3(n6120), .ZN(n8755) );
  AND4_X1 U5600 ( .A1(n6019), .A2(n6018), .A3(n6017), .A4(n6016), .ZN(n6919)
         );
  NAND2_X1 U5601 ( .A1(n4768), .A2(n4769), .ZN(n8364) );
  NAND2_X1 U5602 ( .A1(n7274), .A2(n7273), .ZN(n7277) );
  AND2_X1 U5603 ( .A1(n4413), .A2(n7548), .ZN(n4412) );
  NAND2_X1 U5604 ( .A1(n6076), .A2(n6075), .ZN(n7556) );
  NOR2_X1 U5605 ( .A1(n4416), .A2(n8392), .ZN(n4415) );
  INV_X1 U5606 ( .A(n8274), .ZN(n4416) );
  NAND2_X1 U5607 ( .A1(n8336), .A2(n8274), .ZN(n8393) );
  INV_X1 U5608 ( .A(n8446), .ZN(n7531) );
  NAND2_X1 U5609 ( .A1(n6131), .A2(n6703), .ZN(n4417) );
  OR2_X1 U5610 ( .A1(n5991), .A2(n4419), .ZN(n4418) );
  NAND2_X1 U5611 ( .A1(n6764), .A2(n6761), .ZN(n4761) );
  INV_X1 U5612 ( .A(n4306), .ZN(n4762) );
  NAND2_X1 U5613 ( .A1(n4753), .A2(n4754), .ZN(n8421) );
  INV_X1 U5614 ( .A(n7984), .ZN(n4600) );
  INV_X1 U5615 ( .A(n7271), .ZN(n8448) );
  INV_X1 U5616 ( .A(n6919), .ZN(n8450) );
  INV_X1 U5617 ( .A(n6986), .ZN(n8454) );
  NAND4_X1 U5618 ( .A1(n5974), .A2(n5973), .A3(n5972), .A4(n5971), .ZN(n6849)
         );
  INV_X1 U5619 ( .A(n4399), .ZN(n4398) );
  NAND2_X1 U5620 ( .A1(n4862), .A2(n4861), .ZN(n6596) );
  INV_X1 U5621 ( .A(n4857), .ZN(n4862) );
  NOR2_X1 U5622 ( .A1(n6588), .A2(n4397), .ZN(n6604) );
  AND2_X1 U5623 ( .A1(n5924), .A2(n4431), .ZN(n4397) );
  NAND2_X1 U5624 ( .A1(n6573), .A2(n6572), .ZN(n6571) );
  NAND2_X1 U5625 ( .A1(n6692), .A2(n6693), .ZN(n6691) );
  NOR2_X1 U5626 ( .A1(n7165), .A2(n10099), .ZN(n7164) );
  NAND2_X1 U5627 ( .A1(n4869), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4868) );
  NAND2_X1 U5628 ( .A1(n4317), .A2(n4869), .ZN(n4475) );
  INV_X1 U5629 ( .A(n7312), .ZN(n4869) );
  NAND2_X1 U5630 ( .A1(n7313), .A2(n5936), .ZN(n7347) );
  XNOR2_X1 U5631 ( .A(n4864), .B(n6550), .ZN(n8458) );
  INV_X1 U5632 ( .A(n4742), .ZN(n8494) );
  OAI21_X1 U5633 ( .B1(n4481), .B2(n6965), .A(n5895), .ZN(n8533) );
  NOR2_X1 U5634 ( .A1(n8533), .A2(n8805), .ZN(n8532) );
  XNOR2_X1 U5635 ( .A(n7749), .B(n7959), .ZN(n8587) );
  NAND2_X1 U5636 ( .A1(n6094), .A2(n6093), .ZN(n8253) );
  NAND2_X1 U5637 ( .A1(n6065), .A2(n7880), .ZN(n7493) );
  NAND2_X1 U5638 ( .A1(n6067), .A2(n6066), .ZN(n10071) );
  NAND2_X1 U5639 ( .A1(n4617), .A2(n7866), .ZN(n7286) );
  NAND2_X1 U5640 ( .A1(n6271), .A2(n6270), .ZN(n7070) );
  OAI21_X1 U5641 ( .B1(n7828), .B2(n7822), .A(n7824), .ZN(n6924) );
  INV_X1 U5642 ( .A(n7496), .ZN(n8723) );
  NAND2_X1 U5643 ( .A1(n7746), .A2(n7745), .ZN(n8818) );
  AND2_X1 U5644 ( .A1(n8609), .A2(n8608), .ZN(n8828) );
  NAND2_X1 U5645 ( .A1(n6202), .A2(n6201), .ZN(n8835) );
  NAND2_X1 U5646 ( .A1(n6189), .A2(n6188), .ZN(n8841) );
  NAND2_X1 U5647 ( .A1(n4583), .A2(n4586), .ZN(n8623) );
  OR2_X1 U5648 ( .A1(n8659), .A2(n4589), .ZN(n4583) );
  NAND2_X1 U5649 ( .A1(n6180), .A2(n6179), .ZN(n8847) );
  NAND2_X1 U5650 ( .A1(n4591), .A2(n7927), .ZN(n8636) );
  NAND2_X1 U5651 ( .A1(n8659), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U5652 ( .A1(n6171), .A2(n6170), .ZN(n8853) );
  NAND2_X1 U5653 ( .A1(n8662), .A2(n6291), .ZN(n8652) );
  NAND2_X1 U5654 ( .A1(n8659), .A2(n7807), .ZN(n8650) );
  NAND2_X1 U5655 ( .A1(n6154), .A2(n6153), .ZN(n8996) );
  NAND2_X1 U5656 ( .A1(n8709), .A2(n4620), .ZN(n8674) );
  NAND2_X1 U5657 ( .A1(n6145), .A2(n6144), .ZN(n9002) );
  NAND2_X1 U5658 ( .A1(n8709), .A2(n7812), .ZN(n8688) );
  NAND2_X1 U5659 ( .A1(n6124), .A2(n6123), .ZN(n9012) );
  NAND2_X1 U5660 ( .A1(n6113), .A2(n6112), .ZN(n9018) );
  NAND2_X1 U5661 ( .A1(n8747), .A2(n7901), .ZN(n8730) );
  NAND2_X1 U5662 ( .A1(n9032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5958) );
  INV_X1 U5663 ( .A(n5961), .ZN(n7736) );
  INV_X1 U5664 ( .A(n7767), .ZN(n7821) );
  XNOR2_X1 U5665 ( .A(n5839), .B(n5838), .ZN(n6623) );
  NAND2_X1 U5666 ( .A1(n4432), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5836) );
  INV_X1 U5667 ( .A(n5820), .ZN(n4432) );
  OR2_X1 U5668 ( .A1(n5825), .A2(n5846), .ZN(n5827) );
  NAND2_X1 U5669 ( .A1(n5439), .A2(n5438), .ZN(n9474) );
  OR2_X1 U5670 ( .A1(n5079), .A2(n5616), .ZN(n5080) );
  CLKBUF_X1 U5671 ( .A(n9073), .Z(n9074) );
  INV_X1 U5672 ( .A(n9101), .ZN(n4808) );
  NAND2_X1 U5673 ( .A1(n5147), .A2(n5146), .ZN(n7303) );
  NAND2_X1 U5674 ( .A1(n5349), .A2(n5348), .ZN(n8110) );
  INV_X1 U5675 ( .A(n9084), .ZN(n4784) );
  AND2_X1 U5676 ( .A1(n5623), .A2(n4782), .ZN(n4781) );
  NAND2_X1 U5677 ( .A1(n9084), .A2(n4783), .ZN(n4782) );
  NAND2_X1 U5678 ( .A1(n7619), .A2(n5346), .ZN(n5605) );
  INV_X1 U5679 ( .A(n7238), .ZN(n9178) );
  INV_X1 U5680 ( .A(n7013), .ZN(n9180) );
  INV_X1 U5681 ( .A(n4376), .ZN(n9724) );
  NAND2_X1 U5682 ( .A1(n7697), .A2(n7696), .ZN(n9824) );
  AND2_X1 U5683 ( .A1(n9850), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9852) );
  NOR2_X1 U5684 ( .A1(n9852), .A2(n7707), .ZN(n9871) );
  NAND2_X1 U5685 ( .A1(n9871), .A2(n9872), .ZN(n9870) );
  INV_X1 U5686 ( .A(n4377), .ZN(n7715) );
  OAI211_X1 U5687 ( .C1(n7713), .C2(n9851), .A(n4378), .B(n9898), .ZN(n4377)
         );
  NAND2_X1 U5688 ( .A1(n7714), .A2(n9884), .ZN(n4378) );
  NOR2_X1 U5689 ( .A1(n9255), .A2(n9527), .ZN(n9540) );
  NAND2_X1 U5690 ( .A1(n4669), .A2(n4291), .ZN(n9333) );
  NAND2_X1 U5691 ( .A1(n9357), .A2(n4304), .ZN(n4669) );
  OAI21_X1 U5692 ( .B1(n9357), .B2(n9314), .A(n9313), .ZN(n9352) );
  NAND2_X1 U5693 ( .A1(n5633), .A2(n5632), .ZN(n9556) );
  NAND2_X1 U5694 ( .A1(n7634), .A2(n5346), .ZN(n5633) );
  NAND2_X1 U5695 ( .A1(n4540), .A2(n4545), .ZN(n9391) );
  AND2_X1 U5696 ( .A1(n9438), .A2(n9260), .ZN(n9419) );
  NAND2_X1 U5697 ( .A1(n4647), .A2(n4651), .ZN(n9472) );
  NAND2_X1 U5698 ( .A1(n4654), .A2(n4288), .ZN(n4647) );
  NAND2_X1 U5699 ( .A1(n9484), .A2(n8172), .ZN(n9466) );
  NAND2_X1 U5700 ( .A1(n4653), .A2(n4875), .ZN(n9482) );
  NAND2_X1 U5701 ( .A1(n4654), .A2(n9503), .ZN(n4653) );
  AND2_X1 U5702 ( .A1(n4662), .A2(n4322), .ZN(n9278) );
  NAND2_X1 U5703 ( .A1(n4663), .A2(n4664), .ZN(n4662) );
  OAI21_X1 U5704 ( .B1(n9906), .B2(n8002), .A(n4529), .ZN(n7597) );
  AND2_X1 U5705 ( .A1(n4638), .A2(n4290), .ZN(n7473) );
  NAND2_X1 U5706 ( .A1(n9915), .A2(n9914), .ZN(n4638) );
  NAND2_X1 U5707 ( .A1(n5277), .A2(n5276), .ZN(n9913) );
  INV_X1 U5708 ( .A(n9534), .ZN(n9938) );
  INV_X1 U5709 ( .A(n8213), .ZN(n9636) );
  NAND2_X1 U5710 ( .A1(n4338), .A2(n4551), .ZN(n9637) );
  AOI211_X1 U5711 ( .C1(n9559), .C2(n9958), .A(n9558), .B(n9557), .ZN(n9641)
         );
  INV_X1 U5712 ( .A(n9460), .ZN(n9662) );
  INV_X1 U5713 ( .A(n9512), .ZN(n9674) );
  NAND2_X1 U5714 ( .A1(n7662), .A2(n6238), .ZN(n7741) );
  OR2_X1 U5715 ( .A1(n6237), .A2(SI_29_), .ZN(n6238) );
  NAND2_X1 U5716 ( .A1(n5006), .A2(n4989), .ZN(n4631) );
  OR2_X1 U5717 ( .A1(n5037), .A2(n5036), .ZN(n5038) );
  OR2_X1 U5718 ( .A1(n5015), .A2(n9688), .ZN(n5011) );
  CLKBUF_X1 U5719 ( .A(n5043), .Z(n9350) );
  NAND2_X1 U5720 ( .A1(n4394), .A2(n4392), .ZN(n5098) );
  NAND2_X1 U5721 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4393), .ZN(n4392) );
  NAND2_X1 U5722 ( .A1(n5088), .A2(n5087), .ZN(n6486) );
  CLKBUF_X2 U5723 ( .A(n8455), .Z(P2_U3893) );
  AOI21_X1 U5724 ( .B1(n7976), .B2(n4600), .A(n4459), .ZN(n4597) );
  NAND2_X1 U5725 ( .A1(n9981), .A2(n4398), .ZN(n6635) );
  NAND2_X1 U5726 ( .A1(n4723), .A2(n4725), .ZN(n7157) );
  INV_X1 U5727 ( .A(n4480), .ZN(n7411) );
  INV_X1 U5728 ( .A(n4485), .ZN(n8475) );
  INV_X1 U5729 ( .A(n4482), .ZN(n8513) );
  OR2_X1 U5730 ( .A1(n8570), .A2(n8569), .ZN(n4405) );
  NOR2_X1 U5731 ( .A1(n8568), .A2(n4371), .ZN(n4406) );
  OAI21_X1 U5732 ( .B1(n4745), .B2(n8562), .A(n9990), .ZN(n4744) );
  NAND2_X1 U5733 ( .A1(n4427), .A2(n4425), .ZN(P2_U3201) );
  NOR2_X1 U5734 ( .A1(n5955), .A2(n4426), .ZN(n4425) );
  NAND2_X1 U5735 ( .A1(n4428), .A2(n9990), .ZN(n4427) );
  OAI22_X1 U5736 ( .A1(n6349), .A2(n8810), .B1(n10107), .B2(n6334), .ZN(n6335)
         );
  NAND2_X1 U5737 ( .A1(n8771), .A2(n4871), .ZN(n8773) );
  AOI21_X1 U5738 ( .B1(n8583), .B2(n6352), .A(n6351), .ZN(n6353) );
  NOR2_X1 U5739 ( .A1(n10080), .A2(n6350), .ZN(n6351) );
  OAI21_X1 U5740 ( .B1(n7666), .B2(n6376), .A(n4719), .ZN(P2_U3294) );
  NOR2_X1 U5741 ( .A1(n4721), .A2(n4720), .ZN(n4719) );
  NOR2_X1 U5742 ( .A1(n7734), .A2(n6367), .ZN(n4721) );
  NOR2_X1 U5743 ( .A1(n4506), .A2(n9114), .ZN(n4505) );
  NAND2_X1 U5744 ( .A1(n4574), .A2(n4573), .ZN(P1_U3242) );
  INV_X1 U5745 ( .A(n8242), .ZN(n4573) );
  OAI21_X1 U5746 ( .B1(n4576), .B2(n4575), .A(n8243), .ZN(n4574) );
  INV_X1 U5747 ( .A(n5043), .ZN(n5437) );
  AND2_X1 U5748 ( .A1(n9503), .A2(n4876), .ZN(n4288) );
  OR2_X1 U5749 ( .A1(n4409), .A2(n6998), .ZN(n4289) );
  OR2_X1 U5750 ( .A1(n9913), .A2(n9177), .ZN(n4290) );
  INV_X2 U5751 ( .A(n5148), .ZN(n6404) );
  INV_X1 U5752 ( .A(n9183), .ZN(n4634) );
  AND2_X1 U5753 ( .A1(n4675), .A2(n4674), .ZN(n4291) );
  XNOR2_X1 U5754 ( .A(n8829), .B(n8423), .ZN(n8603) );
  NOR2_X1 U5755 ( .A1(n9144), .A2(n9145), .ZN(n9048) );
  NAND2_X1 U5756 ( .A1(n5128), .A2(n6362), .ZN(n5101) );
  AND2_X1 U5757 ( .A1(n4465), .A2(n9686), .ZN(n4292) );
  AND2_X1 U5758 ( .A1(n7034), .A2(n4468), .ZN(n4293) );
  OR2_X1 U5759 ( .A1(n9556), .A2(n9315), .ZN(n4294) );
  AOI21_X1 U5760 ( .B1(n9986), .B2(n5834), .A(n4431), .ZN(n4732) );
  AND2_X1 U5761 ( .A1(n4637), .A2(n4643), .ZN(n4295) );
  AND2_X1 U5762 ( .A1(n4462), .A2(n4461), .ZN(n4296) );
  AND2_X1 U5763 ( .A1(n6047), .A2(n7866), .ZN(n4297) );
  AND2_X1 U5764 ( .A1(n6074), .A2(n7880), .ZN(n4298) );
  AND2_X1 U5765 ( .A1(n7275), .A2(n7273), .ZN(n4299) );
  XNOR2_X1 U5766 ( .A(n5836), .B(n5835), .ZN(n6381) );
  INV_X1 U5767 ( .A(n6381), .ZN(n4431) );
  OAI21_X1 U5768 ( .B1(n4349), .B2(n7401), .A(n7400), .ZN(n7399) );
  AND2_X1 U5769 ( .A1(n4727), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4301) );
  INV_X1 U5770 ( .A(n9063), .ZN(n4809) );
  NAND3_X1 U5771 ( .A1(n5061), .A2(n5708), .A3(n5060), .ZN(n5078) );
  INV_X2 U5772 ( .A(n5149), .ZN(n5213) );
  AND2_X1 U5773 ( .A1(n4934), .A2(n4933), .ZN(n4302) );
  INV_X1 U5774 ( .A(n6362), .ZN(n4471) );
  OR2_X1 U5775 ( .A1(n8689), .A2(n8690), .ZN(n4303) );
  NAND2_X1 U5776 ( .A1(n6308), .A2(n4471), .ZN(n5990) );
  AND2_X1 U5777 ( .A1(n4294), .A2(n9313), .ZN(n4304) );
  AND2_X1 U5778 ( .A1(n7492), .A2(n7885), .ZN(n4305) );
  AND4_X1 U5779 ( .A1(n5372), .A2(n5368), .A3(n5321), .A4(n4981), .ZN(n4307)
         );
  OR2_X1 U5780 ( .A1(n6308), .A2(n6381), .ZN(n4308) );
  AND2_X1 U5781 ( .A1(n4549), .A2(n9264), .ZN(n4309) );
  NAND2_X1 U5782 ( .A1(n8248), .A2(n8443), .ZN(n4310) );
  NAND2_X1 U5783 ( .A1(n10061), .A2(n8446), .ZN(n4311) );
  NAND2_X1 U5784 ( .A1(n5382), .A2(n5364), .ZN(n4312) );
  NAND2_X1 U5785 ( .A1(n7739), .A2(n5031), .ZN(n5065) );
  INV_X1 U5786 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4404) );
  AND2_X1 U5787 ( .A1(n8203), .A2(n8223), .ZN(n4314) );
  INV_X1 U5788 ( .A(n5993), .ZN(n6242) );
  OR2_X1 U5789 ( .A1(n4450), .A2(n7938), .ZN(n4315) );
  INV_X1 U5790 ( .A(n5206), .ZN(n4919) );
  XNOR2_X1 U5791 ( .A(n4920), .B(SI_7_), .ZN(n5206) );
  AND2_X1 U5792 ( .A1(n9380), .A2(n4464), .ZN(n4316) );
  AND2_X1 U5793 ( .A1(n4477), .A2(n4476), .ZN(n4317) );
  AND2_X1 U5794 ( .A1(n6286), .A2(n4837), .ZN(n4318) );
  NAND2_X1 U5795 ( .A1(n5376), .A2(n5375), .ZN(n8106) );
  INV_X1 U5796 ( .A(n8173), .ZN(n4563) );
  INV_X1 U5797 ( .A(n8204), .ZN(n9318) );
  AND2_X1 U5798 ( .A1(n8206), .A2(n8205), .ZN(n8204) );
  NAND2_X1 U5799 ( .A1(n5325), .A2(n5324), .ZN(n9779) );
  NAND2_X1 U5800 ( .A1(n5302), .A2(n5301), .ZN(n7523) );
  AND2_X1 U5801 ( .A1(n4491), .A2(n4490), .ZN(n9047) );
  NAND2_X1 U5802 ( .A1(n8201), .A2(n9268), .ZN(n9316) );
  OR2_X1 U5803 ( .A1(n8200), .A2(n8209), .ZN(n4319) );
  INV_X1 U5804 ( .A(n7075), .ZN(n4819) );
  AND2_X1 U5805 ( .A1(n10055), .A2(n8447), .ZN(n4320) );
  NAND2_X1 U5806 ( .A1(n5523), .A2(n5524), .ZN(n9144) );
  OR2_X1 U5807 ( .A1(n5792), .A2(n5753), .ZN(n4321) );
  NAND2_X1 U5808 ( .A1(n5760), .A2(n5759), .ZN(n5771) );
  NAND2_X1 U5809 ( .A1(n9686), .A2(n8111), .ZN(n4322) );
  NAND2_X1 U5810 ( .A1(n5234), .A2(n5233), .ZN(n9790) );
  XNOR2_X1 U5811 ( .A(n5042), .B(n5041), .ZN(n5043) );
  AND2_X1 U5812 ( .A1(n8106), .A2(n9174), .ZN(n4323) );
  INV_X1 U5813 ( .A(n8172), .ZN(n4538) );
  AND3_X1 U5814 ( .A1(n8204), .A2(n4884), .A3(n4577), .ZN(n4324) );
  NAND2_X1 U5815 ( .A1(n5658), .A2(n5657), .ZN(n9334) );
  OR2_X1 U5816 ( .A1(n8823), .A2(n8607), .ZN(n4325) );
  NOR2_X1 U5817 ( .A1(n8532), .A2(n5896), .ZN(n4326) );
  INV_X1 U5818 ( .A(n4805), .ZN(n4804) );
  OAI21_X1 U5819 ( .B1(n4807), .B2(n4806), .A(n4809), .ZN(n4805) );
  AND4_X1 U5820 ( .A1(n5285), .A2(n5284), .A3(n5283), .A4(n5282), .ZN(n7449)
         );
  INV_X1 U5821 ( .A(n6272), .ZN(n4822) );
  AND2_X1 U5822 ( .A1(n7853), .A2(n7844), .ZN(n4327) );
  OR2_X1 U5823 ( .A1(n5517), .A2(n7029), .ZN(n4328) );
  AND2_X1 U5824 ( .A1(n6282), .A2(n6281), .ZN(n4329) );
  AND2_X1 U5825 ( .A1(n4742), .A2(n4741), .ZN(n4330) );
  AND2_X1 U5826 ( .A1(n4988), .A2(n4987), .ZN(n4331) );
  NAND2_X1 U5827 ( .A1(n5844), .A2(n6384), .ZN(n4715) );
  NAND2_X1 U5828 ( .A1(n4811), .A2(n4810), .ZN(n9060) );
  AND2_X1 U5829 ( .A1(n5834), .A2(n4431), .ZN(n4332) );
  INV_X1 U5830 ( .A(n9563), .ZN(n9363) );
  NAND2_X1 U5831 ( .A1(n5605), .A2(n5604), .ZN(n9563) );
  NOR2_X1 U5832 ( .A1(n10055), .A2(n8447), .ZN(n4333) );
  NOR2_X1 U5833 ( .A1(n8823), .A2(n7949), .ZN(n4334) );
  NOR2_X1 U5834 ( .A1(n8853), .A2(n8665), .ZN(n4335) );
  NAND2_X1 U5835 ( .A1(n8456), .A2(n6257), .ZN(n7823) );
  INV_X1 U5836 ( .A(n7823), .ZN(n4594) );
  INV_X1 U5837 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4772) );
  AND4_X1 U5838 ( .A1(n5069), .A2(n5068), .A3(n5067), .A4(n5066), .ZN(n5076)
         );
  AND4_X1 U5839 ( .A1(n5186), .A2(n5185), .A3(n5184), .A4(n5183), .ZN(n6976)
         );
  AND2_X1 U5840 ( .A1(n4920), .A2(SI_7_), .ZN(n4336) );
  AND2_X1 U5841 ( .A1(n7800), .A2(n7801), .ZN(n4337) );
  AND2_X1 U5842 ( .A1(n4552), .A2(n9273), .ZN(n4338) );
  AND2_X1 U5843 ( .A1(n9373), .A2(n8189), .ZN(n9390) );
  INV_X1 U5844 ( .A(n9390), .ZN(n4542) );
  OR2_X1 U5845 ( .A1(n8064), .A2(n4643), .ZN(n4339) );
  NAND2_X1 U5846 ( .A1(n8336), .A2(n8335), .ZN(n4340) );
  NAND2_X1 U5847 ( .A1(n8045), .A2(n9328), .ZN(n9351) );
  INV_X1 U5848 ( .A(n9351), .ZN(n4676) );
  NAND2_X1 U5849 ( .A1(n4808), .A2(n4807), .ZN(n4811) );
  INV_X1 U5850 ( .A(n7029), .ZN(n9924) );
  AND3_X1 U5851 ( .A1(n5131), .A2(n5130), .A3(n5129), .ZN(n7029) );
  INV_X1 U5852 ( .A(n8065), .ZN(n4660) );
  AND2_X1 U5853 ( .A1(n8148), .A2(n8138), .ZN(n8065) );
  NOR2_X1 U5854 ( .A1(n7951), .A2(n7949), .ZN(n4341) );
  OAI21_X1 U5855 ( .B1(n4539), .B2(n4538), .A(n9471), .ZN(n4537) );
  OR2_X1 U5856 ( .A1(n9002), .A2(n8706), .ZN(n6288) );
  INV_X1 U5857 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9688) );
  OR2_X1 U5858 ( .A1(n4886), .A2(n4652), .ZN(n4342) );
  OR2_X1 U5859 ( .A1(n6266), .A2(n4832), .ZN(n4343) );
  AND2_X1 U5860 ( .A1(n5876), .A2(n4431), .ZN(n4344) );
  INV_X1 U5861 ( .A(n7848), .ZN(n4610) );
  AND2_X1 U5862 ( .A1(n7941), .A2(n8601), .ZN(n4345) );
  AND2_X1 U5863 ( .A1(n4528), .A2(n8065), .ZN(n4346) );
  INV_X1 U5864 ( .A(n9774), .ZN(n4795) );
  INV_X1 U5865 ( .A(n4651), .ZN(n4650) );
  NAND2_X1 U5866 ( .A1(n4342), .A2(n4876), .ZN(n4651) );
  AND2_X1 U5867 ( .A1(n4627), .A2(n5956), .ZN(n4347) );
  INV_X1 U5868 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4393) );
  INV_X1 U5869 ( .A(n9493), .ZN(n9670) );
  NAND2_X1 U5870 ( .A1(n4994), .A2(n4993), .ZN(n9493) );
  AND2_X1 U5871 ( .A1(n4337), .A2(n4600), .ZN(n4348) );
  INV_X1 U5872 ( .A(n4915), .ZN(n4526) );
  INV_X1 U5873 ( .A(n4621), .ZN(n4620) );
  NAND2_X1 U5874 ( .A1(n6288), .A2(n7812), .ZN(n4621) );
  INV_X1 U5875 ( .A(n5119), .ZN(n5149) );
  OAI21_X1 U5876 ( .B1(n7741), .B2(n5101), .A(n7722), .ZN(n9321) );
  INV_X1 U5877 ( .A(n9321), .ZN(n4461) );
  INV_X1 U5878 ( .A(n5120), .ZN(n5148) );
  AND2_X1 U5879 ( .A1(n5292), .A2(n4792), .ZN(n4349) );
  NOR2_X1 U5880 ( .A1(n5480), .A2(n4703), .ZN(n4702) );
  INV_X1 U5881 ( .A(n4777), .ZN(n5388) );
  INV_X1 U5882 ( .A(n8731), .ZN(n4838) );
  AND3_X1 U5883 ( .A1(n5701), .A2(n9158), .A3(n5700), .ZN(n4350) );
  NAND2_X1 U5884 ( .A1(n4992), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U5885 ( .A1(n4495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5040) );
  INV_X1 U5886 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5321) );
  INV_X1 U5887 ( .A(n7852), .ZN(n4606) );
  NAND2_X1 U5888 ( .A1(n7435), .A2(n7434), .ZN(n7532) );
  NAND2_X1 U5889 ( .A1(n4768), .A2(n4766), .ZN(n8363) );
  NOR2_X1 U5890 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5252) );
  AND2_X1 U5891 ( .A1(n8099), .A2(n8046), .ZN(n4351) );
  AND2_X1 U5892 ( .A1(n8728), .A2(n7814), .ZN(n4352) );
  INV_X1 U5893 ( .A(n7723), .ZN(n9443) );
  NOR2_X1 U5894 ( .A1(n9457), .A2(n9444), .ZN(n7723) );
  NAND2_X1 U5895 ( .A1(n8291), .A2(n8349), .ZN(n4353) );
  AND2_X1 U5896 ( .A1(n8263), .A2(n8262), .ZN(n4354) );
  AND2_X1 U5897 ( .A1(n8278), .A2(n8277), .ZN(n4355) );
  AND2_X1 U5898 ( .A1(n4838), .A2(n7901), .ZN(n4356) );
  OR2_X1 U5899 ( .A1(n4885), .A2(n5730), .ZN(n4357) );
  AND4_X1 U5900 ( .A1(n5310), .A2(n5309), .A3(n5308), .A4(n5307), .ZN(n7450)
         );
  NAND2_X1 U5901 ( .A1(n6241), .A2(n6240), .ZN(n8583) );
  AND2_X1 U5902 ( .A1(n5499), .A2(SI_21_), .ZN(n4358) );
  INV_X1 U5903 ( .A(n4699), .ZN(n4698) );
  NAND2_X1 U5904 ( .A1(n4701), .A2(n5497), .ZN(n4699) );
  OR2_X1 U5905 ( .A1(n6958), .A2(n10097), .ZN(n4359) );
  NAND2_X1 U5906 ( .A1(n5479), .A2(n5478), .ZN(n4360) );
  NAND2_X1 U5907 ( .A1(n5505), .A2(n5504), .ZN(n9424) );
  NOR2_X1 U5908 ( .A1(n7316), .A2(n7380), .ZN(n4361) );
  INV_X1 U5909 ( .A(n5365), .ZN(n4714) );
  AND2_X1 U5910 ( .A1(n4759), .A2(n8344), .ZN(n4362) );
  NAND2_X1 U5911 ( .A1(n6538), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4363) );
  AND2_X1 U5912 ( .A1(n9049), .A2(n4492), .ZN(n4364) );
  INV_X1 U5913 ( .A(n9914), .ZN(n4643) );
  AND2_X1 U5914 ( .A1(n6915), .A2(n6910), .ZN(n4365) );
  AND2_X1 U5915 ( .A1(n7480), .A2(n7589), .ZN(n4366) );
  AOI21_X1 U5916 ( .B1(n8023), .B2(n8022), .A(n8021), .ZN(n4529) );
  NAND2_X1 U5917 ( .A1(n6001), .A2(n7844), .ZN(n6859) );
  NOR2_X1 U5918 ( .A1(n7164), .A2(n4317), .ZN(n4367) );
  NAND2_X1 U5919 ( .A1(n7480), .A2(n4292), .ZN(n4466) );
  INV_X1 U5920 ( .A(n6002), .ZN(n6013) );
  NAND2_X1 U5921 ( .A1(n6538), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4368) );
  AND2_X1 U5922 ( .A1(n7020), .A2(n4293), .ZN(n7182) );
  NAND2_X1 U5923 ( .A1(n4763), .A2(n4306), .ZN(n4369) );
  INV_X1 U5924 ( .A(n4290), .ZN(n4644) );
  XNOR2_X1 U5925 ( .A(n5025), .B(n5028), .ZN(n5723) );
  OR2_X1 U5926 ( .A1(n8519), .A2(n5894), .ZN(n4370) );
  INV_X1 U5927 ( .A(n7263), .ZN(n4468) );
  INV_X1 U5928 ( .A(n6998), .ZN(n4410) );
  OR2_X1 U5929 ( .A1(n8566), .A2(n8567), .ZN(n4371) );
  INV_X1 U5930 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n4738) );
  XNOR2_X1 U5931 ( .A(n5958), .B(n5957), .ZN(n7737) );
  INV_X1 U5932 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4518) );
  NAND3_X1 U5933 ( .A1(n4777), .A2(n4778), .A3(n4331), .ZN(n9687) );
  INV_X1 U5934 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4419) );
  INV_X1 U5935 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n4379) );
  AND2_X1 U5936 ( .A1(n9574), .A2(n4282), .ZN(n4506) );
  OR2_X1 U5937 ( .A1(n5853), .A2(n7161), .ZN(n4727) );
  AND2_X1 U5938 ( .A1(n5853), .A2(n7161), .ZN(n4726) );
  INV_X1 U5939 ( .A(n7161), .ZN(n4476) );
  OR2_X1 U5940 ( .A1(n6947), .A2(n7161), .ZN(n4724) );
  AOI21_X1 U5941 ( .B1(n6947), .B2(n5853), .A(n7161), .ZN(n5854) );
  NOR2_X4 U5942 ( .A1(n6684), .A2(n8644), .ZN(n8762) );
  AND2_X2 U5943 ( .A1(n5290), .A2(n5289), .ZN(n7401) );
  OR2_X1 U5944 ( .A1(n6896), .A2(n6898), .ZN(n5199) );
  NOR2_X1 U5945 ( .A1(n9772), .A2(n5343), .ZN(n7508) );
  AOI21_X1 U5946 ( .B1(n7506), .B2(n4503), .A(n4501), .ZN(n5401) );
  NAND2_X1 U5947 ( .A1(n4489), .A2(n4372), .ZN(n4488) );
  NAND3_X1 U5948 ( .A1(n5096), .A2(n4980), .A3(n4979), .ZN(n5320) );
  OR2_X1 U5949 ( .A1(n5001), .A2(n5000), .ZN(n5005) );
  NAND2_X1 U5950 ( .A1(n9050), .A2(n9049), .ZN(n4491) );
  NOR2_X1 U5951 ( .A1(n5158), .A2(n4500), .ZN(n4498) );
  XNOR2_X1 U5952 ( .A(n4905), .B(SI_3_), .ZN(n4373) );
  XNOR2_X1 U5953 ( .A(n4373), .B(n5126), .ZN(n6380) );
  NAND2_X1 U5954 ( .A1(n5345), .A2(n4951), .ZN(n4387) );
  OAI22_X1 U5955 ( .A1(n4389), .A2(n7751), .B1(SI_30_), .B2(n7750), .ZN(n7754)
         );
  NAND2_X1 U5956 ( .A1(n4390), .A2(n4918), .ZN(n5205) );
  OAI21_X1 U5957 ( .B1(n5086), .B2(n9688), .A(P1_IR_REG_2__SCAN_IN), .ZN(n4394) );
  NAND2_X1 U5958 ( .A1(n4395), .A2(n4934), .ZN(n5273) );
  OAI21_X1 U5959 ( .B1(n6637), .B2(n4400), .A(n6634), .ZN(n4399) );
  NAND2_X1 U5960 ( .A1(n6637), .A2(n4400), .ZN(n6634) );
  AND3_X2 U5961 ( .A1(n4401), .A2(n5794), .A3(n4843), .ZN(n5760) );
  INV_X1 U5962 ( .A(n8557), .ZN(n8554) );
  AND3_X2 U5963 ( .A1(n5826), .A2(n4404), .A3(n4403), .ZN(n5820) );
  NAND3_X1 U5964 ( .A1(n4744), .A2(n4406), .A3(n4405), .ZN(P2_U3200) );
  NAND3_X1 U5965 ( .A1(n4407), .A2(n4289), .A3(n4299), .ZN(n7362) );
  NAND2_X1 U5966 ( .A1(n4411), .A2(n4412), .ZN(n8245) );
  NAND3_X1 U5967 ( .A1(n7435), .A2(n4771), .A3(n7544), .ZN(n4411) );
  NAND2_X2 U5968 ( .A1(n8323), .A2(n8269), .ZN(n8336) );
  NAND3_X1 U5969 ( .A1(n4443), .A2(n4445), .A3(n4345), .ZN(n7946) );
  NAND3_X1 U5970 ( .A1(n7924), .A2(n4446), .A3(n4315), .ZN(n4443) );
  NAND2_X1 U5971 ( .A1(n8615), .A2(n7937), .ZN(n4449) );
  INV_X2 U5972 ( .A(n6308), .ZN(n6131) );
  NAND2_X2 U5973 ( .A1(n6308), .A2(n6362), .ZN(n5991) );
  NAND2_X2 U5974 ( .A1(n5871), .A2(n7657), .ZN(n6308) );
  NOR2_X2 U5975 ( .A1(n4986), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4778) );
  NAND4_X1 U5976 ( .A1(n4985), .A2(n4982), .A3(n4984), .A4(n4983), .ZN(n4986)
         );
  INV_X1 U5977 ( .A(n4466), .ZN(n7640) );
  NAND3_X1 U5978 ( .A1(n7020), .A2(n4293), .A3(n7181), .ZN(n7242) );
  NAND2_X2 U5979 ( .A1(n5128), .A2(n4471), .ZN(n5127) );
  OAI21_X2 U5980 ( .B1(n5128), .B2(n6486), .A(n4469), .ZN(n6666) );
  OAI21_X1 U5981 ( .B1(n7165), .B2(n4868), .A(n4475), .ZN(n7311) );
  OR2_X1 U5982 ( .A1(n5593), .A2(n6541), .ZN(n4489) );
  NAND3_X1 U5983 ( .A1(n4491), .A2(n4490), .A3(n9113), .ZN(n5573) );
  NAND3_X1 U5984 ( .A1(n5523), .A2(n5524), .A3(n4364), .ZN(n4490) );
  NAND2_X1 U5985 ( .A1(n5049), .A2(n4496), .ZN(n4494) );
  OAI21_X1 U5986 ( .B1(n4499), .B2(n4498), .A(n5204), .ZN(n6873) );
  NAND2_X1 U5987 ( .A1(n6646), .A2(n5163), .ZN(n6895) );
  NAND2_X1 U5988 ( .A1(n5158), .A2(n5157), .ZN(n6646) );
  OR2_X1 U5989 ( .A1(n7506), .A2(n4312), .ZN(n9037) );
  OAI21_X1 U5990 ( .B1(n7506), .B2(n4504), .A(n5383), .ZN(n4780) );
  AOI22_X1 U5991 ( .A1(n4312), .A2(n9038), .B1(n4504), .B2(n5383), .ZN(n4502)
         );
  OR2_X1 U5992 ( .A1(n5383), .A2(n9038), .ZN(n4503) );
  NAND2_X1 U5993 ( .A1(n4507), .A2(n4505), .ZN(P1_U3229) );
  NAND2_X1 U5994 ( .A1(n4508), .A2(n9158), .ZN(n4507) );
  NAND2_X1 U5995 ( .A1(n4509), .A2(n9110), .ZN(n4508) );
  NAND2_X1 U5996 ( .A1(n4511), .A2(n4796), .ZN(n9133) );
  NAND2_X1 U5997 ( .A1(n9101), .A2(n4800), .ZN(n4511) );
  NOR2_X1 U5998 ( .A1(n7668), .A2(n5404), .ZN(n9093) );
  NAND2_X1 U5999 ( .A1(n4513), .A2(n4901), .ZN(n5126) );
  NAND2_X1 U6000 ( .A1(n5099), .A2(n5100), .ZN(n4513) );
  INV_X1 U6001 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4516) );
  INV_X1 U6002 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4517) );
  NAND3_X1 U6003 ( .A1(n4519), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4514) );
  NAND3_X1 U6004 ( .A1(n4518), .A2(n4517), .A3(n4516), .ZN(n4515) );
  NAND3_X1 U6005 ( .A1(n4522), .A2(n4919), .A3(n4526), .ZN(n4520) );
  NAND2_X1 U6006 ( .A1(n4527), .A2(n4346), .ZN(n7598) );
  NAND2_X1 U6007 ( .A1(n9906), .A2(n4529), .ZN(n4527) );
  NAND3_X1 U6008 ( .A1(n7451), .A2(n8154), .A3(n8132), .ZN(n4530) );
  NAND2_X1 U6009 ( .A1(n9506), .A2(n4535), .ZN(n4534) );
  AND2_X1 U6010 ( .A1(n9486), .A2(n9483), .ZN(n4539) );
  AOI211_X2 U6011 ( .C1(n9549), .C2(n9917), .A(n9548), .B(n4313), .ZN(n4551)
         );
  AND2_X2 U6012 ( .A1(n8009), .A2(n6776), .ZN(n8051) );
  NAND3_X1 U6013 ( .A1(n4566), .A2(n8173), .A3(n9259), .ZN(n4565) );
  NAND2_X1 U6014 ( .A1(n4567), .A2(n4568), .ZN(n8162) );
  NAND2_X1 U6015 ( .A1(n8150), .A2(n4569), .ZN(n4567) );
  NAND3_X1 U6016 ( .A1(n8199), .A2(n8209), .A3(n8198), .ZN(n4581) );
  NAND2_X1 U6017 ( .A1(n4582), .A2(n4584), .ZN(n6200) );
  NAND2_X1 U6018 ( .A1(n8659), .A2(n4586), .ZN(n4582) );
  NAND2_X1 U6019 ( .A1(n4593), .A2(n7772), .ZN(n6923) );
  INV_X1 U6020 ( .A(n7772), .ZN(n7829) );
  NAND2_X1 U6021 ( .A1(n4595), .A2(n4597), .ZN(P2_U3296) );
  NAND3_X1 U6022 ( .A1(n4596), .A2(n4348), .A3(n7977), .ZN(n4595) );
  NAND2_X1 U6023 ( .A1(n4598), .A2(n4599), .ZN(n4596) );
  INV_X1 U6024 ( .A(n7805), .ZN(n4598) );
  NAND2_X1 U6025 ( .A1(n4603), .A2(n4601), .ZN(n7124) );
  NAND2_X1 U6026 ( .A1(n6001), .A2(n4602), .ZN(n4601) );
  NOR2_X1 U6027 ( .A1(n4608), .A2(n7846), .ZN(n4602) );
  NOR2_X1 U6028 ( .A1(n7846), .A2(n7848), .ZN(n4604) );
  NAND2_X1 U6029 ( .A1(n4609), .A2(n7842), .ZN(n4608) );
  OAI21_X1 U6030 ( .B1(n6001), .B2(n4610), .A(n4607), .ZN(n7041) );
  NAND2_X1 U6031 ( .A1(n4617), .A2(n4297), .ZN(n7285) );
  OAI21_X1 U6032 ( .B1(n8708), .B2(n4621), .A(n4618), .ZN(n6158) );
  NAND4_X1 U6033 ( .A1(n4624), .A2(n4623), .A3(n4772), .A4(n4622), .ZN(n5753)
         );
  NAND2_X1 U6034 ( .A1(n6065), .A2(n4298), .ZN(n7492) );
  AND2_X1 U6035 ( .A1(n5775), .A2(n4627), .ZN(n5959) );
  NAND2_X1 U6036 ( .A1(n5775), .A2(n4347), .ZN(n9032) );
  NAND2_X1 U6037 ( .A1(n4629), .A2(n6801), .ZN(n6803) );
  INV_X1 U6038 ( .A(n6804), .ZN(n4628) );
  NAND2_X1 U6039 ( .A1(n4629), .A2(n6804), .ZN(n6805) );
  NAND2_X1 U6040 ( .A1(n4630), .A2(n8051), .ZN(n6802) );
  INV_X1 U6041 ( .A(n6801), .ZN(n4630) );
  XNOR2_X2 U6042 ( .A(n4631), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6469) );
  OAI22_X2 U6043 ( .A1(n7447), .A2(n7446), .B1(n5265), .B2(n9760), .ZN(n9915)
         );
  INV_X1 U6044 ( .A(n4645), .ZN(n7472) );
  INV_X1 U6045 ( .A(n9501), .ZN(n4654) );
  NAND2_X1 U6046 ( .A1(n4646), .A2(n4648), .ZN(n9289) );
  NAND2_X1 U6047 ( .A1(n9501), .A2(n4651), .ZN(n4646) );
  INV_X1 U6048 ( .A(n4664), .ZN(n4658) );
  INV_X1 U6049 ( .A(n4663), .ZN(n7596) );
  NOR2_X1 U6050 ( .A1(n7596), .A2(n4665), .ZN(n7636) );
  NAND2_X1 U6051 ( .A1(n9311), .A2(n4667), .ZN(n4666) );
  NAND2_X1 U6052 ( .A1(n9311), .A2(n9310), .ZN(n9357) );
  NAND2_X1 U6053 ( .A1(n4666), .A2(n4670), .ZN(n9319) );
  NAND2_X1 U6054 ( .A1(n5576), .A2(n5575), .ZN(n4677) );
  NAND2_X1 U6055 ( .A1(n7967), .A2(n4679), .ZN(n4678) );
  NAND2_X1 U6056 ( .A1(n5294), .A2(n4943), .ZN(n4945) );
  INV_X1 U6057 ( .A(n5272), .ZN(n4683) );
  NAND3_X1 U6058 ( .A1(n4689), .A2(n5206), .A3(n4688), .ZN(n4686) );
  NAND2_X1 U6059 ( .A1(n5627), .A2(n4694), .ZN(n4691) );
  OAI21_X1 U6060 ( .B1(n5627), .B2(n4697), .A(n4694), .ZN(n6234) );
  NAND2_X1 U6061 ( .A1(n4691), .A2(n4692), .ZN(n6236) );
  NAND2_X1 U6062 ( .A1(n5627), .A2(n5626), .ZN(n5651) );
  OAI21_X1 U6063 ( .B1(n5432), .B2(n5431), .A(n5430), .ZN(n5481) );
  NAND2_X1 U6064 ( .A1(n4716), .A2(n5832), .ZN(n6626) );
  NAND2_X1 U6065 ( .A1(n5830), .A2(n4717), .ZN(n4716) );
  NOR2_X1 U6066 ( .A1(n5825), .A2(n5831), .ZN(n4717) );
  INV_X1 U6067 ( .A(n4718), .ZN(n5916) );
  OAI21_X1 U6068 ( .B1(n4718), .B2(n5874), .A(n5875), .ZN(n6624) );
  NAND2_X1 U6069 ( .A1(n6131), .A2(n4718), .ZN(n5970) );
  NOR2_X1 U6070 ( .A1(P2_U3151), .A2(n4718), .ZN(n4720) );
  NAND2_X1 U6071 ( .A1(n5918), .A2(n4718), .ZN(n5919) );
  OAI211_X1 U6072 ( .C1(n9993), .C2(n4718), .A(n6636), .B(n6635), .ZN(P2_U3183) );
  INV_X1 U6073 ( .A(n4729), .ZN(n7156) );
  NAND3_X1 U6074 ( .A1(n4731), .A2(n4730), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n6613) );
  NAND2_X1 U6075 ( .A1(n4332), .A2(n9986), .ZN(n4730) );
  INV_X1 U6076 ( .A(n4732), .ZN(n4731) );
  NAND2_X1 U6077 ( .A1(n6613), .A2(n4731), .ZN(n5840) );
  NAND2_X1 U6078 ( .A1(n7351), .A2(n4737), .ZN(n4733) );
  NAND2_X1 U6079 ( .A1(n4734), .A2(n4733), .ZN(n7415) );
  NAND2_X1 U6080 ( .A1(n5863), .A2(n4743), .ZN(n4739) );
  XNOR2_X1 U6081 ( .A(n5862), .B(n8502), .ZN(n8495) );
  NAND2_X1 U6082 ( .A1(n4743), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4740) );
  INV_X1 U6083 ( .A(n8525), .ZN(n4743) );
  INV_X1 U6084 ( .A(n8564), .ZN(n4747) );
  NAND4_X1 U6085 ( .A1(n4748), .A2(n5798), .A3(n5816), .A4(n5748), .ZN(n5751)
         );
  NAND2_X1 U6086 ( .A1(n8343), .A2(n4362), .ZN(n4753) );
  NAND2_X1 U6087 ( .A1(n4756), .A2(n8344), .ZN(n8419) );
  OR2_X1 U6088 ( .A1(n8343), .A2(n8345), .ZN(n4756) );
  NAND2_X2 U6089 ( .A1(n4763), .A2(n4760), .ZN(n6915) );
  NOR2_X1 U6090 ( .A1(n4762), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U6091 ( .A1(n6741), .A2(n6742), .ZN(n4763) );
  NAND3_X1 U6092 ( .A1(n4306), .A2(n4763), .A3(n6761), .ZN(n6762) );
  NAND2_X1 U6093 ( .A1(n8394), .A2(n8277), .ZN(n4765) );
  AND2_X2 U6094 ( .A1(n4764), .A2(n8280), .ZN(n8313) );
  NAND2_X1 U6095 ( .A1(n4765), .A2(n8279), .ZN(n4764) );
  NAND2_X2 U6096 ( .A1(n6450), .A2(n4774), .ZN(n6714) );
  NAND2_X1 U6097 ( .A1(n5093), .A2(n4776), .ZN(n5094) );
  XNOR2_X1 U6098 ( .A(n4776), .B(n5092), .ZN(n6664) );
  NOR2_X1 U6099 ( .A1(n5388), .A2(n4986), .ZN(n5002) );
  NOR2_X1 U6100 ( .A1(n6875), .A2(n6876), .ZN(n6874) );
  NAND2_X1 U6101 ( .A1(n9110), .A2(n5574), .ZN(n9082) );
  OAI21_X2 U6102 ( .B1(n9110), .B2(n4784), .A(n4781), .ZN(n9157) );
  NAND2_X1 U6103 ( .A1(n9082), .A2(n9084), .ZN(n9083) );
  AND2_X2 U6104 ( .A1(n9157), .A2(n4882), .ZN(n5737) );
  NAND2_X1 U6105 ( .A1(n4785), .A2(n9774), .ZN(n4787) );
  NAND4_X1 U6106 ( .A1(n5291), .A2(n5292), .A3(n4794), .A4(n4786), .ZN(n4790)
         );
  NAND3_X1 U6107 ( .A1(n4790), .A2(n4789), .A3(n4788), .ZN(n9772) );
  NAND2_X1 U6108 ( .A1(n5291), .A2(n5292), .ZN(n9755) );
  INV_X1 U6109 ( .A(n9060), .ZN(n9061) );
  NAND2_X1 U6110 ( .A1(n6271), .A2(n4815), .ZN(n4812) );
  NAND2_X1 U6111 ( .A1(n4812), .A2(n4813), .ZN(n7373) );
  NAND2_X1 U6112 ( .A1(n8663), .A2(n4826), .ZN(n4825) );
  NAND2_X1 U6113 ( .A1(n6887), .A2(n4829), .ZN(n4831) );
  NAND2_X1 U6114 ( .A1(n6284), .A2(n4318), .ZN(n4836) );
  NAND2_X1 U6115 ( .A1(n4842), .A2(n4841), .ZN(n7392) );
  INV_X1 U6116 ( .A(n5753), .ZN(n4843) );
  NAND2_X1 U6117 ( .A1(n5794), .A2(n5752), .ZN(n5792) );
  NAND2_X1 U6118 ( .A1(n4844), .A2(n4845), .ZN(n6299) );
  NAND2_X1 U6119 ( .A1(n8604), .A2(n4846), .ZN(n4844) );
  AND2_X1 U6120 ( .A1(n8604), .A2(n8603), .ZN(n8605) );
  NAND2_X1 U6121 ( .A1(n6692), .A2(n4852), .ZN(n4848) );
  AOI21_X1 U6122 ( .B1(n4856), .B2(n6381), .A(n10087), .ZN(n4860) );
  AOI21_X1 U6123 ( .B1(n9996), .B2(n5876), .A(n4431), .ZN(n4857) );
  INV_X1 U6124 ( .A(n4859), .ZN(n4858) );
  NAND2_X1 U6125 ( .A1(n4344), .A2(n9996), .ZN(n4861) );
  NAND2_X1 U6126 ( .A1(n4863), .A2(n6381), .ZN(n6606) );
  NAND2_X1 U6127 ( .A1(n9996), .A2(n5876), .ZN(n4863) );
  NAND2_X1 U6128 ( .A1(n6608), .A2(n6606), .ZN(n5877) );
  INV_X1 U6129 ( .A(n5535), .ZN(n5532) );
  AOI21_X1 U6130 ( .B1(n9553), .B2(n9958), .A(n9552), .ZN(n9638) );
  XNOR2_X1 U6131 ( .A(n9333), .B(n9332), .ZN(n9553) );
  AOI21_X1 U6132 ( .B1(n8596), .B2(n8752), .A(n8595), .ZN(n8822) );
  NAND2_X1 U6133 ( .A1(n6362), .A2(n6356), .ZN(n4903) );
  OR2_X1 U6134 ( .A1(n6362), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U6135 ( .A1(n4892), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4890) );
  INV_X1 U6136 ( .A(n5990), .ZN(n6028) );
  NAND2_X1 U6137 ( .A1(n5702), .A2(n4350), .ZN(n5733) );
  OR2_X1 U6138 ( .A1(n5290), .A2(n5289), .ZN(n5291) );
  INV_X1 U6139 ( .A(n7737), .ZN(n5962) );
  NAND2_X1 U6140 ( .A1(n7737), .A2(n5961), .ZN(n5992) );
  NAND2_X1 U6141 ( .A1(n4286), .A2(n10085), .ZN(n5873) );
  CLKBUF_X1 U6142 ( .A(n6873), .Z(n6875) );
  INV_X1 U6143 ( .A(n5524), .ZN(n9050) );
  NAND2_X1 U6144 ( .A1(n5879), .A2(n6384), .ZN(n5880) );
  NAND2_X1 U6145 ( .A1(n5401), .A2(n5400), .ZN(n5402) );
  NAND2_X1 U6146 ( .A1(n7362), .A2(n7361), .ZN(n7432) );
  AOI21_X2 U6147 ( .B1(n8252), .B2(n8251), .A(n4873), .ZN(n8430) );
  AND2_X1 U6148 ( .A1(n8799), .A2(n8721), .ZN(n4870) );
  OR2_X1 U6149 ( .A1(n10107), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n4871) );
  INV_X1 U6150 ( .A(n10107), .ZN(n6337) );
  INV_X1 U6151 ( .A(n9023), .ZN(n6352) );
  INV_X1 U6152 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6004) );
  OR2_X1 U6153 ( .A1(n9295), .A2(n9293), .ZN(n4872) );
  AND2_X1 U6154 ( .A1(n8250), .A2(n8249), .ZN(n4873) );
  OR2_X1 U6155 ( .A1(n9276), .A2(n9279), .ZN(n4874) );
  OR2_X1 U6156 ( .A1(n9674), .A2(n9284), .ZN(n4875) );
  OR2_X1 U6157 ( .A1(n9493), .A2(n9286), .ZN(n4876) );
  NOR2_X1 U6158 ( .A1(n8707), .A2(n8700), .ZN(n4877) );
  AND2_X1 U6159 ( .A1(n6253), .A2(n10032), .ZN(n4878) );
  INV_X1 U6160 ( .A(n7947), .ZN(n7959) );
  INV_X1 U6161 ( .A(n9913), .ZN(n9956) );
  OR2_X1 U6162 ( .A1(n7222), .A2(n9180), .ZN(n4879) );
  INV_X1 U6163 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4891) );
  AND2_X1 U6164 ( .A1(n5257), .A2(n9124), .ZN(n4880) );
  AND2_X1 U6165 ( .A1(n8383), .A2(n8331), .ZN(n4881) );
  AND2_X1 U6166 ( .A1(n5734), .A2(n5735), .ZN(n4882) );
  AND2_X1 U6167 ( .A1(n8226), .A2(n8216), .ZN(n4883) );
  INV_X1 U6168 ( .A(n8603), .ZN(n8601) );
  OR2_X1 U6169 ( .A1(n8203), .A2(n8223), .ZN(n4884) );
  AND3_X1 U6170 ( .A1(n5704), .A2(n9158), .A3(n5703), .ZN(n4885) );
  AND2_X1 U6171 ( .A1(n9493), .A2(n9286), .ZN(n4886) );
  INV_X1 U6172 ( .A(n7724), .ZN(n9395) );
  OR2_X1 U6173 ( .A1(n7526), .A2(n8445), .ZN(n4887) );
  INV_X1 U6174 ( .A(n7562), .ZN(n6083) );
  NOR2_X1 U6175 ( .A1(n5560), .A2(n5541), .ZN(n4888) );
  AND2_X1 U6176 ( .A1(n5489), .A2(n5488), .ZN(n9293) );
  INV_X1 U6177 ( .A(n9184), .ZN(n6786) );
  INV_X1 U6178 ( .A(n9444), .ZN(n9295) );
  INV_X1 U6179 ( .A(n9978), .ZN(n9979) );
  AND2_X1 U6180 ( .A1(n6559), .A2(n6855), .ZN(n9971) );
  OR2_X1 U6181 ( .A1(n5708), .A2(n9798), .ZN(n4889) );
  INV_X1 U6182 ( .A(n5593), .ZN(n5125) );
  INV_X1 U6183 ( .A(n8223), .ZN(n8209) );
  AND2_X1 U6184 ( .A1(n8213), .A2(n8209), .ZN(n8210) );
  INV_X1 U6185 ( .A(n7964), .ZN(n7965) );
  AOI21_X1 U6186 ( .B1(n7794), .B2(n7942), .A(n7965), .ZN(n7966) );
  NAND2_X1 U6187 ( .A1(n5247), .A2(n9783), .ZN(n5250) );
  NAND2_X1 U6188 ( .A1(n8217), .A2(n4883), .ZN(n8218) );
  INV_X1 U6189 ( .A(n7278), .ZN(n7275) );
  INV_X1 U6190 ( .A(n5880), .ZN(n5881) );
  NOR2_X1 U6191 ( .A1(n4877), .A2(n4870), .ZN(n6287) );
  NAND2_X1 U6192 ( .A1(n4307), .A2(n4990), .ZN(n4991) );
  INV_X1 U6193 ( .A(n8279), .ZN(n8278) );
  XNOR2_X1 U6194 ( .A(n8467), .B(n5859), .ZN(n8460) );
  INV_X1 U6195 ( .A(n7896), .ZN(n6282) );
  AND2_X1 U6196 ( .A1(n5574), .A2(n5572), .ZN(n9111) );
  NOR2_X1 U6197 ( .A1(n9841), .A2(n9840), .ZN(n9839) );
  INV_X1 U6198 ( .A(n9182), .ZN(n6819) );
  INV_X1 U6199 ( .A(n9790), .ZN(n7181) );
  XNOR2_X1 U6200 ( .A(n9184), .B(n7038), .ZN(n8048) );
  NAND2_X1 U6201 ( .A1(n4910), .A2(SI_4_), .ZN(n4911) );
  AND2_X1 U6202 ( .A1(n6136), .A2(n8409), .ZN(n6138) );
  NAND2_X1 U6203 ( .A1(n6731), .A2(n6987), .ZN(n6739) );
  INV_X1 U6204 ( .A(n6161), .ZN(n6163) );
  NAND2_X1 U6205 ( .A1(n6041), .A2(n6040), .ZN(n6050) );
  INV_X1 U6206 ( .A(n6832), .ZN(n6951) );
  INV_X1 U6207 ( .A(n6205), .ZN(n6204) );
  INV_X1 U6208 ( .A(n6097), .ZN(n6096) );
  INV_X1 U6209 ( .A(n7288), .ZN(n6047) );
  NAND2_X1 U6210 ( .A1(n8592), .A2(n8737), .ZN(n8594) );
  OR2_X1 U6211 ( .A1(n9012), .A2(n8705), .ZN(n7905) );
  NAND2_X1 U6212 ( .A1(n7392), .A2(n7388), .ZN(n7488) );
  INV_X1 U6213 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5957) );
  INV_X1 U6214 ( .A(n5351), .ZN(n5019) );
  AND2_X1 U6215 ( .A1(n5052), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5021) );
  INV_X1 U6216 ( .A(n5127), .ZN(n5191) );
  AND2_X1 U6217 ( .A1(n9159), .A2(n9160), .ZN(n5623) );
  INV_X1 U6218 ( .A(n9334), .ZN(n7725) );
  NAND2_X1 U6219 ( .A1(n9295), .A2(n9293), .ZN(n9296) );
  AND2_X1 U6220 ( .A1(n9460), .A2(n9291), .ZN(n9292) );
  AND2_X1 U6221 ( .A1(n9529), .A2(n9281), .ZN(n9282) );
  NOR2_X1 U6222 ( .A1(n9790), .A2(n9178), .ZN(n7231) );
  OR2_X1 U6223 ( .A1(n7263), .A2(n9179), .ZN(n7172) );
  NAND2_X1 U6224 ( .A1(n5535), .A2(n5534), .ZN(n5553) );
  INV_X1 U6225 ( .A(n5319), .ZN(n4950) );
  NAND2_X1 U6226 ( .A1(n4931), .A2(n4930), .ZN(n4934) );
  NAND2_X1 U6227 ( .A1(n6138), .A2(n6137), .ZN(n6146) );
  AND2_X1 U6228 ( .A1(n6032), .A2(n6031), .ZN(n6041) );
  XNOR2_X1 U6229 ( .A(n6759), .B(n6766), .ZN(n6738) );
  INV_X1 U6230 ( .A(n6763), .ZN(n6764) );
  AOI21_X1 U6231 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n6654), .A(n8485), .ZN(
        n5862) );
  AND2_X1 U6232 ( .A1(n9991), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5903) );
  OR2_X1 U6233 ( .A1(n6215), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U6234 ( .A1(n6117), .A2(n6116), .ZN(n6135) );
  NOR2_X1 U6235 ( .A1(n6020), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U6236 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  AND2_X1 U6237 ( .A1(n7893), .A2(n7894), .ZN(n7892) );
  INV_X1 U6238 ( .A(n8447), .ZN(n7374) );
  NAND2_X1 U6239 ( .A1(n6318), .A2(n6317), .ZN(n6320) );
  NAND2_X1 U6240 ( .A1(n5758), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5769) );
  INV_X1 U6241 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5846) );
  AND2_X1 U6242 ( .A1(n9113), .A2(n5551), .ZN(n9049) );
  INV_X1 U6243 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6900) );
  NOR2_X1 U6244 ( .A1(n5257), .A2(n9124), .ZN(n5278) );
  AND2_X1 U6245 ( .A1(n9774), .A2(n5317), .ZN(n7400) );
  AND2_X1 U6246 ( .A1(n9708), .A2(n9709), .ZN(n9710) );
  INV_X1 U6247 ( .A(n9316), .ZN(n9332) );
  AND2_X1 U6248 ( .A1(n8182), .A2(n8181), .ZN(n9435) );
  NAND2_X1 U6249 ( .A1(n9483), .A2(n8047), .ZN(n9503) );
  INV_X1 U6250 ( .A(n8110), .ZN(n9966) );
  NOR2_X1 U6251 ( .A1(n7236), .A2(n7235), .ZN(n7446) );
  INV_X1 U6252 ( .A(n7182), .ZN(n7184) );
  NOR2_X1 U6253 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5003) );
  NAND2_X1 U6254 ( .A1(n5046), .A2(n5045), .ZN(n5048) );
  INV_X1 U6255 ( .A(n9746), .ZN(n8434) );
  OR2_X1 U6256 ( .A1(n7975), .A2(n7974), .ZN(n7976) );
  AND2_X1 U6257 ( .A1(n6199), .A2(n6198), .ZN(n8287) );
  AND4_X1 U6258 ( .A1(n6082), .A2(n6081), .A3(n6080), .A4(n6079), .ZN(n7575)
         );
  NOR2_X1 U6259 ( .A1(n5890), .A2(n8457), .ZN(n8477) );
  NAND2_X1 U6260 ( .A1(n8553), .A2(n7803), .ZN(n5953) );
  NAND2_X1 U6261 ( .A1(n8822), .A2(n10107), .ZN(n8771) );
  NAND2_X1 U6262 ( .A1(n5303), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5351) );
  AND4_X1 U6263 ( .A1(n5670), .A2(n5669), .A3(n5668), .A4(n5667), .ZN(n7996)
         );
  AND4_X1 U6264 ( .A1(n5398), .A2(n5397), .A3(n5396), .A4(n5395), .ZN(n9279)
         );
  OR2_X1 U6265 ( .A1(n9891), .A2(n9890), .ZN(n9900) );
  XNOR2_X1 U6266 ( .A(n9352), .B(n9351), .ZN(n9559) );
  NOR2_X1 U6267 ( .A1(n5002), .A2(n5003), .ZN(n5004) );
  XNOR2_X1 U6268 ( .A(n4909), .B(SI_4_), .ZN(n5145) );
  AND2_X1 U6269 ( .A1(n6436), .A2(n6435), .ZN(n8391) );
  INV_X1 U6270 ( .A(n8423), .ZN(n8617) );
  INV_X1 U6271 ( .A(n6926), .ZN(n8456) );
  OAI21_X1 U6272 ( .B1(n5954), .B2(n6844), .A(n5953), .ZN(n5955) );
  INV_X1 U6273 ( .A(n6335), .ZN(n6336) );
  INV_X1 U6274 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10085) );
  AND2_X1 U6275 ( .A1(n6348), .A2(n6347), .ZN(n10078) );
  INV_X1 U6276 ( .A(n6585), .ZN(n6384) );
  INV_X1 U6277 ( .A(n9579), .ZN(n9407) );
  INV_X1 U6278 ( .A(n7523), .ZN(n7519) );
  INV_X1 U6279 ( .A(n9158), .ZN(n9792) );
  INV_X1 U6280 ( .A(n9293), .ZN(n9294) );
  AND3_X1 U6281 ( .A1(n5058), .A2(n5057), .A3(n5056), .ZN(n9284) );
  INV_X1 U6282 ( .A(n7580), .ZN(n9175) );
  OR2_X1 U6283 ( .A1(n9938), .A2(n7064), .ZN(n9530) );
  AND2_X1 U6284 ( .A1(n7065), .A2(n9531), .ZN(n9928) );
  INV_X1 U6285 ( .A(n9381), .ZN(n9649) );
  INV_X1 U6286 ( .A(n9424), .ZN(n9655) );
  INV_X1 U6287 ( .A(n6560), .ZN(n9961) );
  NAND2_X1 U6288 ( .A1(n5005), .A2(n5004), .ZN(n7541) );
  XNOR2_X1 U6289 ( .A(n4896), .B(SI_1_), .ZN(n5090) );
  INV_X1 U6290 ( .A(n5090), .ZN(n4895) );
  NAND3_X1 U6291 ( .A1(n4902), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n4894) );
  AND2_X1 U6292 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4893) );
  NAND2_X1 U6293 ( .A1(n4892), .A2(n4893), .ZN(n5977) );
  NAND2_X1 U6294 ( .A1(n4894), .A2(n5977), .ZN(n5089) );
  NAND2_X1 U6295 ( .A1(n4895), .A2(n5089), .ZN(n4898) );
  NAND2_X1 U6296 ( .A1(n4896), .A2(SI_1_), .ZN(n4897) );
  NAND2_X1 U6297 ( .A1(n4898), .A2(n4897), .ZN(n5100) );
  INV_X1 U6298 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6363) );
  INV_X1 U6299 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6378) );
  MUX2_X1 U6300 ( .A(n6363), .B(n6378), .S(n4902), .Z(n4899) );
  XNOR2_X1 U6301 ( .A(n4899), .B(SI_2_), .ZN(n5099) );
  INV_X1 U6302 ( .A(n4899), .ZN(n4900) );
  NAND2_X1 U6303 ( .A1(n4900), .A2(SI_2_), .ZN(n4901) );
  INV_X1 U6304 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6379) );
  INV_X1 U6305 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6356) );
  INV_X1 U6306 ( .A(n4905), .ZN(n4906) );
  NAND2_X1 U6307 ( .A1(n4906), .A2(SI_3_), .ZN(n4907) );
  INV_X1 U6308 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6387) );
  INV_X1 U6309 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4908) );
  MUX2_X1 U6310 ( .A(n6387), .B(n4908), .S(n6362), .Z(n4909) );
  NAND2_X1 U6311 ( .A1(n5144), .A2(n5145), .ZN(n4912) );
  INV_X1 U6312 ( .A(n4909), .ZN(n4910) );
  MUX2_X1 U6313 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6362), .Z(n4914) );
  NAND2_X1 U6314 ( .A1(n4914), .A2(SI_5_), .ZN(n4915) );
  MUX2_X1 U6315 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6362), .Z(n4917) );
  NAND2_X1 U6316 ( .A1(n4917), .A2(SI_6_), .ZN(n4918) );
  MUX2_X1 U6317 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6362), .Z(n4920) );
  INV_X1 U6318 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n4922) );
  INV_X1 U6319 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n4921) );
  MUX2_X1 U6320 ( .A(n4922), .B(n4921), .S(n6362), .Z(n4924) );
  INV_X1 U6321 ( .A(SI_8_), .ZN(n4923) );
  INV_X1 U6322 ( .A(n4924), .ZN(n4925) );
  NAND2_X1 U6323 ( .A1(n4925), .A2(SI_8_), .ZN(n4926) );
  INV_X1 U6324 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n4929) );
  INV_X1 U6325 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4928) );
  MUX2_X1 U6326 ( .A(n4929), .B(n4928), .S(n6362), .Z(n4931) );
  INV_X1 U6327 ( .A(SI_9_), .ZN(n4930) );
  INV_X1 U6328 ( .A(n4931), .ZN(n4932) );
  NAND2_X1 U6329 ( .A1(n4932), .A2(SI_9_), .ZN(n4933) );
  INV_X1 U6330 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n8957) );
  INV_X1 U6331 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n4935) );
  MUX2_X1 U6332 ( .A(n8957), .B(n4935), .S(n6362), .Z(n4940) );
  INV_X1 U6333 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6443) );
  INV_X1 U6334 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6442) );
  MUX2_X1 U6335 ( .A(n6443), .B(n6442), .S(n6362), .Z(n4937) );
  INV_X1 U6336 ( .A(SI_11_), .ZN(n4936) );
  INV_X1 U6337 ( .A(n4937), .ZN(n4938) );
  NAND2_X1 U6338 ( .A1(n4938), .A2(SI_11_), .ZN(n4939) );
  NAND2_X1 U6339 ( .A1(n4944), .A2(n4939), .ZN(n5295) );
  INV_X1 U6340 ( .A(n5295), .ZN(n4942) );
  INV_X1 U6341 ( .A(n4940), .ZN(n4941) );
  NAND2_X1 U6342 ( .A1(n4941), .A2(SI_10_), .ZN(n5293) );
  INV_X1 U6343 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6536) );
  INV_X1 U6344 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n4946) );
  MUX2_X1 U6345 ( .A(n6536), .B(n4946), .S(n6362), .Z(n4947) );
  INV_X1 U6346 ( .A(n4947), .ZN(n4948) );
  NAND2_X1 U6347 ( .A1(n4948), .A2(SI_12_), .ZN(n4949) );
  MUX2_X1 U6348 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6362), .Z(n4952) );
  XNOR2_X1 U6349 ( .A(n4952), .B(SI_13_), .ZN(n5344) );
  INV_X1 U6350 ( .A(n5344), .ZN(n4951) );
  NAND2_X1 U6351 ( .A1(n4952), .A2(SI_13_), .ZN(n4953) );
  INV_X1 U6352 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6653) );
  INV_X1 U6353 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6656) );
  MUX2_X1 U6354 ( .A(n6653), .B(n6656), .S(n6362), .Z(n4955) );
  INV_X1 U6355 ( .A(SI_14_), .ZN(n4954) );
  NAND2_X1 U6356 ( .A1(n4955), .A2(n4954), .ZN(n4958) );
  INV_X1 U6357 ( .A(n4955), .ZN(n4956) );
  NAND2_X1 U6358 ( .A1(n4956), .A2(SI_14_), .ZN(n4957) );
  NAND2_X1 U6359 ( .A1(n4958), .A2(n4957), .ZN(n5365) );
  INV_X1 U6360 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6709) );
  INV_X1 U6361 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n4959) );
  MUX2_X1 U6362 ( .A(n6709), .B(n4959), .S(n6362), .Z(n4960) );
  XNOR2_X1 U6363 ( .A(n4960), .B(SI_15_), .ZN(n5385) );
  INV_X1 U6364 ( .A(n5385), .ZN(n4963) );
  INV_X1 U6365 ( .A(n4960), .ZN(n4961) );
  NAND2_X1 U6366 ( .A1(n4961), .A2(SI_15_), .ZN(n4962) );
  INV_X1 U6367 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6883) );
  INV_X1 U6368 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6882) );
  MUX2_X1 U6369 ( .A(n6883), .B(n6882), .S(n6362), .Z(n4965) );
  INV_X1 U6370 ( .A(SI_16_), .ZN(n4964) );
  NAND2_X1 U6371 ( .A1(n4965), .A2(n4964), .ZN(n4968) );
  INV_X1 U6372 ( .A(n4965), .ZN(n4966) );
  NAND2_X1 U6373 ( .A1(n4966), .A2(SI_16_), .ZN(n4967) );
  NAND2_X1 U6374 ( .A1(n4968), .A2(n4967), .ZN(n5405) );
  INV_X1 U6375 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6963) );
  INV_X1 U6376 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6962) );
  MUX2_X1 U6377 ( .A(n6963), .B(n6962), .S(n6362), .Z(n4970) );
  INV_X1 U6378 ( .A(SI_17_), .ZN(n4969) );
  NAND2_X1 U6379 ( .A1(n4970), .A2(n4969), .ZN(n4973) );
  INV_X1 U6380 ( .A(n4970), .ZN(n4971) );
  NAND2_X1 U6381 ( .A1(n4971), .A2(SI_17_), .ZN(n4972) );
  INV_X1 U6382 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n4974) );
  INV_X1 U6383 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7010) );
  MUX2_X1 U6384 ( .A(n4974), .B(n7010), .S(n6362), .Z(n5428) );
  XNOR2_X1 U6385 ( .A(n5428), .B(SI_18_), .ZN(n5427) );
  XNOR2_X1 U6386 ( .A(n5432), .B(n5427), .ZN(n6966) );
  NOR2_X2 U6387 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5086) );
  AND2_X2 U6388 ( .A1(n5086), .A2(n4393), .ZN(n5096) );
  NOR2_X1 U6389 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4978) );
  NOR2_X1 U6390 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n4984) );
  NOR2_X1 U6391 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4983) );
  NOR2_X1 U6392 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4982) );
  INV_X1 U6393 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4988) );
  INV_X1 U6394 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4987) );
  NAND2_X1 U6395 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n4989) );
  NAND2_X1 U6396 ( .A1(n6966), .A2(n5346), .ZN(n4994) );
  INV_X1 U6397 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4990) );
  INV_X1 U6398 ( .A(n4997), .ZN(n4992) );
  INV_X1 U6399 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4995) );
  XNOR2_X1 U6400 ( .A(n5040), .B(P1_IR_REG_18__SCAN_IN), .ZN(n7709) );
  AOI22_X1 U6401 ( .A1(n5191), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6364), .B2(
        n7709), .ZN(n4993) );
  INV_X1 U6402 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5039) );
  AND3_X1 U6403 ( .A1(n5039), .A2(n4995), .A3(n5041), .ZN(n4996) );
  INV_X1 U6404 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4998) );
  INV_X1 U6405 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5010) );
  NAND2_X1 U6406 ( .A1(n5015), .A2(n5010), .ZN(n5035) );
  INV_X1 U6407 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5036) );
  INV_X1 U6408 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5695) );
  NAND2_X1 U6409 ( .A1(n5036), .A2(n5695), .ZN(n4999) );
  OAI21_X1 U6410 ( .B1(n5035), .B2(n4999), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5001) );
  INV_X1 U6411 ( .A(n5002), .ZN(n5007) );
  XNOR2_X1 U6412 ( .A(n5006), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U6413 ( .A1(n5679), .A2(n7568), .ZN(n5009) );
  INV_X1 U6414 ( .A(n8049), .ZN(n5697) );
  INV_X1 U6415 ( .A(n5012), .ZN(n5013) );
  NAND2_X1 U6416 ( .A1(n5013), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5014) );
  MUX2_X1 U6417 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5014), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5017) );
  INV_X1 U6418 ( .A(n5015), .ZN(n5016) );
  AND2_X2 U6419 ( .A1(n5697), .A2(n7254), .ZN(n6561) );
  NAND2_X4 U6420 ( .A1(n5708), .A2(n6561), .ZN(n5593) );
  NAND2_X1 U6421 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5180) );
  NAND2_X1 U6422 ( .A1(n5182), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5211) );
  INV_X1 U6423 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5210) );
  INV_X1 U6424 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5235) );
  INV_X1 U6425 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9124) );
  NAND2_X1 U6426 ( .A1(n5278), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5305) );
  INV_X1 U6427 ( .A(n5305), .ZN(n5018) );
  NAND2_X1 U6428 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n5020) );
  INV_X1 U6429 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U6430 ( .A1(n5021), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5441) );
  INV_X1 U6431 ( .A(n5021), .ZN(n5055) );
  INV_X1 U6432 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5022) );
  NAND2_X1 U6433 ( .A1(n5055), .A2(n5022), .ZN(n5023) );
  NAND2_X1 U6434 ( .A1(n5441), .A2(n5023), .ZN(n9494) );
  NAND2_X1 U6435 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5024) );
  NAND2_X1 U6436 ( .A1(n5025), .A2(n5024), .ZN(n5026) );
  XNOR2_X2 U6437 ( .A(n5026), .B(P1_IR_REG_29__SCAN_IN), .ZN(n7739) );
  INV_X1 U6438 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6439 ( .A1(n5028), .A2(n5027), .ZN(n9689) );
  AND2_X4 U6440 ( .A1(n5030), .A2(n5031), .ZN(n5666) );
  INV_X1 U6441 ( .A(n5666), .ZN(n5511) );
  OR2_X1 U6442 ( .A1(n9494), .A2(n5511), .ZN(n5034) );
  INV_X1 U6443 ( .A(n5031), .ZN(n7663) );
  AND2_X2 U6444 ( .A1(n5030), .A2(n7663), .ZN(n5119) );
  AND2_X2 U6445 ( .A1(n7663), .A2(n7739), .ZN(n5120) );
  AOI22_X1 U6446 ( .A1(n5213), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6404), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U6447 ( .A1(n7985), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5032) );
  AND3_X1 U6448 ( .A1(n5034), .A2(n5033), .A3(n5032), .ZN(n9287) );
  NAND2_X1 U6449 ( .A1(n5035), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6450 ( .A1(n5037), .A2(n5036), .ZN(n5694) );
  NAND2_X2 U6451 ( .A1(n5694), .A2(n5038), .ZN(n5698) );
  INV_X2 U6452 ( .A(n5698), .ZN(n8237) );
  INV_X1 U6453 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5041) );
  NAND2_X1 U6454 ( .A1(n5043), .A2(n7254), .ZN(n8235) );
  NAND2_X1 U6455 ( .A1(n6561), .A2(n5437), .ZN(n7083) );
  OAI211_X2 U6456 ( .C1(n8237), .C2(n8235), .A(n5708), .B(n7083), .ZN(n5113)
         );
  BUF_X4 U6457 ( .A(n5113), .Z(n5676) );
  NOR2_X1 U6458 ( .A1(n9287), .A2(n5676), .ZN(n5044) );
  AOI21_X1 U6459 ( .B1(n9493), .B2(n5671), .A(n5044), .ZN(n9063) );
  OR2_X1 U6460 ( .A1(n5046), .A2(n5045), .ZN(n5047) );
  NAND2_X1 U6461 ( .A1(n5048), .A2(n5047), .ZN(n6961) );
  NAND2_X1 U6462 ( .A1(n6961), .A2(n5346), .ZN(n5051) );
  XNOR2_X1 U6463 ( .A(n5049), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9882) );
  AOI22_X1 U6464 ( .A1(n5191), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6364), .B2(
        n9882), .ZN(n5050) );
  INV_X1 U6465 ( .A(n5052), .ZN(n5412) );
  INV_X1 U6466 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U6467 ( .A1(n5412), .A2(n5053), .ZN(n5054) );
  AND2_X1 U6468 ( .A1(n5055), .A2(n5054), .ZN(n9513) );
  NAND2_X1 U6469 ( .A1(n9513), .A2(n5666), .ZN(n5058) );
  AOI22_X1 U6470 ( .A1(n5213), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n6404), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U6471 ( .A1(n5105), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5056) );
  NOR2_X1 U6472 ( .A1(n9284), .A2(n5676), .ZN(n5059) );
  AOI21_X1 U6473 ( .B1(n9512), .B2(n5671), .A(n5059), .ZN(n5422) );
  INV_X1 U6474 ( .A(n5422), .ZN(n5425) );
  AND2_X2 U6475 ( .A1(n8237), .A2(n5043), .ZN(n7060) );
  NAND2_X1 U6476 ( .A1(n9512), .A2(n5659), .ZN(n5063) );
  OR2_X1 U6477 ( .A1(n9284), .A2(n5593), .ZN(n5062) );
  NAND2_X1 U6478 ( .A1(n5063), .A2(n5062), .ZN(n5064) );
  XNOR2_X1 U6479 ( .A(n5064), .B(n4287), .ZN(n5423) );
  INV_X1 U6480 ( .A(n5423), .ZN(n5424) );
  NAND2_X1 U6481 ( .A1(n5666), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U6482 ( .A1(n5119), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U6483 ( .A1(n5120), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U6484 ( .A1(n5105), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6485 ( .A1(n9186), .A2(n5125), .ZN(n5074) );
  INV_X1 U6486 ( .A(SI_0_), .ZN(n5070) );
  NOR2_X1 U6487 ( .A1(n4471), .A2(n5070), .ZN(n5072) );
  INV_X1 U6488 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5071) );
  XNOR2_X1 U6489 ( .A(n5072), .B(n5071), .ZN(n9696) );
  MUX2_X1 U6490 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9696), .S(n5128), .Z(n7066) );
  NAND2_X1 U6491 ( .A1(n5104), .A2(n7066), .ZN(n5073) );
  NAND2_X1 U6492 ( .A1(n5074), .A2(n5073), .ZN(n5079) );
  INV_X1 U6493 ( .A(n5079), .ZN(n5075) );
  INV_X1 U6494 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U6495 ( .A1(n5075), .A2(n4889), .ZN(n6467) );
  INV_X1 U6496 ( .A(n5708), .ZN(n6355) );
  AOI22_X1 U6497 ( .A1(n5125), .A2(n7066), .B1(n6355), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5077) );
  OAI21_X1 U6498 ( .B1(n5076), .B2(n5676), .A(n5077), .ZN(n6466) );
  NAND2_X1 U6499 ( .A1(n6467), .A2(n6466), .ZN(n6465) );
  AND2_X1 U6500 ( .A1(n6465), .A2(n5080), .ZN(n6665) );
  NAND2_X1 U6501 ( .A1(n5666), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6502 ( .A1(n5105), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U6503 ( .A1(n5120), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6504 ( .A1(n5119), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5081) );
  AND4_X2 U6505 ( .A1(n5084), .A2(n5083), .A3(n5082), .A4(n5081), .ZN(n6541)
         );
  NAND2_X1 U6506 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5085) );
  MUX2_X1 U6507 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5085), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5088) );
  INV_X1 U6508 ( .A(n5086), .ZN(n5087) );
  XNOR2_X1 U6509 ( .A(n5090), .B(n5089), .ZN(n5967) );
  INV_X1 U6510 ( .A(n5967), .ZN(n6376) );
  OAI22_X1 U6511 ( .A1(n6541), .A2(n5676), .B1(n7025), .B2(n5593), .ZN(n5092)
         );
  NAND2_X1 U6512 ( .A1(n6665), .A2(n6664), .ZN(n5095) );
  INV_X1 U6513 ( .A(n5092), .ZN(n5093) );
  NAND2_X1 U6514 ( .A1(n5095), .A2(n5094), .ZN(n6539) );
  INV_X1 U6515 ( .A(n5096), .ZN(n5097) );
  NAND2_X1 U6516 ( .A1(n5098), .A2(n5097), .ZN(n6507) );
  XNOR2_X1 U6517 ( .A(n5100), .B(n5099), .ZN(n6377) );
  OR2_X1 U6518 ( .A1(n5101), .A2(n6377), .ZN(n5103) );
  OAI211_X2 U6519 ( .C1(n5128), .C2(n6507), .A(n5103), .B(n5102), .ZN(n7038)
         );
  NAND2_X1 U6520 ( .A1(n5104), .A2(n7038), .ZN(n5111) );
  NAND2_X1 U6521 ( .A1(n5666), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U6522 ( .A1(n5119), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6523 ( .A1(n5120), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6524 ( .A1(n5105), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6525 ( .A1(n9184), .A2(n5125), .ZN(n5110) );
  NAND2_X1 U6526 ( .A1(n5111), .A2(n5110), .ZN(n5112) );
  INV_X1 U6527 ( .A(n5113), .ZN(n5415) );
  AOI22_X1 U6528 ( .A1(n9184), .A2(n5415), .B1(n5125), .B2(n7038), .ZN(n5115)
         );
  XNOR2_X1 U6529 ( .A(n5114), .B(n5115), .ZN(n6540) );
  NAND2_X1 U6530 ( .A1(n6539), .A2(n6540), .ZN(n5118) );
  INV_X1 U6531 ( .A(n5114), .ZN(n5116) );
  NAND2_X1 U6532 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  NAND2_X1 U6533 ( .A1(n5118), .A2(n5117), .ZN(n6657) );
  INV_X1 U6534 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U6535 ( .A1(n5666), .A2(n9926), .ZN(n5124) );
  NAND2_X1 U6536 ( .A1(n5105), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6537 ( .A1(n5119), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6538 ( .A1(n5120), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5121) );
  NAND4_X1 U6539 ( .A1(n5124), .A2(n5123), .A3(n5122), .A4(n5121), .ZN(n9183)
         );
  NAND2_X1 U6540 ( .A1(n9183), .A2(n5125), .ZN(n5132) );
  OR2_X1 U6541 ( .A1(n5127), .A2(n6356), .ZN(n5130) );
  OR2_X1 U6542 ( .A1(n5096), .A2(n9688), .ZN(n5141) );
  XNOR2_X1 U6543 ( .A(n5141), .B(n4975), .ZN(n6489) );
  OR2_X1 U6544 ( .A1(n5128), .A2(n6489), .ZN(n5129) );
  NAND2_X1 U6545 ( .A1(n5132), .A2(n4328), .ZN(n5133) );
  NAND2_X1 U6546 ( .A1(n9183), .A2(n5415), .ZN(n5135) );
  NAND2_X1 U6547 ( .A1(n9924), .A2(n5671), .ZN(n5134) );
  NAND2_X1 U6548 ( .A1(n5135), .A2(n5134), .ZN(n5136) );
  XNOR2_X1 U6549 ( .A(n5138), .B(n5136), .ZN(n6658) );
  NAND2_X1 U6550 ( .A1(n6657), .A2(n6658), .ZN(n5140) );
  INV_X1 U6551 ( .A(n5136), .ZN(n5137) );
  NAND2_X1 U6552 ( .A1(n5138), .A2(n5137), .ZN(n5139) );
  NAND2_X1 U6553 ( .A1(n5140), .A2(n5139), .ZN(n6644) );
  INV_X1 U6554 ( .A(n6644), .ZN(n5158) );
  NAND2_X1 U6555 ( .A1(n5141), .A2(n4975), .ZN(n5142) );
  NAND2_X1 U6556 ( .A1(n5142), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5143) );
  XNOR2_X1 U6557 ( .A(n5143), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7210) );
  AOI22_X1 U6558 ( .A1(n5191), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6364), .B2(
        n7210), .ZN(n5147) );
  XNOR2_X1 U6559 ( .A(n5144), .B(n5145), .ZN(n6388) );
  OR2_X1 U6560 ( .A1(n6388), .A2(n5101), .ZN(n5146) );
  NAND2_X1 U6561 ( .A1(n7303), .A2(n5659), .ZN(n5155) );
  NAND2_X1 U6562 ( .A1(n5105), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5153) );
  OAI21_X1 U6563 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5180), .ZN(n6651) );
  INV_X1 U6564 ( .A(n6651), .ZN(n7302) );
  NAND2_X1 U6565 ( .A1(n5666), .A2(n7302), .ZN(n5152) );
  NAND2_X1 U6566 ( .A1(n6404), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U6567 ( .A1(n5213), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5150) );
  NAND4_X1 U6568 ( .A1(n5153), .A2(n5152), .A3(n5151), .A4(n5150), .ZN(n9182)
         );
  NAND2_X1 U6569 ( .A1(n9182), .A2(n5671), .ZN(n5154) );
  NAND2_X1 U6570 ( .A1(n5155), .A2(n5154), .ZN(n5156) );
  AOI22_X1 U6571 ( .A1(n7303), .A2(n5671), .B1(n9182), .B2(n5415), .ZN(n5160)
         );
  INV_X1 U6572 ( .A(n5159), .ZN(n5162) );
  INV_X1 U6573 ( .A(n5160), .ZN(n5161) );
  NAND2_X1 U6574 ( .A1(n5162), .A2(n5161), .ZN(n5163) );
  XNOR2_X1 U6575 ( .A(n5164), .B(n5165), .ZN(n6371) );
  INV_X2 U6576 ( .A(n5101), .ZN(n5346) );
  NAND2_X1 U6577 ( .A1(n6371), .A2(n5346), .ZN(n5169) );
  NOR2_X1 U6578 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5166) );
  NAND2_X1 U6579 ( .A1(n5096), .A2(n5166), .ZN(n5189) );
  NAND2_X1 U6580 ( .A1(n5207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5167) );
  XNOR2_X1 U6581 ( .A(n5167), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9232) );
  AOI22_X1 U6582 ( .A1(n5191), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6364), .B2(
        n9232), .ZN(n5168) );
  NAND2_X1 U6583 ( .A1(n5169), .A2(n5168), .ZN(n7222) );
  NAND2_X1 U6584 ( .A1(n7222), .A2(n5634), .ZN(n5176) );
  NAND2_X1 U6585 ( .A1(n5105), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5174) );
  OR2_X1 U6586 ( .A1(n5182), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5170) );
  AND2_X1 U6587 ( .A1(n5211), .A2(n5170), .ZN(n7223) );
  NAND2_X1 U6588 ( .A1(n5666), .A2(n7223), .ZN(n5173) );
  NAND2_X1 U6589 ( .A1(n6404), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6590 ( .A1(n5213), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6591 ( .A1(n9180), .A2(n5671), .ZN(n5175) );
  NAND2_X1 U6592 ( .A1(n5176), .A2(n5175), .ZN(n5177) );
  XNOR2_X1 U6593 ( .A(n5177), .B(n4287), .ZN(n6973) );
  NAND2_X1 U6594 ( .A1(n7222), .A2(n5671), .ZN(n5179) );
  NAND2_X1 U6595 ( .A1(n9180), .A2(n5415), .ZN(n5178) );
  AND2_X1 U6596 ( .A1(n5179), .A2(n5178), .ZN(n6972) );
  NAND2_X1 U6597 ( .A1(n7985), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5186) );
  AND2_X1 U6598 ( .A1(n5180), .A2(n6900), .ZN(n5181) );
  NOR2_X1 U6599 ( .A1(n5182), .A2(n5181), .ZN(n6894) );
  NAND2_X1 U6600 ( .A1(n5666), .A2(n6894), .ZN(n5185) );
  NAND2_X1 U6601 ( .A1(n6404), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6602 ( .A1(n5213), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5183) );
  INV_X1 U6603 ( .A(n6976), .ZN(n9181) );
  NAND2_X1 U6604 ( .A1(n9181), .A2(n5415), .ZN(n5195) );
  XNOR2_X1 U6605 ( .A(n5187), .B(n5188), .ZN(n6369) );
  NAND2_X1 U6606 ( .A1(n6369), .A2(n5346), .ZN(n5193) );
  NAND2_X1 U6607 ( .A1(n5189), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5190) );
  XNOR2_X1 U6608 ( .A(n5190), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9218) );
  AOI22_X1 U6609 ( .A1(n5191), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6364), .B2(
        n9218), .ZN(n5192) );
  NAND2_X1 U6610 ( .A1(n7012), .A2(n5671), .ZN(n5194) );
  AND2_X1 U6611 ( .A1(n5195), .A2(n5194), .ZN(n6898) );
  NAND2_X1 U6612 ( .A1(n7012), .A2(n5634), .ZN(n5196) );
  OAI21_X1 U6613 ( .B1(n6976), .B2(n5593), .A(n5196), .ZN(n5197) );
  XNOR2_X1 U6614 ( .A(n5197), .B(n4287), .ZN(n6896) );
  AOI22_X1 U6615 ( .A1(n6973), .A2(n6972), .B1(n6898), .B2(n6896), .ZN(n5198)
         );
  INV_X1 U6616 ( .A(n6973), .ZN(n5203) );
  INV_X1 U6617 ( .A(n6896), .ZN(n6971) );
  NAND2_X1 U6618 ( .A1(n5199), .A2(n6972), .ZN(n5202) );
  INV_X1 U6619 ( .A(n5199), .ZN(n5201) );
  INV_X1 U6620 ( .A(n6972), .ZN(n5200) );
  AOI22_X1 U6621 ( .A1(n5203), .A2(n5202), .B1(n5201), .B2(n5200), .ZN(n5204)
         );
  XNOR2_X1 U6622 ( .A(n5205), .B(n5206), .ZN(n6394) );
  NAND2_X1 U6623 ( .A1(n6394), .A2(n5346), .ZN(n5209) );
  NOR2_X1 U6624 ( .A1(n5207), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5253) );
  OR2_X1 U6625 ( .A1(n5253), .A2(n9688), .ZN(n5230) );
  XNOR2_X1 U6626 ( .A(n5230), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9717) );
  AOI22_X1 U6627 ( .A1(n5191), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6364), .B2(
        n9717), .ZN(n5208) );
  NAND2_X1 U6628 ( .A1(n7263), .A2(n5659), .ZN(n5219) );
  NAND2_X1 U6629 ( .A1(n5211), .A2(n5210), .ZN(n5212) );
  AND2_X1 U6630 ( .A1(n5236), .A2(n5212), .ZN(n7101) );
  NAND2_X1 U6631 ( .A1(n5666), .A2(n7101), .ZN(n5217) );
  NAND2_X1 U6632 ( .A1(n5105), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6633 ( .A1(n6404), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U6634 ( .A1(n5213), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5214) );
  INV_X1 U6635 ( .A(n7093), .ZN(n9179) );
  NAND2_X1 U6636 ( .A1(n9179), .A2(n5671), .ZN(n5218) );
  NAND2_X1 U6637 ( .A1(n5219), .A2(n5218), .ZN(n5220) );
  XNOR2_X1 U6638 ( .A(n5220), .B(n4287), .ZN(n5222) );
  NOR2_X1 U6639 ( .A1(n7093), .A2(n5676), .ZN(n5221) );
  AOI21_X1 U6640 ( .B1(n7263), .B2(n5671), .A(n5221), .ZN(n5223) );
  NAND2_X1 U6641 ( .A1(n5222), .A2(n5223), .ZN(n9115) );
  INV_X1 U6642 ( .A(n5222), .ZN(n5225) );
  INV_X1 U6643 ( .A(n5223), .ZN(n5224) );
  NAND2_X1 U6644 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  NAND2_X1 U6645 ( .A1(n9115), .A2(n5226), .ZN(n6876) );
  XNOR2_X1 U6646 ( .A(n5228), .B(n5227), .ZN(n6399) );
  NAND2_X1 U6647 ( .A1(n6399), .A2(n5346), .ZN(n5234) );
  INV_X1 U6648 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6649 ( .A1(n5230), .A2(n5229), .ZN(n5231) );
  NAND2_X1 U6650 ( .A1(n5231), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5232) );
  XNOR2_X1 U6651 ( .A(n5232), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9729) );
  AOI22_X1 U6652 ( .A1(n5191), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6364), .B2(
        n9729), .ZN(n5233) );
  NAND2_X1 U6653 ( .A1(n9790), .A2(n5634), .ZN(n5243) );
  NAND2_X1 U6654 ( .A1(n5236), .A2(n5235), .ZN(n5237) );
  NAND2_X1 U6655 ( .A1(n5257), .A2(n5237), .ZN(n9796) );
  INV_X1 U6656 ( .A(n9796), .ZN(n7185) );
  NAND2_X1 U6657 ( .A1(n5666), .A2(n7185), .ZN(n5241) );
  NAND2_X1 U6658 ( .A1(n7985), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6659 ( .A1(n6404), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6660 ( .A1(n5213), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6661 ( .A1(n9178), .A2(n5671), .ZN(n5242) );
  NAND2_X1 U6662 ( .A1(n5243), .A2(n5242), .ZN(n5244) );
  XNOR2_X1 U6663 ( .A(n5244), .B(n5616), .ZN(n5247) );
  NAND2_X1 U6664 ( .A1(n9790), .A2(n5671), .ZN(n5246) );
  NAND2_X1 U6665 ( .A1(n9178), .A2(n5415), .ZN(n5245) );
  NAND2_X1 U6666 ( .A1(n5246), .A2(n5245), .ZN(n9783) );
  INV_X1 U6667 ( .A(n9115), .ZN(n5249) );
  INV_X1 U6668 ( .A(n5247), .ZN(n9118) );
  INV_X1 U6669 ( .A(n9783), .ZN(n5248) );
  AOI22_X1 U6670 ( .A1(n5250), .A2(n5249), .B1(n9118), .B2(n5248), .ZN(n5267)
         );
  XNOR2_X1 U6671 ( .A(n5251), .B(n4302), .ZN(n6409) );
  NAND2_X1 U6672 ( .A1(n6409), .A2(n5346), .ZN(n5256) );
  NAND2_X1 U6673 ( .A1(n5253), .A2(n5252), .ZN(n5274) );
  NAND2_X1 U6674 ( .A1(n5274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5254) );
  XNOR2_X1 U6675 ( .A(n5254), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9248) );
  AOI22_X1 U6676 ( .A1(n5191), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6364), .B2(
        n9248), .ZN(n5255) );
  NAND2_X1 U6677 ( .A1(n5265), .A2(n5659), .ZN(n5263) );
  NAND2_X1 U6678 ( .A1(n5105), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5261) );
  NOR2_X1 U6679 ( .A1(n5278), .A2(n4880), .ZN(n9127) );
  NAND2_X1 U6680 ( .A1(n5666), .A2(n9127), .ZN(n5260) );
  NAND2_X1 U6681 ( .A1(n6404), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6682 ( .A1(n5213), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6683 ( .A1(n9760), .A2(n5671), .ZN(n5262) );
  NAND2_X1 U6684 ( .A1(n5263), .A2(n5262), .ZN(n5264) );
  NOR2_X1 U6685 ( .A1(n7234), .A2(n5676), .ZN(n5266) );
  AOI21_X1 U6686 ( .B1(n5265), .B2(n5671), .A(n5266), .ZN(n5269) );
  INV_X1 U6687 ( .A(n5268), .ZN(n5270) );
  OR2_X1 U6688 ( .A1(n5270), .A2(n5269), .ZN(n5271) );
  XNOR2_X1 U6689 ( .A(n5273), .B(n5272), .ZN(n6413) );
  NAND2_X1 U6690 ( .A1(n6413), .A2(n5346), .ZN(n5277) );
  OR2_X1 U6691 ( .A1(n5274), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6692 ( .A1(n5275), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5298) );
  XNOR2_X1 U6693 ( .A(n5298), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9705) );
  AOI22_X1 U6694 ( .A1(n5191), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6364), .B2(
        n9705), .ZN(n5276) );
  NAND2_X1 U6695 ( .A1(n9913), .A2(n5634), .ZN(n5287) );
  INV_X1 U6696 ( .A(n5278), .ZN(n5280) );
  INV_X1 U6697 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6698 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  NAND2_X1 U6699 ( .A1(n5305), .A2(n5281), .ZN(n9768) );
  INV_X1 U6700 ( .A(n9768), .ZN(n9912) );
  NAND2_X1 U6701 ( .A1(n5666), .A2(n9912), .ZN(n5285) );
  NAND2_X1 U6702 ( .A1(n7985), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6703 ( .A1(n6404), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6704 ( .A1(n5119), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5282) );
  INV_X1 U6705 ( .A(n7449), .ZN(n9177) );
  NAND2_X1 U6706 ( .A1(n9177), .A2(n5671), .ZN(n5286) );
  NAND2_X1 U6707 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  XNOR2_X1 U6708 ( .A(n5288), .B(n4287), .ZN(n5289) );
  OAI22_X1 U6709 ( .A1(n9956), .A2(n5593), .B1(n7449), .B2(n5676), .ZN(n9756)
         );
  NAND2_X1 U6710 ( .A1(n5294), .A2(n5293), .ZN(n5296) );
  XNOR2_X1 U6711 ( .A(n5296), .B(n5295), .ZN(n6441) );
  NAND2_X1 U6712 ( .A1(n6441), .A2(n5346), .ZN(n5302) );
  NAND2_X1 U6713 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  NAND2_X1 U6714 ( .A1(n5299), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5300) );
  XNOR2_X1 U6715 ( .A(n5300), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7215) );
  AOI22_X1 U6716 ( .A1(n5191), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6364), .B2(
        n7215), .ZN(n5301) );
  NAND2_X1 U6717 ( .A1(n7523), .A2(n5659), .ZN(n5312) );
  INV_X1 U6718 ( .A(n5303), .ZN(n5327) );
  INV_X1 U6719 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6720 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  AND2_X1 U6721 ( .A1(n5327), .A2(n5306), .ZN(n7481) );
  NAND2_X1 U6722 ( .A1(n5666), .A2(n7481), .ZN(n5310) );
  NAND2_X1 U6723 ( .A1(n7985), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6724 ( .A1(n6404), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U6725 ( .A1(n5119), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5307) );
  INV_X1 U6726 ( .A(n7450), .ZN(n9759) );
  NAND2_X1 U6727 ( .A1(n9759), .A2(n5671), .ZN(n5311) );
  NAND2_X1 U6728 ( .A1(n5312), .A2(n5311), .ZN(n5313) );
  XNOR2_X1 U6729 ( .A(n5313), .B(n4287), .ZN(n5316) );
  NOR2_X1 U6730 ( .A1(n7450), .A2(n5676), .ZN(n5314) );
  AOI21_X1 U6731 ( .B1(n7523), .B2(n5671), .A(n5314), .ZN(n5315) );
  NAND2_X1 U6732 ( .A1(n5316), .A2(n5315), .ZN(n9774) );
  OR2_X1 U6733 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  NAND2_X1 U6734 ( .A1(n6527), .A2(n5346), .ZN(n5325) );
  NAND2_X1 U6735 ( .A1(n5320), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5322) );
  MUX2_X1 U6736 ( .A(n5322), .B(P1_IR_REG_31__SCAN_IN), .S(n5321), .Z(n5323)
         );
  OR2_X1 U6737 ( .A1(n5320), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5367) );
  AND2_X1 U6738 ( .A1(n5323), .A2(n5367), .ZN(n7680) );
  AOI22_X1 U6739 ( .A1(n5191), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6364), .B2(
        n7680), .ZN(n5324) );
  NAND2_X1 U6740 ( .A1(n9779), .A2(n5634), .ZN(n5334) );
  INV_X1 U6741 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6742 ( .A1(n5327), .A2(n5326), .ZN(n5328) );
  NAND2_X1 U6743 ( .A1(n5351), .A2(n5328), .ZN(n9781) );
  INV_X1 U6744 ( .A(n9781), .ZN(n7466) );
  NAND2_X1 U6745 ( .A1(n5666), .A2(n7466), .ZN(n5332) );
  NAND2_X1 U6746 ( .A1(n7985), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6747 ( .A1(n6404), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6748 ( .A1(n5213), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6749 ( .A1(n9176), .A2(n5671), .ZN(n5333) );
  NAND2_X1 U6750 ( .A1(n5334), .A2(n5333), .ZN(n5335) );
  XNOR2_X1 U6751 ( .A(n5335), .B(n4287), .ZN(n5337) );
  NOR2_X1 U6752 ( .A1(n7588), .A2(n5676), .ZN(n5336) );
  AOI21_X1 U6753 ( .B1(n9779), .B2(n5671), .A(n5336), .ZN(n5338) );
  NAND2_X1 U6754 ( .A1(n5337), .A2(n5338), .ZN(n5342) );
  INV_X1 U6755 ( .A(n5337), .ZN(n5340) );
  INV_X1 U6756 ( .A(n5338), .ZN(n5339) );
  NAND2_X1 U6757 ( .A1(n5340), .A2(n5339), .ZN(n5341) );
  NAND2_X1 U6758 ( .A1(n5342), .A2(n5341), .ZN(n9773) );
  INV_X1 U6759 ( .A(n5342), .ZN(n5343) );
  XNOR2_X1 U6760 ( .A(n5345), .B(n5344), .ZN(n6546) );
  NAND2_X1 U6761 ( .A1(n6546), .A2(n5346), .ZN(n5349) );
  NAND2_X1 U6762 ( .A1(n5367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5347) );
  XNOR2_X1 U6763 ( .A(n5347), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U6764 ( .A1(n5191), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6364), .B2(
        n9831), .ZN(n5348) );
  NAND2_X1 U6765 ( .A1(n8110), .A2(n5659), .ZN(n5358) );
  NAND2_X1 U6766 ( .A1(n5105), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5356) );
  INV_X1 U6767 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6768 ( .A1(n5351), .A2(n5350), .ZN(n5352) );
  AND2_X1 U6769 ( .A1(n5393), .A2(n5352), .ZN(n7585) );
  NAND2_X1 U6770 ( .A1(n5666), .A2(n7585), .ZN(n5355) );
  NAND2_X1 U6771 ( .A1(n6404), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5354) );
  NAND2_X1 U6772 ( .A1(n5213), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6773 ( .A1(n9175), .A2(n5671), .ZN(n5357) );
  NAND2_X1 U6774 ( .A1(n5358), .A2(n5357), .ZN(n5359) );
  XNOR2_X1 U6775 ( .A(n5359), .B(n5616), .ZN(n5360) );
  OAI22_X1 U6776 ( .A1(n9966), .A2(n5593), .B1(n7580), .B2(n5676), .ZN(n5361)
         );
  XNOR2_X1 U6777 ( .A(n5360), .B(n5361), .ZN(n7507) );
  NOR2_X1 U6778 ( .A1(n7508), .A2(n7507), .ZN(n7506) );
  INV_X1 U6779 ( .A(n5360), .ZN(n5363) );
  INV_X1 U6780 ( .A(n5361), .ZN(n5362) );
  NAND2_X1 U6781 ( .A1(n5363), .A2(n5362), .ZN(n5364) );
  XNOR2_X1 U6782 ( .A(n5366), .B(n5365), .ZN(n6652) );
  NAND2_X1 U6783 ( .A1(n6652), .A2(n5346), .ZN(n5376) );
  INV_X1 U6784 ( .A(n5367), .ZN(n5369) );
  NAND2_X1 U6785 ( .A1(n5369), .A2(n5368), .ZN(n5371) );
  NAND2_X1 U6786 ( .A1(n5371), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5370) );
  MUX2_X1 U6787 ( .A(n5370), .B(P1_IR_REG_31__SCAN_IN), .S(n5372), .Z(n5374)
         );
  INV_X1 U6788 ( .A(n5371), .ZN(n5373) );
  NAND2_X1 U6789 ( .A1(n5373), .A2(n5372), .ZN(n5386) );
  AND2_X1 U6790 ( .A1(n5374), .A2(n5386), .ZN(n7702) );
  AOI22_X1 U6791 ( .A1(n5191), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6364), .B2(
        n7702), .ZN(n5375) );
  NAND2_X1 U6792 ( .A1(n5105), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5380) );
  XNOR2_X1 U6793 ( .A(n5393), .B(P1_REG3_REG_14__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U6794 ( .A1(n5666), .A2(n9044), .ZN(n5379) );
  NAND2_X1 U6795 ( .A1(n6404), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6796 ( .A1(n5213), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5377) );
  AOI22_X1 U6797 ( .A1(n8106), .A2(n5634), .B1(n5671), .B2(n9174), .ZN(n5381)
         );
  XOR2_X1 U6798 ( .A(n5616), .B(n5381), .Z(n5382) );
  AOI22_X1 U6799 ( .A1(n8106), .A2(n5671), .B1(n5415), .B2(n9174), .ZN(n9038)
         );
  INV_X1 U6800 ( .A(n5382), .ZN(n5383) );
  XNOR2_X1 U6801 ( .A(n5384), .B(n5385), .ZN(n6673) );
  NAND2_X1 U6802 ( .A1(n6673), .A2(n5346), .ZN(n5391) );
  NAND2_X1 U6803 ( .A1(n5386), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5387) );
  MUX2_X1 U6804 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5387), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n5389) );
  AND2_X1 U6805 ( .A1(n5389), .A2(n5388), .ZN(n9860) );
  AOI22_X1 U6806 ( .A1(n5191), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6364), .B2(
        n9860), .ZN(n5390) );
  NAND2_X1 U6807 ( .A1(n5105), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5398) );
  INV_X1 U6808 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9040) );
  INV_X1 U6809 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5392) );
  OAI21_X1 U6810 ( .B1(n5393), .B2(n9040), .A(n5392), .ZN(n5394) );
  AND2_X1 U6811 ( .A1(n5394), .A2(n5410), .ZN(n7671) );
  NAND2_X1 U6812 ( .A1(n5666), .A2(n7671), .ZN(n5397) );
  NAND2_X1 U6813 ( .A1(n6404), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6814 ( .A1(n5213), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5395) );
  INV_X1 U6815 ( .A(n9279), .ZN(n9275) );
  AOI22_X1 U6816 ( .A1(n9274), .A2(n5659), .B1(n5671), .B2(n9275), .ZN(n5399)
         );
  XOR2_X1 U6817 ( .A(n5616), .B(n5399), .Z(n5400) );
  NOR2_X1 U6818 ( .A1(n5401), .A2(n5400), .ZN(n5404) );
  INV_X1 U6819 ( .A(n5404), .ZN(n5403) );
  NAND2_X1 U6820 ( .A1(n5403), .A2(n5402), .ZN(n7670) );
  OAI22_X1 U6821 ( .A1(n9276), .A2(n5593), .B1(n9279), .B2(n5676), .ZN(n7669)
         );
  NOR2_X2 U6822 ( .A1(n7670), .A2(n7669), .ZN(n7668) );
  XNOR2_X1 U6823 ( .A(n5406), .B(n5405), .ZN(n6881) );
  NAND2_X1 U6824 ( .A1(n6881), .A2(n5346), .ZN(n5409) );
  NAND2_X1 U6825 ( .A1(n5388), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5407) );
  XNOR2_X1 U6826 ( .A(n5407), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9873) );
  AOI22_X1 U6827 ( .A1(n5191), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6364), .B2(
        n9873), .ZN(n5408) );
  NAND2_X1 U6828 ( .A1(n5410), .A2(n9094), .ZN(n5411) );
  NAND2_X1 U6829 ( .A1(n5412), .A2(n5411), .ZN(n9532) );
  INV_X1 U6830 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9616) );
  OAI22_X1 U6831 ( .A1(n9532), .A2(n5511), .B1(n5149), .B2(n9616), .ZN(n5414)
         );
  INV_X1 U6832 ( .A(n7985), .ZN(n5589) );
  INV_X1 U6833 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9533) );
  INV_X1 U6834 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9676) );
  OAI22_X1 U6835 ( .A1(n5589), .A2(n9533), .B1(n5148), .B2(n9676), .ZN(n5413)
         );
  OR2_X1 U6836 ( .A1(n5414), .A2(n5413), .ZN(n9281) );
  AOI22_X1 U6837 ( .A1(n9529), .A2(n5671), .B1(n5415), .B2(n9281), .ZN(n5419)
         );
  NAND2_X1 U6838 ( .A1(n9529), .A2(n5634), .ZN(n5417) );
  NAND2_X1 U6839 ( .A1(n9281), .A2(n5671), .ZN(n5416) );
  NAND2_X1 U6840 ( .A1(n5417), .A2(n5416), .ZN(n5418) );
  XNOR2_X1 U6841 ( .A(n5418), .B(n5616), .ZN(n5421) );
  XOR2_X1 U6842 ( .A(n5419), .B(n5421), .Z(n9092) );
  INV_X1 U6843 ( .A(n5419), .ZN(n5420) );
  NOR2_X1 U6844 ( .A1(n5421), .A2(n5420), .ZN(n9100) );
  XNOR2_X1 U6845 ( .A(n5423), .B(n5422), .ZN(n9099) );
  OAI22_X1 U6846 ( .A1(n9670), .A2(n5517), .B1(n9287), .B2(n5593), .ZN(n5426)
         );
  XOR2_X1 U6847 ( .A(n5616), .B(n5426), .Z(n9062) );
  INV_X1 U6848 ( .A(n5427), .ZN(n5431) );
  INV_X1 U6849 ( .A(n5428), .ZN(n5429) );
  NAND2_X1 U6850 ( .A1(n5429), .A2(SI_18_), .ZN(n5430) );
  INV_X1 U6851 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7192) );
  INV_X1 U6852 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8956) );
  MUX2_X1 U6853 ( .A(n7192), .B(n8956), .S(n6362), .Z(n5434) );
  INV_X1 U6854 ( .A(SI_19_), .ZN(n5433) );
  NAND2_X1 U6855 ( .A1(n5434), .A2(n5433), .ZN(n5476) );
  INV_X1 U6856 ( .A(n5434), .ZN(n5435) );
  NAND2_X1 U6857 ( .A1(n5435), .A2(SI_19_), .ZN(n5436) );
  NAND2_X1 U6858 ( .A1(n5476), .A2(n5436), .ZN(n5475) );
  XNOR2_X1 U6859 ( .A(n5481), .B(n5475), .ZN(n7191) );
  NAND2_X1 U6860 ( .A1(n7191), .A2(n5346), .ZN(n5439) );
  AOI22_X1 U6861 ( .A1(n5191), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5437), .B2(
        n6364), .ZN(n5438) );
  NAND2_X1 U6862 ( .A1(n9474), .A2(n5634), .ZN(n5449) );
  INV_X1 U6863 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6864 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  NAND2_X1 U6865 ( .A1(n5460), .A2(n5442), .ZN(n9475) );
  OR2_X1 U6866 ( .A1(n9475), .A2(n5511), .ZN(n5447) );
  INV_X1 U6867 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9664) );
  NAND2_X1 U6868 ( .A1(n5105), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6869 ( .A1(n5213), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5443) );
  OAI211_X1 U6870 ( .C1(n5148), .C2(n9664), .A(n5444), .B(n5443), .ZN(n5445)
         );
  INV_X1 U6871 ( .A(n5445), .ZN(n5446) );
  AND2_X1 U6872 ( .A1(n5447), .A2(n5446), .ZN(n9290) );
  INV_X1 U6873 ( .A(n9290), .ZN(n9288) );
  NAND2_X1 U6874 ( .A1(n9288), .A2(n5671), .ZN(n5448) );
  NAND2_X1 U6875 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  XNOR2_X1 U6876 ( .A(n5450), .B(n4287), .ZN(n5468) );
  NOR2_X1 U6877 ( .A1(n9290), .A2(n5676), .ZN(n5451) );
  AOI21_X1 U6878 ( .B1(n9474), .B2(n5671), .A(n5451), .ZN(n5469) );
  NAND2_X1 U6879 ( .A1(n5468), .A2(n5469), .ZN(n9059) );
  OR2_X1 U6880 ( .A1(n5481), .A2(n5475), .ZN(n5452) );
  INV_X1 U6881 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7282) );
  INV_X1 U6882 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7253) );
  MUX2_X1 U6883 ( .A(n7282), .B(n7253), .S(n6362), .Z(n5453) );
  INV_X1 U6884 ( .A(SI_20_), .ZN(n8932) );
  NAND2_X1 U6885 ( .A1(n5453), .A2(n8932), .ZN(n5478) );
  INV_X1 U6886 ( .A(n5453), .ZN(n5454) );
  NAND2_X1 U6887 ( .A1(n5454), .A2(SI_20_), .ZN(n5455) );
  NAND2_X1 U6888 ( .A1(n5478), .A2(n5455), .ZN(n5477) );
  INV_X1 U6889 ( .A(n5477), .ZN(n5456) );
  NAND2_X1 U6890 ( .A1(n7252), .A2(n5346), .ZN(n5459) );
  OR2_X1 U6891 ( .A1(n5127), .A2(n7253), .ZN(n5458) );
  INV_X1 U6892 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9138) );
  NAND2_X1 U6893 ( .A1(n5460), .A2(n9138), .ZN(n5461) );
  AND2_X1 U6894 ( .A1(n5508), .A2(n5461), .ZN(n9454) );
  INV_X1 U6895 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U6896 ( .A1(n6404), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6897 ( .A1(n5213), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5462) );
  OAI211_X1 U6898 ( .C1(n5589), .C2(n9461), .A(n5463), .B(n5462), .ZN(n5464)
         );
  AOI21_X1 U6899 ( .B1(n9454), .B2(n5666), .A(n5464), .ZN(n9173) );
  OAI22_X1 U6900 ( .A1(n9662), .A2(n5517), .B1(n9173), .B2(n5593), .ZN(n5465)
         );
  XNOR2_X1 U6901 ( .A(n5465), .B(n5616), .ZN(n5467) );
  OAI22_X1 U6902 ( .A1(n9662), .A2(n5593), .B1(n9173), .B2(n5676), .ZN(n5466)
         );
  NOR2_X1 U6903 ( .A1(n5467), .A2(n5466), .ZN(n5473) );
  AOI21_X1 U6904 ( .B1(n5467), .B2(n5466), .A(n5473), .ZN(n9134) );
  INV_X1 U6905 ( .A(n5468), .ZN(n5471) );
  INV_X1 U6906 ( .A(n5469), .ZN(n5470) );
  NAND2_X1 U6907 ( .A1(n5471), .A2(n5470), .ZN(n9135) );
  NAND2_X1 U6908 ( .A1(n9133), .A2(n5472), .ZN(n9132) );
  INV_X1 U6909 ( .A(n5473), .ZN(n5474) );
  NAND2_X1 U6910 ( .A1(n9132), .A2(n5474), .ZN(n9072) );
  OR2_X1 U6911 ( .A1(n5475), .A2(n5477), .ZN(n5480) );
  OR2_X1 U6912 ( .A1(n5477), .A2(n5476), .ZN(n5479) );
  INV_X1 U6913 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7342) );
  INV_X1 U6914 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7331) );
  MUX2_X1 U6915 ( .A(n7342), .B(n7331), .S(n6362), .Z(n5498) );
  XNOR2_X1 U6916 ( .A(n5498), .B(SI_21_), .ZN(n5497) );
  XNOR2_X1 U6917 ( .A(n5496), .B(n5497), .ZN(n7330) );
  NAND2_X1 U6918 ( .A1(n7330), .A2(n5346), .ZN(n5483) );
  OR2_X1 U6919 ( .A1(n5127), .A2(n7331), .ZN(n5482) );
  XNOR2_X1 U6920 ( .A(n5508), .B(P1_REG3_REG_21__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U6921 ( .A1(n9445), .A2(n5666), .ZN(n5489) );
  INV_X1 U6922 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6923 ( .A1(n6404), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U6924 ( .A1(n5213), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5484) );
  OAI211_X1 U6925 ( .C1(n5589), .C2(n5486), .A(n5485), .B(n5484), .ZN(n5487)
         );
  INV_X1 U6926 ( .A(n5487), .ZN(n5488) );
  NAND2_X1 U6927 ( .A1(n9444), .A2(n5659), .ZN(n5491) );
  NAND2_X1 U6928 ( .A1(n9294), .A2(n5671), .ZN(n5490) );
  NAND2_X1 U6929 ( .A1(n5491), .A2(n5490), .ZN(n5492) );
  XOR2_X1 U6930 ( .A(n5493), .B(n5494), .Z(n9075) );
  NAND2_X1 U6931 ( .A1(n9072), .A2(n9075), .ZN(n9073) );
  NAND2_X1 U6932 ( .A1(n9073), .A2(n5495), .ZN(n5522) );
  INV_X1 U6933 ( .A(n5522), .ZN(n5520) );
  INV_X1 U6934 ( .A(n5498), .ZN(n5499) );
  INV_X1 U6935 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7385) );
  INV_X1 U6936 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7387) );
  MUX2_X1 U6937 ( .A(n7385), .B(n7387), .S(n6362), .Z(n5501) );
  INV_X1 U6938 ( .A(SI_22_), .ZN(n5500) );
  NAND2_X1 U6939 ( .A1(n5501), .A2(n5500), .ZN(n5525) );
  INV_X1 U6940 ( .A(n5501), .ZN(n5502) );
  NAND2_X1 U6941 ( .A1(n5502), .A2(SI_22_), .ZN(n5503) );
  NAND2_X1 U6942 ( .A1(n5525), .A2(n5503), .ZN(n5526) );
  XNOR2_X1 U6943 ( .A(n5527), .B(n5526), .ZN(n7384) );
  NAND2_X1 U6944 ( .A1(n7384), .A2(n5346), .ZN(n5505) );
  OR2_X1 U6945 ( .A1(n5127), .A2(n7387), .ZN(n5504) );
  NAND2_X1 U6946 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n5506) );
  INV_X1 U6947 ( .A(n5540), .ZN(n5510) );
  INV_X1 U6948 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9078) );
  INV_X1 U6949 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5507) );
  OAI21_X1 U6950 ( .B1(n5508), .B2(n9078), .A(n5507), .ZN(n5509) );
  NAND2_X1 U6951 ( .A1(n5510), .A2(n5509), .ZN(n9425) );
  OR2_X1 U6952 ( .A1(n9425), .A2(n5511), .ZN(n5516) );
  INV_X1 U6953 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9586) );
  NAND2_X1 U6954 ( .A1(n5105), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U6955 ( .A1(n6404), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5512) );
  OAI211_X1 U6956 ( .C1(n9586), .C2(n5149), .A(n5513), .B(n5512), .ZN(n5514)
         );
  INV_X1 U6957 ( .A(n5514), .ZN(n5515) );
  OAI22_X1 U6958 ( .A1(n9655), .A2(n5517), .B1(n9299), .B2(n5593), .ZN(n5518)
         );
  XOR2_X1 U6959 ( .A(n5616), .B(n5518), .Z(n5521) );
  INV_X1 U6960 ( .A(n5521), .ZN(n5519) );
  NAND2_X1 U6961 ( .A1(n5520), .A2(n5519), .ZN(n5523) );
  OAI22_X1 U6962 ( .A1(n9655), .A2(n5593), .B1(n9299), .B2(n5676), .ZN(n9145)
         );
  INV_X1 U6963 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7431) );
  INV_X1 U6964 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5537) );
  MUX2_X1 U6965 ( .A(n7431), .B(n5537), .S(n6362), .Z(n5529) );
  INV_X1 U6966 ( .A(SI_23_), .ZN(n5528) );
  NAND2_X1 U6967 ( .A1(n5529), .A2(n5528), .ZN(n5552) );
  INV_X1 U6968 ( .A(n5529), .ZN(n5530) );
  NAND2_X1 U6969 ( .A1(n5530), .A2(SI_23_), .ZN(n5531) );
  NAND2_X1 U6970 ( .A1(n5552), .A2(n5531), .ZN(n5533) );
  NAND2_X1 U6971 ( .A1(n5532), .A2(n5533), .ZN(n5536) );
  INV_X1 U6972 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U6973 ( .A1(n5536), .A2(n5553), .ZN(n7429) );
  NAND2_X1 U6974 ( .A1(n7429), .A2(n5346), .ZN(n5539) );
  OR2_X1 U6975 ( .A1(n5127), .A2(n5537), .ZN(n5538) );
  NAND2_X1 U6976 ( .A1(n9579), .A2(n5634), .ZN(n5546) );
  NOR2_X1 U6977 ( .A1(n5540), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5541) );
  INV_X1 U6978 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9406) );
  NAND2_X1 U6979 ( .A1(n5213), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U6980 ( .A1(n6404), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5542) );
  OAI211_X1 U6981 ( .C1(n5589), .C2(n9406), .A(n5543), .B(n5542), .ZN(n5544)
         );
  AOI21_X1 U6982 ( .B1(n4888), .B2(n5666), .A(n5544), .ZN(n9301) );
  OR2_X1 U6983 ( .A1(n9301), .A2(n5593), .ZN(n5545) );
  NAND2_X1 U6984 ( .A1(n5546), .A2(n5545), .ZN(n5547) );
  XNOR2_X1 U6985 ( .A(n5547), .B(n4287), .ZN(n5550) );
  NOR2_X1 U6986 ( .A1(n9301), .A2(n5676), .ZN(n5548) );
  AOI21_X1 U6987 ( .B1(n9579), .B2(n5671), .A(n5548), .ZN(n5549) );
  NAND2_X1 U6988 ( .A1(n5550), .A2(n5549), .ZN(n9113) );
  OR2_X1 U6989 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  INV_X1 U6990 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7664) );
  INV_X1 U6991 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7540) );
  MUX2_X1 U6992 ( .A(n7664), .B(n7540), .S(n6362), .Z(n5555) );
  INV_X1 U6993 ( .A(SI_24_), .ZN(n5554) );
  NAND2_X1 U6994 ( .A1(n5555), .A2(n5554), .ZN(n5577) );
  INV_X1 U6995 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U6996 ( .A1(n5556), .A2(SI_24_), .ZN(n5557) );
  AND2_X1 U6997 ( .A1(n5577), .A2(n5557), .ZN(n5575) );
  XNOR2_X1 U6998 ( .A(n5576), .B(n5575), .ZN(n7539) );
  NAND2_X1 U6999 ( .A1(n7539), .A2(n5346), .ZN(n5559) );
  OR2_X1 U7000 ( .A1(n5127), .A2(n7540), .ZN(n5558) );
  NAND2_X1 U7001 ( .A1(n9574), .A2(n5659), .ZN(n5567) );
  NOR2_X1 U7002 ( .A1(n5560), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5561) );
  OR2_X1 U7003 ( .A1(n5584), .A2(n5561), .ZN(n9109) );
  INV_X1 U7004 ( .A(n9109), .ZN(n9396) );
  INV_X1 U7005 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7006 ( .A1(n5213), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U7007 ( .A1(n5120), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5562) );
  OAI211_X1 U7008 ( .C1(n5589), .C2(n5564), .A(n5563), .B(n5562), .ZN(n5565)
         );
  AOI21_X1 U7009 ( .B1(n9396), .B2(n5666), .A(n5565), .ZN(n9172) );
  OR2_X1 U7010 ( .A1(n9172), .A2(n5593), .ZN(n5566) );
  NAND2_X1 U7011 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  XNOR2_X1 U7012 ( .A(n5568), .B(n4287), .ZN(n5571) );
  NOR2_X1 U7013 ( .A1(n9172), .A2(n5676), .ZN(n5569) );
  AOI21_X1 U7014 ( .B1(n9574), .B2(n5671), .A(n5569), .ZN(n5570) );
  NAND2_X1 U7015 ( .A1(n5571), .A2(n5570), .ZN(n5574) );
  OR2_X1 U7016 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  NAND2_X1 U7017 ( .A1(n5573), .A2(n9111), .ZN(n9110) );
  INV_X1 U7018 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8905) );
  INV_X1 U7019 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7569) );
  MUX2_X1 U7020 ( .A(n8905), .B(n7569), .S(n6362), .Z(n5579) );
  INV_X1 U7021 ( .A(SI_25_), .ZN(n5578) );
  NAND2_X1 U7022 ( .A1(n5579), .A2(n5578), .ZN(n5599) );
  INV_X1 U7023 ( .A(n5579), .ZN(n5580) );
  NAND2_X1 U7024 ( .A1(n5580), .A2(SI_25_), .ZN(n5581) );
  AND2_X1 U7025 ( .A1(n5599), .A2(n5581), .ZN(n5597) );
  XNOR2_X1 U7026 ( .A(n5598), .B(n5597), .ZN(n7567) );
  NAND2_X1 U7027 ( .A1(n7567), .A2(n5346), .ZN(n5583) );
  OR2_X1 U7028 ( .A1(n5127), .A2(n7569), .ZN(n5582) );
  OR2_X1 U7029 ( .A1(n5584), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7030 ( .A1(n5584), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5607) );
  AND2_X1 U7031 ( .A1(n5585), .A2(n5607), .ZN(n9382) );
  NAND2_X1 U7032 ( .A1(n9382), .A2(n5666), .ZN(n5592) );
  INV_X1 U7033 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7034 ( .A1(n5213), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7035 ( .A1(n5120), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5586) );
  OAI211_X1 U7036 ( .C1(n5589), .C2(n5588), .A(n5587), .B(n5586), .ZN(n5590)
         );
  INV_X1 U7037 ( .A(n5590), .ZN(n5591) );
  OAI22_X1 U7038 ( .A1(n9649), .A2(n5593), .B1(n9307), .B2(n5676), .ZN(n5620)
         );
  NAND2_X1 U7039 ( .A1(n9381), .A2(n5634), .ZN(n5595) );
  INV_X1 U7040 ( .A(n9307), .ZN(n9309) );
  NAND2_X1 U7041 ( .A1(n9309), .A2(n5671), .ZN(n5594) );
  NAND2_X1 U7042 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  XNOR2_X1 U7043 ( .A(n5596), .B(n5616), .ZN(n5619) );
  XOR2_X1 U7044 ( .A(n5620), .B(n5619), .Z(n9084) );
  INV_X1 U7045 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7622) );
  INV_X1 U7046 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7620) );
  MUX2_X1 U7047 ( .A(n7622), .B(n7620), .S(n6362), .Z(n5601) );
  INV_X1 U7048 ( .A(SI_26_), .ZN(n5600) );
  NAND2_X1 U7049 ( .A1(n5601), .A2(n5600), .ZN(n5626) );
  INV_X1 U7050 ( .A(n5601), .ZN(n5602) );
  NAND2_X1 U7051 ( .A1(n5602), .A2(SI_26_), .ZN(n5603) );
  AND2_X1 U7052 ( .A1(n5626), .A2(n5603), .ZN(n5624) );
  OR2_X1 U7053 ( .A1(n5127), .A2(n7620), .ZN(n5604) );
  NAND2_X1 U7054 ( .A1(n9563), .A2(n5659), .ZN(n5615) );
  NAND2_X1 U7055 ( .A1(n5105), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5613) );
  INV_X1 U7056 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7057 ( .A1(n5606), .A2(n5607), .ZN(n5609) );
  INV_X1 U7058 ( .A(n5607), .ZN(n5608) );
  NAND2_X1 U7059 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n5608), .ZN(n5664) );
  AND2_X1 U7060 ( .A1(n5609), .A2(n5664), .ZN(n9361) );
  NAND2_X1 U7061 ( .A1(n5666), .A2(n9361), .ZN(n5612) );
  NAND2_X1 U7062 ( .A1(n5120), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U7063 ( .A1(n5119), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5610) );
  INV_X1 U7064 ( .A(n9312), .ZN(n9171) );
  NAND2_X1 U7065 ( .A1(n9171), .A2(n5671), .ZN(n5614) );
  NAND2_X1 U7066 ( .A1(n5615), .A2(n5614), .ZN(n5617) );
  XNOR2_X1 U7067 ( .A(n5617), .B(n5616), .ZN(n5649) );
  NOR2_X1 U7068 ( .A1(n9312), .A2(n5676), .ZN(n5618) );
  AOI21_X1 U7069 ( .B1(n9563), .B2(n5671), .A(n5618), .ZN(n5647) );
  XNOR2_X1 U7070 ( .A(n5649), .B(n5647), .ZN(n9159) );
  INV_X1 U7071 ( .A(n5619), .ZN(n5622) );
  INV_X1 U7072 ( .A(n5620), .ZN(n5621) );
  NAND2_X1 U7073 ( .A1(n5622), .A2(n5621), .ZN(n9160) );
  INV_X1 U7074 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7635) );
  INV_X1 U7075 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7653) );
  MUX2_X1 U7076 ( .A(n7635), .B(n7653), .S(n6362), .Z(n5629) );
  INV_X1 U7077 ( .A(SI_27_), .ZN(n5628) );
  NAND2_X1 U7078 ( .A1(n5629), .A2(n5628), .ZN(n5652) );
  INV_X1 U7079 ( .A(n5629), .ZN(n5630) );
  NAND2_X1 U7080 ( .A1(n5630), .A2(SI_27_), .ZN(n5631) );
  AND2_X1 U7081 ( .A1(n5652), .A2(n5631), .ZN(n5650) );
  OR2_X1 U7082 ( .A1(n5127), .A2(n7653), .ZN(n5632) );
  NAND2_X1 U7083 ( .A1(n9556), .A2(n5634), .ZN(n5640) );
  XNOR2_X1 U7084 ( .A(n5664), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U7085 ( .A1(n5666), .A2(n9342), .ZN(n5638) );
  NAND2_X1 U7086 ( .A1(n7985), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7087 ( .A1(n5120), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7088 ( .A1(n5119), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5635) );
  INV_X1 U7089 ( .A(n9162), .ZN(n9315) );
  NAND2_X1 U7090 ( .A1(n9315), .A2(n5671), .ZN(n5639) );
  NAND2_X1 U7091 ( .A1(n5640), .A2(n5639), .ZN(n5641) );
  XNOR2_X1 U7092 ( .A(n5641), .B(n4287), .ZN(n5644) );
  INV_X1 U7093 ( .A(n5644), .ZN(n5646) );
  NOR2_X1 U7094 ( .A1(n9162), .A2(n5676), .ZN(n5642) );
  AOI21_X1 U7095 ( .B1(n9556), .B2(n5671), .A(n5642), .ZN(n5643) );
  INV_X1 U7096 ( .A(n5643), .ZN(n5645) );
  AOI21_X1 U7097 ( .B1(n5646), .B2(n5645), .A(n5703), .ZN(n5734) );
  INV_X1 U7098 ( .A(n5647), .ZN(n5648) );
  NAND2_X1 U7099 ( .A1(n5649), .A2(n5648), .ZN(n5735) );
  INV_X1 U7100 ( .A(n5737), .ZN(n5702) );
  INV_X1 U7101 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7656) );
  INV_X1 U7102 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7732) );
  MUX2_X1 U7103 ( .A(n7656), .B(n7732), .S(n6362), .Z(n5654) );
  INV_X1 U7104 ( .A(SI_28_), .ZN(n5653) );
  NAND2_X1 U7105 ( .A1(n5654), .A2(n5653), .ZN(n6235) );
  INV_X1 U7106 ( .A(n5654), .ZN(n5655) );
  NAND2_X1 U7107 ( .A1(n5655), .A2(SI_28_), .ZN(n5656) );
  AND2_X1 U7108 ( .A1(n6235), .A2(n5656), .ZN(n6233) );
  NAND2_X1 U7109 ( .A1(n7655), .A2(n5346), .ZN(n5658) );
  OR2_X1 U7110 ( .A1(n5127), .A2(n7732), .ZN(n5657) );
  NAND2_X1 U7111 ( .A1(n9334), .A2(n5659), .ZN(n5673) );
  NAND2_X1 U7112 ( .A1(n5105), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5670) );
  INV_X1 U7113 ( .A(n5664), .ZN(n5661) );
  AND2_X1 U7114 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5660) );
  NAND2_X1 U7115 ( .A1(n5661), .A2(n5660), .ZN(n5718) );
  INV_X1 U7116 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5663) );
  INV_X1 U7117 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5662) );
  OAI21_X1 U7118 ( .B1(n5664), .B2(n5663), .A(n5662), .ZN(n5665) );
  AND2_X1 U7119 ( .A1(n5718), .A2(n5665), .ZN(n9336) );
  NAND2_X1 U7120 ( .A1(n5666), .A2(n9336), .ZN(n5669) );
  NAND2_X1 U7121 ( .A1(n5120), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7122 ( .A1(n5119), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5667) );
  INV_X1 U7123 ( .A(n7996), .ZN(n9317) );
  NAND2_X1 U7124 ( .A1(n9317), .A2(n5671), .ZN(n5672) );
  NAND2_X1 U7125 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  XNOR2_X1 U7126 ( .A(n5674), .B(n4287), .ZN(n5678) );
  NAND2_X1 U7127 ( .A1(n9334), .A2(n5671), .ZN(n5675) );
  OAI21_X1 U7128 ( .B1(n7996), .B2(n5676), .A(n5675), .ZN(n5677) );
  XNOR2_X1 U7129 ( .A(n5678), .B(n5677), .ZN(n5704) );
  INV_X1 U7130 ( .A(n5704), .ZN(n5701) );
  INV_X1 U7131 ( .A(P1_B_REG_SCAN_IN), .ZN(n7726) );
  OR2_X1 U7132 ( .A1(n7568), .A2(n7726), .ZN(n5680) );
  MUX2_X1 U7133 ( .A(P1_B_REG_SCAN_IN), .B(n5680), .S(n7541), .Z(n5681) );
  AND2_X1 U7134 ( .A1(n5679), .A2(n5681), .ZN(n6389) );
  INV_X1 U7135 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5682) );
  INV_X1 U7136 ( .A(n5679), .ZN(n7621) );
  AND2_X1 U7137 ( .A1(n7541), .A2(n7621), .ZN(n6393) );
  AOI21_X1 U7138 ( .B1(n6389), .B2(n5682), .A(n6393), .ZN(n6853) );
  INV_X1 U7139 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5683) );
  NOR2_X1 U7140 ( .A1(n5679), .A2(n7568), .ZN(n6391) );
  AOI21_X1 U7141 ( .B1(n6389), .B2(n5683), .A(n6391), .ZN(n7054) );
  NOR4_X1 U7142 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5687) );
  NOR4_X1 U7143 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5686) );
  NOR4_X1 U7144 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5685) );
  NOR4_X1 U7145 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5684) );
  NAND4_X1 U7146 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .ZN(n5693)
         );
  NOR2_X1 U7147 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n5691) );
  NOR4_X1 U7148 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5690) );
  NOR4_X1 U7149 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5689) );
  NOR4_X1 U7150 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5688) );
  NAND4_X1 U7151 ( .A1(n5691), .A2(n5690), .A3(n5689), .A4(n5688), .ZN(n5692)
         );
  OAI21_X1 U7152 ( .B1(n5693), .B2(n5692), .A(n6389), .ZN(n6556) );
  NAND3_X1 U7153 ( .A1(n6853), .A2(n7054), .A3(n6556), .ZN(n5713) );
  NAND2_X1 U7154 ( .A1(n5694), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5696) );
  XNOR2_X1 U7155 ( .A(n5696), .B(n5695), .ZN(n6365) );
  AND2_X1 U7156 ( .A1(n6365), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6531) );
  NAND2_X1 U7157 ( .A1(n6531), .A2(n5708), .ZN(n6554) );
  OR2_X1 U7158 ( .A1(n5713), .A2(n6554), .ZN(n5717) );
  AND2_X1 U7159 ( .A1(n8237), .A2(n8225), .ZN(n8093) );
  INV_X1 U7160 ( .A(n8093), .ZN(n5706) );
  AND2_X1 U7161 ( .A1(n5698), .A2(n8049), .ZN(n5705) );
  NAND2_X1 U7162 ( .A1(n5705), .A2(n8235), .ZN(n9965) );
  NAND2_X1 U7163 ( .A1(n5706), .A2(n9965), .ZN(n5699) );
  NOR2_X2 U7164 ( .A1(n5717), .A2(n5699), .ZN(n9158) );
  INV_X1 U7165 ( .A(n5703), .ZN(n5700) );
  AND2_X1 U7166 ( .A1(n5704), .A2(n9158), .ZN(n5731) );
  INV_X1 U7167 ( .A(n5705), .ZN(n7056) );
  OR2_X1 U7168 ( .A1(n7056), .A2(n7254), .ZN(n7064) );
  AND2_X1 U7169 ( .A1(n5705), .A2(n7254), .ZN(n9917) );
  NAND2_X1 U7170 ( .A1(n9917), .A2(n5437), .ZN(n6557) );
  OR2_X1 U7171 ( .A1(n6554), .A2(n6557), .ZN(n9531) );
  INV_X1 U7172 ( .A(n8235), .ZN(n6562) );
  NAND2_X1 U7173 ( .A1(n5713), .A2(n9965), .ZN(n5707) );
  MUX2_X1 U7174 ( .A(n6562), .B(n5707), .S(n5706), .Z(n5709) );
  NAND2_X1 U7175 ( .A1(n5709), .A2(n5708), .ZN(n6529) );
  NAND2_X1 U7176 ( .A1(n6529), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5716) );
  NAND2_X1 U7177 ( .A1(n7060), .A2(n6561), .ZN(n5710) );
  NOR2_X1 U7178 ( .A1(n6554), .A2(n5710), .ZN(n8241) );
  NOR2_X1 U7179 ( .A1(n7064), .A2(P1_U3086), .ZN(n5711) );
  OR2_X1 U7180 ( .A1(n8241), .A2(n5711), .ZN(n5712) );
  NAND2_X1 U7181 ( .A1(n5713), .A2(n5712), .ZN(n6530) );
  INV_X1 U7182 ( .A(n6365), .ZN(n5714) );
  NAND2_X1 U7183 ( .A1(n5714), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8238) );
  AND2_X1 U7184 ( .A1(n6530), .A2(n8238), .ZN(n5715) );
  AND2_X1 U7185 ( .A1(n5716), .A2(n5715), .ZN(n9797) );
  INV_X1 U7186 ( .A(n9336), .ZN(n5727) );
  NOR2_X2 U7187 ( .A1(n5717), .A2(n8235), .ZN(n9164) );
  INV_X1 U7188 ( .A(n5718), .ZN(n9322) );
  NAND2_X1 U7189 ( .A1(n5666), .A2(n9322), .ZN(n5722) );
  NAND2_X1 U7190 ( .A1(n7985), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7191 ( .A1(n5120), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7192 ( .A1(n5119), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5719) );
  AND4_X1 U7193 ( .A1(n5722), .A2(n5721), .A3(n5720), .A4(n5719), .ZN(n7988)
         );
  NAND2_X1 U7194 ( .A1(n8093), .A2(n4285), .ZN(n9161) );
  NOR2_X1 U7195 ( .A1(n7988), .A2(n9161), .ZN(n5725) );
  INV_X1 U7196 ( .A(n4285), .ZN(n6495) );
  NAND2_X1 U7197 ( .A1(n8093), .A2(n6495), .ZN(n9163) );
  NOR2_X1 U7198 ( .A1(n9162), .A2(n9163), .ZN(n5724) );
  OR2_X1 U7199 ( .A1(n5725), .A2(n5724), .ZN(n9330) );
  AOI22_X1 U7200 ( .A1(n9164), .A2(n9330), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5726) );
  OAI21_X1 U7201 ( .B1(n9797), .B2(n5727), .A(n5726), .ZN(n5728) );
  AOI21_X1 U7202 ( .B1(n9334), .B2(n4282), .A(n5728), .ZN(n5729) );
  INV_X1 U7203 ( .A(n5729), .ZN(n5730) );
  AOI21_X1 U7204 ( .B1(n5737), .B2(n5731), .A(n4357), .ZN(n5732) );
  NAND2_X1 U7205 ( .A1(n5733), .A2(n5732), .ZN(P1_U3220) );
  AOI21_X1 U7206 ( .B1(n9157), .B2(n5735), .A(n5734), .ZN(n5736) );
  OAI21_X1 U7207 ( .B1(n5737), .B2(n5736), .A(n9158), .ZN(n5744) );
  NAND2_X1 U7208 ( .A1(n9556), .A2(n4282), .ZN(n5743) );
  NOR2_X1 U7209 ( .A1(n7996), .A2(n9161), .ZN(n5739) );
  NOR2_X1 U7210 ( .A1(n9312), .A2(n9163), .ZN(n5738) );
  OR2_X1 U7211 ( .A1(n5739), .A2(n5738), .ZN(n9346) );
  AOI22_X1 U7212 ( .A1(n9164), .A2(n9346), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n5741) );
  INV_X1 U7213 ( .A(n9797), .ZN(n9140) );
  NAND2_X1 U7214 ( .A1(n9140), .A2(n9342), .ZN(n5740) );
  AND2_X1 U7215 ( .A1(n5741), .A2(n5740), .ZN(n5742) );
  NAND3_X1 U7216 ( .A1(n5744), .A2(n5743), .A3(n5742), .ZN(P1_U3214) );
  NOR2_X1 U7217 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5746) );
  NOR2_X1 U7218 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5745) );
  AND2_X1 U7219 ( .A1(n5746), .A2(n5745), .ZN(n5747) );
  AND2_X2 U7220 ( .A1(n5820), .A2(n5747), .ZN(n5794) );
  INV_X1 U7221 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5749) );
  NAND4_X1 U7222 ( .A1(n5803), .A2(n5808), .A3(n5796), .A4(n5749), .ZN(n5750)
         );
  INV_X1 U7223 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U7224 ( .A1(n5769), .A2(n5768), .ZN(n5754) );
  INV_X1 U7225 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7226 ( .A1(n5763), .A2(n5762), .ZN(n5755) );
  INV_X1 U7227 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5756) );
  NOR3_X1 U7228 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U7229 ( .A1(n5771), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5761) );
  XNOR2_X1 U7230 ( .A(n5761), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6317) );
  INV_X1 U7231 ( .A(n6317), .ZN(n7624) );
  OR3_X1 U7232 ( .A1(n7731), .A2(n7624), .A3(n7667), .ZN(n6423) );
  NOR2_X1 U7233 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5764) );
  INV_X1 U7234 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7235 ( .A1(n6248), .A2(n5765), .ZN(n6251) );
  NAND2_X1 U7236 ( .A1(n6251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5766) );
  XNOR2_X1 U7237 ( .A(n5766), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U7238 ( .A1(n4321), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5767) );
  XNOR2_X1 U7239 ( .A(n5767), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U7240 ( .A1(n7767), .A2(n7982), .ZN(n7942) );
  NAND2_X1 U7241 ( .A1(n6423), .A2(n7942), .ZN(n5770) );
  XNOR2_X1 U7242 ( .A(n5769), .B(n5768), .ZN(n6712) );
  NAND2_X1 U7243 ( .A1(n5770), .A2(n6712), .ZN(n5870) );
  INV_X1 U7244 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5772) );
  INV_X1 U7245 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U7246 ( .A1(n5779), .A2(n5778), .ZN(n5871) );
  NAND2_X1 U7247 ( .A1(n5870), .A2(n6308), .ZN(n5780) );
  NAND2_X1 U7248 ( .A1(n5780), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  AND2_X1 U7249 ( .A1(n6712), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6429) );
  INV_X1 U7250 ( .A(n6429), .ZN(n5781) );
  NOR2_X1 U7251 ( .A1(n6423), .A2(n5781), .ZN(n8455) );
  INV_X1 U7252 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5786) );
  INV_X1 U7253 ( .A(n5782), .ZN(n5783) );
  NAND2_X1 U7254 ( .A1(n5783), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7255 ( .A1(n5788), .A2(n5787), .ZN(n5790) );
  INV_X1 U7256 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5784) );
  MUX2_X1 U7257 ( .A(n5786), .B(P2_REG2_REG_19__SCAN_IN), .S(n7193), .Z(n5947)
         );
  OR2_X1 U7258 ( .A1(n5788), .A2(n5787), .ZN(n5789) );
  AND2_X1 U7259 ( .A1(n5790), .A2(n5789), .ZN(n6968) );
  INV_X1 U7260 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8724) );
  OR2_X1 U7261 ( .A1(n6968), .A2(n8724), .ZN(n5868) );
  NAND2_X1 U7262 ( .A1(n6968), .A2(n8724), .ZN(n5791) );
  NAND2_X1 U7263 ( .A1(n5868), .A2(n5791), .ZN(n8563) );
  NAND2_X1 U7264 ( .A1(n5792), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5793) );
  XNOR2_X1 U7265 ( .A(n5793), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8519) );
  INV_X1 U7266 ( .A(n8519), .ZN(n6885) );
  INV_X1 U7267 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7268 ( .A1(n5794), .A2(n5795), .ZN(n5850) );
  OR2_X1 U7269 ( .A1(n5850), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7270 ( .A1(n5816), .A2(n5796), .ZN(n5797) );
  NOR2_X1 U7271 ( .A1(n5815), .A2(n5797), .ZN(n5810) );
  NAND2_X1 U7272 ( .A1(n5810), .A2(n5798), .ZN(n5812) );
  OR2_X1 U7273 ( .A1(n5812), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7274 ( .A1(n5799), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5807) );
  INV_X1 U7275 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U7276 ( .A1(n5807), .A2(n5800), .ZN(n5801) );
  NAND2_X1 U7277 ( .A1(n5801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7278 ( .A1(n5804), .A2(n5803), .ZN(n5806) );
  NAND2_X1 U7279 ( .A1(n5806), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5802) );
  XNOR2_X1 U7280 ( .A(n5802), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8502) );
  OR2_X1 U7281 ( .A1(n5804), .A2(n5803), .ZN(n5805) );
  NAND2_X1 U7282 ( .A1(n5806), .A2(n5805), .ZN(n6654) );
  XNOR2_X1 U7283 ( .A(n5807), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U7284 ( .A1(n5812), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5809) );
  XNOR2_X1 U7285 ( .A(n5809), .B(n5808), .ZN(n6538) );
  NOR2_X1 U7286 ( .A1(n5810), .A2(n5846), .ZN(n5811) );
  MUX2_X1 U7287 ( .A(n5846), .B(n5811), .S(P2_IR_REG_11__SCAN_IN), .Z(n5814)
         );
  INV_X1 U7288 ( .A(n5812), .ZN(n5813) );
  OR2_X1 U7289 ( .A1(n5814), .A2(n5813), .ZN(n6445) );
  INV_X1 U7290 ( .A(n6445), .ZN(n7349) );
  NAND2_X1 U7291 ( .A1(n5815), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U7292 ( .A1(n5819), .A2(n5816), .ZN(n5817) );
  NAND2_X1 U7293 ( .A1(n5817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5818) );
  XNOR2_X1 U7294 ( .A(n5818), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7316) );
  INV_X1 U7295 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7380) );
  INV_X1 U7296 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7294) );
  XNOR2_X1 U7297 ( .A(n5819), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7161) );
  INV_X1 U7298 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5824) );
  OR2_X1 U7299 ( .A1(n5837), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5842) );
  OAI21_X1 U7300 ( .B1(n5842), .B2(P2_IR_REG_5__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5821) );
  MUX2_X1 U7301 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5821), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5823) );
  INV_X1 U7302 ( .A(n5794), .ZN(n5822) );
  MUX2_X1 U7303 ( .A(n5824), .B(P2_REG2_REG_6__SCAN_IN), .S(n6703), .Z(n6696)
         );
  INV_X1 U7304 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5828) );
  MUX2_X1 U7305 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n5828), .S(n5833), .Z(n9988)
         );
  INV_X1 U7306 ( .A(n5825), .ZN(n5829) );
  INV_X1 U7307 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5917) );
  NOR2_X1 U7308 ( .A1(n5917), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U7309 ( .A1(n5825), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5832) );
  INV_X1 U7310 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6625) );
  OR2_X1 U7311 ( .A1(n6626), .A2(n6625), .ZN(n6628) );
  NAND2_X1 U7312 ( .A1(n6628), .A2(n5832), .ZN(n9987) );
  NAND2_X1 U7313 ( .A1(n9988), .A2(n9987), .ZN(n9986) );
  NAND2_X1 U7314 ( .A1(n4286), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5834) );
  INV_X1 U7315 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6993) );
  NAND2_X1 U7316 ( .A1(n5837), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5839) );
  INV_X1 U7317 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5838) );
  INV_X1 U7318 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6889) );
  XNOR2_X1 U7319 ( .A(n6623), .B(n6889), .ZN(n6611) );
  NAND2_X1 U7320 ( .A1(n5840), .A2(n6611), .ZN(n6615) );
  NAND2_X1 U7321 ( .A1(n6623), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U7322 ( .A1(n6615), .A2(n5841), .ZN(n5844) );
  NAND2_X1 U7323 ( .A1(n5842), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5843) );
  XNOR2_X1 U7324 ( .A(n5843), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6585) );
  INV_X1 U7325 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6869) );
  NAND2_X1 U7326 ( .A1(n6574), .A2(n4715), .ZN(n6695) );
  NAND2_X1 U7327 ( .A1(n6696), .A2(n6695), .ZN(n6694) );
  INV_X1 U7328 ( .A(n6703), .ZN(n6386) );
  NAND2_X1 U7329 ( .A1(n6386), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7330 ( .A1(n6694), .A2(n5845), .ZN(n5848) );
  OR2_X1 U7331 ( .A1(n5794), .A2(n5846), .ZN(n5847) );
  XNOR2_X1 U7332 ( .A(n5847), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6842) );
  INV_X1 U7333 ( .A(n6842), .ZN(n6398) );
  NAND2_X1 U7334 ( .A1(n5848), .A2(n6398), .ZN(n5849) );
  OAI21_X1 U7335 ( .B1(n5848), .B2(n6398), .A(n5849), .ZN(n6835) );
  INV_X1 U7336 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7132) );
  INV_X1 U7337 ( .A(n5849), .ZN(n6944) );
  INV_X1 U7338 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U7339 ( .A1(n5850), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5851) );
  XNOR2_X1 U7340 ( .A(n5851), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6958) );
  MUX2_X1 U7341 ( .A(n5852), .B(P2_REG2_REG_8__SCAN_IN), .S(n6958), .Z(n6943)
         );
  INV_X1 U7342 ( .A(n6958), .ZN(n5915) );
  NAND2_X1 U7343 ( .A1(n5915), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5853) );
  MUX2_X1 U7344 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7380), .S(n7316), .Z(n7322)
         );
  NAND2_X1 U7345 ( .A1(n5855), .A2(n6445), .ZN(n5856) );
  OR2_X1 U7346 ( .A1(n6538), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7347 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6538), .ZN(n5857) );
  NAND2_X1 U7348 ( .A1(n5858), .A2(n5857), .ZN(n7416) );
  NOR2_X1 U7349 ( .A1(n8467), .A2(n5859), .ZN(n5860) );
  INV_X1 U7350 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8958) );
  NOR2_X1 U7351 ( .A1(n8958), .A2(n8460), .ZN(n8459) );
  NAND2_X1 U7352 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6654), .ZN(n5861) );
  OAI21_X1 U7353 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n6654), .A(n5861), .ZN(
        n8486) );
  NOR2_X1 U7354 ( .A1(n8502), .A2(n5862), .ZN(n5863) );
  INV_X1 U7355 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8917) );
  INV_X1 U7356 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8937) );
  NOR2_X1 U7357 ( .A1(n6885), .A2(n8937), .ZN(n5864) );
  AOI21_X1 U7358 ( .B1(n8937), .B2(n6885), .A(n5864), .ZN(n8525) );
  NAND2_X1 U7359 ( .A1(n5865), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5866) );
  XNOR2_X1 U7360 ( .A(n5866), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8543) );
  INV_X1 U7361 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8537) );
  NOR2_X1 U7362 ( .A1(n5867), .A2(n8535), .ZN(n8564) );
  INV_X1 U7363 ( .A(n5868), .ZN(n5869) );
  NAND2_X1 U7364 ( .A1(n5870), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5950) );
  INV_X1 U7365 ( .A(n7657), .ZN(n7979) );
  INV_X1 U7366 ( .A(n5871), .ZN(n5900) );
  NAND2_X1 U7367 ( .A1(n7979), .A2(n5900), .ZN(n6302) );
  OR2_X1 U7368 ( .A1(n5950), .A2(n6302), .ZN(n8565) );
  INV_X1 U7369 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8802) );
  OR2_X1 U7370 ( .A1(n6968), .A2(n8802), .ZN(n5897) );
  NAND2_X1 U7371 ( .A1(n6968), .A2(n8802), .ZN(n5872) );
  NAND2_X1 U7372 ( .A1(n5897), .A2(n5872), .ZN(n8556) );
  OAI21_X1 U7373 ( .B1(n4286), .B2(n10085), .A(n5873), .ZN(n9998) );
  AND2_X1 U7374 ( .A1(n4404), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7375 ( .A1(n5825), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5875) );
  INV_X1 U7376 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U7377 ( .A1(n4286), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5876) );
  INV_X1 U7378 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10087) );
  XNOR2_X1 U7379 ( .A(n6623), .B(n10089), .ZN(n6605) );
  NAND2_X1 U7380 ( .A1(n5877), .A2(n6605), .ZN(n6610) );
  NAND2_X1 U7381 ( .A1(n6623), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7382 ( .A1(n6610), .A2(n5878), .ZN(n5879) );
  OAI21_X1 U7383 ( .B1(n5879), .B2(n6384), .A(n5880), .ZN(n6579) );
  INV_X1 U7384 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10091) );
  NOR2_X1 U7385 ( .A1(n6579), .A2(n10091), .ZN(n6578) );
  INV_X1 U7386 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10093) );
  MUX2_X1 U7387 ( .A(n10093), .B(P2_REG1_REG_6__SCAN_IN), .S(n6703), .Z(n6693)
         );
  NAND2_X1 U7388 ( .A1(n6386), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5882) );
  INV_X1 U7389 ( .A(n6833), .ZN(n5883) );
  INV_X1 U7390 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10095) );
  NAND2_X1 U7391 ( .A1(n5883), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6832) );
  INV_X1 U7392 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10097) );
  MUX2_X1 U7393 ( .A(n10097), .B(P2_REG1_REG_8__SCAN_IN), .S(n6958), .Z(n6950)
         );
  INV_X1 U7394 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10099) );
  INV_X1 U7395 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10101) );
  INV_X1 U7396 ( .A(n7316), .ZN(n6416) );
  AOI22_X1 U7397 ( .A1(n7316), .A2(P2_REG1_REG_10__SCAN_IN), .B1(n10101), .B2(
        n6416), .ZN(n7312) );
  NOR2_X1 U7398 ( .A1(n7316), .A2(n10101), .ZN(n5884) );
  INV_X1 U7399 ( .A(n5885), .ZN(n5887) );
  INV_X1 U7400 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10103) );
  OAI21_X1 U7401 ( .B1(n5886), .B2(n6445), .A(n5885), .ZN(n7345) );
  NAND2_X1 U7402 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6538), .ZN(n5888) );
  OAI21_X1 U7403 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n6538), .A(n5888), .ZN(
        n7410) );
  NOR2_X1 U7404 ( .A1(n8467), .A2(n5889), .ZN(n5890) );
  INV_X1 U7405 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9752) );
  INV_X1 U7406 ( .A(n8467), .ZN(n6550) );
  NAND2_X1 U7407 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6654), .ZN(n5891) );
  OAI21_X1 U7408 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n6654), .A(n5891), .ZN(
        n8476) );
  NOR2_X1 U7409 ( .A1(n8502), .A2(n5892), .ZN(n5893) );
  INV_X1 U7410 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8498) );
  INV_X1 U7411 ( .A(n8502), .ZN(n6711) );
  INV_X1 U7412 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n5894) );
  AOI22_X1 U7413 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8519), .B1(n6885), .B2(
        n5894), .ZN(n8514) );
  INV_X1 U7414 ( .A(n8543), .ZN(n6965) );
  INV_X1 U7415 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8805) );
  INV_X1 U7416 ( .A(n5895), .ZN(n5896) );
  INV_X1 U7417 ( .A(n5897), .ZN(n5898) );
  XNOR2_X1 U7418 ( .A(n7193), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n5946) );
  XNOR2_X1 U7419 ( .A(n5899), .B(n5946), .ZN(n5904) );
  NOR2_X1 U7420 ( .A1(n5950), .A2(n7657), .ZN(n6640) );
  INV_X2 U7421 ( .A(n5900), .ZN(n7978) );
  NAND2_X1 U7422 ( .A1(n6640), .A2(n7978), .ZN(n8559) );
  INV_X1 U7423 ( .A(n8559), .ZN(n10000) );
  INV_X1 U7424 ( .A(n6712), .ZN(n5901) );
  NOR2_X1 U7425 ( .A1(n6423), .A2(n5901), .ZN(n5902) );
  OR2_X1 U7426 ( .A1(P2_U3150), .A2(n5902), .ZN(n8561) );
  INV_X1 U7427 ( .A(n8561), .ZN(n9991) );
  NAND2_X1 U7428 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8325) );
  MUX2_X1 U7429 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n7978), .Z(n5943) );
  XNOR2_X1 U7430 ( .A(n5943), .B(n8543), .ZN(n8546) );
  MUX2_X1 U7431 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n7978), .Z(n5906) );
  OR2_X1 U7432 ( .A1(n5906), .A2(n6885), .ZN(n5942) );
  XNOR2_X1 U7433 ( .A(n5906), .B(n8519), .ZN(n8518) );
  MUX2_X1 U7434 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n7978), .Z(n5907) );
  OR2_X1 U7435 ( .A1(n5907), .A2(n6711), .ZN(n5941) );
  XNOR2_X1 U7436 ( .A(n8502), .B(n5907), .ZN(n8505) );
  MUX2_X1 U7437 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n7978), .Z(n5908) );
  OR2_X1 U7438 ( .A1(n5908), .A2(n6654), .ZN(n5940) );
  INV_X1 U7439 ( .A(n6654), .ZN(n8481) );
  XNOR2_X1 U7440 ( .A(n5908), .B(n8481), .ZN(n8480) );
  MUX2_X1 U7441 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n7978), .Z(n5909) );
  OR2_X1 U7442 ( .A1(n5909), .A2(n6550), .ZN(n5939) );
  XNOR2_X1 U7443 ( .A(n5909), .B(n8467), .ZN(n8470) );
  MUX2_X1 U7444 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n7978), .Z(n5910) );
  OR2_X1 U7445 ( .A1(n5910), .A2(n6538), .ZN(n5938) );
  INV_X1 U7446 ( .A(n6538), .ZN(n7418) );
  XNOR2_X1 U7447 ( .A(n5910), .B(n7418), .ZN(n7414) );
  MUX2_X1 U7448 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n7978), .Z(n5911) );
  OR2_X1 U7449 ( .A1(n5911), .A2(n6445), .ZN(n5937) );
  XNOR2_X1 U7450 ( .A(n5911), .B(n7349), .ZN(n7348) );
  MUX2_X1 U7451 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n7978), .Z(n5912) );
  OR2_X1 U7452 ( .A1(n5912), .A2(n6416), .ZN(n5936) );
  XNOR2_X1 U7453 ( .A(n5912), .B(n7316), .ZN(n7315) );
  MUX2_X1 U7454 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n7978), .Z(n5914) );
  INV_X1 U7455 ( .A(n5914), .ZN(n5913) );
  NAND2_X1 U7456 ( .A1(n7161), .A2(n5913), .ZN(n5935) );
  XNOR2_X1 U7457 ( .A(n5914), .B(n7161), .ZN(n7160) );
  MUX2_X1 U7458 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n7978), .Z(n5933) );
  OR2_X1 U7459 ( .A1(n5933), .A2(n5915), .ZN(n5934) );
  MUX2_X1 U7460 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n7978), .Z(n5930) );
  INV_X1 U7461 ( .A(n5930), .ZN(n5931) );
  MUX2_X1 U7462 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n7978), .Z(n5928) );
  INV_X1 U7463 ( .A(n5928), .ZN(n5929) );
  INV_X1 U7464 ( .A(n6623), .ZN(n5927) );
  MUX2_X1 U7465 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n7978), .Z(n5925) );
  INV_X1 U7466 ( .A(n5925), .ZN(n5926) );
  MUX2_X1 U7467 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n7978), .Z(n5923) );
  INV_X1 U7468 ( .A(n5923), .ZN(n5924) );
  INV_X1 U7469 ( .A(n4286), .ZN(n5922) );
  MUX2_X1 U7470 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n7978), .Z(n5920) );
  INV_X1 U7471 ( .A(n5920), .ZN(n5921) );
  MUX2_X1 U7472 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n7978), .Z(n5918) );
  INV_X1 U7473 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10081) );
  MUX2_X1 U7474 ( .A(n5917), .B(n10081), .S(n7978), .Z(n6638) );
  NAND2_X1 U7475 ( .A1(n6638), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6637) );
  NAND2_X1 U7476 ( .A1(n6634), .A2(n5919), .ZN(n9984) );
  XNOR2_X1 U7477 ( .A(n5920), .B(n5922), .ZN(n9983) );
  NAND2_X1 U7478 ( .A1(n9984), .A2(n9983), .ZN(n9982) );
  OAI21_X1 U7479 ( .B1(n5922), .B2(n5921), .A(n9982), .ZN(n6589) );
  XNOR2_X1 U7480 ( .A(n5923), .B(n6381), .ZN(n6590) );
  NOR2_X1 U7481 ( .A1(n6589), .A2(n6590), .ZN(n6588) );
  XOR2_X1 U7482 ( .A(n6623), .B(n5925), .Z(n6603) );
  XNOR2_X1 U7483 ( .A(n5928), .B(n6585), .ZN(n6572) );
  OAI21_X1 U7484 ( .B1(n6585), .B2(n5929), .A(n6571), .ZN(n6689) );
  XOR2_X1 U7485 ( .A(n6703), .B(n5930), .Z(n6690) );
  NOR2_X1 U7486 ( .A1(n6689), .A2(n6690), .ZN(n6688) );
  AOI21_X1 U7487 ( .B1(n6703), .B2(n5931), .A(n6688), .ZN(n6830) );
  MUX2_X1 U7488 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n7978), .Z(n5932) );
  XOR2_X1 U7489 ( .A(n6842), .B(n5932), .Z(n6831) );
  OAI22_X1 U7490 ( .A1(n6830), .A2(n6831), .B1(n5932), .B2(n6398), .ZN(n6941)
         );
  XNOR2_X1 U7491 ( .A(n5933), .B(n6958), .ZN(n6940) );
  NAND2_X1 U7492 ( .A1(n6941), .A2(n6940), .ZN(n6939) );
  NAND2_X1 U7493 ( .A1(n5934), .A2(n6939), .ZN(n7159) );
  NAND2_X1 U7494 ( .A1(n7348), .A2(n7347), .ZN(n7346) );
  NAND2_X1 U7495 ( .A1(n5937), .A2(n7346), .ZN(n7413) );
  NAND2_X1 U7496 ( .A1(n8480), .A2(n8479), .ZN(n8478) );
  NAND2_X1 U7497 ( .A1(n5940), .A2(n8478), .ZN(n8504) );
  NAND2_X1 U7498 ( .A1(n8546), .A2(n8545), .ZN(n8544) );
  OAI21_X1 U7499 ( .B1(n5943), .B2(n6965), .A(n8544), .ZN(n5945) );
  MUX2_X1 U7500 ( .A(n8724), .B(n8802), .S(n7978), .Z(n5944) );
  INV_X1 U7501 ( .A(n6968), .ZN(n8569) );
  NAND2_X1 U7502 ( .A1(n5945), .A2(n5944), .ZN(n8552) );
  OAI21_X1 U7503 ( .B1(n8551), .B2(n8569), .A(n8552), .ZN(n5949) );
  MUX2_X1 U7504 ( .A(n5947), .B(n5946), .S(n7978), .Z(n5948) );
  XNOR2_X1 U7505 ( .A(n5949), .B(n5948), .ZN(n5954) );
  AND2_X1 U7506 ( .A1(n7657), .A2(P2_U3893), .ZN(n9981) );
  INV_X1 U7507 ( .A(n9981), .ZN(n6844) );
  INV_X1 U7508 ( .A(n5950), .ZN(n5951) );
  MUX2_X1 U7509 ( .A(n5951), .B(P2_U3893), .S(n7979), .Z(n5952) );
  AND2_X1 U7510 ( .A1(n5952), .A2(n6308), .ZN(n8553) );
  INV_X1 U7511 ( .A(n7193), .ZN(n7803) );
  INV_X1 U7512 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7513 ( .A1(n5985), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7514 ( .A1(n6002), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5963) );
  OR2_X1 U7515 ( .A1(n5991), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5969) );
  OR2_X1 U7516 ( .A1(n5990), .A2(n5967), .ZN(n5968) );
  INV_X1 U7518 ( .A(n6459), .ZN(n6257) );
  NAND2_X1 U7519 ( .A1(n6926), .A2(n6459), .ZN(n7824) );
  NAND2_X1 U7520 ( .A1(n6002), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5974) );
  OR2_X1 U7521 ( .A1(n5992), .A2(n10081), .ZN(n5973) );
  NAND2_X1 U7522 ( .A1(n6125), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7523 ( .A1(n5993), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5971) );
  INV_X1 U7524 ( .A(n6849), .ZN(n6460) );
  NAND2_X1 U7525 ( .A1(n4471), .A2(SI_0_), .ZN(n5976) );
  INV_X1 U7526 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7527 ( .A1(n5976), .A2(n5975), .ZN(n5978) );
  AND2_X1 U7528 ( .A1(n5978), .A2(n5977), .ZN(n9036) );
  MUX2_X1 U7529 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9036), .S(n6308), .Z(n10007)
         );
  NAND2_X1 U7530 ( .A1(n5993), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7531 ( .A1(n5985), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7532 ( .A1(n6125), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7533 ( .A1(n6002), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5979) );
  OR2_X1 U7534 ( .A1(n5991), .A2(n6363), .ZN(n5984) );
  OR2_X1 U7535 ( .A1(n5990), .A2(n6377), .ZN(n5983) );
  OAI211_X1 U7536 ( .C1(n6308), .C2(n4286), .A(n5984), .B(n5983), .ZN(n6521)
         );
  NAND2_X1 U7537 ( .A1(n6986), .A2(n6521), .ZN(n7832) );
  NAND2_X1 U7538 ( .A1(n5985), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7539 ( .A1(n6125), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5988) );
  INV_X1 U7540 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U7541 ( .A1(n5993), .A2(n6990), .ZN(n5987) );
  NAND2_X1 U7542 ( .A1(n6002), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7543 ( .A1(n6925), .A2(n6991), .ZN(n7847) );
  NAND2_X1 U7544 ( .A1(n7847), .A2(n7841), .ZN(n6258) );
  NAND2_X1 U7545 ( .A1(n6989), .A2(n6259), .ZN(n6988) );
  NAND2_X1 U7546 ( .A1(n6988), .A2(n7847), .ZN(n6886) );
  NAND2_X1 U7547 ( .A1(n6002), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7548 ( .A1(n7758), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5997) );
  AND2_X1 U7549 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5994) );
  OR2_X1 U7550 ( .A1(n5994), .A2(n6003), .ZN(n6890) );
  NAND2_X1 U7551 ( .A1(n6227), .A2(n6890), .ZN(n5996) );
  NAND2_X1 U7552 ( .A1(n6125), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5995) );
  OR2_X1 U7553 ( .A1(n5990), .A2(n6388), .ZN(n6000) );
  OR2_X1 U7554 ( .A1(n5991), .A2(n6387), .ZN(n5999) );
  INV_X1 U7555 ( .A(n6891), .ZN(n6264) );
  NAND2_X1 U7556 ( .A1(n8452), .A2(n6264), .ZN(n7849) );
  NAND2_X1 U7557 ( .A1(n6886), .A2(n7849), .ZN(n6001) );
  NAND2_X1 U7558 ( .A1(n6987), .A2(n6891), .ZN(n7844) );
  NAND2_X1 U7559 ( .A1(n7758), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7560 ( .A1(n6243), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7561 ( .A1(n6003), .A2(n6004), .ZN(n6014) );
  OR2_X1 U7562 ( .A1(n6004), .A2(n6003), .ZN(n6005) );
  NAND2_X1 U7563 ( .A1(n6014), .A2(n6005), .ZN(n6730) );
  NAND2_X1 U7564 ( .A1(n5993), .A2(n6730), .ZN(n6007) );
  NAND2_X1 U7565 ( .A1(n6125), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6006) );
  NAND4_X1 U7566 ( .A1(n6009), .A2(n6008), .A3(n6007), .A4(n6006), .ZN(n8451)
         );
  INV_X1 U7567 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U7568 ( .A1(n6369), .A2(n6028), .ZN(n6011) );
  NAND2_X1 U7569 ( .A1(n6131), .A2(n6585), .ZN(n6010) );
  OAI211_X1 U7570 ( .C1(n5991), .C2(n6382), .A(n6011), .B(n6010), .ZN(n6744)
         );
  INV_X1 U7571 ( .A(n6744), .ZN(n6867) );
  NAND2_X1 U7572 ( .A1(n8451), .A2(n6867), .ZN(n7848) );
  NAND2_X1 U7573 ( .A1(n6766), .A2(n6744), .ZN(n7842) );
  NAND2_X1 U7574 ( .A1(n6371), .A2(n6028), .ZN(n6012) );
  NAND2_X1 U7575 ( .A1(n7758), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6019) );
  INV_X2 U7576 ( .A(n6013), .ZN(n7759) );
  NAND2_X1 U7577 ( .A1(n7759), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7578 ( .A1(n6014), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7579 ( .A1(n6020), .A2(n6015), .ZN(n7049) );
  NAND2_X1 U7580 ( .A1(n6227), .A2(n7049), .ZN(n6017) );
  NAND2_X1 U7581 ( .A1(n6125), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6016) );
  NOR2_X1 U7582 ( .A1(n10039), .A2(n8450), .ZN(n7846) );
  NAND2_X1 U7583 ( .A1(n10039), .A2(n8450), .ZN(n7852) );
  NAND2_X1 U7584 ( .A1(n7758), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6025) );
  NAND2_X1 U7585 ( .A1(n6243), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6024) );
  AND2_X1 U7586 ( .A1(n6020), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6021) );
  OR2_X1 U7587 ( .A1(n6021), .A2(n6032), .ZN(n7131) );
  NAND2_X1 U7588 ( .A1(n6227), .A2(n7131), .ZN(n6023) );
  NAND2_X1 U7589 ( .A1(n6125), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7590 ( .A1(n6394), .A2(n6028), .ZN(n6027) );
  AOI22_X1 U7591 ( .A1(n6132), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6131), .B2(
        n6842), .ZN(n6026) );
  NAND2_X1 U7592 ( .A1(n6027), .A2(n6026), .ZN(n6905) );
  OR2_X1 U7593 ( .A1(n7072), .A2(n6905), .ZN(n7074) );
  NAND2_X1 U7594 ( .A1(n6905), .A2(n7072), .ZN(n7865) );
  NAND2_X1 U7595 ( .A1(n7124), .A2(n7778), .ZN(n7073) );
  NAND2_X1 U7596 ( .A1(n6399), .A2(n7755), .ZN(n6030) );
  AOI22_X1 U7597 ( .A1(n6132), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6131), .B2(
        n6958), .ZN(n6029) );
  NAND2_X1 U7598 ( .A1(n6030), .A2(n6029), .ZN(n6997) );
  NAND2_X1 U7599 ( .A1(n7758), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7600 ( .A1(n7759), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6036) );
  INV_X1 U7601 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6031) );
  NOR2_X1 U7602 ( .A1(n6032), .A2(n6031), .ZN(n6033) );
  OR2_X1 U7603 ( .A1(n6041), .A2(n6033), .ZN(n7077) );
  NAND2_X1 U7604 ( .A1(n6227), .A2(n7077), .ZN(n6035) );
  NAND2_X1 U7605 ( .A1(n6125), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6034) );
  OR2_X1 U7606 ( .A1(n6997), .A2(n7271), .ZN(n7856) );
  AND2_X1 U7607 ( .A1(n7856), .A2(n7074), .ZN(n7864) );
  NAND2_X1 U7608 ( .A1(n6997), .A2(n7271), .ZN(n7866) );
  NAND2_X1 U7609 ( .A1(n6409), .A2(n7755), .ZN(n6039) );
  AOI22_X1 U7610 ( .A1(n6132), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6131), .B2(
        n7161), .ZN(n6038) );
  NAND2_X1 U7611 ( .A1(n6039), .A2(n6038), .ZN(n10055) );
  NAND2_X1 U7612 ( .A1(n7758), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7613 ( .A1(n6243), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6045) );
  INV_X2 U7614 ( .A(n6242), .ZN(n6227) );
  INV_X1 U7615 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6040) );
  OR2_X1 U7616 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  NAND2_X1 U7617 ( .A1(n6050), .A2(n6042), .ZN(n7267) );
  NAND2_X1 U7618 ( .A1(n6227), .A2(n7267), .ZN(n6044) );
  NAND2_X1 U7619 ( .A1(n6125), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6043) );
  NAND4_X1 U7620 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n8447)
         );
  OR2_X1 U7621 ( .A1(n10055), .A2(n7374), .ZN(n7859) );
  NAND2_X1 U7622 ( .A1(n10055), .A2(n7374), .ZN(n7867) );
  NAND2_X1 U7623 ( .A1(n7859), .A2(n7867), .ZN(n7288) );
  NAND2_X1 U7624 ( .A1(n6413), .A2(n7755), .ZN(n6049) );
  AOI22_X1 U7625 ( .A1(n6132), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6131), .B2(
        n7316), .ZN(n6048) );
  NAND2_X1 U7626 ( .A1(n6049), .A2(n6048), .ZN(n10061) );
  NAND2_X1 U7627 ( .A1(n7758), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7628 ( .A1(n7759), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7629 ( .A1(n6050), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7630 ( .A1(n6059), .A2(n6051), .ZN(n7378) );
  NAND2_X1 U7631 ( .A1(n6227), .A2(n7378), .ZN(n6053) );
  NAND2_X1 U7632 ( .A1(n6125), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6052) );
  NAND4_X1 U7633 ( .A1(n6055), .A2(n6054), .A3(n6053), .A4(n6052), .ZN(n8446)
         );
  OR2_X1 U7634 ( .A1(n10061), .A2(n7531), .ZN(n7878) );
  AND2_X1 U7635 ( .A1(n7878), .A2(n7859), .ZN(n7863) );
  NAND2_X1 U7636 ( .A1(n7285), .A2(n7863), .ZN(n6056) );
  NAND2_X1 U7637 ( .A1(n10061), .A2(n7531), .ZN(n7875) );
  NAND2_X1 U7638 ( .A1(n6056), .A2(n7875), .ZN(n7395) );
  NAND2_X1 U7639 ( .A1(n6441), .A2(n7755), .ZN(n6058) );
  AOI22_X1 U7640 ( .A1(n6132), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6131), .B2(
        n7349), .ZN(n6057) );
  NAND2_X1 U7641 ( .A1(n7759), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7642 ( .A1(n6125), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7643 ( .A1(n6059), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7644 ( .A1(n6068), .A2(n6060), .ZN(n7527) );
  NAND2_X1 U7645 ( .A1(n6227), .A2(n7527), .ZN(n6062) );
  NAND2_X1 U7646 ( .A1(n7758), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6061) );
  NAND4_X1 U7647 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n8445)
         );
  XNOR2_X1 U7648 ( .A(n7526), .B(n8445), .ZN(n7771) );
  NAND2_X1 U7649 ( .A1(n7395), .A2(n7771), .ZN(n6065) );
  INV_X1 U7650 ( .A(n8445), .ZN(n7489) );
  NAND2_X1 U7651 ( .A1(n7526), .A2(n7489), .ZN(n7880) );
  NAND2_X1 U7652 ( .A1(n6527), .A2(n7755), .ZN(n6067) );
  AOI22_X1 U7653 ( .A1(n6132), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6131), .B2(
        n7418), .ZN(n6066) );
  NAND2_X1 U7654 ( .A1(n7759), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7655 ( .A1(n6125), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6072) );
  AND2_X1 U7656 ( .A1(n6068), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6069) );
  OR2_X1 U7657 ( .A1(n6069), .A2(n6077), .ZN(n7491) );
  NAND2_X1 U7658 ( .A1(n6227), .A2(n7491), .ZN(n6071) );
  NAND2_X1 U7659 ( .A1(n7758), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6070) );
  NAND4_X1 U7660 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(n8444)
         );
  INV_X1 U7661 ( .A(n8444), .ZN(n7559) );
  NAND2_X1 U7662 ( .A1(n10071), .A2(n7559), .ZN(n7886) );
  NAND2_X1 U7663 ( .A1(n7885), .A2(n7886), .ZN(n7888) );
  INV_X1 U7664 ( .A(n7888), .ZN(n6074) );
  NAND2_X1 U7665 ( .A1(n6546), .A2(n7755), .ZN(n6076) );
  AOI22_X1 U7666 ( .A1(n6132), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6131), .B2(
        n8467), .ZN(n6075) );
  INV_X1 U7667 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7550) );
  NAND2_X1 U7668 ( .A1(n6077), .A2(n7550), .ZN(n6086) );
  OR2_X1 U7669 ( .A1(n6077), .A2(n7550), .ZN(n6078) );
  NAND2_X1 U7670 ( .A1(n6086), .A2(n6078), .ZN(n7561) );
  NAND2_X1 U7671 ( .A1(n6227), .A2(n7561), .ZN(n6082) );
  NAND2_X1 U7672 ( .A1(n7759), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7673 ( .A1(n6125), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7674 ( .A1(n7758), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6079) );
  XNOR2_X1 U7675 ( .A(n7556), .B(n7575), .ZN(n7562) );
  NAND2_X1 U7676 ( .A1(n7556), .A2(n7575), .ZN(n7890) );
  NAND2_X1 U7677 ( .A1(n7563), .A2(n7890), .ZN(n7571) );
  NAND2_X1 U7678 ( .A1(n6652), .A2(n7755), .ZN(n6085) );
  AOI22_X1 U7679 ( .A1(n6132), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6131), .B2(
        n8481), .ZN(n6084) );
  NAND2_X1 U7680 ( .A1(n7759), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7681 ( .A1(n7758), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7682 ( .A1(n6125), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7683 ( .A1(n6086), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6087) );
  AND2_X1 U7684 ( .A1(n6097), .A2(n6087), .ZN(n9747) );
  INV_X1 U7685 ( .A(n9747), .ZN(n7577) );
  NAND2_X1 U7686 ( .A1(n6227), .A2(n7577), .ZN(n6088) );
  NAND4_X1 U7687 ( .A1(n6091), .A2(n6090), .A3(n6089), .A4(n6088), .ZN(n8443)
         );
  INV_X1 U7688 ( .A(n8443), .ZN(n8249) );
  OR2_X1 U7689 ( .A1(n8248), .A2(n8249), .ZN(n7893) );
  NAND2_X1 U7690 ( .A1(n8248), .A2(n8249), .ZN(n7894) );
  INV_X1 U7691 ( .A(n7894), .ZN(n6092) );
  NAND2_X1 U7692 ( .A1(n6673), .A2(n7755), .ZN(n6094) );
  AOI22_X1 U7693 ( .A1(n6132), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8502), .B2(
        n6131), .ZN(n6093) );
  NAND2_X1 U7694 ( .A1(n6243), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7695 ( .A1(n7758), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6101) );
  INV_X1 U7696 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7697 ( .A1(n6097), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7698 ( .A1(n6106), .A2(n6098), .ZN(n8435) );
  NAND2_X1 U7699 ( .A1(n6227), .A2(n8435), .ZN(n6100) );
  NAND2_X1 U7700 ( .A1(n6125), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7701 ( .A1(n8253), .A2(n9733), .ZN(n6103) );
  NAND2_X1 U7702 ( .A1(n7626), .A2(n7896), .ZN(n7625) );
  NAND2_X1 U7703 ( .A1(n7625), .A2(n7899), .ZN(n8745) );
  NAND2_X1 U7704 ( .A1(n6881), .A2(n7755), .ZN(n6105) );
  AOI22_X1 U7705 ( .A1(n6132), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6131), .B2(
        n8519), .ZN(n6104) );
  NAND2_X1 U7706 ( .A1(n7759), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7707 ( .A1(n7758), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6110) );
  OR2_X2 U7708 ( .A1(n6106), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7709 ( .A1(n6106), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7710 ( .A1(n6118), .A2(n6107), .ZN(n8760) );
  NAND2_X1 U7711 ( .A1(n6227), .A2(n8760), .ZN(n6109) );
  NAND2_X1 U7712 ( .A1(n6125), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7713 ( .A1(n8809), .A2(n8432), .ZN(n7902) );
  NAND2_X1 U7714 ( .A1(n7901), .A2(n7902), .ZN(n7785) );
  INV_X1 U7715 ( .A(n7785), .ZN(n8749) );
  NAND2_X1 U7716 ( .A1(n8745), .A2(n8749), .ZN(n8747) );
  NAND2_X1 U7717 ( .A1(n6961), .A2(n7755), .ZN(n6113) );
  AOI22_X1 U7718 ( .A1(n6132), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6131), .B2(
        n8543), .ZN(n6112) );
  NAND2_X1 U7719 ( .A1(n7759), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7720 ( .A1(n6125), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6114) );
  AND2_X1 U7721 ( .A1(n6115), .A2(n6114), .ZN(n6122) );
  INV_X1 U7722 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7723 ( .A1(n6118), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7724 ( .A1(n6135), .A2(n6119), .ZN(n8732) );
  NAND2_X1 U7725 ( .A1(n8732), .A2(n6227), .ZN(n6121) );
  NAND2_X1 U7726 ( .A1(n7758), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6120) );
  OR2_X1 U7727 ( .A1(n9018), .A2(n8755), .ZN(n7904) );
  NAND2_X1 U7728 ( .A1(n9018), .A2(n8755), .ZN(n7814) );
  NAND2_X1 U7729 ( .A1(n7904), .A2(n7814), .ZN(n8731) );
  NAND2_X1 U7730 ( .A1(n6966), .A2(n7755), .ZN(n6124) );
  AOI22_X1 U7731 ( .A1(n6132), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6131), .B2(
        n6968), .ZN(n6123) );
  XNOR2_X1 U7732 ( .A(n6135), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U7733 ( .A1(n8725), .A2(n6227), .ZN(n6130) );
  INV_X1 U7734 ( .A(n6125), .ZN(n6305) );
  NAND2_X1 U7735 ( .A1(n7759), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7736 ( .A1(n7758), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6126) );
  OAI211_X1 U7737 ( .C1(n8724), .C2(n6305), .A(n6127), .B(n6126), .ZN(n6128)
         );
  INV_X1 U7738 ( .A(n6128), .ZN(n6129) );
  NAND2_X1 U7739 ( .A1(n6130), .A2(n6129), .ZN(n8738) );
  INV_X1 U7740 ( .A(n8738), .ZN(n8705) );
  NAND2_X1 U7741 ( .A1(n9012), .A2(n8705), .ZN(n7912) );
  NAND2_X1 U7742 ( .A1(n7905), .A2(n7912), .ZN(n7770) );
  NAND2_X1 U7743 ( .A1(n8717), .A2(n7905), .ZN(n8708) );
  NAND2_X1 U7744 ( .A1(n7191), .A2(n7755), .ZN(n6134) );
  AOI22_X1 U7745 ( .A1(n6132), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7803), .B2(
        n6131), .ZN(n6133) );
  INV_X1 U7746 ( .A(n6135), .ZN(n6136) );
  INV_X1 U7747 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8409) );
  INV_X1 U7748 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6137) );
  INV_X1 U7749 ( .A(n6138), .ZN(n6139) );
  NAND2_X1 U7750 ( .A1(n6139), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7751 ( .A1(n6146), .A2(n6140), .ZN(n8711) );
  NAND2_X1 U7752 ( .A1(n8711), .A2(n6227), .ZN(n6143) );
  AOI22_X1 U7753 ( .A1(n7758), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n7759), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7754 ( .A1(n6125), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7755 ( .A1(n8799), .A2(n8386), .ZN(n7815) );
  NAND2_X1 U7756 ( .A1(n7812), .A2(n7815), .ZN(n8702) );
  INV_X1 U7757 ( .A(n8702), .ZN(n8707) );
  NAND2_X1 U7758 ( .A1(n7252), .A2(n7755), .ZN(n6145) );
  OR2_X1 U7759 ( .A1(n5991), .A2(n7282), .ZN(n6144) );
  NAND2_X1 U7760 ( .A1(n6146), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7761 ( .A1(n6161), .A2(n6147), .ZN(n8696) );
  NAND2_X1 U7762 ( .A1(n8696), .A2(n6227), .ZN(n6152) );
  INV_X1 U7763 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U7764 ( .A1(n7758), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7765 ( .A1(n6243), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6148) );
  OAI211_X1 U7766 ( .C1(n8695), .C2(n6305), .A(n6149), .B(n6148), .ZN(n6150)
         );
  INV_X1 U7767 ( .A(n6150), .ZN(n6151) );
  INV_X1 U7768 ( .A(n6288), .ZN(n7914) );
  NAND2_X1 U7769 ( .A1(n7330), .A2(n7755), .ZN(n6154) );
  OR2_X1 U7770 ( .A1(n5991), .A2(n7342), .ZN(n6153) );
  XNOR2_X1 U7771 ( .A(n6161), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8685) );
  INV_X1 U7772 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U7773 ( .A1(n7758), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7774 ( .A1(n7759), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6155) );
  OAI211_X1 U7775 ( .C1(n8684), .C2(n6305), .A(n6156), .B(n6155), .ZN(n6157)
         );
  AOI21_X1 U7776 ( .B1(n8685), .B2(n6227), .A(n6157), .ZN(n8270) );
  NAND2_X1 U7777 ( .A1(n8996), .A2(n8270), .ZN(n7922) );
  NAND2_X1 U7778 ( .A1(n9002), .A2(n8706), .ZN(n8673) );
  AND2_X1 U7779 ( .A1(n7922), .A2(n8673), .ZN(n7917) );
  NAND2_X1 U7780 ( .A1(n6158), .A2(n7921), .ZN(n8661) );
  NAND2_X1 U7781 ( .A1(n7384), .A2(n7755), .ZN(n6160) );
  OR2_X1 U7782 ( .A1(n5991), .A2(n7385), .ZN(n6159) );
  OAI21_X1 U7783 ( .B1(n6161), .B2(P2_REG3_REG_21__SCAN_IN), .A(
        P2_REG3_REG_22__SCAN_IN), .ZN(n6164) );
  NOR2_X1 U7784 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n6162) );
  NAND2_X1 U7785 ( .A1(n6163), .A2(n6162), .ZN(n6172) );
  NAND2_X1 U7786 ( .A1(n6164), .A2(n6172), .ZN(n8667) );
  NAND2_X1 U7787 ( .A1(n8667), .A2(n6227), .ZN(n6169) );
  INV_X1 U7788 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U7789 ( .A1(n7759), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7790 ( .A1(n7758), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6165) );
  OAI211_X1 U7791 ( .C1(n6305), .C2(n8669), .A(n6166), .B(n6165), .ZN(n6167)
         );
  INV_X1 U7792 ( .A(n6167), .ZN(n6168) );
  XNOR2_X1 U7793 ( .A(n8788), .B(n8316), .ZN(n8664) );
  INV_X1 U7794 ( .A(n8664), .ZN(n8660) );
  NAND2_X1 U7795 ( .A1(n8661), .A2(n8660), .ZN(n8659) );
  OR2_X1 U7796 ( .A1(n8788), .A2(n8316), .ZN(n7807) );
  NAND2_X1 U7797 ( .A1(n7429), .A2(n7755), .ZN(n6171) );
  OR2_X1 U7798 ( .A1(n5991), .A2(n7431), .ZN(n6170) );
  INV_X1 U7799 ( .A(n8853), .ZN(n8320) );
  NAND2_X1 U7800 ( .A1(n6172), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7801 ( .A1(n6181), .A2(n6173), .ZN(n8656) );
  NAND2_X1 U7802 ( .A1(n8656), .A2(n6227), .ZN(n6178) );
  INV_X1 U7803 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U7804 ( .A1(n7758), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7805 ( .A1(n6243), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6174) );
  OAI211_X1 U7806 ( .C1(n8655), .C2(n6305), .A(n6175), .B(n6174), .ZN(n6176)
         );
  INV_X1 U7807 ( .A(n6176), .ZN(n6177) );
  NAND2_X1 U7808 ( .A1(n6178), .A2(n6177), .ZN(n8665) );
  INV_X1 U7809 ( .A(n8665), .ZN(n8397) );
  NAND2_X1 U7810 ( .A1(n8853), .A2(n8397), .ZN(n7927) );
  NAND2_X1 U7811 ( .A1(n7539), .A2(n7755), .ZN(n6180) );
  OR2_X1 U7812 ( .A1(n5991), .A2(n7664), .ZN(n6179) );
  NAND2_X1 U7813 ( .A1(n6181), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7814 ( .A1(n6192), .A2(n6182), .ZN(n8641) );
  NAND2_X1 U7815 ( .A1(n8641), .A2(n6227), .ZN(n6187) );
  INV_X1 U7816 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U7817 ( .A1(n6125), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7818 ( .A1(n6243), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6183) );
  OAI211_X1 U7819 ( .C1(n5992), .C2(n8899), .A(n6184), .B(n6183), .ZN(n6185)
         );
  INV_X1 U7820 ( .A(n6185), .ZN(n6186) );
  NAND2_X1 U7821 ( .A1(n6187), .A2(n6186), .ZN(n8653) );
  INV_X1 U7822 ( .A(n8653), .ZN(n8282) );
  NAND2_X1 U7823 ( .A1(n7567), .A2(n7755), .ZN(n6189) );
  OR2_X1 U7824 ( .A1(n5991), .A2(n8905), .ZN(n6188) );
  INV_X1 U7825 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7826 ( .A1(n6192), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7827 ( .A1(n6205), .A2(n6193), .ZN(n8631) );
  NAND2_X1 U7828 ( .A1(n8631), .A2(n6227), .ZN(n6199) );
  INV_X1 U7829 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7830 ( .A1(n7758), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7831 ( .A1(n6243), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6194) );
  OAI211_X1 U7832 ( .C1(n6196), .C2(n6305), .A(n6195), .B(n6194), .ZN(n6197)
         );
  INV_X1 U7833 ( .A(n6197), .ZN(n6198) );
  NAND2_X1 U7834 ( .A1(n8841), .A2(n8287), .ZN(n7936) );
  NAND2_X1 U7835 ( .A1(n6200), .A2(n7935), .ZN(n8614) );
  NAND2_X1 U7836 ( .A1(n7619), .A2(n7755), .ZN(n6202) );
  OR2_X1 U7837 ( .A1(n5991), .A2(n7622), .ZN(n6201) );
  INV_X1 U7838 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7839 ( .A1(n6204), .A2(n6203), .ZN(n6215) );
  NAND2_X1 U7840 ( .A1(n6205), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7841 ( .A1(n6215), .A2(n6206), .ZN(n8620) );
  NAND2_X1 U7842 ( .A1(n8620), .A2(n6227), .ZN(n6211) );
  INV_X1 U7843 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U7844 ( .A1(n7758), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7845 ( .A1(n7759), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6207) );
  OAI211_X1 U7846 ( .C1(n8619), .C2(n6305), .A(n6208), .B(n6207), .ZN(n6209)
         );
  INV_X1 U7847 ( .A(n6209), .ZN(n6210) );
  NAND2_X1 U7848 ( .A1(n6211), .A2(n6210), .ZN(n8629) );
  NAND2_X1 U7849 ( .A1(n8835), .A2(n8349), .ZN(n7940) );
  NAND2_X1 U7850 ( .A1(n8614), .A2(n8615), .ZN(n6212) );
  NAND2_X1 U7851 ( .A1(n7634), .A2(n7755), .ZN(n6214) );
  OR2_X1 U7852 ( .A1(n5991), .A2(n7635), .ZN(n6213) );
  NAND2_X1 U7853 ( .A1(n6215), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7854 ( .A1(n6225), .A2(n6216), .ZN(n8611) );
  NAND2_X1 U7855 ( .A1(n8611), .A2(n6227), .ZN(n6221) );
  INV_X1 U7856 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U7857 ( .A1(n7758), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7858 ( .A1(n7759), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6217) );
  OAI211_X1 U7859 ( .C1(n8610), .C2(n6305), .A(n6218), .B(n6217), .ZN(n6219)
         );
  INV_X1 U7860 ( .A(n6219), .ZN(n6220) );
  NAND2_X1 U7861 ( .A1(n7655), .A2(n7755), .ZN(n6223) );
  OR2_X1 U7862 ( .A1(n5991), .A2(n7656), .ZN(n6222) );
  INV_X1 U7863 ( .A(n6225), .ZN(n6224) );
  INV_X1 U7864 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U7865 ( .A1(n6224), .A2(n8296), .ZN(n8573) );
  NAND2_X1 U7866 ( .A1(n6225), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7867 ( .A1(n8573), .A2(n6226), .ZN(n8598) );
  NAND2_X1 U7868 ( .A1(n8598), .A2(n6227), .ZN(n6232) );
  INV_X1 U7869 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8970) );
  NAND2_X1 U7870 ( .A1(n7758), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6229) );
  NAND2_X1 U7871 ( .A1(n6125), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6228) );
  OAI211_X1 U7872 ( .C1(n6013), .C2(n8970), .A(n6229), .B(n6228), .ZN(n6230)
         );
  INV_X1 U7873 ( .A(n6230), .ZN(n6231) );
  NAND2_X1 U7874 ( .A1(n6232), .A2(n6231), .ZN(n8607) );
  INV_X1 U7875 ( .A(n8607), .ZN(n7949) );
  MUX2_X1 U7876 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6362), .Z(n7658) );
  INV_X1 U7877 ( .A(n7741), .ZN(n6239) );
  INV_X1 U7878 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7735) );
  OR2_X1 U7879 ( .A1(n5991), .A2(n7735), .ZN(n6240) );
  OR2_X1 U7880 ( .A1(n8573), .A2(n6242), .ZN(n7764) );
  INV_X1 U7881 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U7882 ( .A1(n7758), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7883 ( .A1(n6243), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6244) );
  OAI211_X1 U7884 ( .C1(n8580), .C2(n6305), .A(n6245), .B(n6244), .ZN(n6246)
         );
  INV_X1 U7885 ( .A(n6246), .ZN(n6247) );
  INV_X1 U7886 ( .A(n8587), .ZN(n6253) );
  NAND2_X1 U7887 ( .A1(n6249), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6250) );
  MUX2_X1 U7888 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6250), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6252) );
  NAND2_X1 U7889 ( .A1(n6252), .A2(n6251), .ZN(n7284) );
  AND2_X1 U7890 ( .A1(n7284), .A2(n7803), .ZN(n6935) );
  INV_X1 U7891 ( .A(n7982), .ZN(n7820) );
  NAND2_X1 U7892 ( .A1(n6935), .A2(n7820), .ZN(n10057) );
  INV_X1 U7893 ( .A(n10057), .ZN(n10032) );
  NAND2_X1 U7894 ( .A1(n7963), .A2(n6449), .ZN(n6425) );
  NAND2_X1 U7895 ( .A1(n7821), .A2(n7820), .ZN(n10072) );
  OAI21_X1 U7896 ( .B1(n7284), .B2(n7982), .A(n7193), .ZN(n6254) );
  INV_X1 U7897 ( .A(n6254), .ZN(n6255) );
  AND2_X1 U7898 ( .A1(n10072), .A2(n6255), .ZN(n6256) );
  NAND2_X1 U7899 ( .A1(n6425), .A2(n6256), .ZN(n7610) );
  NAND2_X1 U7900 ( .A1(n6849), .A2(n10007), .ZN(n6848) );
  NAND2_X1 U7901 ( .A1(n6926), .A2(n6257), .ZN(n6928) );
  NAND2_X1 U7902 ( .A1(n6929), .A2(n6928), .ZN(n6927) );
  AND2_X1 U7903 ( .A1(n7829), .A2(n6258), .ZN(n6261) );
  INV_X1 U7904 ( .A(n6258), .ZN(n6259) );
  NAND2_X1 U7905 ( .A1(n6986), .A2(n6515), .ZN(n6981) );
  NOR2_X1 U7906 ( .A1(n6259), .A2(n6981), .ZN(n6260) );
  NAND2_X1 U7907 ( .A1(n6925), .A2(n10020), .ZN(n6262) );
  NAND2_X1 U7908 ( .A1(n6984), .A2(n6262), .ZN(n6887) );
  NAND2_X1 U7909 ( .A1(n8452), .A2(n6891), .ZN(n6263) );
  NAND2_X1 U7910 ( .A1(n6987), .A2(n6264), .ZN(n6265) );
  NOR2_X1 U7911 ( .A1(n8451), .A2(n6744), .ZN(n7043) );
  NAND2_X1 U7912 ( .A1(n6919), .A2(n10039), .ZN(n7042) );
  INV_X1 U7913 ( .A(n7042), .ZN(n6267) );
  OR2_X1 U7914 ( .A1(n7043), .A2(n6267), .ZN(n6266) );
  NAND2_X1 U7915 ( .A1(n8451), .A2(n6744), .ZN(n7045) );
  OR2_X1 U7916 ( .A1(n6267), .A2(n7045), .ZN(n6268) );
  INV_X1 U7917 ( .A(n10039), .ZN(n7050) );
  NAND2_X1 U7918 ( .A1(n8450), .A2(n7050), .ZN(n7125) );
  INV_X1 U7919 ( .A(n7778), .ZN(n7862) );
  AND2_X1 U7920 ( .A1(n7125), .A2(n7862), .ZN(n6269) );
  NAND2_X1 U7921 ( .A1(n7126), .A2(n6269), .ZN(n6271) );
  INV_X1 U7922 ( .A(n7072), .ZN(n8449) );
  OR2_X1 U7923 ( .A1(n8449), .A2(n6905), .ZN(n6270) );
  NAND2_X1 U7924 ( .A1(n7856), .A2(n7866), .ZN(n7075) );
  NOR2_X1 U7925 ( .A1(n6997), .A2(n8448), .ZN(n6272) );
  INV_X1 U7926 ( .A(n7373), .ZN(n6273) );
  OR2_X1 U7927 ( .A1(n10061), .A2(n8446), .ZN(n6274) );
  NAND2_X1 U7928 ( .A1(n7526), .A2(n8445), .ZN(n7388) );
  OR2_X1 U7929 ( .A1(n10071), .A2(n8444), .ZN(n6275) );
  NAND2_X1 U7930 ( .A1(n7488), .A2(n6275), .ZN(n6277) );
  NAND2_X1 U7931 ( .A1(n10071), .A2(n8444), .ZN(n6276) );
  NAND2_X1 U7932 ( .A1(n6277), .A2(n6276), .ZN(n7557) );
  NAND2_X1 U7933 ( .A1(n7557), .A2(n7562), .ZN(n6279) );
  INV_X1 U7934 ( .A(n7575), .ZN(n9736) );
  NAND2_X1 U7935 ( .A1(n7556), .A2(n9736), .ZN(n6278) );
  NAND2_X1 U7936 ( .A1(n6279), .A2(n6278), .ZN(n7573) );
  INV_X1 U7937 ( .A(n7573), .ZN(n6280) );
  OR2_X1 U7938 ( .A1(n8248), .A2(n8443), .ZN(n6281) );
  INV_X1 U7939 ( .A(n9733), .ZN(n8442) );
  NAND2_X1 U7940 ( .A1(n8253), .A2(n8442), .ZN(n8748) );
  NAND2_X1 U7941 ( .A1(n8750), .A2(n8748), .ZN(n6283) );
  NAND2_X1 U7942 ( .A1(n6283), .A2(n7785), .ZN(n8733) );
  INV_X1 U7943 ( .A(n8432), .ZN(n8740) );
  NAND2_X1 U7944 ( .A1(n8809), .A2(n8740), .ZN(n8734) );
  NAND2_X1 U7945 ( .A1(n8733), .A2(n8734), .ZN(n6284) );
  INV_X1 U7946 ( .A(n8755), .ZN(n8720) );
  NAND2_X1 U7947 ( .A1(n9018), .A2(n8720), .ZN(n6285) );
  OR2_X1 U7948 ( .A1(n9012), .A2(n8738), .ZN(n8699) );
  AND2_X1 U7949 ( .A1(n8699), .A2(n8702), .ZN(n6286) );
  NAND2_X1 U7950 ( .A1(n9012), .A2(n8738), .ZN(n8700) );
  INV_X1 U7951 ( .A(n8386), .ZN(n8721) );
  INV_X1 U7952 ( .A(n8706), .ZN(n8681) );
  OR2_X1 U7953 ( .A1(n9002), .A2(n8681), .ZN(n8677) );
  NAND2_X1 U7954 ( .A1(n4303), .A2(n8677), .ZN(n6289) );
  NAND2_X1 U7955 ( .A1(n7921), .A2(n7922), .ZN(n8676) );
  NAND2_X1 U7956 ( .A1(n6289), .A2(n8676), .ZN(n8680) );
  INV_X1 U7957 ( .A(n8270), .ZN(n8693) );
  OR2_X1 U7958 ( .A1(n8996), .A2(n8693), .ZN(n6290) );
  NAND2_X1 U7959 ( .A1(n8680), .A2(n6290), .ZN(n8663) );
  INV_X1 U7960 ( .A(n8316), .ZN(n8682) );
  OR2_X1 U7961 ( .A1(n8682), .A2(n8788), .ZN(n6291) );
  NAND2_X1 U7962 ( .A1(n8853), .A2(n8665), .ZN(n6292) );
  NOR2_X1 U7963 ( .A1(n8847), .A2(n8653), .ZN(n6294) );
  NAND2_X1 U7964 ( .A1(n8847), .A2(n8653), .ZN(n6293) );
  OAI21_X1 U7965 ( .B1(n8637), .B2(n6294), .A(n6293), .ZN(n8624) );
  INV_X1 U7966 ( .A(n8287), .ZN(n8639) );
  OR2_X1 U7967 ( .A1(n8841), .A2(n8639), .ZN(n6295) );
  NAND2_X1 U7968 ( .A1(n8626), .A2(n6295), .ZN(n8616) );
  NAND2_X1 U7969 ( .A1(n8835), .A2(n8629), .ZN(n6297) );
  NOR2_X1 U7970 ( .A1(n8835), .A2(n8629), .ZN(n6296) );
  AOI21_X1 U7971 ( .B1(n8616), .B2(n6297), .A(n6296), .ZN(n8604) );
  INV_X1 U7972 ( .A(n8823), .ZN(n7951) );
  XNOR2_X1 U7973 ( .A(n6299), .B(n7959), .ZN(n6301) );
  INV_X1 U7974 ( .A(n7284), .ZN(n7801) );
  NAND2_X1 U7975 ( .A1(n7767), .A2(n7801), .ZN(n6300) );
  NAND2_X1 U7976 ( .A1(n7803), .A2(n7982), .ZN(n6340) );
  NAND2_X1 U7977 ( .A1(n6301), .A2(n8752), .ZN(n6311) );
  NAND2_X1 U7978 ( .A1(n6308), .A2(n6302), .ZN(n6457) );
  INV_X1 U7979 ( .A(n6457), .ZN(n6438) );
  INV_X1 U7980 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U7981 ( .A1(n7758), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7982 ( .A1(n7759), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6303) );
  OAI211_X1 U7983 ( .C1(n8986), .C2(n6305), .A(n6304), .B(n6303), .ZN(n6306)
         );
  INV_X1 U7984 ( .A(n6306), .ZN(n6307) );
  NAND2_X1 U7985 ( .A1(n7764), .A2(n6307), .ZN(n8440) );
  NAND2_X1 U7986 ( .A1(n6457), .A2(n7963), .ZN(n8754) );
  AND2_X1 U7987 ( .A1(n6308), .A2(P2_B_REG_SCAN_IN), .ZN(n6309) );
  NOR2_X1 U7988 ( .A1(n8754), .A2(n6309), .ZN(n8571) );
  AOI22_X1 U7989 ( .A1(n8607), .A2(n8739), .B1(n8440), .B2(n8571), .ZN(n6310)
         );
  NAND2_X1 U7990 ( .A1(n7667), .A2(P2_B_REG_SCAN_IN), .ZN(n6315) );
  INV_X1 U7991 ( .A(n7667), .ZN(n6313) );
  INV_X1 U7992 ( .A(P2_B_REG_SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7993 ( .A1(n6313), .A2(n6312), .ZN(n6314) );
  NAND2_X1 U7994 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  NAND2_X1 U7995 ( .A1(n6316), .A2(n7731), .ZN(n6318) );
  OR2_X1 U7996 ( .A1(n6320), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7997 ( .A1(n7731), .A2(n7624), .ZN(n6360) );
  NAND2_X1 U7998 ( .A1(n6319), .A2(n6360), .ZN(n6338) );
  NAND2_X1 U7999 ( .A1(n7667), .A2(n7624), .ZN(n6357) );
  OAI21_X1 U8000 ( .B1(n6320), .B2(P2_D_REG_0__SCAN_IN), .A(n6357), .ZN(n6447)
         );
  NAND3_X1 U8001 ( .A1(n7801), .A2(n7982), .A3(n7193), .ZN(n6321) );
  NAND2_X1 U8002 ( .A1(n7942), .A2(n6321), .ZN(n6322) );
  MUX2_X1 U8003 ( .A(n6338), .B(n6447), .S(n6322), .Z(n6682) );
  NOR4_X1 U8004 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6326) );
  NOR4_X1 U8005 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6325) );
  NOR4_X1 U8006 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6324) );
  NOR4_X1 U8007 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6323) );
  NAND4_X1 U8008 ( .A1(n6326), .A2(n6325), .A3(n6324), .A4(n6323), .ZN(n6331)
         );
  NOR2_X1 U8009 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n8967) );
  NOR4_X1 U8010 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6329) );
  NOR4_X1 U8011 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6328) );
  NOR4_X1 U8012 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6327) );
  NAND4_X1 U8013 ( .A1(n8967), .A2(n6329), .A3(n6328), .A4(n6327), .ZN(n6330)
         );
  NOR2_X1 U8014 ( .A1(n6331), .A2(n6330), .ZN(n6332) );
  OR2_X1 U8015 ( .A1(n6320), .A2(n6332), .ZN(n6339) );
  AND2_X1 U8016 ( .A1(n6423), .A2(n6429), .ZN(n6675) );
  NAND2_X1 U8017 ( .A1(n7963), .A2(n6448), .ZN(n6421) );
  NAND3_X1 U8018 ( .A1(n6339), .A2(n6675), .A3(n6421), .ZN(n6678) );
  NOR2_X1 U8019 ( .A1(n10057), .A2(n7767), .ZN(n6676) );
  NOR2_X1 U8020 ( .A1(n6678), .A2(n6676), .ZN(n6333) );
  NAND2_X1 U8021 ( .A1(n6447), .A2(n6338), .ZN(n6344) );
  AND3_X2 U8022 ( .A1(n6682), .A2(n6333), .A3(n6344), .ZN(n10107) );
  INV_X1 U8023 ( .A(n8583), .ZN(n6349) );
  INV_X1 U8024 ( .A(n10072), .ZN(n10062) );
  NAND2_X1 U8025 ( .A1(n10107), .A2(n10062), .ZN(n8810) );
  INV_X1 U8026 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6334) );
  OAI21_X1 U8027 ( .B1(n6354), .B2(n6337), .A(n6336), .ZN(P2_U3488) );
  OR2_X1 U8028 ( .A1(n6447), .A2(n6338), .ZN(n6679) );
  INV_X1 U8029 ( .A(n6339), .ZN(n6343) );
  OR2_X1 U8030 ( .A1(n6679), .A2(n6343), .ZN(n6419) );
  INV_X1 U8031 ( .A(n6675), .ZN(n6345) );
  NOR2_X1 U8032 ( .A1(n6419), .A2(n6345), .ZN(n6433) );
  NOR2_X1 U8033 ( .A1(n7767), .A2(n7284), .ZN(n6446) );
  INV_X1 U8034 ( .A(n6340), .ZN(n6341) );
  NAND2_X1 U8035 ( .A1(n6446), .A2(n6341), .ZN(n6420) );
  NAND2_X1 U8036 ( .A1(n6425), .A2(n6420), .ZN(n6342) );
  NAND2_X1 U8037 ( .A1(n6433), .A2(n6342), .ZN(n6348) );
  OR2_X1 U8038 ( .A1(n6344), .A2(n6343), .ZN(n6426) );
  NOR2_X1 U8039 ( .A1(n6426), .A2(n6345), .ZN(n6437) );
  AND2_X1 U8040 ( .A1(n7942), .A2(n10072), .ZN(n6346) );
  NAND2_X1 U8041 ( .A1(n6420), .A2(n6346), .ZN(n6431) );
  INV_X1 U8042 ( .A(n6935), .ZN(n7972) );
  NAND2_X1 U8043 ( .A1(n10062), .A2(n7972), .ZN(n8644) );
  NAND2_X1 U8044 ( .A1(n6431), .A2(n8644), .ZN(n6418) );
  NAND2_X1 U8045 ( .A1(n6437), .A2(n6418), .ZN(n6347) );
  INV_X2 U8046 ( .A(n10078), .ZN(n10080) );
  OR2_X1 U8047 ( .A1(n10078), .A2(n10072), .ZN(n9023) );
  INV_X1 U8048 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6350) );
  OAI21_X1 U8049 ( .B1(n6354), .B2(n10078), .A(n6353), .ZN(P2_U3456) );
  AND2_X2 U8050 ( .A1(n6531), .A2(n6355), .ZN(P1_U3973) );
  NAND2_X1 U8051 ( .A1(n4471), .A2(P1_U3086), .ZN(n8303) );
  NAND2_X1 U8052 ( .A1(n6362), .A2(P1_U3086), .ZN(n9694) );
  OAI222_X1 U8053 ( .A1(n8303), .A2(n6356), .B1(n9694), .B2(n6380), .C1(
        P1_U3086), .C2(n6489), .ZN(P1_U3352) );
  NAND2_X1 U8054 ( .A1(n6320), .A2(n6429), .ZN(n6373) );
  INV_X1 U8055 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6359) );
  INV_X1 U8056 ( .A(n6357), .ZN(n6358) );
  AOI22_X1 U8057 ( .A1(n6373), .A2(n6359), .B1(n6429), .B2(n6358), .ZN(
        P2_U3376) );
  INV_X1 U8058 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8963) );
  INV_X1 U8059 ( .A(n6360), .ZN(n6361) );
  AOI22_X1 U8060 ( .A1(n6373), .A2(n8963), .B1(n6429), .B2(n6361), .ZN(
        P2_U3377) );
  AND2_X1 U8061 ( .A1(n6373), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8062 ( .A1(n6373), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8063 ( .A1(n6373), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8064 ( .A1(n6373), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8065 ( .A1(n6373), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8066 ( .A1(n6373), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8067 ( .A1(n6373), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8068 ( .A1(n6373), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8069 ( .A1(n6373), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8070 ( .A1(n6373), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8071 ( .A1(n6373), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8072 ( .A1(n6373), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8073 ( .A1(n6373), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8074 ( .A1(n6373), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8075 ( .A1(n6373), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8076 ( .A1(n6373), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8077 ( .A1(n6373), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8078 ( .A1(n6373), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8079 ( .A1(n6373), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8080 ( .A1(n6373), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8081 ( .A1(n6373), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8082 ( .A1(n6373), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8083 ( .A1(n6373), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8084 ( .A1(n6373), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8085 ( .A1(n6373), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8086 ( .A1(n6373), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  NAND2_X1 U8087 ( .A1(n6362), .A2(P2_U3151), .ZN(n7734) );
  INV_X1 U8088 ( .A(n7734), .ZN(n6967) );
  INV_X1 U8089 ( .A(n6967), .ZN(n9030) );
  NAND2_X1 U8090 ( .A1(n4471), .A2(P2_U3151), .ZN(n9035) );
  OAI222_X1 U8091 ( .A1(n9030), .A2(n6363), .B1(n9035), .B2(n6377), .C1(n4286), 
        .C2(P2_U3151), .ZN(P2_U3293) );
  AOI21_X1 U8092 ( .B1(n8093), .B2(n6365), .A(n6364), .ZN(n6481) );
  INV_X1 U8093 ( .A(n6481), .ZN(n6366) );
  NAND2_X1 U8094 ( .A1(n6554), .A2(n8238), .ZN(n6482) );
  AND2_X1 U8095 ( .A1(n6366), .A2(n6482), .ZN(n9869) );
  NOR2_X1 U8096 ( .A1(n9869), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8097 ( .A(n9035), .ZN(n7428) );
  INV_X1 U8098 ( .A(n7428), .ZN(n7666) );
  INV_X1 U8099 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6367) );
  INV_X1 U8100 ( .A(n8303), .ZN(n9690) );
  AOI22_X1 U8101 ( .A1(n7210), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n9690), .ZN(n6368) );
  OAI21_X1 U8102 ( .B1(n6388), .B2(n9694), .A(n6368), .ZN(P1_U3351) );
  INV_X1 U8103 ( .A(n6369), .ZN(n6383) );
  AOI22_X1 U8104 ( .A1(n9218), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9690), .ZN(n6370) );
  OAI21_X1 U8105 ( .B1(n6383), .B2(n9694), .A(n6370), .ZN(P1_U3350) );
  INV_X1 U8106 ( .A(n6371), .ZN(n6385) );
  AOI22_X1 U8107 ( .A1(n9232), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9690), .ZN(n6372) );
  OAI21_X1 U8108 ( .B1(n6385), .B2(n9694), .A(n6372), .ZN(P1_U3349) );
  INV_X1 U8109 ( .A(n6373), .ZN(n6375) );
  INV_X1 U8110 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n8909) );
  NOR2_X1 U8111 ( .A1(n6375), .A2(n8909), .ZN(P2_U3251) );
  INV_X1 U8112 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n8947) );
  NOR2_X1 U8113 ( .A1(n6375), .A2(n8947), .ZN(P2_U3234) );
  INV_X1 U8114 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6374) );
  NOR2_X1 U8115 ( .A1(n6375), .A2(n6374), .ZN(P2_U3259) );
  INV_X1 U8116 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n8918) );
  NOR2_X1 U8117 ( .A1(n6375), .A2(n8918), .ZN(P2_U3260) );
  INV_X1 U8118 ( .A(n9694), .ZN(n7426) );
  INV_X1 U8119 ( .A(n7426), .ZN(n7742) );
  OAI222_X1 U8120 ( .A1(n8303), .A2(n4891), .B1(n7742), .B2(n6376), .C1(
        P1_U3086), .C2(n6486), .ZN(P1_U3354) );
  OAI222_X1 U8121 ( .A1(n8303), .A2(n6378), .B1(n7742), .B2(n6377), .C1(
        P1_U3086), .C2(n6507), .ZN(P1_U3353) );
  OAI222_X1 U8122 ( .A1(n6381), .A2(P2_U3151), .B1(n9035), .B2(n6380), .C1(
        n6379), .C2(n9030), .ZN(P2_U3292) );
  OAI222_X1 U8123 ( .A1(n6384), .A2(P2_U3151), .B1(n9035), .B2(n6383), .C1(
        n6382), .C2(n9030), .ZN(P2_U3290) );
  OAI222_X1 U8124 ( .A1(n6386), .A2(P2_U3151), .B1(n9035), .B2(n6385), .C1(
        n4419), .C2(n9030), .ZN(P2_U3289) );
  OAI222_X1 U8125 ( .A1(n6623), .A2(P2_U3151), .B1(n9035), .B2(n6388), .C1(
        n6387), .C2(n9030), .ZN(P2_U3291) );
  NOR2_X1 U8126 ( .A1(n6389), .A2(n6554), .ZN(n9940) );
  NAND2_X1 U8127 ( .A1(n9941), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6390) );
  OAI21_X1 U8128 ( .B1(n9941), .B2(n6391), .A(n6390), .ZN(P1_U3440) );
  NAND2_X1 U8129 ( .A1(n9941), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6392) );
  OAI21_X1 U8130 ( .B1(n9941), .B2(n6393), .A(n6392), .ZN(P1_U3439) );
  INV_X1 U8131 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8862) );
  INV_X1 U8132 ( .A(n6394), .ZN(n6397) );
  INV_X1 U8133 ( .A(n9717), .ZN(n6395) );
  OAI222_X1 U8134 ( .A1(n8303), .A2(n8862), .B1(n7742), .B2(n6397), .C1(
        P1_U3086), .C2(n6395), .ZN(P1_U3348) );
  INV_X1 U8135 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6396) );
  OAI222_X1 U8136 ( .A1(n6398), .A2(P2_U3151), .B1(n9035), .B2(n6397), .C1(
        n6396), .C2(n9030), .ZN(P2_U3288) );
  INV_X1 U8137 ( .A(n6399), .ZN(n6402) );
  AOI22_X1 U8138 ( .A1(n9729), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9690), .ZN(n6400) );
  OAI21_X1 U8139 ( .B1(n6402), .B2(n9694), .A(n6400), .ZN(P1_U3347) );
  AOI22_X1 U8140 ( .A1(n6958), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n6967), .ZN(n6401) );
  OAI21_X1 U8141 ( .B1(n6402), .B2(n9035), .A(n6401), .ZN(P2_U3287) );
  INV_X1 U8142 ( .A(P1_U3973), .ZN(n6708) );
  NAND2_X1 U8143 ( .A1(n6708), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n6403) );
  OAI21_X1 U8144 ( .B1(n9284), .B2(n6708), .A(n6403), .ZN(P1_U3571) );
  INV_X1 U8145 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8894) );
  NAND2_X1 U8146 ( .A1(n7985), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8147 ( .A1(n5119), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U8148 ( .A1(n6404), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6405) );
  AND3_X1 U8149 ( .A1(n6407), .A2(n6406), .A3(n6405), .ZN(n8043) );
  INV_X1 U8150 ( .A(n8043), .ZN(n8215) );
  NAND2_X1 U8151 ( .A1(n8215), .A2(P1_U3973), .ZN(n6408) );
  OAI21_X1 U8152 ( .B1(P1_U3973), .B2(n8894), .A(n6408), .ZN(P1_U3585) );
  INV_X1 U8153 ( .A(n6409), .ZN(n6412) );
  AOI22_X1 U8154 ( .A1(n9248), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9690), .ZN(n6410) );
  OAI21_X1 U8155 ( .B1(n6412), .B2(n7742), .A(n6410), .ZN(P1_U3346) );
  AOI22_X1 U8156 ( .A1(n7161), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n6967), .ZN(n6411) );
  OAI21_X1 U8157 ( .B1(n6412), .B2(n7666), .A(n6411), .ZN(P2_U3286) );
  INV_X1 U8158 ( .A(n6413), .ZN(n6415) );
  AOI22_X1 U8159 ( .A1(n9705), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9690), .ZN(n6414) );
  OAI21_X1 U8160 ( .B1(n6415), .B2(n9694), .A(n6414), .ZN(P1_U3345) );
  OAI222_X1 U8161 ( .A1(P2_U3151), .A2(n6416), .B1(n9035), .B2(n6415), .C1(
        n8957), .C2(n9030), .ZN(P2_U3285) );
  NAND2_X1 U8162 ( .A1(n6849), .A2(P2_U3893), .ZN(n6417) );
  OAI21_X1 U8163 ( .B1(P2_U3893), .B2(n5071), .A(n6417), .ZN(P2_U3491) );
  NAND2_X1 U8164 ( .A1(n6419), .A2(n6418), .ZN(n6424) );
  INV_X1 U8165 ( .A(n6420), .ZN(n6434) );
  NAND2_X1 U8166 ( .A1(n6426), .A2(n6434), .ZN(n6422) );
  NAND4_X1 U8167 ( .A1(n6424), .A2(n6423), .A3(n6422), .A4(n6421), .ZN(n6428)
         );
  INV_X1 U8168 ( .A(n6425), .ZN(n6677) );
  AND2_X1 U8169 ( .A1(n6677), .A2(n6675), .ZN(n7980) );
  AND2_X1 U8170 ( .A1(n6426), .A2(n7980), .ZN(n6427) );
  AOI21_X1 U8171 ( .B1(n6428), .B2(P2_STATE_REG_SCAN_IN), .A(n6427), .ZN(n6713) );
  AND2_X1 U8172 ( .A1(n6713), .A2(n6429), .ZN(n6526) );
  INV_X1 U8173 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6687) );
  AND2_X1 U8174 ( .A1(n6675), .A2(n6935), .ZN(n6430) );
  OR2_X1 U8175 ( .A1(n6433), .A2(n6430), .ZN(n9740) );
  AND2_X1 U8176 ( .A1(n9740), .A2(n10062), .ZN(n8369) );
  INV_X1 U8177 ( .A(n6431), .ZN(n6432) );
  NAND2_X1 U8178 ( .A1(n6433), .A2(n6432), .ZN(n6436) );
  NAND2_X1 U8179 ( .A1(n6437), .A2(n6434), .ZN(n6435) );
  AND2_X1 U8180 ( .A1(n7822), .A2(n7826), .ZN(n10003) );
  NAND2_X1 U8181 ( .A1(n6437), .A2(n6677), .ZN(n6458) );
  OR2_X1 U8182 ( .A1(n6458), .A2(n6438), .ZN(n9734) );
  OAI22_X1 U8183 ( .A1(n8391), .A2(n10003), .B1(n9734), .B2(n6926), .ZN(n6439)
         );
  AOI21_X1 U8184 ( .B1(n10007), .B2(n8369), .A(n6439), .ZN(n6440) );
  OAI21_X1 U8185 ( .B1(n6526), .B2(n6687), .A(n6440), .ZN(P2_U3172) );
  INV_X1 U8186 ( .A(n6441), .ZN(n6444) );
  INV_X1 U8187 ( .A(n7215), .ZN(n9818) );
  OAI222_X1 U8188 ( .A1(n8303), .A2(n6442), .B1(n9694), .B2(n6444), .C1(
        P1_U3086), .C2(n9818), .ZN(P1_U3344) );
  OAI222_X1 U8189 ( .A1(n6445), .A2(P2_U3151), .B1(n7666), .B2(n6444), .C1(
        n6443), .C2(n9030), .ZN(P2_U3284) );
  INV_X1 U8190 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6464) );
  INV_X1 U8191 ( .A(n6448), .ZN(n6449) );
  NAND2_X1 U8192 ( .A1(n6451), .A2(n6926), .ZN(n6516) );
  INV_X1 U8193 ( .A(n6451), .ZN(n6452) );
  NAND2_X1 U8194 ( .A1(n6452), .A2(n8456), .ZN(n6453) );
  OAI21_X1 U8195 ( .B1(n10007), .B2(n6714), .A(n7822), .ZN(n6454) );
  OAI21_X1 U8196 ( .B1(n6455), .B2(n6454), .A(n6517), .ZN(n6456) );
  INV_X1 U8197 ( .A(n8391), .ZN(n9742) );
  NAND2_X1 U8198 ( .A1(n6456), .A2(n9742), .ZN(n6463) );
  INV_X1 U8199 ( .A(n9734), .ZN(n8410) );
  OR2_X1 U8200 ( .A1(n6458), .A2(n6457), .ZN(n8412) );
  INV_X1 U8201 ( .A(n9740), .ZN(n7008) );
  NAND2_X1 U8202 ( .A1(n6459), .A2(n10062), .ZN(n10009) );
  OAI22_X1 U8203 ( .A1(n6460), .A2(n8412), .B1(n7008), .B2(n10009), .ZN(n6461)
         );
  AOI21_X1 U8204 ( .B1(n8410), .B2(n8454), .A(n6461), .ZN(n6462) );
  OAI211_X1 U8205 ( .C1(n6526), .C2(n6464), .A(n6463), .B(n6462), .ZN(P2_U3162) );
  OAI21_X1 U8206 ( .B1(n6467), .B2(n6466), .A(n6465), .ZN(n6468) );
  INV_X1 U8207 ( .A(n6468), .ZN(n6533) );
  INV_X1 U8208 ( .A(n6469), .ZN(n6491) );
  NOR3_X1 U8209 ( .A1(n6533), .A2(n6491), .A3(n4285), .ZN(n6473) );
  NAND2_X1 U8210 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6477) );
  AND2_X1 U8211 ( .A1(n6495), .A2(n6491), .ZN(n8240) );
  INV_X1 U8212 ( .A(n8240), .ZN(n6483) );
  OR2_X1 U8213 ( .A1(n6469), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U8214 ( .A1(n6495), .A2(n6470), .ZN(n9799) );
  INV_X1 U8215 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U8216 ( .A1(n9799), .A2(n6471), .ZN(n9803) );
  OAI211_X1 U8217 ( .C1(n6477), .C2(n6483), .A(P1_U3973), .B(n9803), .ZN(n6472) );
  NOR2_X1 U8218 ( .A1(n6473), .A2(n6472), .ZN(n6514) );
  INV_X1 U8219 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6474) );
  MUX2_X1 U8220 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6474), .S(n7210), .Z(n6485)
         );
  INV_X1 U8221 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6475) );
  MUX2_X1 U8222 ( .A(n6475), .B(P1_REG2_REG_2__SCAN_IN), .S(n6507), .Z(n6503)
         );
  INV_X1 U8223 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6476) );
  MUX2_X1 U8224 ( .A(n6476), .B(P1_REG2_REG_1__SCAN_IN), .S(n6486), .Z(n9189)
         );
  INV_X1 U8225 ( .A(n6477), .ZN(n9188) );
  NAND2_X1 U8226 ( .A1(n9189), .A2(n9188), .ZN(n9187) );
  INV_X1 U8227 ( .A(n6486), .ZN(n9193) );
  NAND2_X1 U8228 ( .A1(n9193), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8229 ( .A1(n9187), .A2(n6478), .ZN(n6502) );
  NAND2_X1 U8230 ( .A1(n6503), .A2(n6502), .ZN(n6501) );
  OR2_X1 U8231 ( .A1(n6507), .A2(n6475), .ZN(n6479) );
  NAND2_X1 U8232 ( .A1(n6501), .A2(n6479), .ZN(n9203) );
  XNOR2_X1 U8233 ( .A(n6489), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U8234 ( .A1(n9203), .A2(n9204), .ZN(n9202) );
  INV_X1 U8235 ( .A(n6489), .ZN(n9201) );
  NAND2_X1 U8236 ( .A1(n9201), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U8237 ( .A1(n9202), .A2(n6480), .ZN(n6484) );
  NAND2_X1 U8238 ( .A1(n6482), .A2(n6481), .ZN(n9807) );
  OR2_X1 U8239 ( .A1(n9807), .A2(n6483), .ZN(n9889) );
  INV_X1 U8240 ( .A(n9889), .ZN(n9884) );
  NAND2_X1 U8241 ( .A1(n6484), .A2(n6485), .ZN(n7197) );
  OAI211_X1 U8242 ( .C1(n6485), .C2(n6484), .A(n9884), .B(n7197), .ZN(n6499)
         );
  INV_X1 U8243 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9972) );
  MUX2_X1 U8244 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9972), .S(n7210), .Z(n6493)
         );
  INV_X1 U8245 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6490) );
  INV_X1 U8246 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6488) );
  INV_X1 U8247 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6487) );
  MUX2_X1 U8248 ( .A(n6487), .B(P1_REG1_REG_1__SCAN_IN), .S(n6486), .Z(n9192)
         );
  NAND3_X1 U8249 ( .A1(n9192), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9190) );
  OAI21_X1 U8250 ( .B1(n6487), .B2(n6486), .A(n9190), .ZN(n6505) );
  MUX2_X1 U8251 ( .A(n6488), .B(P1_REG1_REG_2__SCAN_IN), .S(n6507), .Z(n6506)
         );
  NAND2_X1 U8252 ( .A1(n6505), .A2(n6506), .ZN(n6504) );
  OAI21_X1 U8253 ( .B1(n6488), .B2(n6507), .A(n6504), .ZN(n9206) );
  XNOR2_X1 U8254 ( .A(n6489), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U8255 ( .A1(n9206), .A2(n9207), .ZN(n9205) );
  OAI21_X1 U8256 ( .B1(n6490), .B2(n6489), .A(n9205), .ZN(n6492) );
  OR2_X1 U8257 ( .A1(n9807), .A2(n6491), .ZN(n9851) );
  INV_X1 U8258 ( .A(n9851), .ZN(n9892) );
  OAI211_X1 U8259 ( .C1(n6493), .C2(n6492), .A(n9892), .B(n7209), .ZN(n6498)
         );
  INV_X1 U8260 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8935) );
  NOR2_X1 U8261 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8935), .ZN(n6494) );
  AOI21_X1 U8262 ( .B1(n9869), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6494), .ZN(
        n6497) );
  OR2_X1 U8263 ( .A1(n9807), .A2(n6495), .ZN(n9898) );
  INV_X1 U8264 ( .A(n9898), .ZN(n9881) );
  NAND2_X1 U8265 ( .A1(n9881), .A2(n7210), .ZN(n6496) );
  NAND4_X1 U8266 ( .A1(n6499), .A2(n6498), .A3(n6497), .A4(n6496), .ZN(n6500)
         );
  OR2_X1 U8267 ( .A1(n6514), .A2(n6500), .ZN(P1_U3247) );
  OAI211_X1 U8268 ( .C1(n6503), .C2(n6502), .A(n9884), .B(n6501), .ZN(n6512)
         );
  OAI211_X1 U8269 ( .C1(n6506), .C2(n6505), .A(n9892), .B(n6504), .ZN(n6511)
         );
  AOI22_X1 U8270 ( .A1(n9869), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6510) );
  INV_X1 U8271 ( .A(n6507), .ZN(n6508) );
  NAND2_X1 U8272 ( .A1(n9881), .A2(n6508), .ZN(n6509) );
  NAND4_X1 U8273 ( .A1(n6512), .A2(n6511), .A3(n6510), .A4(n6509), .ZN(n6513)
         );
  OR2_X1 U8274 ( .A1(n6514), .A2(n6513), .ZN(P1_U3245) );
  INV_X1 U8275 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6525) );
  XNOR2_X1 U8276 ( .A(n6515), .B(n6714), .ZN(n6716) );
  XNOR2_X1 U8277 ( .A(n6716), .B(n6986), .ZN(n6519) );
  NAND2_X1 U8278 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  NAND2_X1 U8279 ( .A1(n6518), .A2(n6519), .ZN(n6719) );
  OAI21_X1 U8280 ( .B1(n6519), .B2(n6518), .A(n6719), .ZN(n6520) );
  NAND2_X1 U8281 ( .A1(n6520), .A2(n9742), .ZN(n6524) );
  NAND2_X1 U8282 ( .A1(n6521), .A2(n10062), .ZN(n10014) );
  OAI22_X1 U8283 ( .A1(n6926), .A2(n8412), .B1(n7008), .B2(n10014), .ZN(n6522)
         );
  AOI21_X1 U8284 ( .B1(n8410), .B2(n8453), .A(n6522), .ZN(n6523) );
  OAI211_X1 U8285 ( .C1(n6526), .C2(n6525), .A(n6524), .B(n6523), .ZN(P2_U3177) );
  INV_X1 U8286 ( .A(n6527), .ZN(n6537) );
  AOI22_X1 U8287 ( .A1(n7680), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9690), .ZN(n6528) );
  OAI21_X1 U8288 ( .B1(n6537), .B2(n9694), .A(n6528), .ZN(P1_U3343) );
  INV_X1 U8289 ( .A(n4282), .ZN(n9143) );
  INV_X1 U8290 ( .A(n7066), .ZN(n6568) );
  INV_X1 U8291 ( .A(n6529), .ZN(n6532) );
  NAND3_X1 U8292 ( .A1(n6532), .A2(n6531), .A3(n6530), .ZN(n6668) );
  NAND2_X1 U8293 ( .A1(n6668), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6535) );
  NOR2_X1 U8294 ( .A1(n6541), .A2(n9161), .ZN(n7058) );
  AOI22_X1 U8295 ( .A1(n9158), .A2(n6533), .B1(n9164), .B2(n7058), .ZN(n6534)
         );
  OAI211_X1 U8296 ( .C1(n9143), .C2(n6568), .A(n6535), .B(n6534), .ZN(P1_U3232) );
  OAI222_X1 U8297 ( .A1(P2_U3151), .A2(n6538), .B1(n7666), .B2(n6537), .C1(
        n6536), .C2(n7734), .ZN(P2_U3283) );
  XOR2_X1 U8298 ( .A(n6540), .B(n6539), .Z(n6545) );
  INV_X1 U8299 ( .A(n6541), .ZN(n9185) );
  INV_X1 U8300 ( .A(n9163), .ZN(n9761) );
  INV_X1 U8301 ( .A(n9161), .ZN(n9758) );
  AOI22_X1 U8302 ( .A1(n9185), .A2(n9761), .B1(n9758), .B2(n9183), .ZN(n6779)
         );
  INV_X1 U8303 ( .A(n6779), .ZN(n6542) );
  AOI22_X1 U8304 ( .A1(n4282), .A2(n7038), .B1(n9164), .B2(n6542), .ZN(n6544)
         );
  NAND2_X1 U8305 ( .A1(n6668), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6543) );
  OAI211_X1 U8306 ( .C1(n6545), .C2(n9792), .A(n6544), .B(n6543), .ZN(P1_U3237) );
  INV_X1 U8307 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6547) );
  INV_X1 U8308 ( .A(n6546), .ZN(n6549) );
  INV_X1 U8309 ( .A(n9831), .ZN(n7678) );
  OAI222_X1 U8310 ( .A1(n8303), .A2(n6547), .B1(n9694), .B2(n6549), .C1(
        P1_U3086), .C2(n7678), .ZN(P1_U3342) );
  INV_X1 U8311 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6548) );
  OAI222_X1 U8312 ( .A1(n6550), .A2(P2_U3151), .B1(n7666), .B2(n6549), .C1(
        n6548), .C2(n9030), .ZN(P2_U3282) );
  INV_X1 U8313 ( .A(n9301), .ZN(n6551) );
  NAND2_X1 U8314 ( .A1(n6551), .A2(P1_U3973), .ZN(n6552) );
  OAI21_X1 U8315 ( .B1(P1_U3973), .B2(n7431), .A(n6552), .ZN(P1_U3577) );
  INV_X1 U8316 ( .A(n6853), .ZN(n7055) );
  AND2_X1 U8317 ( .A1(n8093), .A2(n8235), .ZN(n6553) );
  NOR2_X1 U8318 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  AND2_X1 U8319 ( .A1(n6556), .A2(n6555), .ZN(n7053) );
  AND2_X1 U8320 ( .A1(n7055), .A2(n7053), .ZN(n6559) );
  INV_X1 U8321 ( .A(n6557), .ZN(n6558) );
  NOR2_X1 U8322 ( .A1(n7054), .A2(n6558), .ZN(n6855) );
  INV_X1 U8323 ( .A(n9971), .ZN(n6560) );
  INV_X1 U8324 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6570) );
  MUX2_X1 U8325 ( .A(n6562), .B(n5060), .S(n7060), .Z(n6563) );
  NAND2_X1 U8326 ( .A1(n6563), .A2(n7056), .ZN(n7478) );
  NAND2_X1 U8327 ( .A1(n5698), .A2(n5437), .ZN(n8223) );
  OR2_X1 U8328 ( .A1(n8223), .A2(n8232), .ZN(n7514) );
  NAND2_X1 U8329 ( .A1(n7478), .A2(n7514), .ZN(n9958) );
  OR2_X1 U8330 ( .A1(n5698), .A2(n9350), .ZN(n6565) );
  NAND2_X1 U8331 ( .A1(n8225), .A2(n8232), .ZN(n6564) );
  AND2_X1 U8332 ( .A1(n6565), .A2(n6564), .ZN(n9469) );
  INV_X1 U8333 ( .A(n9469), .ZN(n9910) );
  NAND2_X1 U8334 ( .A1(n5076), .A2(n7066), .ZN(n6804) );
  INV_X1 U8335 ( .A(n5076), .ZN(n9186) );
  NAND2_X1 U8336 ( .A1(n9186), .A2(n6568), .ZN(n8008) );
  AND2_X1 U8337 ( .A1(n6804), .A2(n8008), .ZN(n8050) );
  INV_X1 U8338 ( .A(n8050), .ZN(n7057) );
  OAI21_X1 U8339 ( .B1(n9958), .B2(n9910), .A(n7057), .ZN(n6567) );
  INV_X1 U8340 ( .A(n7058), .ZN(n6566) );
  OAI211_X1 U8341 ( .C1(n7056), .C2(n6568), .A(n6567), .B(n6566), .ZN(n9628)
         );
  NAND2_X1 U8342 ( .A1(n9628), .A2(n9961), .ZN(n6569) );
  OAI21_X1 U8343 ( .B1(n9961), .B2(n6570), .A(n6569), .ZN(P1_U3453) );
  OAI211_X1 U8344 ( .C1(n6573), .C2(n6572), .A(n6571), .B(n9981), .ZN(n6587)
         );
  INV_X1 U8345 ( .A(n6574), .ZN(n6575) );
  AOI21_X1 U8346 ( .B1(n6576), .B2(n6869), .A(n6575), .ZN(n6577) );
  NOR2_X1 U8347 ( .A1(n6577), .A2(n8565), .ZN(n6584) );
  AOI21_X1 U8348 ( .B1(n6579), .B2(n10091), .A(n6578), .ZN(n6582) );
  NAND2_X1 U8349 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3151), .ZN(n6581) );
  NAND2_X1 U8350 ( .A1(n9991), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n6580) );
  OAI211_X1 U8351 ( .C1(n8559), .C2(n6582), .A(n6581), .B(n6580), .ZN(n6583)
         );
  AOI211_X1 U8352 ( .C1(n8553), .C2(n6585), .A(n6584), .B(n6583), .ZN(n6586)
         );
  NAND2_X1 U8353 ( .A1(n6587), .A2(n6586), .ZN(P2_U3187) );
  AOI21_X1 U8354 ( .B1(n6590), .B2(n6589), .A(n6588), .ZN(n6601) );
  INV_X1 U8355 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U8356 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6725) );
  INV_X1 U8357 ( .A(n6613), .ZN(n6591) );
  AOI21_X1 U8358 ( .B1(n6993), .B2(n6592), .A(n6591), .ZN(n6593) );
  OR2_X1 U8359 ( .A1(n8565), .A2(n6593), .ZN(n6594) );
  OAI211_X1 U8360 ( .C1(n8561), .C2(n6595), .A(n6725), .B(n6594), .ZN(n6599)
         );
  NAND2_X1 U8361 ( .A1(n6596), .A2(n10087), .ZN(n6597) );
  AOI21_X1 U8362 ( .B1(n6608), .B2(n6597), .A(n8559), .ZN(n6598) );
  AOI211_X1 U8363 ( .C1(n8553), .C2(n4431), .A(n6599), .B(n6598), .ZN(n6600)
         );
  OAI21_X1 U8364 ( .B1(n6601), .B2(n6844), .A(n6600), .ZN(P2_U3185) );
  INV_X1 U8365 ( .A(n8553), .ZN(n9993) );
  OAI211_X1 U8366 ( .C1(n6604), .C2(n6603), .A(n6602), .B(n9981), .ZN(n6622)
         );
  INV_X1 U8367 ( .A(n6605), .ZN(n6607) );
  NAND3_X1 U8368 ( .A1(n6608), .A2(n6607), .A3(n6606), .ZN(n6609) );
  AOI21_X1 U8369 ( .B1(n6610), .B2(n6609), .A(n8559), .ZN(n6620) );
  INV_X1 U8370 ( .A(n6611), .ZN(n6612) );
  NAND3_X1 U8371 ( .A1(n6613), .A2(n6612), .A3(n4731), .ZN(n6614) );
  AOI21_X1 U8372 ( .B1(n6615), .B2(n6614), .A(n8565), .ZN(n6619) );
  INV_X1 U8373 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6616) );
  NOR2_X1 U8374 ( .A1(n8561), .A2(n6616), .ZN(n6618) );
  NAND2_X1 U8375 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6749) );
  INV_X1 U8376 ( .A(n6749), .ZN(n6617) );
  NOR4_X1 U8377 ( .A1(n6620), .A2(n6619), .A3(n6618), .A4(n6617), .ZN(n6621)
         );
  OAI211_X1 U8378 ( .C1(n9993), .C2(n6623), .A(n6622), .B(n6621), .ZN(P2_U3186) );
  XNOR2_X1 U8379 ( .A(n6624), .B(n10083), .ZN(n6633) );
  INV_X1 U8380 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10112) );
  INV_X1 U8381 ( .A(n8565), .ZN(n9990) );
  NAND2_X1 U8382 ( .A1(n6626), .A2(n6625), .ZN(n6627) );
  NAND2_X1 U8383 ( .A1(n6628), .A2(n6627), .ZN(n6629) );
  NAND2_X1 U8384 ( .A1(n9990), .A2(n6629), .ZN(n6631) );
  NAND2_X1 U8385 ( .A1(P2_U3151), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6630) );
  OAI211_X1 U8386 ( .C1(n8561), .C2(n10112), .A(n6631), .B(n6630), .ZN(n6632)
         );
  AOI21_X1 U8387 ( .B1(n10000), .B2(n6633), .A(n6632), .ZN(n6636) );
  OAI21_X1 U8388 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6638), .A(n6637), .ZN(n6639) );
  OAI21_X1 U8389 ( .B1(n6640), .B2(n9981), .A(n6639), .ZN(n6641) );
  OAI21_X1 U8390 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6687), .A(n6641), .ZN(n6642) );
  AOI21_X1 U8391 ( .B1(n9991), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6642), .ZN(
        n6643) );
  OAI21_X1 U8392 ( .B1(n4404), .B2(n9993), .A(n6643), .ZN(P2_U3182) );
  AOI21_X1 U8393 ( .B1(n6644), .B2(n6645), .A(n9792), .ZN(n6647) );
  NAND2_X1 U8394 ( .A1(n6647), .A2(n6646), .ZN(n6650) );
  INV_X1 U8395 ( .A(n9164), .ZN(n9787) );
  AOI22_X1 U8396 ( .A1(n9181), .A2(n9758), .B1(n9761), .B2(n9183), .ZN(n7306)
         );
  OAI22_X1 U8397 ( .A1(n9787), .A2(n7306), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8935), .ZN(n6648) );
  AOI21_X1 U8398 ( .B1(n7303), .B2(n4282), .A(n6648), .ZN(n6649) );
  OAI211_X1 U8399 ( .C1(n9797), .C2(n6651), .A(n6650), .B(n6649), .ZN(P1_U3230) );
  INV_X1 U8400 ( .A(n6652), .ZN(n6655) );
  OAI222_X1 U8401 ( .A1(n6654), .A2(P2_U3151), .B1(n7666), .B2(n6655), .C1(
        n6653), .C2(n7734), .ZN(P2_U3281) );
  INV_X1 U8402 ( .A(n7702), .ZN(n9845) );
  OAI222_X1 U8403 ( .A1(n8303), .A2(n6656), .B1(n9694), .B2(n6655), .C1(
        P1_U3086), .C2(n9845), .ZN(P1_U3341) );
  XOR2_X1 U8404 ( .A(n6658), .B(n6657), .Z(n6663) );
  NAND2_X1 U8405 ( .A1(n9184), .A2(n9761), .ZN(n6660) );
  NAND2_X1 U8406 ( .A1(n9182), .A2(n9758), .ZN(n6659) );
  NAND2_X1 U8407 ( .A1(n6660), .A2(n6659), .ZN(n6793) );
  AOI22_X1 U8408 ( .A1(n9924), .A2(n4282), .B1(n9164), .B2(n6793), .ZN(n6662)
         );
  MUX2_X1 U8409 ( .A(n9797), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6661) );
  OAI211_X1 U8410 ( .C1(n6663), .C2(n9792), .A(n6662), .B(n6661), .ZN(P1_U3218) );
  XOR2_X1 U8411 ( .A(n6665), .B(n6664), .Z(n6671) );
  NAND2_X1 U8412 ( .A1(n9184), .A2(n9758), .ZN(n6667) );
  OAI21_X1 U8413 ( .B1(n5076), .B2(n9163), .A(n6667), .ZN(n6807) );
  AOI22_X1 U8414 ( .A1(n6666), .A2(n4282), .B1(n9164), .B2(n6807), .ZN(n6670)
         );
  NAND2_X1 U8415 ( .A1(n6668), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6669) );
  OAI211_X1 U8416 ( .C1(n6671), .C2(n9792), .A(n6670), .B(n6669), .ZN(P1_U3222) );
  NAND2_X1 U8417 ( .A1(n8665), .A2(P2_U3893), .ZN(n6672) );
  OAI21_X1 U8418 ( .B1(P2_U3893), .B2(n5537), .A(n6672), .ZN(P2_U3514) );
  INV_X1 U8419 ( .A(n6673), .ZN(n6710) );
  AOI22_X1 U8420 ( .A1(n9860), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n9690), .ZN(n6674) );
  OAI21_X1 U8421 ( .B1(n6710), .B2(n9694), .A(n6674), .ZN(P1_U3340) );
  NAND2_X1 U8422 ( .A1(n6676), .A2(n6675), .ZN(n8642) );
  NOR3_X1 U8423 ( .A1(n10003), .A2(n10062), .A3(n6677), .ZN(n6683) );
  NOR2_X1 U8424 ( .A1(n6926), .A2(n8754), .ZN(n10006) );
  INV_X1 U8425 ( .A(n6678), .ZN(n6680) );
  NAND2_X1 U8426 ( .A1(n6680), .A2(n6679), .ZN(n6681) );
  OR2_X1 U8427 ( .A1(n6682), .A2(n6681), .ZN(n6684) );
  NAND2_X1 U8428 ( .A1(n6684), .A2(n8642), .ZN(n8715) );
  INV_X1 U8429 ( .A(n8715), .ZN(n7496) );
  OAI21_X1 U8430 ( .B1(n6683), .B2(n10006), .A(n8723), .ZN(n6686) );
  AOI22_X1 U8431 ( .A1(n10007), .A2(n8762), .B1(n7496), .B2(
        P2_REG2_REG_0__SCAN_IN), .ZN(n6685) );
  OAI211_X1 U8432 ( .C1(n8642), .C2(n6687), .A(n6686), .B(n6685), .ZN(P2_U3233) );
  AOI21_X1 U8433 ( .B1(n6690), .B2(n6689), .A(n6688), .ZN(n6706) );
  OAI21_X1 U8434 ( .B1(n6693), .B2(n6692), .A(n6691), .ZN(n6702) );
  INV_X1 U8435 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6700) );
  OAI21_X1 U8436 ( .B1(n6696), .B2(n6695), .A(n6694), .ZN(n6697) );
  NAND2_X1 U8437 ( .A1(n9990), .A2(n6697), .ZN(n6699) );
  INV_X1 U8438 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6698) );
  OR2_X1 U8439 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6698), .ZN(n6767) );
  OAI211_X1 U8440 ( .C1(n8561), .C2(n6700), .A(n6699), .B(n6767), .ZN(n6701)
         );
  AOI21_X1 U8441 ( .B1(n10000), .B2(n6702), .A(n6701), .ZN(n6705) );
  NAND2_X1 U8442 ( .A1(n8553), .A2(n6703), .ZN(n6704) );
  OAI211_X1 U8443 ( .C1(n6706), .C2(n6844), .A(n6705), .B(n6704), .ZN(P2_U3188) );
  NAND2_X1 U8444 ( .A1(n6708), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6707) );
  OAI21_X1 U8445 ( .B1(n6708), .B2(n7988), .A(n6707), .ZN(P1_U3583) );
  OAI222_X1 U8446 ( .A1(P2_U3151), .A2(n6711), .B1(n7666), .B2(n6710), .C1(
        n6709), .C2(n7734), .ZN(P2_U3280) );
  OR2_X1 U8447 ( .A1(n6712), .A2(P2_U3151), .ZN(n7984) );
  AND2_X1 U8448 ( .A1(n6713), .A2(n7984), .ZN(n9746) );
  INV_X1 U8449 ( .A(n6714), .ZN(n6715) );
  XNOR2_X1 U8450 ( .A(n6714), .B(n10020), .ZN(n6734) );
  XNOR2_X1 U8451 ( .A(n6734), .B(n8453), .ZN(n6723) );
  INV_X1 U8452 ( .A(n6716), .ZN(n6717) );
  NAND2_X1 U8453 ( .A1(n6717), .A2(n6986), .ZN(n6718) );
  NAND2_X1 U8454 ( .A1(n6719), .A2(n6718), .ZN(n6722) );
  INV_X1 U8455 ( .A(n6722), .ZN(n6721) );
  NAND2_X1 U8456 ( .A1(n6721), .A2(n6720), .ZN(n6742) );
  INV_X1 U8457 ( .A(n6742), .ZN(n6753) );
  AOI211_X1 U8458 ( .C1(n6723), .C2(n6722), .A(n8391), .B(n6753), .ZN(n6724)
         );
  INV_X1 U8459 ( .A(n6724), .ZN(n6729) );
  INV_X1 U8460 ( .A(n6725), .ZN(n6727) );
  INV_X1 U8461 ( .A(n8369), .ZN(n8438) );
  OAI22_X1 U8462 ( .A1(n8438), .A2(n10020), .B1(n6986), .B2(n8412), .ZN(n6726)
         );
  AOI211_X1 U8463 ( .C1(n8410), .C2(n8452), .A(n6727), .B(n6726), .ZN(n6728)
         );
  OAI211_X1 U8464 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9746), .A(n6729), .B(
        n6728), .ZN(P2_U3158) );
  INV_X1 U8465 ( .A(n6730), .ZN(n6868) );
  INV_X1 U8466 ( .A(n6731), .ZN(n6732) );
  NAND2_X1 U8467 ( .A1(n6732), .A2(n8452), .ZN(n6733) );
  NAND2_X1 U8468 ( .A1(n6739), .A2(n6733), .ZN(n6751) );
  AND2_X1 U8469 ( .A1(n6734), .A2(n8453), .ZN(n6752) );
  NOR2_X1 U8470 ( .A1(n6751), .A2(n6752), .ZN(n6737) );
  NAND2_X1 U8471 ( .A1(n6742), .A2(n6737), .ZN(n6754) );
  INV_X1 U8472 ( .A(n6754), .ZN(n6736) );
  INV_X1 U8473 ( .A(n6739), .ZN(n6735) );
  XNOR2_X1 U8474 ( .A(n6714), .B(n6867), .ZN(n6759) );
  NOR3_X1 U8475 ( .A1(n6736), .A2(n6735), .A3(n6738), .ZN(n6743) );
  AND2_X1 U8476 ( .A1(n6737), .A2(n6738), .ZN(n6741) );
  INV_X1 U8477 ( .A(n6738), .ZN(n6740) );
  OAI21_X1 U8478 ( .B1(n6743), .B2(n4369), .A(n9742), .ZN(n6748) );
  AND2_X1 U8479 ( .A1(n6744), .A2(n10062), .ZN(n10031) );
  NOR2_X1 U8480 ( .A1(n8412), .A2(n6987), .ZN(n6746) );
  OAI22_X1 U8481 ( .A1(n9734), .A2(n6919), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6004), .ZN(n6745) );
  AOI211_X1 U8482 ( .C1(n10031), .C2(n9740), .A(n6746), .B(n6745), .ZN(n6747)
         );
  OAI211_X1 U8483 ( .C1(n6868), .C2(n9746), .A(n6748), .B(n6747), .ZN(P2_U3167) );
  NAND2_X1 U8484 ( .A1(n6891), .A2(n10062), .ZN(n10025) );
  INV_X1 U8485 ( .A(n8412), .ZN(n9737) );
  AOI22_X1 U8486 ( .A1(n9737), .A2(n8453), .B1(n8410), .B2(n8451), .ZN(n6750)
         );
  OAI211_X1 U8487 ( .C1(n7008), .C2(n10025), .A(n6750), .B(n6749), .ZN(n6757)
         );
  OAI21_X1 U8488 ( .B1(n6753), .B2(n6752), .A(n6751), .ZN(n6755) );
  AOI21_X1 U8489 ( .B1(n6755), .B2(n6754), .A(n8391), .ZN(n6756) );
  AOI211_X1 U8490 ( .C1(n6890), .C2(n8434), .A(n6757), .B(n6756), .ZN(n6758)
         );
  INV_X1 U8491 ( .A(n6758), .ZN(P2_U3170) );
  INV_X1 U8492 ( .A(n6759), .ZN(n6760) );
  NAND2_X1 U8493 ( .A1(n6760), .A2(n6766), .ZN(n6761) );
  XNOR2_X1 U8494 ( .A(n6909), .B(n8450), .ZN(n6763) );
  AOI21_X1 U8495 ( .B1(n6762), .B2(n6763), .A(n8391), .ZN(n6765) );
  NAND2_X1 U8496 ( .A1(n6765), .A2(n6915), .ZN(n6771) );
  OR2_X1 U8497 ( .A1(n8412), .A2(n6766), .ZN(n6768) );
  OAI211_X1 U8498 ( .C1(n9734), .C2(n7072), .A(n6768), .B(n6767), .ZN(n6769)
         );
  AOI21_X1 U8499 ( .B1(n8434), .B2(n7049), .A(n6769), .ZN(n6770) );
  OAI211_X1 U8500 ( .C1(n10039), .C2(n8438), .A(n6771), .B(n6770), .ZN(
        P2_U3179) );
  INV_X1 U8501 ( .A(n7514), .ZN(n6782) );
  NAND2_X1 U8502 ( .A1(n9185), .A2(n7025), .ZN(n8009) );
  NAND2_X1 U8503 ( .A1(n6541), .A2(n6666), .ZN(n6776) );
  NAND2_X1 U8504 ( .A1(n9186), .A2(n7066), .ZN(n6801) );
  NAND2_X1 U8505 ( .A1(n6541), .A2(n7025), .ZN(n6772) );
  NAND2_X1 U8506 ( .A1(n6803), .A2(n6772), .ZN(n6774) );
  INV_X1 U8507 ( .A(n8048), .ZN(n6773) );
  NAND2_X1 U8508 ( .A1(n6774), .A2(n6773), .ZN(n6788) );
  OR2_X1 U8509 ( .A1(n6774), .A2(n6773), .ZN(n6775) );
  NAND2_X1 U8510 ( .A1(n6788), .A2(n6775), .ZN(n7121) );
  OR2_X1 U8511 ( .A1(n6666), .A2(n7066), .ZN(n6814) );
  INV_X1 U8512 ( .A(n9917), .ZN(n9527) );
  AOI211_X1 U8513 ( .C1(n7038), .C2(n6814), .A(n9527), .B(n6796), .ZN(n7116)
         );
  NAND2_X1 U8514 ( .A1(n6777), .A2(n8048), .ZN(n6792) );
  OAI21_X1 U8515 ( .B1(n6777), .B2(n8048), .A(n6792), .ZN(n6778) );
  NAND2_X1 U8516 ( .A1(n6778), .A2(n9910), .ZN(n6781) );
  INV_X1 U8517 ( .A(n7478), .ZN(n6809) );
  NAND2_X1 U8518 ( .A1(n7121), .A2(n6809), .ZN(n6780) );
  NAND3_X1 U8519 ( .A1(n6781), .A2(n6780), .A3(n6779), .ZN(n7118) );
  AOI211_X1 U8520 ( .C1(n6782), .C2(n7121), .A(n7116), .B(n7118), .ZN(n7040)
         );
  INV_X1 U8521 ( .A(n9965), .ZN(n9580) );
  NAND2_X1 U8522 ( .A1(n9961), .A2(n9580), .ZN(n9685) );
  INV_X1 U8523 ( .A(n7038), .ZN(n8006) );
  INV_X1 U8524 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6783) );
  OAI22_X1 U8525 ( .A1(n9685), .A2(n8006), .B1(n9961), .B2(n6783), .ZN(n6784)
         );
  INV_X1 U8526 ( .A(n6784), .ZN(n6785) );
  OAI21_X1 U8527 ( .B1(n7040), .B2(n6560), .A(n6785), .ZN(P1_U3459) );
  NAND2_X1 U8528 ( .A1(n6786), .A2(n8006), .ZN(n6787) );
  XNOR2_X1 U8529 ( .A(n9183), .B(n9924), .ZN(n8054) );
  INV_X1 U8530 ( .A(n8054), .ZN(n6789) );
  OAI21_X1 U8531 ( .B1(n6790), .B2(n6789), .A(n6818), .ZN(n9934) );
  INV_X1 U8532 ( .A(n9934), .ZN(n6797) );
  INV_X1 U8533 ( .A(n9958), .ZN(n9962) );
  NAND2_X1 U8534 ( .A1(n6786), .A2(n7038), .ZN(n6791) );
  NAND2_X1 U8535 ( .A1(n6792), .A2(n6791), .ZN(n6823) );
  XNOR2_X1 U8536 ( .A(n6823), .B(n8054), .ZN(n6794) );
  AOI21_X1 U8537 ( .B1(n6794), .B2(n9910), .A(n6793), .ZN(n9937) );
  AND2_X1 U8538 ( .A1(n6796), .A2(n7029), .ZN(n7301) );
  INV_X1 U8539 ( .A(n7301), .ZN(n6795) );
  OAI211_X1 U8540 ( .C1(n7029), .C2(n6796), .A(n6795), .B(n9917), .ZN(n9932)
         );
  OAI211_X1 U8541 ( .C1(n6797), .C2(n9962), .A(n9937), .B(n9932), .ZN(n7031)
         );
  INV_X1 U8542 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6798) );
  OAI22_X1 U8543 ( .A1(n9685), .A2(n7029), .B1(n9961), .B2(n6798), .ZN(n6799)
         );
  AOI21_X1 U8544 ( .B1(n7031), .B2(n9961), .A(n6799), .ZN(n6800) );
  INV_X1 U8545 ( .A(n6800), .ZN(P1_U3462) );
  NAND2_X1 U8546 ( .A1(n6803), .A2(n6802), .ZN(n6810) );
  INV_X1 U8547 ( .A(n6810), .ZN(n7090) );
  NAND2_X1 U8548 ( .A1(n6806), .A2(n6805), .ZN(n6808) );
  AOI21_X1 U8549 ( .B1(n6808), .B2(n9910), .A(n6807), .ZN(n6812) );
  NAND2_X1 U8550 ( .A1(n6810), .A2(n6809), .ZN(n6811) );
  AND2_X1 U8551 ( .A1(n6812), .A2(n6811), .ZN(n7087) );
  NAND2_X1 U8552 ( .A1(n6666), .A2(n7066), .ZN(n6813) );
  NAND3_X1 U8553 ( .A1(n6814), .A2(n9917), .A3(n6813), .ZN(n7085) );
  OAI211_X1 U8554 ( .C1(n7090), .C2(n7514), .A(n7087), .B(n7085), .ZN(n7027)
         );
  INV_X1 U8555 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6815) );
  OAI22_X1 U8556 ( .A1(n9685), .A2(n7025), .B1(n9961), .B2(n6815), .ZN(n6816)
         );
  AOI21_X1 U8557 ( .B1(n9961), .B2(n7027), .A(n6816), .ZN(n6817) );
  INV_X1 U8558 ( .A(n6817), .ZN(P1_U3456) );
  INV_X1 U8559 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U8560 ( .A1(n6819), .A2(n7303), .ZN(n8003) );
  NAND2_X1 U8561 ( .A1(n9182), .A2(n9943), .ZN(n8010) );
  NAND2_X1 U8562 ( .A1(n8003), .A2(n8010), .ZN(n8052) );
  NAND2_X1 U8563 ( .A1(n9943), .A2(n6819), .ZN(n6820) );
  NAND2_X1 U8564 ( .A1(n7298), .A2(n6820), .ZN(n6821) );
  INV_X1 U8565 ( .A(n7012), .ZN(n7110) );
  NAND2_X1 U8566 ( .A1(n7110), .A2(n9181), .ZN(n8118) );
  NAND2_X1 U8567 ( .A1(n6976), .A2(n7012), .ZN(n8115) );
  AND2_X1 U8568 ( .A1(n8118), .A2(n8115), .ZN(n8056) );
  INV_X1 U8569 ( .A(n8056), .ZN(n7015) );
  NAND2_X1 U8570 ( .A1(n6821), .A2(n7015), .ZN(n7011) );
  OAI21_X1 U8571 ( .B1(n6821), .B2(n7015), .A(n7011), .ZN(n6822) );
  INV_X1 U8572 ( .A(n6822), .ZN(n7115) );
  NAND2_X1 U8573 ( .A1(n9183), .A2(n7029), .ZN(n8011) );
  NAND2_X1 U8574 ( .A1(n6823), .A2(n8011), .ZN(n6825) );
  NAND2_X1 U8575 ( .A1(n4634), .A2(n9924), .ZN(n6824) );
  NAND2_X1 U8576 ( .A1(n6825), .A2(n6824), .ZN(n7305) );
  NAND2_X1 U8577 ( .A1(n7305), .A2(n8010), .ZN(n8005) );
  NAND2_X1 U8578 ( .A1(n8005), .A2(n8003), .ZN(n8117) );
  XNOR2_X1 U8579 ( .A(n8117), .B(n8056), .ZN(n6827) );
  AOI22_X1 U8580 ( .A1(n9180), .A2(n9758), .B1(n9761), .B2(n9182), .ZN(n6901)
         );
  INV_X1 U8581 ( .A(n6901), .ZN(n6826) );
  AOI21_X1 U8582 ( .B1(n6827), .B2(n9910), .A(n6826), .ZN(n7107) );
  NAND2_X1 U8583 ( .A1(n7301), .A2(n9943), .ZN(n7300) );
  AOI21_X1 U8584 ( .B1(n7012), .B2(n7300), .A(n7020), .ZN(n7112) );
  AOI22_X1 U8585 ( .A1(n7112), .A2(n9917), .B1(n9580), .B2(n7012), .ZN(n6828)
         );
  OAI211_X1 U8586 ( .C1(n7115), .C2(n9962), .A(n7107), .B(n6828), .ZN(n6856)
         );
  NAND2_X1 U8587 ( .A1(n6856), .A2(n9961), .ZN(n6829) );
  OAI21_X1 U8588 ( .B1(n9961), .B2(n8907), .A(n6829), .ZN(P1_U3468) );
  XOR2_X1 U8589 ( .A(n6831), .B(n6830), .Z(n6845) );
  AOI21_X1 U8590 ( .B1(n10095), .B2(n6833), .A(n6951), .ZN(n6834) );
  NOR2_X1 U8591 ( .A1(n6834), .A2(n8559), .ZN(n6841) );
  AOI21_X1 U8592 ( .B1(n7132), .B2(n6835), .A(n6945), .ZN(n6839) );
  INV_X1 U8593 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8933) );
  NOR2_X1 U8594 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8933), .ZN(n6917) );
  INV_X1 U8595 ( .A(n6917), .ZN(n6838) );
  INV_X1 U8596 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6836) );
  OR2_X1 U8597 ( .A1(n8561), .A2(n6836), .ZN(n6837) );
  OAI211_X1 U8598 ( .C1(n6839), .C2(n8565), .A(n6838), .B(n6837), .ZN(n6840)
         );
  AOI211_X1 U8599 ( .C1(n8553), .C2(n6842), .A(n6841), .B(n6840), .ZN(n6843)
         );
  OAI21_X1 U8600 ( .B1(n6845), .B2(n6844), .A(n6843), .ZN(P2_U3189) );
  INV_X1 U8601 ( .A(n7828), .ZN(n7773) );
  XNOR2_X1 U8602 ( .A(n7773), .B(n7822), .ZN(n10011) );
  AND2_X1 U8603 ( .A1(n6935), .A2(n7767), .ZN(n6866) );
  INV_X1 U8604 ( .A(n6866), .ZN(n6846) );
  NAND2_X1 U8605 ( .A1(n7610), .A2(n6846), .ZN(n6847) );
  NAND2_X1 U8606 ( .A1(n8723), .A2(n6847), .ZN(n8765) );
  OAI21_X1 U8607 ( .B1(n6848), .B2(n7828), .A(n6929), .ZN(n6850) );
  INV_X1 U8608 ( .A(n8754), .ZN(n8737) );
  AOI222_X1 U8609 ( .A1(n8752), .A2(n6850), .B1(n8454), .B2(n8737), .C1(n6849), 
        .C2(n8739), .ZN(n10010) );
  MUX2_X1 U8610 ( .A(n6625), .B(n10010), .S(n8723), .Z(n6852) );
  INV_X1 U8611 ( .A(n8642), .ZN(n8761) );
  AOI22_X1 U8612 ( .A1(n8762), .A2(n6459), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8761), .ZN(n6851) );
  OAI211_X1 U8613 ( .C1(n10011), .C2(n8765), .A(n6852), .B(n6851), .ZN(
        P2_U3232) );
  AND2_X1 U8614 ( .A1(n7053), .A2(n6853), .ZN(n6854) );
  AND2_X2 U8615 ( .A1(n6855), .A2(n6854), .ZN(n9978) );
  INV_X1 U8616 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6858) );
  NAND2_X1 U8617 ( .A1(n6856), .A2(n9978), .ZN(n6857) );
  OAI21_X1 U8618 ( .B1(n9978), .B2(n6858), .A(n6857), .ZN(P1_U3527) );
  XNOR2_X1 U8619 ( .A(n8451), .B(n6867), .ZN(n7774) );
  INV_X1 U8620 ( .A(n7774), .ZN(n6860) );
  XNOR2_X1 U8621 ( .A(n6859), .B(n6860), .ZN(n10033) );
  INV_X1 U8622 ( .A(n7610), .ZN(n6933) );
  NAND2_X1 U8623 ( .A1(n10033), .A2(n6933), .ZN(n6865) );
  XNOR2_X1 U8624 ( .A(n7044), .B(n7774), .ZN(n6863) );
  NAND2_X1 U8625 ( .A1(n8452), .A2(n8739), .ZN(n6861) );
  OAI21_X1 U8626 ( .B1(n6919), .B2(n8754), .A(n6861), .ZN(n6862) );
  AOI21_X1 U8627 ( .B1(n6863), .B2(n8752), .A(n6862), .ZN(n6864) );
  AND2_X1 U8628 ( .A1(n6865), .A2(n6864), .ZN(n10035) );
  NAND2_X1 U8629 ( .A1(n8723), .A2(n6866), .ZN(n8586) );
  INV_X1 U8630 ( .A(n8586), .ZN(n7134) );
  INV_X1 U8631 ( .A(n8762), .ZN(n8575) );
  NOR2_X1 U8632 ( .A1(n8575), .A2(n6867), .ZN(n6871) );
  OAI22_X1 U8633 ( .A1(n8723), .A2(n6869), .B1(n6868), .B2(n8642), .ZN(n6870)
         );
  AOI211_X1 U8634 ( .C1(n10033), .C2(n7134), .A(n6871), .B(n6870), .ZN(n6872)
         );
  OAI21_X1 U8635 ( .B1(n10035), .B2(n7496), .A(n6872), .ZN(P2_U3228) );
  AOI21_X1 U8636 ( .B1(n6876), .B2(n6875), .A(n6874), .ZN(n6880) );
  AOI22_X1 U8637 ( .A1(n9761), .A2(n9180), .B1(n9178), .B2(n9758), .ZN(n7095)
         );
  NAND2_X1 U8638 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9718) );
  NAND2_X1 U8639 ( .A1(n4282), .A2(n7263), .ZN(n6877) );
  OAI211_X1 U8640 ( .C1(n9787), .C2(n7095), .A(n9718), .B(n6877), .ZN(n6878)
         );
  AOI21_X1 U8641 ( .B1(n9140), .B2(n7101), .A(n6878), .ZN(n6879) );
  OAI21_X1 U8642 ( .B1(n6880), .B2(n9792), .A(n6879), .ZN(P1_U3213) );
  INV_X1 U8643 ( .A(n6881), .ZN(n6884) );
  INV_X1 U8644 ( .A(n9873), .ZN(n7693) );
  OAI222_X1 U8645 ( .A1(n8303), .A2(n6882), .B1(n9694), .B2(n6884), .C1(
        P1_U3086), .C2(n7693), .ZN(P1_U3339) );
  OAI222_X1 U8646 ( .A1(n6885), .A2(P2_U3151), .B1(n7666), .B2(n6884), .C1(
        n6883), .C2(n7734), .ZN(P2_U3279) );
  NAND2_X1 U8647 ( .A1(n7844), .A2(n7849), .ZN(n7839) );
  XNOR2_X1 U8648 ( .A(n6886), .B(n7839), .ZN(n10027) );
  XNOR2_X1 U8649 ( .A(n6887), .B(n7839), .ZN(n6888) );
  AOI222_X1 U8650 ( .A1(n8752), .A2(n6888), .B1(n8451), .B2(n8737), .C1(n8453), 
        .C2(n8739), .ZN(n10026) );
  MUX2_X1 U8651 ( .A(n6889), .B(n10026), .S(n8723), .Z(n6893) );
  AOI22_X1 U8652 ( .A1(n8762), .A2(n6891), .B1(n8761), .B2(n6890), .ZN(n6892)
         );
  OAI211_X1 U8653 ( .C1(n8765), .C2(n10027), .A(n6893), .B(n6892), .ZN(
        P2_U3229) );
  INV_X1 U8654 ( .A(n6894), .ZN(n7109) );
  XNOR2_X1 U8655 ( .A(n6895), .B(n6896), .ZN(n6897) );
  NAND2_X1 U8656 ( .A1(n6897), .A2(n6898), .ZN(n6970) );
  OAI21_X1 U8657 ( .B1(n6898), .B2(n6897), .A(n6970), .ZN(n6899) );
  NAND2_X1 U8658 ( .A1(n6899), .A2(n9158), .ZN(n6904) );
  OAI22_X1 U8659 ( .A1(n9787), .A2(n6901), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6900), .ZN(n6902) );
  AOI21_X1 U8660 ( .B1(n7012), .B2(n4282), .A(n6902), .ZN(n6903) );
  OAI211_X1 U8661 ( .C1(n9797), .C2(n7109), .A(n6904), .B(n6903), .ZN(P1_U3227) );
  INV_X1 U8662 ( .A(n6905), .ZN(n10043) );
  XNOR2_X1 U8663 ( .A(n6905), .B(n6714), .ZN(n6906) );
  NAND2_X1 U8664 ( .A1(n6906), .A2(n7072), .ZN(n6998) );
  INV_X1 U8665 ( .A(n6906), .ZN(n6907) );
  NAND2_X1 U8666 ( .A1(n6907), .A2(n8449), .ZN(n6908) );
  NAND2_X1 U8667 ( .A1(n6998), .A2(n6908), .ZN(n6912) );
  AND2_X1 U8668 ( .A1(n6909), .A2(n8450), .ZN(n6911) );
  NOR2_X1 U8669 ( .A1(n6912), .A2(n6911), .ZN(n6910) );
  INV_X1 U8670 ( .A(n6911), .ZN(n6914) );
  INV_X1 U8671 ( .A(n6912), .ZN(n6913) );
  AOI21_X1 U8672 ( .B1(n6915), .B2(n6914), .A(n6913), .ZN(n6916) );
  OAI21_X1 U8673 ( .B1(n4365), .B2(n6916), .A(n9742), .ZN(n6922) );
  AOI21_X1 U8674 ( .B1(n8410), .B2(n8448), .A(n6917), .ZN(n6918) );
  OAI21_X1 U8675 ( .B1(n6919), .B2(n8412), .A(n6918), .ZN(n6920) );
  AOI21_X1 U8676 ( .B1(n7131), .B2(n8434), .A(n6920), .ZN(n6921) );
  OAI211_X1 U8677 ( .C1(n10043), .C2(n8438), .A(n6922), .B(n6921), .ZN(
        P2_U3153) );
  OAI21_X1 U8678 ( .B1(n6924), .B2(n7772), .A(n6923), .ZN(n10018) );
  INV_X1 U8679 ( .A(n8739), .ZN(n8753) );
  OAI22_X1 U8680 ( .A1(n6926), .A2(n8753), .B1(n6925), .B2(n8754), .ZN(n6932)
         );
  NAND2_X1 U8681 ( .A1(n6927), .A2(n7829), .ZN(n6982) );
  NAND3_X1 U8682 ( .A1(n6929), .A2(n7772), .A3(n6928), .ZN(n6930) );
  INV_X1 U8683 ( .A(n8752), .ZN(n10004) );
  AOI21_X1 U8684 ( .B1(n6982), .B2(n6930), .A(n10004), .ZN(n6931) );
  AOI211_X1 U8685 ( .C1(n6933), .C2(n10018), .A(n6932), .B(n6931), .ZN(n10015)
         );
  NAND2_X1 U8686 ( .A1(n8761), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6934) );
  OAI211_X1 U8687 ( .C1(n6935), .C2(n10014), .A(n10015), .B(n6934), .ZN(n6936)
         );
  MUX2_X1 U8688 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6936), .S(n8723), .Z(n6937)
         );
  AOI21_X1 U8689 ( .B1(n7134), .B2(n10018), .A(n6937), .ZN(n6938) );
  INV_X1 U8690 ( .A(n6938), .ZN(P2_U3231) );
  OAI21_X1 U8691 ( .B1(n6941), .B2(n6940), .A(n6939), .ZN(n6942) );
  NAND2_X1 U8692 ( .A1(n6942), .A2(n9981), .ZN(n6960) );
  OR3_X1 U8693 ( .A1(n6945), .A2(n6944), .A3(n6943), .ZN(n6946) );
  AOI21_X1 U8694 ( .B1(n6947), .B2(n6946), .A(n8565), .ZN(n6957) );
  INV_X1 U8695 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6955) );
  INV_X1 U8696 ( .A(n6948), .ZN(n6949) );
  NOR3_X1 U8697 ( .A1(n6951), .A2(n6950), .A3(n6949), .ZN(n6952) );
  OAI21_X1 U8698 ( .B1(n6953), .B2(n6952), .A(n10000), .ZN(n6954) );
  NAND2_X1 U8699 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7002) );
  OAI211_X1 U8700 ( .C1(n8561), .C2(n6955), .A(n6954), .B(n7002), .ZN(n6956)
         );
  AOI211_X1 U8701 ( .C1(n8553), .C2(n6958), .A(n6957), .B(n6956), .ZN(n6959)
         );
  NAND2_X1 U8702 ( .A1(n6960), .A2(n6959), .ZN(P2_U3190) );
  INV_X1 U8703 ( .A(n6961), .ZN(n6964) );
  INV_X1 U8704 ( .A(n9882), .ZN(n7708) );
  OAI222_X1 U8705 ( .A1(n8303), .A2(n6962), .B1(n7742), .B2(n6964), .C1(
        P1_U3086), .C2(n7708), .ZN(P1_U3338) );
  OAI222_X1 U8706 ( .A1(n6965), .A2(P2_U3151), .B1(n7666), .B2(n6964), .C1(
        n6963), .C2(n7734), .ZN(P2_U3278) );
  INV_X1 U8707 ( .A(n6966), .ZN(n7009) );
  AOI22_X1 U8708 ( .A1(n6968), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n6967), .ZN(n6969) );
  OAI21_X1 U8709 ( .B1(n7009), .B2(n9035), .A(n6969), .ZN(P2_U3277) );
  OAI21_X1 U8710 ( .B1(n6971), .B2(n6895), .A(n6970), .ZN(n6975) );
  XNOR2_X1 U8711 ( .A(n6973), .B(n6972), .ZN(n6974) );
  XNOR2_X1 U8712 ( .A(n6975), .B(n6974), .ZN(n6980) );
  INV_X1 U8713 ( .A(n7222), .ZN(n7034) );
  OAI22_X1 U8714 ( .A1(n6976), .A2(n9163), .B1(n7093), .B2(n9161), .ZN(n7018)
         );
  AOI22_X1 U8715 ( .A1(n9164), .A2(n7018), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n6977) );
  OAI21_X1 U8716 ( .B1(n9143), .B2(n7034), .A(n6977), .ZN(n6978) );
  AOI21_X1 U8717 ( .B1(n9140), .B2(n7223), .A(n6978), .ZN(n6979) );
  OAI21_X1 U8718 ( .B1(n6980), .B2(n9792), .A(n6979), .ZN(P1_U3239) );
  NAND3_X1 U8719 ( .A1(n6982), .A2(n6259), .A3(n6981), .ZN(n6983) );
  AND2_X1 U8720 ( .A1(n6984), .A2(n6983), .ZN(n6985) );
  OAI222_X1 U8721 ( .A1(n8754), .A2(n6987), .B1(n8753), .B2(n6986), .C1(n10004), .C2(n6985), .ZN(n10021) );
  INV_X1 U8722 ( .A(n10021), .ZN(n6996) );
  OAI21_X1 U8723 ( .B1(n6989), .B2(n6259), .A(n6988), .ZN(n10023) );
  INV_X1 U8724 ( .A(n8765), .ZN(n7564) );
  AOI22_X1 U8725 ( .A1(n8762), .A2(n6991), .B1(n8761), .B2(n6990), .ZN(n6992)
         );
  OAI21_X1 U8726 ( .B1(n6993), .B2(n8715), .A(n6992), .ZN(n6994) );
  AOI21_X1 U8727 ( .B1(n10023), .B2(n7564), .A(n6994), .ZN(n6995) );
  OAI21_X1 U8728 ( .B1(n6996), .B2(n7496), .A(n6995), .ZN(P2_U3230) );
  INV_X1 U8729 ( .A(n6997), .ZN(n7079) );
  NOR2_X1 U8730 ( .A1(n7079), .A2(n10072), .ZN(n10049) );
  INV_X1 U8731 ( .A(n10049), .ZN(n7007) );
  XNOR2_X1 U8732 ( .A(n6997), .B(n6714), .ZN(n7272) );
  XNOR2_X1 U8733 ( .A(n7272), .B(n8448), .ZN(n6999) );
  NOR3_X1 U8734 ( .A1(n4365), .A2(n4410), .A3(n6999), .ZN(n7001) );
  INV_X1 U8735 ( .A(n7274), .ZN(n7000) );
  OAI21_X1 U8736 ( .B1(n7001), .B2(n7000), .A(n9742), .ZN(n7006) );
  NAND2_X1 U8737 ( .A1(n9737), .A2(n8449), .ZN(n7003) );
  OAI211_X1 U8738 ( .C1(n7374), .C2(n9734), .A(n7003), .B(n7002), .ZN(n7004)
         );
  AOI21_X1 U8739 ( .B1(n7077), .B2(n8434), .A(n7004), .ZN(n7005) );
  OAI211_X1 U8740 ( .C1(n7008), .C2(n7007), .A(n7006), .B(n7005), .ZN(P2_U3161) );
  INV_X1 U8741 ( .A(n7709), .ZN(n9897) );
  OAI222_X1 U8742 ( .A1(n8303), .A2(n7010), .B1(n9897), .B2(P1_U3086), .C1(
        n7742), .C2(n7009), .ZN(P1_U3337) );
  OR2_X1 U8743 ( .A1(n7222), .A2(n7013), .ZN(n8124) );
  NAND2_X1 U8744 ( .A1(n7222), .A2(n7013), .ZN(n8120) );
  AND2_X1 U8745 ( .A1(n8124), .A2(n8120), .ZN(n8055) );
  INV_X1 U8746 ( .A(n8055), .ZN(n7017) );
  OAI21_X1 U8747 ( .B1(n7014), .B2(n7017), .A(n7097), .ZN(n7228) );
  INV_X1 U8748 ( .A(n7228), .ZN(n7021) );
  OR2_X1 U8749 ( .A1(n8117), .A2(n7015), .ZN(n7016) );
  NAND2_X1 U8750 ( .A1(n7016), .A2(n8118), .ZN(n7452) );
  XNOR2_X1 U8751 ( .A(n7452), .B(n7017), .ZN(n7019) );
  AOI21_X1 U8752 ( .B1(n7019), .B2(n9910), .A(n7018), .ZN(n7230) );
  OAI211_X1 U8753 ( .C1(n7020), .C2(n7034), .A(n7100), .B(n9917), .ZN(n7226)
         );
  OAI211_X1 U8754 ( .C1(n7021), .C2(n9962), .A(n7230), .B(n7226), .ZN(n7036)
         );
  INV_X1 U8755 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7022) );
  OAI22_X1 U8756 ( .A1(n9685), .A2(n7034), .B1(n9961), .B2(n7022), .ZN(n7023)
         );
  AOI21_X1 U8757 ( .B1(n7036), .B2(n9961), .A(n7023), .ZN(n7024) );
  INV_X1 U8758 ( .A(n7024), .ZN(P1_U3471) );
  NAND2_X1 U8759 ( .A1(n9978), .A2(n9580), .ZN(n9627) );
  OAI22_X1 U8760 ( .A1(n9627), .A2(n7025), .B1(n9978), .B2(n6487), .ZN(n7026)
         );
  AOI21_X1 U8761 ( .B1(n9978), .B2(n7027), .A(n7026), .ZN(n7028) );
  INV_X1 U8762 ( .A(n7028), .ZN(P1_U3523) );
  OAI22_X1 U8763 ( .A1(n9627), .A2(n7029), .B1(n9978), .B2(n6490), .ZN(n7030)
         );
  AOI21_X1 U8764 ( .B1(n7031), .B2(n9978), .A(n7030), .ZN(n7032) );
  INV_X1 U8765 ( .A(n7032), .ZN(P1_U3525) );
  INV_X1 U8766 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7033) );
  OAI22_X1 U8767 ( .A1(n9627), .A2(n7034), .B1(n9978), .B2(n7033), .ZN(n7035)
         );
  AOI21_X1 U8768 ( .B1(n7036), .B2(n9978), .A(n7035), .ZN(n7037) );
  INV_X1 U8769 ( .A(n7037), .ZN(P1_U3528) );
  INV_X1 U8770 ( .A(n9627), .ZN(n7522) );
  AOI22_X1 U8771 ( .A1(n7522), .A2(n7038), .B1(n9979), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n7039) );
  OAI21_X1 U8772 ( .B1(n7040), .B2(n9979), .A(n7039), .ZN(P1_U3524) );
  AND2_X1 U8773 ( .A1(n7042), .A2(n7125), .ZN(n7775) );
  XNOR2_X1 U8774 ( .A(n7041), .B(n7775), .ZN(n10037) );
  OR2_X1 U8775 ( .A1(n7044), .A2(n7043), .ZN(n7046) );
  NAND2_X1 U8776 ( .A1(n7046), .A2(n7045), .ZN(n7047) );
  XOR2_X1 U8777 ( .A(n7775), .B(n7047), .Z(n7048) );
  AOI222_X1 U8778 ( .A1(n8752), .A2(n7048), .B1(n8449), .B2(n8737), .C1(n8451), 
        .C2(n8739), .ZN(n10038) );
  MUX2_X1 U8779 ( .A(n5824), .B(n10038), .S(n8723), .Z(n7052) );
  AOI22_X1 U8780 ( .A1(n8762), .A2(n7050), .B1(n8761), .B2(n7049), .ZN(n7051)
         );
  OAI211_X1 U8781 ( .C1(n10037), .C2(n8765), .A(n7052), .B(n7051), .ZN(
        P2_U3227) );
  NAND3_X1 U8782 ( .A1(n7055), .A2(n7054), .A3(n7053), .ZN(n7065) );
  NAND2_X1 U8783 ( .A1(n7057), .A2(n7056), .ZN(n7061) );
  INV_X1 U8784 ( .A(n7061), .ZN(n7063) );
  INV_X1 U8785 ( .A(n9531), .ZN(n9927) );
  INV_X1 U8786 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n8920) );
  AOI21_X1 U8787 ( .B1(n9927), .B2(P1_REG3_REG_0__SCAN_IN), .A(n7058), .ZN(
        n7059) );
  OAI21_X1 U8788 ( .B1(n7061), .B2(n7060), .A(n7059), .ZN(n7062) );
  AOI21_X1 U8789 ( .B1(n7063), .B2(n5060), .A(n7062), .ZN(n7069) );
  INV_X1 U8790 ( .A(n9530), .ZN(n9925) );
  OR2_X1 U8791 ( .A1(n7065), .A2(n5437), .ZN(n9931) );
  NOR2_X1 U8792 ( .A1(n9931), .A2(n9527), .ZN(n9325) );
  OAI21_X1 U8793 ( .B1(n9925), .B2(n9325), .A(n7066), .ZN(n7068) );
  NAND2_X1 U8794 ( .A1(n9928), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7067) );
  OAI211_X1 U8795 ( .C1(n9938), .C2(n7069), .A(n7068), .B(n7067), .ZN(P1_U3293) );
  XNOR2_X1 U8796 ( .A(n7070), .B(n4819), .ZN(n7071) );
  OAI222_X1 U8797 ( .A1(n8754), .A2(n7374), .B1(n8753), .B2(n7072), .C1(n10004), .C2(n7071), .ZN(n10048) );
  INV_X1 U8798 ( .A(n10048), .ZN(n7082) );
  NAND2_X1 U8799 ( .A1(n7073), .A2(n7074), .ZN(n7076) );
  XNOR2_X1 U8800 ( .A(n7076), .B(n7075), .ZN(n10050) );
  AOI22_X1 U8801 ( .A1(n7496), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8761), .B2(
        n7077), .ZN(n7078) );
  OAI21_X1 U8802 ( .B1(n7079), .B2(n8575), .A(n7078), .ZN(n7080) );
  AOI21_X1 U8803 ( .B1(n10050), .B2(n7564), .A(n7080), .ZN(n7081) );
  OAI21_X1 U8804 ( .B1(n7082), .B2(n7496), .A(n7081), .ZN(P2_U3225) );
  OR2_X1 U8805 ( .A1(n9938), .A2(n7083), .ZN(n7487) );
  INV_X1 U8806 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7084) );
  OAI22_X1 U8807 ( .A1(n9931), .A2(n7085), .B1(n7084), .B2(n9531), .ZN(n7086)
         );
  AOI21_X1 U8808 ( .B1(n9925), .B2(n6666), .A(n7086), .ZN(n7089) );
  MUX2_X1 U8809 ( .A(n7087), .B(n6476), .S(n9938), .Z(n7088) );
  OAI211_X1 U8810 ( .C1(n7090), .C2(n7487), .A(n7089), .B(n7088), .ZN(P1_U3292) );
  INV_X1 U8811 ( .A(n7452), .ZN(n7092) );
  INV_X1 U8812 ( .A(n8120), .ZN(n7091) );
  AOI21_X1 U8813 ( .B1(n7092), .B2(n8124), .A(n7091), .ZN(n7094) );
  OR2_X1 U8814 ( .A1(n7263), .A2(n7093), .ZN(n7453) );
  NAND2_X1 U8815 ( .A1(n7263), .A2(n7093), .ZN(n7237) );
  AND2_X1 U8816 ( .A1(n7453), .A2(n7237), .ZN(n8125) );
  NOR2_X1 U8817 ( .A1(n7094), .A2(n7098), .ZN(n7239) );
  AOI21_X1 U8818 ( .B1(n7094), .B2(n7098), .A(n7239), .ZN(n7096) );
  OAI21_X1 U8819 ( .B1(n7096), .B2(n9469), .A(n7095), .ZN(n7255) );
  INV_X1 U8820 ( .A(n7255), .ZN(n7106) );
  OAI21_X1 U8821 ( .B1(n7099), .B2(n7098), .A(n7173), .ZN(n7257) );
  OAI21_X2 U8822 ( .B1(n9938), .B2(n7478), .A(n7487), .ZN(n9935) );
  AOI211_X1 U8823 ( .C1(n7263), .C2(n7100), .A(n9527), .B(n7182), .ZN(n7256)
         );
  INV_X1 U8824 ( .A(n9931), .ZN(n9921) );
  NAND2_X1 U8825 ( .A1(n7256), .A2(n9921), .ZN(n7103) );
  AOI22_X1 U8826 ( .A1(n9928), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7101), .B2(
        n9927), .ZN(n7102) );
  OAI211_X1 U8827 ( .C1(n4468), .C2(n9530), .A(n7103), .B(n7102), .ZN(n7104)
         );
  AOI21_X1 U8828 ( .B1(n7257), .B2(n9935), .A(n7104), .ZN(n7105) );
  OAI21_X1 U8829 ( .B1(n7106), .B2(n9928), .A(n7105), .ZN(P1_U3286) );
  INV_X1 U8830 ( .A(n9935), .ZN(n9518) );
  INV_X1 U8831 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7108) );
  INV_X1 U8832 ( .A(n9928), .ZN(n9534) );
  MUX2_X1 U8833 ( .A(n7108), .B(n7107), .S(n9534), .Z(n7114) );
  OAI22_X1 U8834 ( .A1(n9530), .A2(n7110), .B1(n7109), .B2(n9531), .ZN(n7111)
         );
  AOI21_X1 U8835 ( .B1(n9325), .B2(n7112), .A(n7111), .ZN(n7113) );
  OAI211_X1 U8836 ( .C1(n9518), .C2(n7115), .A(n7114), .B(n7113), .ZN(P1_U3288) );
  INV_X1 U8837 ( .A(n7487), .ZN(n7122) );
  AOI22_X1 U8838 ( .A1(n9921), .A2(n7116), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9927), .ZN(n7117) );
  OAI21_X1 U8839 ( .B1(n8006), .B2(n9530), .A(n7117), .ZN(n7120) );
  MUX2_X1 U8840 ( .A(n7118), .B(P1_REG2_REG_2__SCAN_IN), .S(n9938), .Z(n7119)
         );
  AOI211_X1 U8841 ( .C1(n7122), .C2(n7121), .A(n7120), .B(n7119), .ZN(n7123)
         );
  INV_X1 U8842 ( .A(n7123), .ZN(P1_U3291) );
  OAI21_X1 U8843 ( .B1(n7124), .B2(n7778), .A(n7073), .ZN(n10044) );
  AOI22_X1 U8844 ( .A1(n8739), .A2(n8450), .B1(n8448), .B2(n8737), .ZN(n7130)
         );
  NAND2_X1 U8845 ( .A1(n7126), .A2(n7125), .ZN(n7127) );
  XNOR2_X1 U8846 ( .A(n7127), .B(n7778), .ZN(n7128) );
  NAND2_X1 U8847 ( .A1(n7128), .A2(n8752), .ZN(n7129) );
  OAI211_X1 U8848 ( .C1(n10044), .C2(n7610), .A(n7130), .B(n7129), .ZN(n10046)
         );
  AOI21_X1 U8849 ( .B1(n8761), .B2(n7131), .A(n10046), .ZN(n7137) );
  INV_X1 U8850 ( .A(n10044), .ZN(n7135) );
  OAI22_X1 U8851 ( .A1(n8575), .A2(n10043), .B1(n7132), .B2(n8715), .ZN(n7133)
         );
  AOI21_X1 U8852 ( .B1(n7135), .B2(n7134), .A(n7133), .ZN(n7136) );
  OAI21_X1 U8853 ( .B1(n7137), .B2(n7496), .A(n7136), .ZN(P2_U3226) );
  INV_X1 U8854 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10114) );
  INV_X1 U8855 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9888) );
  INV_X1 U8856 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8534) );
  AOI22_X1 U8857 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n9888), .B2(n8534), .ZN(n10120) );
  NOR2_X1 U8858 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7138) );
  AOI21_X1 U8859 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7138), .ZN(n10123) );
  NOR2_X1 U8860 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7139) );
  AOI21_X1 U8861 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7139), .ZN(n10126) );
  NOR2_X1 U8862 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7140) );
  AOI21_X1 U8863 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7140), .ZN(n10129) );
  INV_X1 U8864 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8465) );
  INV_X1 U8865 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9834) );
  AOI22_X1 U8866 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .B1(n8465), .B2(n9834), .ZN(n10132) );
  NOR2_X1 U8867 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7141) );
  AOI21_X1 U8868 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7141), .ZN(n10135) );
  NOR2_X1 U8869 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7142) );
  AOI21_X1 U8870 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7142), .ZN(n10138) );
  NOR2_X1 U8871 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7143) );
  AOI21_X1 U8872 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7143), .ZN(n10141) );
  NOR2_X1 U8873 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7144) );
  AOI21_X1 U8874 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7144), .ZN(n10150) );
  NOR2_X1 U8875 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7145) );
  AOI21_X1 U8876 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7145), .ZN(n10156) );
  NOR2_X1 U8877 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7146) );
  AOI21_X1 U8878 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7146), .ZN(n10153) );
  NOR2_X1 U8879 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7147) );
  AOI21_X1 U8880 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7147), .ZN(n10144) );
  NOR2_X1 U8881 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n7148) );
  AOI21_X1 U8882 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n7148), .ZN(n10147) );
  AND2_X1 U8883 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7149) );
  NOR2_X1 U8884 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7149), .ZN(n10109) );
  INV_X1 U8885 ( .A(n10109), .ZN(n10110) );
  NAND3_X1 U8886 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10111) );
  NAND2_X1 U8887 ( .A1(n10112), .A2(n10111), .ZN(n10108) );
  NAND2_X1 U8888 ( .A1(n10110), .A2(n10108), .ZN(n10159) );
  NAND2_X1 U8889 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7150) );
  OAI21_X1 U8890 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7150), .ZN(n10158) );
  NOR2_X1 U8891 ( .A1(n10159), .A2(n10158), .ZN(n10157) );
  AOI21_X1 U8892 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10157), .ZN(n10162) );
  NAND2_X1 U8893 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7151) );
  OAI21_X1 U8894 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7151), .ZN(n10161) );
  NOR2_X1 U8895 ( .A1(n10162), .A2(n10161), .ZN(n10160) );
  AOI21_X1 U8896 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10160), .ZN(n10165) );
  NOR2_X1 U8897 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7152) );
  AOI21_X1 U8898 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7152), .ZN(n10164) );
  NAND2_X1 U8899 ( .A1(n10165), .A2(n10164), .ZN(n10163) );
  OAI21_X1 U8900 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10163), .ZN(n10146) );
  NAND2_X1 U8901 ( .A1(n10147), .A2(n10146), .ZN(n10145) );
  OAI21_X1 U8902 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10145), .ZN(n10143) );
  NAND2_X1 U8903 ( .A1(n10144), .A2(n10143), .ZN(n10142) );
  OAI21_X1 U8904 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10142), .ZN(n10152) );
  NAND2_X1 U8905 ( .A1(n10153), .A2(n10152), .ZN(n10151) );
  OAI21_X1 U8906 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10151), .ZN(n10155) );
  NAND2_X1 U8907 ( .A1(n10156), .A2(n10155), .ZN(n10154) );
  OAI21_X1 U8908 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10154), .ZN(n10149) );
  NAND2_X1 U8909 ( .A1(n10150), .A2(n10149), .ZN(n10148) );
  OAI21_X1 U8910 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10148), .ZN(n10140) );
  NAND2_X1 U8911 ( .A1(n10141), .A2(n10140), .ZN(n10139) );
  OAI21_X1 U8912 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10139), .ZN(n10137) );
  NAND2_X1 U8913 ( .A1(n10138), .A2(n10137), .ZN(n10136) );
  OAI21_X1 U8914 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10136), .ZN(n10134) );
  NAND2_X1 U8915 ( .A1(n10135), .A2(n10134), .ZN(n10133) );
  OAI21_X1 U8916 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10133), .ZN(n10131) );
  NAND2_X1 U8917 ( .A1(n10132), .A2(n10131), .ZN(n10130) );
  OAI21_X1 U8918 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10130), .ZN(n10128) );
  NAND2_X1 U8919 ( .A1(n10129), .A2(n10128), .ZN(n10127) );
  OAI21_X1 U8920 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10127), .ZN(n10125) );
  NAND2_X1 U8921 ( .A1(n10126), .A2(n10125), .ZN(n10124) );
  OAI21_X1 U8922 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10124), .ZN(n10122) );
  NAND2_X1 U8923 ( .A1(n10123), .A2(n10122), .ZN(n10121) );
  OAI21_X1 U8924 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10121), .ZN(n10119) );
  NAND2_X1 U8925 ( .A1(n10120), .A2(n10119), .ZN(n10118) );
  OAI21_X1 U8926 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10118), .ZN(n10115) );
  NAND2_X1 U8927 ( .A1(n10114), .A2(n10115), .ZN(n7153) );
  NOR2_X1 U8928 ( .A1(n10114), .A2(n10115), .ZN(n10113) );
  AOI21_X1 U8929 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7153), .A(n10113), .ZN(
        n7155) );
  XNOR2_X1 U8930 ( .A(n4518), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7154) );
  XNOR2_X1 U8931 ( .A(n7155), .B(n7154), .ZN(ADD_1068_U4) );
  AOI21_X1 U8932 ( .B1(n7294), .B2(n7157), .A(n7156), .ZN(n7171) );
  OAI21_X1 U8933 ( .B1(n7160), .B2(n7159), .A(n7158), .ZN(n7169) );
  NAND2_X1 U8934 ( .A1(n8553), .A2(n7161), .ZN(n7163) );
  AND2_X1 U8935 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7268) );
  AOI21_X1 U8936 ( .B1(n9991), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7268), .ZN(
        n7162) );
  NAND2_X1 U8937 ( .A1(n7163), .A2(n7162), .ZN(n7168) );
  AOI21_X1 U8938 ( .B1(n10099), .B2(n7165), .A(n7164), .ZN(n7166) );
  NOR2_X1 U8939 ( .A1(n7166), .A2(n8559), .ZN(n7167) );
  AOI211_X1 U8940 ( .C1(n9981), .C2(n7169), .A(n7168), .B(n7167), .ZN(n7170)
         );
  OAI21_X1 U8941 ( .B1(n7171), .B2(n8565), .A(n7170), .ZN(P2_U3191) );
  NAND2_X1 U8942 ( .A1(n7173), .A2(n7172), .ZN(n7233) );
  XNOR2_X1 U8943 ( .A(n9790), .B(n9178), .ZN(n7176) );
  INV_X1 U8944 ( .A(n7176), .ZN(n7174) );
  XNOR2_X1 U8945 ( .A(n7233), .B(n7174), .ZN(n7334) );
  INV_X1 U8946 ( .A(n7334), .ZN(n7190) );
  INV_X1 U8947 ( .A(n7237), .ZN(n7175) );
  NOR2_X1 U8948 ( .A1(n7239), .A2(n7175), .ZN(n7177) );
  XNOR2_X1 U8949 ( .A(n7177), .B(n7176), .ZN(n7180) );
  NAND2_X1 U8950 ( .A1(n9179), .A2(n9761), .ZN(n7179) );
  NAND2_X1 U8951 ( .A1(n9760), .A2(n9758), .ZN(n7178) );
  AND2_X1 U8952 ( .A1(n7179), .A2(n7178), .ZN(n9786) );
  OAI21_X1 U8953 ( .B1(n7180), .B2(n9469), .A(n9786), .ZN(n7332) );
  INV_X1 U8954 ( .A(n7242), .ZN(n7183) );
  AOI211_X1 U8955 ( .C1(n9790), .C2(n7184), .A(n9527), .B(n7183), .ZN(n7333)
         );
  NAND2_X1 U8956 ( .A1(n7333), .A2(n9921), .ZN(n7187) );
  AOI22_X1 U8957 ( .A1(n9938), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7185), .B2(
        n9927), .ZN(n7186) );
  OAI211_X1 U8958 ( .C1(n7181), .C2(n9530), .A(n7187), .B(n7186), .ZN(n7188)
         );
  AOI21_X1 U8959 ( .B1(n7332), .B2(n9534), .A(n7188), .ZN(n7189) );
  OAI21_X1 U8960 ( .B1(n9518), .B2(n7190), .A(n7189), .ZN(P1_U3285) );
  INV_X1 U8961 ( .A(n7191), .ZN(n8302) );
  OAI222_X1 U8962 ( .A1(P2_U3151), .A2(n7193), .B1(n7666), .B2(n8302), .C1(
        n7192), .C2(n7734), .ZN(P2_U3276) );
  INV_X1 U8963 ( .A(n7680), .ZN(n7695) );
  NAND2_X1 U8964 ( .A1(n9705), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7194) );
  OAI21_X1 U8965 ( .B1(n9705), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7194), .ZN(
        n9701) );
  NOR2_X1 U8966 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n9248), .ZN(n7195) );
  AOI21_X1 U8967 ( .B1(n9248), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7195), .ZN(
        n9241) );
  NAND2_X1 U8968 ( .A1(n7210), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U8969 ( .A1(n7197), .A2(n7196), .ZN(n9220) );
  MUX2_X1 U8970 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7108), .S(n9218), .Z(n9221)
         );
  NAND2_X1 U8971 ( .A1(n9220), .A2(n9221), .ZN(n9219) );
  NAND2_X1 U8972 ( .A1(n9218), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7198) );
  NAND2_X1 U8973 ( .A1(n9219), .A2(n7198), .ZN(n9234) );
  INV_X1 U8974 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7199) );
  XNOR2_X1 U8975 ( .A(n9232), .B(n7199), .ZN(n9235) );
  NAND2_X1 U8976 ( .A1(n9234), .A2(n9235), .ZN(n9233) );
  NAND2_X1 U8977 ( .A1(n9232), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7200) );
  NAND2_X1 U8978 ( .A1(n9233), .A2(n7200), .ZN(n9708) );
  INV_X1 U8979 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n8981) );
  MUX2_X1 U8980 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n8981), .S(n9717), .Z(n9709)
         );
  AOI21_X1 U8981 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n9717), .A(n9710), .ZN(
        n9723) );
  NAND2_X1 U8982 ( .A1(n9729), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7201) );
  OAI21_X1 U8983 ( .B1(n9729), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7201), .ZN(
        n9722) );
  NOR2_X1 U8984 ( .A1(n9723), .A2(n9722), .ZN(n9721) );
  AOI21_X1 U8985 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9729), .A(n9721), .ZN(
        n9240) );
  NAND2_X1 U8986 ( .A1(n9241), .A2(n9240), .ZN(n9239) );
  OAI21_X1 U8987 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9248), .A(n9239), .ZN(
        n9702) );
  NOR2_X1 U8988 ( .A1(n9701), .A2(n9702), .ZN(n9700) );
  AOI21_X1 U8989 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9705), .A(n9700), .ZN(
        n9809) );
  INV_X1 U8990 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7202) );
  AOI22_X1 U8991 ( .A1(n7215), .A2(n7202), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n9818), .ZN(n9810) );
  NOR2_X1 U8992 ( .A1(n9809), .A2(n9810), .ZN(n9808) );
  AOI21_X1 U8993 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7215), .A(n9808), .ZN(
        n7206) );
  INV_X1 U8994 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7203) );
  MUX2_X1 U8995 ( .A(n7203), .B(P1_REG2_REG_12__SCAN_IN), .S(n7680), .Z(n7204)
         );
  INV_X1 U8996 ( .A(n7204), .ZN(n7205) );
  NAND2_X1 U8997 ( .A1(n7205), .A2(n7206), .ZN(n7679) );
  OAI21_X1 U8998 ( .B1(n7206), .B2(n7205), .A(n7679), .ZN(n7219) );
  NAND2_X1 U8999 ( .A1(n9705), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7207) );
  OAI21_X1 U9000 ( .B1(n9705), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7207), .ZN(
        n9698) );
  NOR2_X1 U9001 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9248), .ZN(n7208) );
  AOI21_X1 U9002 ( .B1(n9248), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7208), .ZN(
        n9246) );
  XNOR2_X1 U9003 ( .A(n9218), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9212) );
  AOI21_X1 U9004 ( .B1(n9218), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9211), .ZN(
        n9227) );
  XNOR2_X1 U9005 ( .A(n9232), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9226) );
  NOR2_X1 U9006 ( .A1(n9227), .A2(n9226), .ZN(n9225) );
  AOI21_X1 U9007 ( .B1(n9232), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9225), .ZN(
        n9714) );
  OR2_X1 U9008 ( .A1(n9717), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7212) );
  NAND2_X1 U9009 ( .A1(n9717), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7211) );
  NAND2_X1 U9010 ( .A1(n7212), .A2(n7211), .ZN(n9713) );
  NOR2_X1 U9011 ( .A1(n9714), .A2(n9713), .ZN(n9712) );
  AOI21_X1 U9012 ( .B1(n9717), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9712), .ZN(
        n9726) );
  NAND2_X1 U9013 ( .A1(n9729), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7213) );
  OAI21_X1 U9014 ( .B1(n9729), .B2(P1_REG1_REG_8__SCAN_IN), .A(n7213), .ZN(
        n9725) );
  NOR2_X1 U9015 ( .A1(n9698), .A2(n9699), .ZN(n9697) );
  AOI21_X1 U9016 ( .B1(n9705), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9697), .ZN(
        n9813) );
  INV_X1 U9017 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7214) );
  MUX2_X1 U9018 ( .A(n7214), .B(P1_REG1_REG_11__SCAN_IN), .S(n7215), .Z(n9814)
         );
  NOR2_X1 U9019 ( .A1(n9813), .A2(n9814), .ZN(n9812) );
  INV_X1 U9020 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7694) );
  MUX2_X1 U9021 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7694), .S(n7680), .Z(n7216)
         );
  OAI21_X1 U9022 ( .B1(n7217), .B2(n7216), .A(n7697), .ZN(n7218) );
  AOI22_X1 U9023 ( .A1(n9884), .A2(n7219), .B1(n9892), .B2(n7218), .ZN(n7221)
         );
  AND2_X1 U9024 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9769) );
  AOI21_X1 U9025 ( .B1(n9869), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n9769), .ZN(
        n7220) );
  OAI211_X1 U9026 ( .C1(n7695), .C2(n9898), .A(n7221), .B(n7220), .ZN(P1_U3255) );
  NAND2_X1 U9027 ( .A1(n9925), .A2(n7222), .ZN(n7225) );
  AOI22_X1 U9028 ( .A1(n9928), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7223), .B2(
        n9927), .ZN(n7224) );
  OAI211_X1 U9029 ( .C1(n7226), .C2(n9931), .A(n7225), .B(n7224), .ZN(n7227)
         );
  AOI21_X1 U9030 ( .B1(n7228), .B2(n9935), .A(n7227), .ZN(n7229) );
  OAI21_X1 U9031 ( .B1(n9938), .B2(n7230), .A(n7229), .ZN(P1_U3287) );
  NAND2_X1 U9032 ( .A1(n9790), .A2(n9178), .ZN(n7232) );
  AOI21_X2 U9033 ( .B1(n7233), .B2(n7232), .A(n7231), .ZN(n7447) );
  OR2_X1 U9034 ( .A1(n5265), .A2(n7234), .ZN(n8154) );
  INV_X1 U9035 ( .A(n8154), .ZN(n7236) );
  NAND2_X1 U9036 ( .A1(n5265), .A2(n7234), .ZN(n8151) );
  INV_X1 U9037 ( .A(n8151), .ZN(n7235) );
  XNOR2_X1 U9038 ( .A(n7447), .B(n7446), .ZN(n9952) );
  INV_X1 U9039 ( .A(n9952), .ZN(n7251) );
  NAND2_X1 U9040 ( .A1(n9790), .A2(n7238), .ZN(n8134) );
  AND2_X1 U9041 ( .A1(n8134), .A2(n7237), .ZN(n8129) );
  INV_X1 U9042 ( .A(n8129), .ZN(n7451) );
  OR2_X1 U9043 ( .A1(n9790), .A2(n7238), .ZN(n8132) );
  OAI21_X1 U9044 ( .B1(n7239), .B2(n7451), .A(n8132), .ZN(n7240) );
  XNOR2_X1 U9045 ( .A(n7240), .B(n7446), .ZN(n7241) );
  NAND2_X1 U9046 ( .A1(n9178), .A2(n9761), .ZN(n9123) );
  OAI21_X1 U9047 ( .B1(n7241), .B2(n9469), .A(n9123), .ZN(n9950) );
  AOI211_X1 U9048 ( .C1(n5265), .C2(n7242), .A(n9527), .B(n9919), .ZN(n7244)
         );
  NAND2_X1 U9049 ( .A1(n9177), .A2(n9758), .ZN(n9122) );
  INV_X1 U9050 ( .A(n9122), .ZN(n7243) );
  NOR2_X1 U9051 ( .A1(n7244), .A2(n7243), .ZN(n9948) );
  INV_X1 U9052 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7246) );
  INV_X1 U9053 ( .A(n9127), .ZN(n7245) );
  OAI22_X1 U9054 ( .A1(n9534), .A2(n7246), .B1(n7245), .B2(n9531), .ZN(n7247)
         );
  AOI21_X1 U9055 ( .B1(n9925), .B2(n5265), .A(n7247), .ZN(n7248) );
  OAI21_X1 U9056 ( .B1(n9948), .B2(n9931), .A(n7248), .ZN(n7249) );
  AOI21_X1 U9057 ( .B1(n9950), .B2(n9534), .A(n7249), .ZN(n7250) );
  OAI21_X1 U9058 ( .B1(n7251), .B2(n9518), .A(n7250), .ZN(P1_U3284) );
  INV_X1 U9059 ( .A(n7252), .ZN(n7283) );
  OAI222_X1 U9060 ( .A1(n7742), .A2(n7283), .B1(n7254), .B2(P1_U3086), .C1(
        n7253), .C2(n8303), .ZN(P1_U3335) );
  AOI211_X1 U9061 ( .C1(n9958), .C2(n7257), .A(n7256), .B(n7255), .ZN(n7266)
         );
  INV_X1 U9062 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7258) );
  NOR2_X1 U9063 ( .A1(n9978), .A2(n7258), .ZN(n7259) );
  AOI21_X1 U9064 ( .B1(n7522), .B2(n7263), .A(n7259), .ZN(n7260) );
  OAI21_X1 U9065 ( .B1(n7266), .B2(n9979), .A(n7260), .ZN(P1_U3529) );
  INV_X1 U9066 ( .A(n9685), .ZN(n7264) );
  INV_X1 U9067 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7261) );
  NOR2_X1 U9068 ( .A1(n9961), .A2(n7261), .ZN(n7262) );
  AOI21_X1 U9069 ( .B1(n7264), .B2(n7263), .A(n7262), .ZN(n7265) );
  OAI21_X1 U9070 ( .B1(n7266), .B2(n6560), .A(n7265), .ZN(P1_U3474) );
  INV_X1 U9071 ( .A(n7267), .ZN(n7293) );
  AOI21_X1 U9072 ( .B1(n8410), .B2(n8446), .A(n7268), .ZN(n7270) );
  OR2_X1 U9073 ( .A1(n8412), .A2(n7271), .ZN(n7269) );
  OAI211_X1 U9074 ( .C1(n7293), .C2(n9746), .A(n7270), .B(n7269), .ZN(n7280)
         );
  XNOR2_X1 U9075 ( .A(n10055), .B(n8293), .ZN(n7359) );
  XNOR2_X1 U9076 ( .A(n7359), .B(n7374), .ZN(n7278) );
  NAND2_X1 U9077 ( .A1(n7272), .A2(n7271), .ZN(n7273) );
  INV_X1 U9078 ( .A(n7362), .ZN(n7276) );
  AOI211_X1 U9079 ( .C1(n7278), .C2(n7277), .A(n8391), .B(n7276), .ZN(n7279)
         );
  AOI211_X1 U9080 ( .C1(n8369), .C2(n10055), .A(n7280), .B(n7279), .ZN(n7281)
         );
  INV_X1 U9081 ( .A(n7281), .ZN(P2_U3171) );
  OAI222_X1 U9082 ( .A1(n7284), .A2(P2_U3151), .B1(n7666), .B2(n7283), .C1(
        n7282), .C2(n7734), .ZN(P2_U3275) );
  NAND2_X1 U9083 ( .A1(n7286), .A2(n7288), .ZN(n7287) );
  NAND2_X1 U9084 ( .A1(n7285), .A2(n7287), .ZN(n10052) );
  XNOR2_X1 U9085 ( .A(n7289), .B(n6047), .ZN(n7290) );
  NAND2_X1 U9086 ( .A1(n7290), .A2(n8752), .ZN(n7292) );
  AOI22_X1 U9087 ( .A1(n8448), .A2(n8739), .B1(n8737), .B2(n8446), .ZN(n7291)
         );
  OAI211_X1 U9088 ( .C1(n7610), .C2(n10052), .A(n7292), .B(n7291), .ZN(n10053)
         );
  NAND2_X1 U9089 ( .A1(n10053), .A2(n8715), .ZN(n7297) );
  OAI22_X1 U9090 ( .A1(n8723), .A2(n7294), .B1(n7293), .B2(n8642), .ZN(n7295)
         );
  AOI21_X1 U9091 ( .B1(n10055), .B2(n8762), .A(n7295), .ZN(n7296) );
  OAI211_X1 U9092 ( .C1(n10052), .C2(n8586), .A(n7297), .B(n7296), .ZN(
        P2_U3224) );
  OAI21_X1 U9093 ( .B1(n7299), .B2(n8052), .A(n7298), .ZN(n9946) );
  OAI211_X1 U9094 ( .C1(n7301), .C2(n9943), .A(n9917), .B(n7300), .ZN(n9942)
         );
  AOI22_X1 U9095 ( .A1(n9925), .A2(n7303), .B1(n9927), .B2(n7302), .ZN(n7304)
         );
  OAI21_X1 U9096 ( .B1(n9931), .B2(n9942), .A(n7304), .ZN(n7309) );
  XNOR2_X1 U9097 ( .A(n7305), .B(n8052), .ZN(n7307) );
  OAI21_X1 U9098 ( .B1(n7307), .B2(n9469), .A(n7306), .ZN(n9944) );
  MUX2_X1 U9099 ( .A(n9944), .B(P1_REG2_REG_4__SCAN_IN), .S(n9938), .Z(n7308)
         );
  AOI211_X1 U9100 ( .C1(n9935), .C2(n9946), .A(n7309), .B(n7308), .ZN(n7310)
         );
  INV_X1 U9101 ( .A(n7310), .ZN(P1_U3289) );
  AOI21_X1 U9102 ( .B1(n4367), .B2(n7312), .A(n7311), .ZN(n7329) );
  OAI21_X1 U9103 ( .B1(n7315), .B2(n7314), .A(n7313), .ZN(n7327) );
  INV_X1 U9104 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7320) );
  NAND2_X1 U9105 ( .A1(n8553), .A2(n7316), .ZN(n7319) );
  INV_X1 U9106 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7317) );
  NOR2_X1 U9107 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7317), .ZN(n7366) );
  INV_X1 U9108 ( .A(n7366), .ZN(n7318) );
  OAI211_X1 U9109 ( .C1(n7320), .C2(n8561), .A(n7319), .B(n7318), .ZN(n7326)
         );
  AOI21_X1 U9110 ( .B1(n7323), .B2(n7322), .A(n7321), .ZN(n7324) );
  NOR2_X1 U9111 ( .A1(n7324), .A2(n8565), .ZN(n7325) );
  AOI211_X1 U9112 ( .C1(n9981), .C2(n7327), .A(n7326), .B(n7325), .ZN(n7328)
         );
  OAI21_X1 U9113 ( .B1(n7329), .B2(n8559), .A(n7328), .ZN(P2_U3192) );
  INV_X1 U9114 ( .A(n7330), .ZN(n7343) );
  OAI222_X1 U9115 ( .A1(n7742), .A2(n7343), .B1(n8049), .B2(P1_U3086), .C1(
        n7331), .C2(n8303), .ZN(P1_U3334) );
  AOI211_X1 U9116 ( .C1(n7334), .C2(n9958), .A(n7333), .B(n7332), .ZN(n7341)
         );
  INV_X1 U9117 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7335) );
  OAI22_X1 U9118 ( .A1(n9627), .A2(n7181), .B1(n9978), .B2(n7335), .ZN(n7336)
         );
  INV_X1 U9119 ( .A(n7336), .ZN(n7337) );
  OAI21_X1 U9120 ( .B1(n7341), .B2(n9979), .A(n7337), .ZN(P1_U3530) );
  INV_X1 U9121 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7338) );
  OAI22_X1 U9122 ( .A1(n9685), .A2(n7181), .B1(n9961), .B2(n7338), .ZN(n7339)
         );
  INV_X1 U9123 ( .A(n7339), .ZN(n7340) );
  OAI21_X1 U9124 ( .B1(n7341), .B2(n6560), .A(n7340), .ZN(P1_U3477) );
  OAI222_X1 U9125 ( .A1(n7821), .A2(P2_U3151), .B1(n7666), .B2(n7343), .C1(
        n7342), .C2(n7734), .ZN(P2_U3274) );
  AOI21_X1 U9126 ( .B1(n7345), .B2(n10103), .A(n7344), .ZN(n7358) );
  OAI21_X1 U9127 ( .B1(n7348), .B2(n7347), .A(n7346), .ZN(n7356) );
  INV_X1 U9128 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U9129 ( .A1(n8553), .A2(n7349), .ZN(n7354) );
  OAI21_X1 U9130 ( .B1(n7351), .B2(P2_REG2_REG_11__SCAN_IN), .A(n7350), .ZN(
        n7352) );
  INV_X1 U9131 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8859) );
  NOR2_X1 U9132 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8859), .ZN(n7528) );
  AOI21_X1 U9133 ( .B1(n9990), .B2(n7352), .A(n7528), .ZN(n7353) );
  OAI211_X1 U9134 ( .C1(n8922), .C2(n8561), .A(n7354), .B(n7353), .ZN(n7355)
         );
  AOI21_X1 U9135 ( .B1(n9981), .B2(n7356), .A(n7355), .ZN(n7357) );
  OAI21_X1 U9136 ( .B1(n7358), .B2(n8559), .A(n7357), .ZN(P2_U3193) );
  INV_X1 U9137 ( .A(n10061), .ZN(n7371) );
  INV_X1 U9138 ( .A(n7359), .ZN(n7360) );
  NAND2_X1 U9139 ( .A1(n7360), .A2(n8447), .ZN(n7361) );
  XNOR2_X1 U9140 ( .A(n7432), .B(n7531), .ZN(n7364) );
  XNOR2_X1 U9141 ( .A(n10061), .B(n6714), .ZN(n7363) );
  NAND2_X1 U9142 ( .A1(n7364), .A2(n7363), .ZN(n7435) );
  OAI21_X1 U9143 ( .B1(n7364), .B2(n7363), .A(n7435), .ZN(n7365) );
  NAND2_X1 U9144 ( .A1(n7365), .A2(n9742), .ZN(n7370) );
  AOI21_X1 U9145 ( .B1(n8410), .B2(n8445), .A(n7366), .ZN(n7367) );
  OAI21_X1 U9146 ( .B1(n7374), .B2(n8412), .A(n7367), .ZN(n7368) );
  AOI21_X1 U9147 ( .B1(n7378), .B2(n8434), .A(n7368), .ZN(n7369) );
  OAI211_X1 U9148 ( .C1(n7371), .C2(n8438), .A(n7370), .B(n7369), .ZN(P2_U3157) );
  XNOR2_X1 U9149 ( .A(n10061), .B(n7531), .ZN(n7779) );
  NAND2_X1 U9150 ( .A1(n7285), .A2(n7859), .ZN(n7372) );
  XOR2_X1 U9151 ( .A(n7779), .B(n7372), .Z(n10058) );
  XOR2_X1 U9152 ( .A(n7373), .B(n7779), .Z(n7376) );
  OAI22_X1 U9153 ( .A1(n7374), .A2(n8753), .B1(n7489), .B2(n8754), .ZN(n7375)
         );
  AOI21_X1 U9154 ( .B1(n7376), .B2(n8752), .A(n7375), .ZN(n7377) );
  OAI21_X1 U9155 ( .B1(n10058), .B2(n7610), .A(n7377), .ZN(n10059) );
  NAND2_X1 U9156 ( .A1(n10059), .A2(n8715), .ZN(n7383) );
  INV_X1 U9157 ( .A(n7378), .ZN(n7379) );
  OAI22_X1 U9158 ( .A1(n8723), .A2(n7380), .B1(n7379), .B2(n8642), .ZN(n7381)
         );
  AOI21_X1 U9159 ( .B1(n10061), .B2(n8762), .A(n7381), .ZN(n7382) );
  OAI211_X1 U9160 ( .C1(n10058), .C2(n8586), .A(n7383), .B(n7382), .ZN(
        P2_U3223) );
  INV_X1 U9161 ( .A(n7384), .ZN(n7386) );
  OAI222_X1 U9162 ( .A1(P2_U3151), .A2(n7820), .B1(n7666), .B2(n7386), .C1(
        n7385), .C2(n9030), .ZN(P2_U3273) );
  OAI222_X1 U9163 ( .A1(n8303), .A2(n7387), .B1(n7742), .B2(n7386), .C1(
        P1_U3086), .C2(n5698), .ZN(P1_U3333) );
  INV_X1 U9164 ( .A(n7388), .ZN(n7391) );
  AOI21_X1 U9165 ( .B1(n7389), .B2(n7771), .A(n10004), .ZN(n7390) );
  OAI21_X1 U9166 ( .B1(n7392), .B2(n7391), .A(n7390), .ZN(n7394) );
  AOI22_X1 U9167 ( .A1(n8737), .A2(n8444), .B1(n8446), .B2(n8739), .ZN(n7393)
         );
  NAND2_X1 U9168 ( .A1(n7394), .A2(n7393), .ZN(n10067) );
  AOI21_X1 U9169 ( .B1(n8761), .B2(n7527), .A(n10067), .ZN(n7398) );
  XNOR2_X1 U9170 ( .A(n7395), .B(n7771), .ZN(n10064) );
  INV_X1 U9171 ( .A(n7526), .ZN(n7876) );
  OAI22_X1 U9172 ( .A1(n7876), .A2(n8575), .B1(n4738), .B2(n8715), .ZN(n7396)
         );
  AOI21_X1 U9173 ( .B1(n10064), .B2(n7564), .A(n7396), .ZN(n7397) );
  OAI21_X1 U9174 ( .B1(n7398), .B2(n7496), .A(n7397), .ZN(P2_U3222) );
  INV_X1 U9175 ( .A(n7399), .ZN(n7403) );
  NOR3_X1 U9176 ( .A1(n4349), .A2(n7401), .A3(n7400), .ZN(n7402) );
  OAI21_X1 U9177 ( .B1(n7403), .B2(n7402), .A(n9158), .ZN(n7408) );
  NAND2_X1 U9178 ( .A1(n9176), .A2(n9758), .ZN(n7405) );
  NAND2_X1 U9179 ( .A1(n9177), .A2(n9761), .ZN(n7404) );
  AND2_X1 U9180 ( .A1(n7405), .A2(n7404), .ZN(n7477) );
  NAND2_X1 U9181 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9820) );
  OAI21_X1 U9182 ( .B1(n9787), .B2(n7477), .A(n9820), .ZN(n7406) );
  AOI21_X1 U9183 ( .B1(n9140), .B2(n7481), .A(n7406), .ZN(n7407) );
  OAI211_X1 U9184 ( .C1(n7519), .C2(n9143), .A(n7408), .B(n7407), .ZN(P1_U3236) );
  AOI21_X1 U9185 ( .B1(n7411), .B2(n7410), .A(n7409), .ZN(n7425) );
  OAI21_X1 U9186 ( .B1(n7414), .B2(n7413), .A(n7412), .ZN(n7423) );
  AOI21_X1 U9187 ( .B1(n7417), .B2(n7416), .A(n7415), .ZN(n7421) );
  NAND2_X1 U9188 ( .A1(n8553), .A2(n7418), .ZN(n7420) );
  AND2_X1 U9189 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7440) );
  AOI21_X1 U9190 ( .B1(n9991), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7440), .ZN(
        n7419) );
  OAI211_X1 U9191 ( .C1(n7421), .C2(n8565), .A(n7420), .B(n7419), .ZN(n7422)
         );
  AOI21_X1 U9192 ( .B1(n9981), .B2(n7423), .A(n7422), .ZN(n7424) );
  OAI21_X1 U9193 ( .B1(n7425), .B2(n8559), .A(n7424), .ZN(P2_U3194) );
  NAND2_X1 U9194 ( .A1(n7429), .A2(n7426), .ZN(n7427) );
  OAI211_X1 U9195 ( .C1(n5537), .C2(n8303), .A(n7427), .B(n8238), .ZN(P1_U3332) );
  NAND2_X1 U9196 ( .A1(n7429), .A2(n7428), .ZN(n7430) );
  OAI211_X1 U9197 ( .C1(n7431), .C2(n9030), .A(n7430), .B(n7984), .ZN(P2_U3272) );
  INV_X1 U9198 ( .A(n7432), .ZN(n7433) );
  NAND2_X1 U9199 ( .A1(n7433), .A2(n7531), .ZN(n7434) );
  XNOR2_X1 U9200 ( .A(n7526), .B(n6714), .ZN(n7437) );
  XNOR2_X1 U9201 ( .A(n7437), .B(n7489), .ZN(n7535) );
  INV_X1 U9202 ( .A(n7535), .ZN(n7436) );
  INV_X1 U9203 ( .A(n7437), .ZN(n7438) );
  NAND2_X1 U9204 ( .A1(n7438), .A2(n8445), .ZN(n7439) );
  XNOR2_X1 U9205 ( .A(n10071), .B(n8293), .ZN(n7546) );
  XNOR2_X1 U9206 ( .A(n7546), .B(n8444), .ZN(n7544) );
  XNOR2_X1 U9207 ( .A(n7545), .B(n7544), .ZN(n7445) );
  NAND2_X1 U9208 ( .A1(n8434), .A2(n7491), .ZN(n7442) );
  AOI21_X1 U9209 ( .B1(n8410), .B2(n9736), .A(n7440), .ZN(n7441) );
  OAI211_X1 U9210 ( .C1(n7489), .C2(n8412), .A(n7442), .B(n7441), .ZN(n7443)
         );
  AOI21_X1 U9211 ( .B1(n10071), .B2(n8369), .A(n7443), .ZN(n7444) );
  OAI21_X1 U9212 ( .B1(n7445), .B2(n8391), .A(n7444), .ZN(P2_U3164) );
  NOR2_X1 U9213 ( .A1(n9913), .A2(n7449), .ZN(n8001) );
  INV_X1 U9214 ( .A(n8001), .ZN(n7448) );
  NAND2_X1 U9215 ( .A1(n9913), .A2(n7449), .ZN(n8152) );
  NAND2_X1 U9216 ( .A1(n7448), .A2(n8152), .ZN(n9914) );
  OR2_X1 U9217 ( .A1(n7523), .A2(n7450), .ZN(n7581) );
  NAND2_X1 U9218 ( .A1(n7523), .A2(n7450), .ZN(n8157) );
  XNOR2_X1 U9219 ( .A(n9779), .B(n9176), .ZN(n8062) );
  XNOR2_X1 U9220 ( .A(n7591), .B(n8062), .ZN(n7500) );
  INV_X1 U9221 ( .A(n7500), .ZN(n7471) );
  NAND2_X1 U9222 ( .A1(n8019), .A2(n7452), .ZN(n7457) );
  AND2_X1 U9223 ( .A1(n8132), .A2(n7453), .ZN(n8128) );
  NAND2_X1 U9224 ( .A1(n8154), .A2(n8128), .ZN(n8059) );
  INV_X1 U9225 ( .A(n8124), .ZN(n7454) );
  OR2_X1 U9226 ( .A1(n8059), .A2(n7454), .ZN(n7455) );
  NAND2_X1 U9227 ( .A1(n7456), .A2(n7455), .ZN(n8016) );
  NAND2_X1 U9228 ( .A1(n7457), .A2(n8016), .ZN(n9905) );
  OR2_X1 U9229 ( .A1(n9905), .A2(n9914), .ZN(n9906) );
  NAND2_X1 U9230 ( .A1(n8157), .A2(n8152), .ZN(n8022) );
  INV_X1 U9231 ( .A(n8022), .ZN(n7458) );
  NAND2_X1 U9232 ( .A1(n7582), .A2(n7581), .ZN(n7460) );
  INV_X1 U9233 ( .A(n8062), .ZN(n7459) );
  XNOR2_X1 U9234 ( .A(n7460), .B(n7459), .ZN(n7461) );
  NAND2_X1 U9235 ( .A1(n7461), .A2(n9910), .ZN(n7464) );
  NAND2_X1 U9236 ( .A1(n9175), .A2(n9758), .ZN(n7463) );
  NAND2_X1 U9237 ( .A1(n9759), .A2(n9761), .ZN(n7462) );
  AND2_X1 U9238 ( .A1(n7463), .A2(n7462), .ZN(n9771) );
  NAND2_X1 U9239 ( .A1(n7464), .A2(n9771), .ZN(n7498) );
  INV_X1 U9240 ( .A(n9779), .ZN(n7589) );
  INV_X1 U9241 ( .A(n7480), .ZN(n7465) );
  AOI211_X1 U9242 ( .C1(n9779), .C2(n7465), .A(n9527), .B(n4366), .ZN(n7499)
         );
  NAND2_X1 U9243 ( .A1(n7499), .A2(n9921), .ZN(n7468) );
  AOI22_X1 U9244 ( .A1(n9928), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7466), .B2(
        n9927), .ZN(n7467) );
  OAI211_X1 U9245 ( .C1(n7589), .C2(n9530), .A(n7468), .B(n7467), .ZN(n7469)
         );
  AOI21_X1 U9246 ( .B1(n9534), .B2(n7498), .A(n7469), .ZN(n7470) );
  OAI21_X1 U9247 ( .B1(n7471), .B2(n9518), .A(n7470), .ZN(P1_U3281) );
  AOI21_X1 U9248 ( .B1(n7473), .B2(n8064), .A(n7472), .ZN(n7515) );
  NAND2_X1 U9249 ( .A1(n9906), .A2(n8152), .ZN(n7474) );
  XNOR2_X1 U9250 ( .A(n7474), .B(n8064), .ZN(n7475) );
  NAND2_X1 U9251 ( .A1(n7475), .A2(n9910), .ZN(n7476) );
  OAI211_X1 U9252 ( .C1(n7515), .C2(n7478), .A(n7477), .B(n7476), .ZN(n7517)
         );
  NAND2_X1 U9253 ( .A1(n7517), .A2(n9534), .ZN(n7486) );
  OAI21_X1 U9254 ( .B1(n9916), .B2(n7519), .A(n9917), .ZN(n7479) );
  OR2_X1 U9255 ( .A1(n7480), .A2(n7479), .ZN(n7513) );
  INV_X1 U9256 ( .A(n7513), .ZN(n7484) );
  AOI22_X1 U9257 ( .A1(n9928), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7481), .B2(
        n9927), .ZN(n7482) );
  OAI21_X1 U9258 ( .B1(n7519), .B2(n9530), .A(n7482), .ZN(n7483) );
  AOI21_X1 U9259 ( .B1(n7484), .B2(n9921), .A(n7483), .ZN(n7485) );
  OAI211_X1 U9260 ( .C1(n7515), .C2(n7487), .A(n7486), .B(n7485), .ZN(P1_U3282) );
  NOR2_X1 U9261 ( .A1(n7575), .A2(n8754), .ZN(n10075) );
  XNOR2_X1 U9262 ( .A(n7488), .B(n7888), .ZN(n7490) );
  OAI22_X1 U9263 ( .A1(n7490), .A2(n10004), .B1(n7489), .B2(n8753), .ZN(n10077) );
  AOI211_X1 U9264 ( .C1(n8761), .C2(n7491), .A(n10075), .B(n10077), .ZN(n7497)
         );
  AOI22_X1 U9265 ( .A1(n10071), .A2(n8762), .B1(P2_REG2_REG_12__SCAN_IN), .B2(
        n7496), .ZN(n7495) );
  NAND2_X1 U9266 ( .A1(n7493), .A2(n7888), .ZN(n10069) );
  NAND3_X1 U9267 ( .A1(n7492), .A2(n10069), .A3(n7564), .ZN(n7494) );
  OAI211_X1 U9268 ( .C1(n7497), .C2(n7496), .A(n7495), .B(n7494), .ZN(P2_U3221) );
  AOI211_X1 U9269 ( .C1(n7500), .C2(n9958), .A(n7499), .B(n7498), .ZN(n7505)
         );
  INV_X1 U9270 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7501) );
  OAI22_X1 U9271 ( .A1(n7589), .A2(n9685), .B1(n9971), .B2(n7501), .ZN(n7502)
         );
  INV_X1 U9272 ( .A(n7502), .ZN(n7503) );
  OAI21_X1 U9273 ( .B1(n7505), .B2(n6560), .A(n7503), .ZN(P1_U3489) );
  AOI22_X1 U9274 ( .A1(n9779), .A2(n7522), .B1(n9979), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7504) );
  OAI21_X1 U9275 ( .B1(n7505), .B2(n9979), .A(n7504), .ZN(P1_U3534) );
  AOI21_X1 U9276 ( .B1(n7508), .B2(n7507), .A(n7506), .ZN(n7512) );
  AOI22_X1 U9277 ( .A1(n9761), .A2(n9176), .B1(n9174), .B2(n9758), .ZN(n7583)
         );
  NAND2_X1 U9278 ( .A1(n9140), .A2(n7585), .ZN(n7509) );
  NAND2_X1 U9279 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9832) );
  OAI211_X1 U9280 ( .C1(n7583), .C2(n9787), .A(n7509), .B(n9832), .ZN(n7510)
         );
  AOI21_X1 U9281 ( .B1(n8110), .B2(n4282), .A(n7510), .ZN(n7511) );
  OAI21_X1 U9282 ( .B1(n7512), .B2(n9792), .A(n7511), .ZN(P1_U3234) );
  OAI21_X1 U9283 ( .B1(n7515), .B2(n7514), .A(n7513), .ZN(n7516) );
  NOR2_X1 U9284 ( .A1(n7517), .A2(n7516), .ZN(n7525) );
  INV_X1 U9285 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7518) );
  OAI22_X1 U9286 ( .A1(n7519), .A2(n9685), .B1(n9971), .B2(n7518), .ZN(n7520)
         );
  INV_X1 U9287 ( .A(n7520), .ZN(n7521) );
  OAI21_X1 U9288 ( .B1(n7525), .B2(n6560), .A(n7521), .ZN(P1_U3486) );
  AOI22_X1 U9289 ( .A1(n7523), .A2(n7522), .B1(n9979), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7524) );
  OAI21_X1 U9290 ( .B1(n7525), .B2(n9979), .A(n7524), .ZN(P1_U3533) );
  AND2_X1 U9291 ( .A1(n7526), .A2(n10062), .ZN(n10066) );
  NAND2_X1 U9292 ( .A1(n8434), .A2(n7527), .ZN(n7530) );
  AOI21_X1 U9293 ( .B1(n8410), .B2(n8444), .A(n7528), .ZN(n7529) );
  OAI211_X1 U9294 ( .C1(n7531), .C2(n8412), .A(n7530), .B(n7529), .ZN(n7537)
         );
  INV_X1 U9295 ( .A(n7533), .ZN(n7534) );
  AOI211_X1 U9296 ( .C1(n7535), .C2(n7532), .A(n8391), .B(n7534), .ZN(n7536)
         );
  AOI211_X1 U9297 ( .C1(n10066), .C2(n9740), .A(n7537), .B(n7536), .ZN(n7538)
         );
  INV_X1 U9298 ( .A(n7538), .ZN(P2_U3176) );
  INV_X1 U9299 ( .A(n7539), .ZN(n7665) );
  OAI222_X1 U9300 ( .A1(n7742), .A2(n7665), .B1(P1_U3086), .B2(n7541), .C1(
        n7540), .C2(n8303), .ZN(P1_U3331) );
  INV_X2 U9301 ( .A(n6715), .ZN(n8293) );
  XNOR2_X1 U9302 ( .A(n7556), .B(n8293), .ZN(n7543) );
  INV_X1 U9303 ( .A(n7543), .ZN(n7542) );
  NAND2_X1 U9304 ( .A1(n7542), .A2(n9736), .ZN(n8246) );
  NAND2_X1 U9305 ( .A1(n7543), .A2(n7575), .ZN(n8244) );
  NAND2_X1 U9306 ( .A1(n8246), .A2(n8244), .ZN(n7549) );
  INV_X1 U9307 ( .A(n7546), .ZN(n7547) );
  NAND2_X1 U9308 ( .A1(n7547), .A2(n8444), .ZN(n7548) );
  XOR2_X1 U9309 ( .A(n7549), .B(n8245), .Z(n7555) );
  NAND2_X1 U9310 ( .A1(n8434), .A2(n7561), .ZN(n7552) );
  NOR2_X1 U9311 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7550), .ZN(n8462) );
  AOI21_X1 U9312 ( .B1(n8410), .B2(n8443), .A(n8462), .ZN(n7551) );
  OAI211_X1 U9313 ( .C1(n7559), .C2(n8412), .A(n7552), .B(n7551), .ZN(n7553)
         );
  AOI21_X1 U9314 ( .B1(n7556), .B2(n8369), .A(n7553), .ZN(n7554) );
  OAI21_X1 U9315 ( .B1(n7555), .B2(n8391), .A(n7554), .ZN(P2_U3174) );
  INV_X1 U9316 ( .A(n7556), .ZN(n9748) );
  NOR2_X1 U9317 ( .A1(n9748), .A2(n8644), .ZN(n7560) );
  XNOR2_X1 U9318 ( .A(n7557), .B(n7562), .ZN(n7558) );
  OAI222_X1 U9319 ( .A1(n8754), .A2(n8249), .B1(n8753), .B2(n7559), .C1(n10004), .C2(n7558), .ZN(n9749) );
  AOI211_X1 U9320 ( .C1(n8761), .C2(n7561), .A(n7560), .B(n9749), .ZN(n7566)
         );
  OAI21_X1 U9321 ( .B1(n4305), .B2(n6083), .A(n7563), .ZN(n9751) );
  AOI22_X1 U9322 ( .A1(n9751), .A2(n7564), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7496), .ZN(n7565) );
  OAI21_X1 U9323 ( .B1(n7566), .B2(n7496), .A(n7565), .ZN(P2_U3220) );
  INV_X1 U9324 ( .A(n7567), .ZN(n7730) );
  INV_X1 U9325 ( .A(n7568), .ZN(n7570) );
  OAI222_X1 U9326 ( .A1(n7742), .A2(n7730), .B1(P1_U3086), .B2(n7570), .C1(
        n7569), .C2(n8303), .ZN(P1_U3330) );
  INV_X1 U9327 ( .A(n7892), .ZN(n7572) );
  XNOR2_X1 U9328 ( .A(n7571), .B(n7572), .ZN(n7618) );
  XOR2_X1 U9329 ( .A(n7573), .B(n7892), .Z(n7574) );
  OAI222_X1 U9330 ( .A1(n8754), .A2(n9733), .B1(n8753), .B2(n7575), .C1(n7574), 
        .C2(n10004), .ZN(n7612) );
  INV_X1 U9331 ( .A(n8248), .ZN(n7611) );
  NOR2_X1 U9332 ( .A1(n7611), .A2(n8644), .ZN(n7576) );
  OAI21_X1 U9333 ( .B1(n7612), .B2(n7576), .A(n8723), .ZN(n7579) );
  AOI22_X1 U9334 ( .A1(n7496), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8761), .B2(
        n7577), .ZN(n7578) );
  OAI211_X1 U9335 ( .C1(n7618), .C2(n8765), .A(n7579), .B(n7578), .ZN(P2_U3219) );
  OR2_X1 U9336 ( .A1(n8110), .A2(n7580), .ZN(n8148) );
  NAND2_X1 U9337 ( .A1(n8110), .A2(n7580), .ZN(n8138) );
  OR2_X1 U9338 ( .A1(n9779), .A2(n7588), .ZN(n8156) );
  NAND2_X1 U9339 ( .A1(n8156), .A2(n7581), .ZN(n8002) );
  INV_X1 U9340 ( .A(n8002), .ZN(n8023) );
  AND2_X1 U9341 ( .A1(n9779), .A2(n7588), .ZN(n8021) );
  INV_X1 U9342 ( .A(n8021), .ZN(n8158) );
  XOR2_X1 U9343 ( .A(n8065), .B(n7597), .Z(n7584) );
  OAI21_X1 U9344 ( .B1(n7584), .B2(n9469), .A(n7583), .ZN(n9968) );
  OAI211_X1 U9345 ( .C1(n4366), .C2(n9966), .A(n9917), .B(n7604), .ZN(n9964)
         );
  AOI22_X1 U9346 ( .A1(n9938), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7585), .B2(
        n9927), .ZN(n7587) );
  NAND2_X1 U9347 ( .A1(n8110), .A2(n9925), .ZN(n7586) );
  OAI211_X1 U9348 ( .C1(n9964), .C2(n9931), .A(n7587), .B(n7586), .ZN(n7594)
         );
  NOR2_X1 U9349 ( .A1(n7589), .A2(n7588), .ZN(n7590) );
  AND2_X1 U9350 ( .A1(n7592), .A2(n8065), .ZN(n9963) );
  NOR3_X1 U9351 ( .A1(n7596), .A2(n9963), .A3(n9518), .ZN(n7593) );
  AOI211_X1 U9352 ( .C1(n9534), .C2(n9968), .A(n7594), .B(n7593), .ZN(n7595)
         );
  INV_X1 U9353 ( .A(n7595), .ZN(P1_U3280) );
  OR2_X1 U9354 ( .A1(n8106), .A2(n8111), .ZN(n8149) );
  NAND2_X1 U9355 ( .A1(n8106), .A2(n8111), .ZN(n8139) );
  NAND2_X1 U9356 ( .A1(n8149), .A2(n8139), .ZN(n8067) );
  XNOR2_X1 U9357 ( .A(n7636), .B(n8067), .ZN(n9624) );
  INV_X1 U9358 ( .A(n9624), .ZN(n7609) );
  NAND2_X1 U9359 ( .A1(n7598), .A2(n8138), .ZN(n7599) );
  NAND2_X1 U9360 ( .A1(n7599), .A2(n8067), .ZN(n7600) );
  NAND3_X1 U9361 ( .A1(n7637), .A2(n9910), .A3(n7600), .ZN(n7603) );
  NAND2_X1 U9362 ( .A1(n9275), .A2(n9758), .ZN(n7602) );
  NAND2_X1 U9363 ( .A1(n9175), .A2(n9761), .ZN(n7601) );
  AND2_X1 U9364 ( .A1(n7602), .A2(n7601), .ZN(n9041) );
  NAND2_X1 U9365 ( .A1(n7603), .A2(n9041), .ZN(n9622) );
  AOI211_X1 U9366 ( .C1(n8106), .C2(n7604), .A(n9527), .B(n7640), .ZN(n9623)
         );
  NAND2_X1 U9367 ( .A1(n9623), .A2(n9921), .ZN(n7606) );
  AOI22_X1 U9368 ( .A1(n9928), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9044), .B2(
        n9927), .ZN(n7605) );
  OAI211_X1 U9369 ( .C1(n9686), .C2(n9530), .A(n7606), .B(n7605), .ZN(n7607)
         );
  AOI21_X1 U9370 ( .B1(n9534), .B2(n9622), .A(n7607), .ZN(n7608) );
  OAI21_X1 U9371 ( .B1(n7609), .B2(n9518), .A(n7608), .ZN(P1_U3279) );
  NAND2_X1 U9372 ( .A1(n7610), .A2(n10057), .ZN(n10070) );
  INV_X1 U9373 ( .A(n10070), .ZN(n10028) );
  OR2_X1 U9374 ( .A1(n10078), .A2(n10028), .ZN(n9025) );
  INV_X1 U9375 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7613) );
  NOR2_X1 U9376 ( .A1(n7611), .A2(n10072), .ZN(n9741) );
  NOR2_X1 U9377 ( .A1(n7612), .A2(n9741), .ZN(n7615) );
  MUX2_X1 U9378 ( .A(n7613), .B(n7615), .S(n10080), .Z(n7614) );
  OAI21_X1 U9379 ( .B1(n7618), .B2(n9025), .A(n7614), .ZN(P2_U3432) );
  NAND2_X1 U9380 ( .A1(n10107), .A2(n10070), .ZN(n8811) );
  INV_X1 U9381 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7616) );
  MUX2_X1 U9382 ( .A(n7616), .B(n7615), .S(n10107), .Z(n7617) );
  OAI21_X1 U9383 ( .B1(n8811), .B2(n7618), .A(n7617), .ZN(P2_U3473) );
  INV_X1 U9384 ( .A(n7619), .ZN(n7623) );
  OAI222_X1 U9385 ( .A1(n7742), .A2(n7623), .B1(P1_U3086), .B2(n7621), .C1(
        n7620), .C2(n8303), .ZN(P1_U3329) );
  OAI222_X1 U9386 ( .A1(n7624), .A2(P2_U3151), .B1(n7666), .B2(n7623), .C1(
        n7622), .C2(n9030), .ZN(P2_U3269) );
  OAI21_X1 U9387 ( .B1(n7626), .B2(n7896), .A(n7625), .ZN(n7650) );
  NAND2_X1 U9388 ( .A1(n7627), .A2(n7896), .ZN(n7628) );
  NAND3_X1 U9389 ( .A1(n8750), .A2(n8752), .A3(n7628), .ZN(n7630) );
  AOI22_X1 U9390 ( .A1(n8740), .A2(n8737), .B1(n8739), .B2(n8443), .ZN(n7629)
         );
  NAND2_X1 U9391 ( .A1(n7630), .A2(n7629), .ZN(n7649) );
  INV_X1 U9392 ( .A(n7649), .ZN(n7631) );
  MUX2_X1 U9393 ( .A(n7631), .B(n8917), .S(n7496), .Z(n7633) );
  AOI22_X1 U9394 ( .A1(n8253), .A2(n8762), .B1(n8761), .B2(n8435), .ZN(n7632)
         );
  OAI211_X1 U9395 ( .C1(n7650), .C2(n8765), .A(n7633), .B(n7632), .ZN(P2_U3218) );
  INV_X1 U9396 ( .A(n7634), .ZN(n7654) );
  OAI222_X1 U9397 ( .A1(P2_U3151), .A2(n7978), .B1(n9035), .B2(n7654), .C1(
        n7635), .C2(n9030), .ZN(P2_U3268) );
  XNOR2_X1 U9398 ( .A(n9274), .B(n9275), .ZN(n8068) );
  XNOR2_X1 U9399 ( .A(n9278), .B(n8068), .ZN(n9620) );
  INV_X1 U9400 ( .A(n9620), .ZN(n7646) );
  INV_X1 U9401 ( .A(n8068), .ZN(n8080) );
  XNOR2_X1 U9402 ( .A(n8080), .B(n8081), .ZN(n7638) );
  NAND2_X1 U9403 ( .A1(n7638), .A2(n9910), .ZN(n7639) );
  AOI22_X1 U9404 ( .A1(n9174), .A2(n9761), .B1(n9758), .B2(n9281), .ZN(n7673)
         );
  NAND2_X1 U9405 ( .A1(n7639), .A2(n7673), .ZN(n9618) );
  INV_X1 U9406 ( .A(n9528), .ZN(n7641) );
  AOI211_X1 U9407 ( .C1(n9274), .C2(n4466), .A(n9527), .B(n7641), .ZN(n9619)
         );
  NAND2_X1 U9408 ( .A1(n9619), .A2(n9921), .ZN(n7643) );
  AOI22_X1 U9409 ( .A1(n9928), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7671), .B2(
        n9927), .ZN(n7642) );
  OAI211_X1 U9410 ( .C1(n9276), .C2(n9530), .A(n7643), .B(n7642), .ZN(n7644)
         );
  AOI21_X1 U9411 ( .B1(n9534), .B2(n9618), .A(n7644), .ZN(n7645) );
  OAI21_X1 U9412 ( .B1(n7646), .B2(n9518), .A(n7645), .ZN(P1_U3278) );
  MUX2_X1 U9413 ( .A(n7649), .B(P2_REG0_REG_15__SCAN_IN), .S(n10078), .Z(n7648) );
  INV_X1 U9414 ( .A(n8253), .ZN(n8439) );
  OAI22_X1 U9415 ( .A1(n7650), .A2(n9025), .B1(n8439), .B2(n9023), .ZN(n7647)
         );
  OR2_X1 U9416 ( .A1(n7648), .A2(n7647), .ZN(P2_U3435) );
  MUX2_X1 U9417 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n7649), .S(n10107), .Z(n7652) );
  OAI22_X1 U9418 ( .A1(n7650), .A2(n8811), .B1(n8439), .B2(n8810), .ZN(n7651)
         );
  OR2_X1 U9419 ( .A1(n7652), .A2(n7651), .ZN(P2_U3474) );
  OAI222_X1 U9420 ( .A1(n7742), .A2(n7654), .B1(P1_U3086), .B2(n6469), .C1(
        n7653), .C2(n8303), .ZN(P1_U3328) );
  INV_X1 U9421 ( .A(n7655), .ZN(n7733) );
  OAI222_X1 U9422 ( .A1(P2_U3151), .A2(n7657), .B1(n9035), .B2(n7733), .C1(
        n7656), .C2(n9030), .ZN(P2_U3267) );
  INV_X1 U9423 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7719) );
  INV_X1 U9424 ( .A(n7658), .ZN(n7659) );
  MUX2_X1 U9425 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4471), .Z(n7750) );
  XNOR2_X1 U9426 ( .A(n7750), .B(SI_30_), .ZN(n7751) );
  INV_X1 U9427 ( .A(n7743), .ZN(n7738) );
  OAI222_X1 U9428 ( .A1(n8303), .A2(n7719), .B1(n7742), .B2(n7738), .C1(
        P1_U3086), .C2(n7663), .ZN(P1_U3325) );
  OAI222_X1 U9429 ( .A1(n7667), .A2(P2_U3151), .B1(n7666), .B2(n7665), .C1(
        n7664), .C2(n7734), .ZN(P2_U3271) );
  AOI21_X1 U9430 ( .B1(n7670), .B2(n7669), .A(n7668), .ZN(n7676) );
  NAND2_X1 U9431 ( .A1(n9140), .A2(n7671), .ZN(n7672) );
  NAND2_X1 U9432 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9861) );
  OAI211_X1 U9433 ( .C1(n7673), .C2(n9787), .A(n7672), .B(n9861), .ZN(n7674)
         );
  AOI21_X1 U9434 ( .B1(n9274), .B2(n4282), .A(n7674), .ZN(n7675) );
  OAI21_X1 U9435 ( .B1(n7676), .B2(n9792), .A(n7675), .ZN(P1_U3241) );
  INV_X1 U9436 ( .A(n9869), .ZN(n9904) );
  NAND2_X1 U9437 ( .A1(n7702), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7683) );
  INV_X1 U9438 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7677) );
  AOI22_X1 U9439 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7678), .B1(n9831), .B2(
        n7677), .ZN(n9828) );
  OAI21_X1 U9440 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7680), .A(n7679), .ZN(
        n9827) );
  NOR2_X1 U9441 ( .A1(n9828), .A2(n9827), .ZN(n9826) );
  AOI21_X1 U9442 ( .B1(n9831), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9826), .ZN(
        n9836) );
  INV_X1 U9443 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7681) );
  AOI22_X1 U9444 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9845), .B1(n7702), .B2(
        n7681), .ZN(n9837) );
  NOR2_X1 U9445 ( .A1(n9836), .A2(n9837), .ZN(n9835) );
  INV_X1 U9446 ( .A(n9835), .ZN(n7682) );
  NAND2_X1 U9447 ( .A1(n7683), .A2(n7682), .ZN(n7685) );
  INV_X1 U9448 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9857) );
  INV_X1 U9449 ( .A(n7686), .ZN(n7684) );
  OAI21_X1 U9450 ( .B1(n9860), .B2(n7685), .A(n7684), .ZN(n9856) );
  NOR2_X1 U9451 ( .A1(n9857), .A2(n9856), .ZN(n9855) );
  NOR2_X1 U9452 ( .A1(n7686), .A2(n9855), .ZN(n9866) );
  AOI22_X1 U9453 ( .A1(n9873), .A2(n9533), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n7693), .ZN(n9865) );
  NOR2_X1 U9454 ( .A1(n9866), .A2(n9865), .ZN(n9864) );
  AOI21_X1 U9455 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9873), .A(n9864), .ZN(
        n9878) );
  INV_X1 U9456 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7687) );
  XNOR2_X1 U9457 ( .A(n9882), .B(n7687), .ZN(n9877) );
  NAND2_X1 U9458 ( .A1(n9878), .A2(n9877), .ZN(n7689) );
  OR2_X1 U9459 ( .A1(n9882), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U9460 ( .A1(n7689), .A2(n7688), .ZN(n9891) );
  NAND2_X1 U9461 ( .A1(n7709), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7691) );
  OR2_X1 U9462 ( .A1(n7709), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7690) );
  NAND2_X1 U9463 ( .A1(n7691), .A2(n7690), .ZN(n9890) );
  NAND2_X1 U9464 ( .A1(n9900), .A2(n7691), .ZN(n7692) );
  INV_X1 U9465 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9476) );
  XNOR2_X1 U9466 ( .A(n7692), .B(n9476), .ZN(n7712) );
  AOI22_X1 U9467 ( .A1(n9873), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9616), .B2(
        n7693), .ZN(n9872) );
  NAND2_X1 U9468 ( .A1(n7702), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7704) );
  NAND2_X1 U9469 ( .A1(n7695), .A2(n7694), .ZN(n7696) );
  INV_X1 U9470 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7698) );
  OR2_X1 U9471 ( .A1(n9831), .A2(n7698), .ZN(n7700) );
  NAND2_X1 U9472 ( .A1(n9831), .A2(n7698), .ZN(n7699) );
  AND2_X1 U9473 ( .A1(n7700), .A2(n7699), .ZN(n9825) );
  AND2_X1 U9474 ( .A1(n9831), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7701) );
  XNOR2_X1 U9475 ( .A(n7702), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9840) );
  INV_X1 U9476 ( .A(n9839), .ZN(n7703) );
  NAND2_X1 U9477 ( .A1(n7704), .A2(n7703), .ZN(n7705) );
  NOR2_X1 U9478 ( .A1(n7705), .A2(n9860), .ZN(n7706) );
  OAI21_X1 U9479 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9873), .A(n9870), .ZN(
        n9880) );
  INV_X1 U9480 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9610) );
  XNOR2_X1 U9481 ( .A(n9882), .B(n9610), .ZN(n9879) );
  AOI22_X1 U9482 ( .A1(n9880), .A2(n9879), .B1(n9610), .B2(n7708), .ZN(n9895)
         );
  INV_X1 U9483 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9605) );
  AND2_X1 U9484 ( .A1(n7709), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7710) );
  AOI21_X1 U9485 ( .B1(n9897), .B2(n9605), .A(n7710), .ZN(n9894) );
  NAND2_X1 U9486 ( .A1(n9895), .A2(n9894), .ZN(n9893) );
  INV_X1 U9487 ( .A(n7710), .ZN(n7711) );
  AOI22_X1 U9488 ( .A1(n7712), .A2(n9884), .B1(n9892), .B2(n7713), .ZN(n7716)
         );
  INV_X1 U9489 ( .A(n7712), .ZN(n7714) );
  MUX2_X1 U9490 ( .A(n7716), .B(n7715), .S(n5437), .Z(n7718) );
  NAND2_X1 U9491 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n7717) );
  OAI211_X1 U9492 ( .C1(n4518), .C2(n9904), .A(n7718), .B(n7717), .ZN(P1_U3262) );
  NAND2_X1 U9493 ( .A1(n7743), .A2(n5346), .ZN(n7721) );
  OR2_X1 U9494 ( .A1(n5127), .A2(n7719), .ZN(n7720) );
  INV_X1 U9495 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7740) );
  OR2_X1 U9496 ( .A1(n5127), .A2(n7740), .ZN(n7722) );
  NAND2_X1 U9497 ( .A1(n9662), .A2(n9473), .ZN(n9457) );
  NOR2_X2 U9498 ( .A1(n9395), .A2(n9381), .ZN(n9380) );
  NAND2_X1 U9499 ( .A1(n9636), .A2(n9320), .ZN(n9254) );
  OAI211_X1 U9500 ( .C1(n9636), .C2(n9320), .A(n9917), .B(n9254), .ZN(n9544)
         );
  NOR2_X1 U9501 ( .A1(n6469), .A2(n7726), .ZN(n7727) );
  NOR2_X1 U9502 ( .A1(n9161), .A2(n7727), .ZN(n9272) );
  AND2_X1 U9503 ( .A1(n8215), .A2(n9272), .ZN(n9539) );
  INV_X1 U9504 ( .A(n9539), .ZN(n9543) );
  NOR2_X1 U9505 ( .A1(n9938), .A2(n9543), .ZN(n9256) );
  NOR2_X1 U9506 ( .A1(n9636), .A2(n9530), .ZN(n7728) );
  AOI211_X1 U9507 ( .C1(n9928), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9256), .B(
        n7728), .ZN(n7729) );
  OAI21_X1 U9508 ( .B1(n9544), .B2(n9931), .A(n7729), .ZN(P1_U3264) );
  OAI222_X1 U9509 ( .A1(n7731), .A2(P2_U3151), .B1(n9035), .B2(n7730), .C1(
        n8905), .C2(n7734), .ZN(P2_U3270) );
  OAI222_X1 U9510 ( .A1(n7742), .A2(n7733), .B1(n4285), .B2(P1_U3086), .C1(
        n7732), .C2(n8303), .ZN(P1_U3327) );
  OAI222_X1 U9511 ( .A1(P2_U3151), .A2(n7736), .B1(n9035), .B2(n7741), .C1(
        n7735), .C2(n7734), .ZN(P2_U3266) );
  INV_X1 U9512 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7744) );
  OAI222_X1 U9513 ( .A1(n7737), .A2(P2_U3151), .B1(n9035), .B2(n7738), .C1(
        n7744), .C2(n9030), .ZN(P2_U3265) );
  OAI222_X1 U9514 ( .A1(n7742), .A2(n7741), .B1(P1_U3086), .B2(n7739), .C1(
        n7740), .C2(n8303), .ZN(P1_U3326) );
  INV_X1 U9515 ( .A(n7790), .ZN(n7748) );
  NAND2_X1 U9516 ( .A1(n7743), .A2(n7755), .ZN(n7746) );
  OR2_X1 U9517 ( .A1(n5991), .A2(n7744), .ZN(n7745) );
  INV_X1 U9518 ( .A(n8440), .ZN(n7766) );
  INV_X1 U9519 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8039) );
  MUX2_X1 U9520 ( .A(n8039), .B(n8894), .S(n4471), .Z(n7752) );
  XNOR2_X1 U9521 ( .A(n7752), .B(SI_31_), .ZN(n7753) );
  NAND2_X1 U9522 ( .A1(n9029), .A2(n7755), .ZN(n7757) );
  OR2_X1 U9523 ( .A1(n5991), .A2(n8894), .ZN(n7756) );
  NAND2_X1 U9524 ( .A1(n6125), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7762) );
  NAND2_X1 U9525 ( .A1(n7758), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7761) );
  NAND2_X1 U9526 ( .A1(n7759), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7760) );
  AND3_X1 U9527 ( .A1(n7762), .A2(n7761), .A3(n7760), .ZN(n7763) );
  NAND2_X1 U9528 ( .A1(n8814), .A2(n7795), .ZN(n7968) );
  NAND2_X1 U9529 ( .A1(n7765), .A2(n7968), .ZN(n7805) );
  INV_X1 U9530 ( .A(n8814), .ZN(n8576) );
  OAI211_X1 U9531 ( .C1(n8576), .C2(n7794), .A(n7767), .B(n7803), .ZN(n7802)
         );
  NOR2_X1 U9532 ( .A1(n8814), .A2(n7795), .ZN(n7969) );
  INV_X1 U9533 ( .A(n7968), .ZN(n7792) );
  INV_X1 U9534 ( .A(n8588), .ZN(n8590) );
  INV_X1 U9535 ( .A(n7769), .ZN(n7932) );
  INV_X1 U9536 ( .A(n7927), .ZN(n7809) );
  INV_X1 U9537 ( .A(n7770), .ZN(n8718) );
  INV_X1 U9538 ( .A(n7771), .ZN(n7782) );
  NAND4_X1 U9539 ( .A1(n7773), .A2(n6259), .A3(n7772), .A4(n10003), .ZN(n7776)
         );
  NOR4_X1 U9540 ( .A1(n7776), .A2(n7775), .A3(n7839), .A4(n7774), .ZN(n7777)
         );
  NAND4_X1 U9541 ( .A1(n6047), .A2(n7778), .A3(n7777), .A4(n4819), .ZN(n7780)
         );
  OR2_X1 U9542 ( .A1(n7780), .A2(n7779), .ZN(n7781) );
  NOR3_X1 U9543 ( .A1(n7888), .A2(n7782), .A3(n7781), .ZN(n7783) );
  NAND4_X1 U9544 ( .A1(n7896), .A2(n7892), .A3(n7783), .A4(n6083), .ZN(n7784)
         );
  NOR3_X1 U9545 ( .A1(n8731), .A2(n7785), .A3(n7784), .ZN(n7786) );
  NAND4_X1 U9546 ( .A1(n8690), .A2(n8707), .A3(n8718), .A4(n7786), .ZN(n7787)
         );
  NOR4_X1 U9547 ( .A1(n8651), .A2(n8664), .A3(n8676), .A4(n7787), .ZN(n7788)
         );
  NAND4_X1 U9548 ( .A1(n8615), .A2(n8625), .A3(n8638), .A4(n7788), .ZN(n7789)
         );
  NAND2_X1 U9549 ( .A1(n7794), .A2(n7790), .ZN(n7950) );
  XNOR2_X1 U9550 ( .A(n7793), .B(n7803), .ZN(n7799) );
  XNOR2_X1 U9551 ( .A(n8814), .B(n7803), .ZN(n7797) );
  INV_X1 U9552 ( .A(n7794), .ZN(n7962) );
  NOR2_X1 U9553 ( .A1(n7962), .A2(n7803), .ZN(n7796) );
  INV_X1 U9554 ( .A(n7795), .ZN(n8572) );
  NOR2_X1 U9555 ( .A1(n8818), .A2(n8572), .ZN(n7806) );
  NOR4_X1 U9556 ( .A1(n7797), .A2(n7796), .A3(n7806), .A4(n7821), .ZN(n7798)
         );
  AOI21_X1 U9557 ( .B1(n7799), .B2(n7821), .A(n7798), .ZN(n7800) );
  NOR2_X1 U9558 ( .A1(n7821), .A2(n7803), .ZN(n7804) );
  OAI211_X1 U9559 ( .C1(n7806), .C2(n8814), .A(n7805), .B(n7804), .ZN(n7977)
         );
  MUX2_X1 U9560 ( .A(n7949), .B(n7951), .S(n7942), .Z(n7956) );
  INV_X1 U9561 ( .A(n7807), .ZN(n7808) );
  NOR2_X1 U9562 ( .A1(n7925), .A2(n7808), .ZN(n7811) );
  AOI21_X1 U9563 ( .B1(n8316), .B2(n8788), .A(n7809), .ZN(n7810) );
  MUX2_X1 U9564 ( .A(n7811), .B(n7810), .S(n7942), .Z(n7931) );
  NAND2_X1 U9565 ( .A1(n8690), .A2(n7812), .ZN(n7818) );
  AND2_X1 U9566 ( .A1(n7812), .A2(n7905), .ZN(n7813) );
  OAI21_X1 U9567 ( .B1(n7813), .B2(n7942), .A(n7815), .ZN(n7819) );
  AND2_X1 U9568 ( .A1(n7912), .A2(n7814), .ZN(n7816) );
  OAI211_X1 U9569 ( .C1(n7819), .C2(n7816), .A(n8673), .B(n7815), .ZN(n7817)
         );
  MUX2_X1 U9570 ( .A(n7818), .B(n7817), .S(n7963), .Z(n7920) );
  INV_X1 U9571 ( .A(n7819), .ZN(n7913) );
  OAI21_X1 U9572 ( .B1(n7830), .B2(n4594), .A(n7824), .ZN(n7825) );
  MUX2_X1 U9573 ( .A(n7825), .B(n7824), .S(n7963), .Z(n7838) );
  INV_X1 U9574 ( .A(n7826), .ZN(n7827) );
  NOR2_X1 U9575 ( .A1(n7828), .A2(n7827), .ZN(n7831) );
  AOI21_X1 U9576 ( .B1(n7831), .B2(n7830), .A(n7829), .ZN(n7837) );
  NAND2_X1 U9577 ( .A1(n7847), .A2(n7832), .ZN(n7835) );
  NAND2_X1 U9578 ( .A1(n7841), .A2(n7833), .ZN(n7834) );
  MUX2_X1 U9579 ( .A(n7835), .B(n7834), .S(n7963), .Z(n7836) );
  AOI21_X1 U9580 ( .B1(n7838), .B2(n7837), .A(n7836), .ZN(n7840) );
  INV_X1 U9581 ( .A(n7841), .ZN(n7845) );
  INV_X1 U9582 ( .A(n7842), .ZN(n7843) );
  NOR2_X1 U9583 ( .A1(n7843), .A2(n7846), .ZN(n7853) );
  INV_X1 U9584 ( .A(n7847), .ZN(n7850) );
  OAI211_X1 U9585 ( .C1(n7851), .C2(n7850), .A(n7849), .B(n7848), .ZN(n7854)
         );
  AOI21_X1 U9586 ( .B1(n7854), .B2(n7853), .A(n4606), .ZN(n7855) );
  INV_X1 U9587 ( .A(n7856), .ZN(n7858) );
  NAND2_X1 U9588 ( .A1(n7867), .A2(n7866), .ZN(n7857) );
  MUX2_X1 U9589 ( .A(n7858), .B(n7857), .S(n7942), .Z(n7861) );
  INV_X1 U9590 ( .A(n7859), .ZN(n7860) );
  OR2_X1 U9591 ( .A1(n7861), .A2(n7860), .ZN(n7869) );
  NOR2_X1 U9592 ( .A1(n7869), .A2(n7862), .ZN(n7873) );
  OAI21_X1 U9593 ( .B1(n7869), .B2(n7864), .A(n7863), .ZN(n7871) );
  AND2_X1 U9594 ( .A1(n7866), .A2(n7865), .ZN(n7868) );
  OAI211_X1 U9595 ( .C1(n7869), .C2(n7868), .A(n7867), .B(n7875), .ZN(n7870)
         );
  MUX2_X1 U9596 ( .A(n7871), .B(n7870), .S(n7963), .Z(n7872) );
  AOI21_X1 U9597 ( .B1(n7874), .B2(n7873), .A(n7872), .ZN(n7882) );
  NAND2_X1 U9598 ( .A1(n7880), .A2(n7875), .ZN(n7877) );
  NAND2_X1 U9599 ( .A1(n7876), .A2(n8445), .ZN(n7879) );
  OAI21_X1 U9600 ( .B1(n7882), .B2(n7877), .A(n7879), .ZN(n7884) );
  NAND2_X1 U9601 ( .A1(n7879), .A2(n7878), .ZN(n7881) );
  OAI21_X1 U9602 ( .B1(n7882), .B2(n7881), .A(n7880), .ZN(n7883) );
  MUX2_X1 U9603 ( .A(n7886), .B(n7885), .S(n7963), .Z(n7887) );
  NAND2_X1 U9604 ( .A1(n9748), .A2(n9736), .ZN(n7889) );
  MUX2_X1 U9605 ( .A(n7890), .B(n7889), .S(n7942), .Z(n7891) );
  MUX2_X1 U9606 ( .A(n7894), .B(n7893), .S(n7963), .Z(n7895) );
  NAND3_X1 U9607 ( .A1(n8253), .A2(n9733), .A3(n7963), .ZN(n7897) );
  NAND3_X1 U9608 ( .A1(n7898), .A2(n8749), .A3(n7897), .ZN(n7907) );
  INV_X1 U9609 ( .A(n7899), .ZN(n7900) );
  NOR2_X1 U9610 ( .A1(n7907), .A2(n7900), .ZN(n7906) );
  MUX2_X1 U9611 ( .A(n7902), .B(n7901), .S(n7963), .Z(n7903) );
  NAND2_X1 U9612 ( .A1(n4838), .A2(n7903), .ZN(n7908) );
  OAI211_X1 U9613 ( .C1(n7906), .C2(n7908), .A(n7905), .B(n7904), .ZN(n7911)
         );
  INV_X1 U9614 ( .A(n7907), .ZN(n7909) );
  OAI21_X1 U9615 ( .B1(n7909), .B2(n7908), .A(n7963), .ZN(n7910) );
  AND4_X1 U9616 ( .A1(n7913), .A2(n7912), .A3(n7911), .A4(n7910), .ZN(n7919)
         );
  INV_X1 U9617 ( .A(n7921), .ZN(n7915) );
  NOR2_X1 U9618 ( .A1(n7915), .A2(n7914), .ZN(n7916) );
  MUX2_X1 U9619 ( .A(n7917), .B(n7916), .S(n7963), .Z(n7918) );
  OAI21_X1 U9620 ( .B1(n7920), .B2(n7919), .A(n7918), .ZN(n7924) );
  MUX2_X1 U9621 ( .A(n7922), .B(n7921), .S(n7942), .Z(n7923) );
  INV_X1 U9622 ( .A(n7925), .ZN(n7926) );
  NAND2_X1 U9623 ( .A1(n7933), .A2(n7926), .ZN(n7929) );
  NAND2_X1 U9624 ( .A1(n7932), .A2(n7927), .ZN(n7928) );
  MUX2_X1 U9625 ( .A(n7929), .B(n7928), .S(n7963), .Z(n7930) );
  MUX2_X1 U9626 ( .A(n7933), .B(n7932), .S(n7942), .Z(n7934) );
  NAND2_X1 U9627 ( .A1(n8625), .A2(n7934), .ZN(n7938) );
  MUX2_X1 U9628 ( .A(n7936), .B(n7935), .S(n7942), .Z(n7937) );
  MUX2_X1 U9629 ( .A(n7940), .B(n7939), .S(n7963), .Z(n7941) );
  NAND2_X1 U9630 ( .A1(n8829), .A2(n8423), .ZN(n7944) );
  MUX2_X1 U9631 ( .A(n7944), .B(n7943), .S(n7942), .Z(n7945) );
  NAND2_X1 U9632 ( .A1(n7946), .A2(n7945), .ZN(n7955) );
  AOI21_X1 U9633 ( .B1(n7952), .B2(n7949), .A(n7948), .ZN(n7954) );
  AOI21_X1 U9634 ( .B1(n7952), .B2(n7951), .A(n7950), .ZN(n7953) );
  MUX2_X1 U9635 ( .A(n7954), .B(n7953), .S(n7963), .Z(n7961) );
  INV_X1 U9636 ( .A(n7955), .ZN(n7958) );
  INV_X1 U9637 ( .A(n7956), .ZN(n7957) );
  NAND3_X1 U9638 ( .A1(n7959), .A2(n7958), .A3(n7957), .ZN(n7960) );
  NAND2_X1 U9639 ( .A1(n7961), .A2(n7960), .ZN(n7967) );
  INV_X1 U9640 ( .A(n7969), .ZN(n7970) );
  NOR2_X1 U9641 ( .A1(n7971), .A2(n6448), .ZN(n7975) );
  NOR2_X1 U9642 ( .A1(n7973), .A2(n7972), .ZN(n7974) );
  NAND3_X1 U9643 ( .A1(n7980), .A2(n7979), .A3(n7978), .ZN(n7981) );
  OAI211_X1 U9644 ( .C1(n7982), .C2(n7984), .A(n7981), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7983) );
  INV_X1 U9645 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U9646 ( .A1(n7985), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7987) );
  NAND2_X1 U9647 ( .A1(n5120), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7986) );
  OAI211_X1 U9648 ( .C1(n5149), .C2(n9545), .A(n7987), .B(n7986), .ZN(n9271)
         );
  INV_X1 U9649 ( .A(n9271), .ZN(n8036) );
  NAND2_X1 U9650 ( .A1(n8213), .A2(n8036), .ZN(n8076) );
  NAND2_X1 U9651 ( .A1(n9321), .A2(n7988), .ZN(n8205) );
  AND2_X1 U9652 ( .A1(n8076), .A2(n8205), .ZN(n8088) );
  INV_X1 U9653 ( .A(n8088), .ZN(n8038) );
  NAND2_X1 U9654 ( .A1(n8206), .A2(n8201), .ZN(n8086) );
  NAND2_X1 U9655 ( .A1(n9563), .A2(n9312), .ZN(n9266) );
  NAND2_X1 U9656 ( .A1(n9381), .A2(n9307), .ZN(n9265) );
  AND2_X1 U9657 ( .A1(n9266), .A2(n9265), .ZN(n8195) );
  OR2_X1 U9658 ( .A1(n9381), .A2(n9307), .ZN(n8193) );
  OR2_X1 U9659 ( .A1(n9574), .A2(n9172), .ZN(n9373) );
  OR2_X1 U9660 ( .A1(n9579), .A2(n9301), .ZN(n8185) );
  OR2_X1 U9661 ( .A1(n9424), .A2(n9299), .ZN(n9261) );
  NAND2_X1 U9662 ( .A1(n8185), .A2(n9261), .ZN(n8098) );
  NAND2_X1 U9663 ( .A1(n9579), .A2(n9301), .ZN(n9264) );
  NAND2_X1 U9664 ( .A1(n8098), .A2(n9264), .ZN(n7989) );
  NAND2_X1 U9665 ( .A1(n9373), .A2(n7989), .ZN(n7990) );
  NAND2_X1 U9666 ( .A1(n9574), .A2(n9172), .ZN(n8189) );
  NAND2_X1 U9667 ( .A1(n7990), .A2(n8189), .ZN(n7991) );
  AND2_X1 U9668 ( .A1(n8193), .A2(n7991), .ZN(n7998) );
  NAND2_X1 U9669 ( .A1(n9424), .A2(n9299), .ZN(n9262) );
  NAND2_X1 U9670 ( .A1(n9264), .A2(n9262), .ZN(n8097) );
  INV_X1 U9671 ( .A(n8097), .ZN(n7992) );
  NAND2_X1 U9672 ( .A1(n9444), .A2(n9293), .ZN(n8181) );
  NAND2_X1 U9673 ( .A1(n9460), .A2(n9173), .ZN(n9259) );
  NAND2_X1 U9674 ( .A1(n8181), .A2(n9259), .ZN(n8177) );
  OR2_X1 U9675 ( .A1(n9444), .A2(n9293), .ZN(n8182) );
  NAND2_X1 U9676 ( .A1(n8177), .A2(n8182), .ZN(n9260) );
  NAND3_X1 U9677 ( .A1(n8189), .A2(n7992), .A3(n9260), .ZN(n7993) );
  NAND2_X1 U9678 ( .A1(n7998), .A2(n7993), .ZN(n7994) );
  AND2_X1 U9679 ( .A1(n8195), .A2(n7994), .ZN(n7995) );
  NAND2_X1 U9680 ( .A1(n8045), .A2(n8198), .ZN(n8000) );
  NOR2_X1 U9681 ( .A1(n7995), .A2(n8000), .ZN(n7997) );
  NAND2_X1 U9682 ( .A1(n9334), .A2(n7996), .ZN(n9268) );
  NAND2_X1 U9683 ( .A1(n9268), .A2(n9328), .ZN(n9267) );
  OR2_X1 U9684 ( .A1(n7997), .A2(n9267), .ZN(n8084) );
  INV_X1 U9685 ( .A(n7998), .ZN(n7999) );
  OR2_X1 U9686 ( .A1(n9460), .A2(n9173), .ZN(n9433) );
  NAND2_X1 U9687 ( .A1(n8182), .A2(n9433), .ZN(n8176) );
  OR3_X1 U9688 ( .A1(n8000), .A2(n7999), .A3(n8176), .ZN(n8082) );
  OR2_X1 U9689 ( .A1(n9474), .A2(n9290), .ZN(n8099) );
  OR2_X1 U9690 ( .A1(n9493), .A2(n9287), .ZN(n8046) );
  OR2_X1 U9691 ( .A1(n9512), .A2(n9284), .ZN(n9483) );
  NAND2_X1 U9692 ( .A1(n8046), .A2(n9483), .ZN(n8174) );
  INV_X1 U9693 ( .A(n9281), .ZN(n9103) );
  NAND2_X1 U9694 ( .A1(n9529), .A2(n9103), .ZN(n9502) );
  NAND2_X1 U9695 ( .A1(n9274), .A2(n9279), .ZN(n8079) );
  NAND2_X1 U9696 ( .A1(n9502), .A2(n8079), .ZN(n8100) );
  NOR2_X1 U9697 ( .A1(n8002), .A2(n8001), .ZN(n8155) );
  AND2_X1 U9698 ( .A1(n8115), .A2(n8003), .ZN(n8004) );
  NAND2_X1 U9699 ( .A1(n8005), .A2(n8004), .ZN(n8119) );
  NAND2_X1 U9700 ( .A1(n9184), .A2(n8006), .ZN(n8007) );
  NAND4_X1 U9701 ( .A1(n8009), .A2(n8008), .A3(n8225), .A4(n8007), .ZN(n8014)
         );
  INV_X1 U9702 ( .A(n8010), .ZN(n8013) );
  INV_X1 U9703 ( .A(n8011), .ZN(n8012) );
  NOR3_X1 U9704 ( .A1(n8014), .A2(n8013), .A3(n8012), .ZN(n8015) );
  OAI21_X1 U9705 ( .B1(n8119), .B2(n8015), .A(n8118), .ZN(n8018) );
  INV_X1 U9706 ( .A(n8016), .ZN(n8017) );
  AOI21_X1 U9707 ( .B1(n8019), .B2(n8018), .A(n8017), .ZN(n8020) );
  NAND2_X1 U9708 ( .A1(n8155), .A2(n8020), .ZN(n8024) );
  AOI21_X1 U9709 ( .B1(n8023), .B2(n8022), .A(n8021), .ZN(n8141) );
  NAND3_X1 U9710 ( .A1(n8024), .A2(n8141), .A3(n8138), .ZN(n8025) );
  NAND3_X1 U9711 ( .A1(n8025), .A2(n8148), .A3(n8149), .ZN(n8026) );
  NAND2_X1 U9712 ( .A1(n8026), .A2(n8139), .ZN(n8029) );
  OR2_X1 U9713 ( .A1(n9274), .A2(n9279), .ZN(n8145) );
  NAND2_X1 U9714 ( .A1(n8164), .A2(n8145), .ZN(n8027) );
  NAND2_X1 U9715 ( .A1(n8027), .A2(n9502), .ZN(n8028) );
  OAI21_X1 U9716 ( .B1(n8100), .B2(n8029), .A(n8028), .ZN(n8031) );
  NAND2_X1 U9717 ( .A1(n9493), .A2(n9287), .ZN(n8172) );
  NAND2_X1 U9718 ( .A1(n9512), .A2(n9284), .ZN(n8047) );
  NAND2_X1 U9719 ( .A1(n8172), .A2(n8047), .ZN(n8171) );
  INV_X1 U9720 ( .A(n8171), .ZN(n8030) );
  OAI21_X1 U9721 ( .B1(n8174), .B2(n8031), .A(n8030), .ZN(n8032) );
  NAND2_X1 U9722 ( .A1(n9474), .A2(n9290), .ZN(n8173) );
  AOI21_X1 U9723 ( .B1(n4351), .B2(n8032), .A(n4563), .ZN(n8033) );
  NOR2_X1 U9724 ( .A1(n8082), .A2(n8033), .ZN(n8034) );
  NOR2_X1 U9725 ( .A1(n8084), .A2(n8034), .ZN(n8035) );
  NOR2_X1 U9726 ( .A1(n8086), .A2(n8035), .ZN(n8037) );
  OR2_X1 U9727 ( .A1(n8213), .A2(n8036), .ZN(n8090) );
  OAI21_X1 U9728 ( .B1(n8038), .B2(n8037), .A(n8090), .ZN(n8042) );
  NAND2_X1 U9729 ( .A1(n9029), .A2(n5346), .ZN(n8041) );
  OR2_X1 U9730 ( .A1(n5127), .A2(n8039), .ZN(n8040) );
  OR2_X1 U9731 ( .A1(n9253), .A2(n8043), .ZN(n8226) );
  NAND2_X1 U9732 ( .A1(n8042), .A2(n8226), .ZN(n8044) );
  AND2_X1 U9733 ( .A1(n9253), .A2(n8043), .ZN(n8211) );
  INV_X1 U9734 ( .A(n8211), .ZN(n8224) );
  NAND2_X1 U9735 ( .A1(n8044), .A2(n8224), .ZN(n8236) );
  NAND2_X1 U9736 ( .A1(n8236), .A2(n5437), .ZN(n8234) );
  OR2_X1 U9737 ( .A1(n9316), .A2(n9351), .ZN(n8202) );
  NAND2_X1 U9738 ( .A1(n8198), .A2(n9266), .ZN(n9356) );
  NAND2_X1 U9739 ( .A1(n9433), .A2(n9259), .ZN(n9455) );
  NAND2_X1 U9740 ( .A1(n8164), .A2(n9502), .ZN(n9283) );
  NAND4_X1 U9741 ( .A1(n8051), .A2(n8050), .A3(n8049), .A4(n8048), .ZN(n8053)
         );
  NOR2_X1 U9742 ( .A1(n8053), .A2(n8052), .ZN(n8057) );
  NAND4_X1 U9743 ( .A1(n8057), .A2(n8056), .A3(n8055), .A4(n8054), .ZN(n8058)
         );
  OR3_X1 U9744 ( .A1(n8060), .A2(n8059), .A3(n8058), .ZN(n8061) );
  NOR2_X1 U9745 ( .A1(n8061), .A2(n9914), .ZN(n8063) );
  NAND4_X1 U9746 ( .A1(n8065), .A2(n8064), .A3(n8063), .A4(n8062), .ZN(n8066)
         );
  NOR4_X1 U9747 ( .A1(n9503), .A2(n9283), .A3(n8067), .A4(n8066), .ZN(n8069)
         );
  NAND4_X1 U9748 ( .A1(n9471), .A2(n9486), .A3(n8069), .A4(n8068), .ZN(n8070)
         );
  NOR2_X1 U9749 ( .A1(n9455), .A2(n8070), .ZN(n8071) );
  XNOR2_X1 U9750 ( .A(n9424), .B(n9299), .ZN(n9416) );
  INV_X1 U9751 ( .A(n9416), .ZN(n9418) );
  NAND4_X1 U9752 ( .A1(n9409), .A2(n9435), .A3(n8071), .A4(n9418), .ZN(n8072)
         );
  NOR2_X1 U9753 ( .A1(n4542), .A2(n8072), .ZN(n8073) );
  NAND2_X1 U9754 ( .A1(n9379), .A2(n8073), .ZN(n8074) );
  OR3_X1 U9755 ( .A1(n8202), .A2(n9356), .A3(n8074), .ZN(n8075) );
  NOR2_X1 U9756 ( .A1(n9318), .A2(n8075), .ZN(n8077) );
  AND3_X1 U9757 ( .A1(n8077), .A2(n8090), .A3(n8076), .ZN(n8078) );
  AND3_X1 U9758 ( .A1(n8226), .A2(n8078), .A3(n8224), .ZN(n8221) );
  INV_X1 U9759 ( .A(n8221), .ZN(n8096) );
  NOR2_X1 U9760 ( .A1(n8213), .A2(n8215), .ZN(n8089) );
  INV_X1 U9761 ( .A(n9283), .ZN(n9524) );
  INV_X1 U9762 ( .A(n9503), .ZN(n9285) );
  NAND3_X1 U9763 ( .A1(n9520), .A2(n9285), .A3(n9502), .ZN(n9506) );
  NOR2_X1 U9764 ( .A1(n8082), .A2(n9451), .ZN(n8083) );
  NOR2_X1 U9765 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  OR2_X1 U9766 ( .A1(n8086), .A2(n8085), .ZN(n8087) );
  OAI211_X1 U9767 ( .C1(n9253), .C2(n8089), .A(n8088), .B(n8087), .ZN(n8094)
         );
  INV_X1 U9768 ( .A(n8090), .ZN(n8091) );
  NAND2_X1 U9769 ( .A1(n8091), .A2(n9253), .ZN(n8092) );
  NAND4_X1 U9770 ( .A1(n8094), .A2(n8093), .A3(n8224), .A4(n8092), .ZN(n8095)
         );
  NAND2_X1 U9771 ( .A1(n8096), .A2(n8095), .ZN(n8222) );
  MUX2_X1 U9772 ( .A(n8098), .B(n8097), .S(n8223), .Z(n8188) );
  AOI21_X1 U9773 ( .B1(n9433), .B2(n8099), .A(n8223), .ZN(n8180) );
  NAND2_X1 U9774 ( .A1(n8100), .A2(n8164), .ZN(n8168) );
  OAI21_X1 U9775 ( .B1(n8223), .B2(n9274), .A(n8168), .ZN(n8103) );
  NAND2_X1 U9776 ( .A1(n9502), .A2(n9275), .ZN(n8101) );
  NAND2_X1 U9777 ( .A1(n8101), .A2(n8209), .ZN(n8102) );
  NAND2_X1 U9778 ( .A1(n8103), .A2(n8102), .ZN(n8170) );
  INV_X1 U9779 ( .A(n8164), .ZN(n8104) );
  NAND2_X1 U9780 ( .A1(n8104), .A2(n8223), .ZN(n8167) );
  NOR2_X1 U9781 ( .A1(n9175), .A2(n8223), .ZN(n8105) );
  NAND2_X1 U9782 ( .A1(n8110), .A2(n8105), .ZN(n8109) );
  OAI21_X1 U9783 ( .B1(n8223), .B2(n9174), .A(n8109), .ZN(n8107) );
  NAND2_X1 U9784 ( .A1(n8107), .A2(n8106), .ZN(n8108) );
  OAI21_X1 U9785 ( .B1(n8109), .B2(n9174), .A(n8108), .ZN(n8147) );
  NAND2_X1 U9786 ( .A1(n9175), .A2(n8223), .ZN(n8112) );
  OAI22_X1 U9787 ( .A1(n8110), .A2(n8112), .B1(n8111), .B2(n8209), .ZN(n8114)
         );
  NOR2_X1 U9788 ( .A1(n8112), .A2(n8111), .ZN(n8113) );
  AOI22_X1 U9789 ( .A1(n9686), .A2(n8114), .B1(n9966), .B2(n8113), .ZN(n8144)
         );
  NAND2_X1 U9790 ( .A1(n8120), .A2(n8115), .ZN(n8116) );
  AOI21_X1 U9791 ( .B1(n8117), .B2(n8118), .A(n8116), .ZN(n8123) );
  NAND3_X1 U9792 ( .A1(n8119), .A2(n8124), .A3(n8118), .ZN(n8121) );
  NAND2_X1 U9793 ( .A1(n8121), .A2(n8120), .ZN(n8122) );
  MUX2_X1 U9794 ( .A(n8123), .B(n8122), .S(n8223), .Z(n8127) );
  NOR2_X1 U9795 ( .A1(n8124), .A2(n8223), .ZN(n8126) );
  OAI21_X1 U9796 ( .B1(n8127), .B2(n8126), .A(n8125), .ZN(n8131) );
  MUX2_X1 U9797 ( .A(n8129), .B(n8128), .S(n8209), .Z(n8130) );
  NAND2_X1 U9798 ( .A1(n8131), .A2(n8130), .ZN(n8136) );
  AND2_X1 U9799 ( .A1(n8154), .A2(n8132), .ZN(n8133) );
  MUX2_X1 U9800 ( .A(n8134), .B(n8133), .S(n8223), .Z(n8135) );
  NAND2_X1 U9801 ( .A1(n8136), .A2(n8135), .ZN(n8150) );
  NAND2_X1 U9802 ( .A1(n8150), .A2(n8151), .ZN(n8137) );
  NAND2_X1 U9803 ( .A1(n8137), .A2(n8155), .ZN(n8142) );
  AND2_X1 U9804 ( .A1(n8138), .A2(n8223), .ZN(n8140) );
  NAND4_X1 U9805 ( .A1(n8142), .A2(n8141), .A3(n8140), .A4(n8139), .ZN(n8143)
         );
  NAND3_X1 U9806 ( .A1(n8145), .A2(n8144), .A3(n8143), .ZN(n8146) );
  AOI21_X1 U9807 ( .B1(n8164), .B2(n8147), .A(n8146), .ZN(n8166) );
  AND3_X1 U9808 ( .A1(n8149), .A2(n8209), .A3(n8148), .ZN(n8163) );
  INV_X1 U9809 ( .A(n8152), .ZN(n8153) );
  INV_X1 U9810 ( .A(n8155), .ZN(n8161) );
  INV_X1 U9811 ( .A(n8156), .ZN(n8160) );
  AND2_X1 U9812 ( .A1(n8158), .A2(n8157), .ZN(n8159) );
  NAND3_X1 U9813 ( .A1(n8164), .A2(n8163), .A3(n8162), .ZN(n8165) );
  NAND4_X1 U9814 ( .A1(n8168), .A2(n8167), .A3(n8166), .A4(n8165), .ZN(n8169)
         );
  AOI21_X1 U9815 ( .B1(n8170), .B2(n8169), .A(n9503), .ZN(n8175) );
  MUX2_X1 U9816 ( .A(n8177), .B(n8176), .S(n8223), .Z(n8178) );
  INV_X1 U9817 ( .A(n8178), .ZN(n8179) );
  MUX2_X1 U9818 ( .A(n8182), .B(n8181), .S(n8223), .Z(n8183) );
  AOI21_X1 U9819 ( .B1(n8184), .B2(n8183), .A(n9416), .ZN(n8187) );
  MUX2_X1 U9820 ( .A(n9264), .B(n8185), .S(n8223), .Z(n8186) );
  OAI211_X1 U9821 ( .C1(n8188), .C2(n8187), .A(n9390), .B(n8186), .ZN(n8191)
         );
  MUX2_X1 U9822 ( .A(n9373), .B(n8189), .S(n8223), .Z(n8190) );
  NAND2_X1 U9823 ( .A1(n8198), .A2(n8193), .ZN(n8192) );
  AOI22_X1 U9824 ( .A1(n8195), .A2(n8194), .B1(n8192), .B2(n9266), .ZN(n8200)
         );
  INV_X1 U9825 ( .A(n8193), .ZN(n8197) );
  INV_X1 U9826 ( .A(n8194), .ZN(n8196) );
  OAI21_X1 U9827 ( .B1(n8197), .B2(n8196), .A(n8195), .ZN(n8199) );
  NAND2_X1 U9828 ( .A1(n9267), .A2(n8201), .ZN(n8203) );
  MUX2_X1 U9829 ( .A(n8206), .B(n8205), .S(n8223), .Z(n8207) );
  NAND2_X1 U9830 ( .A1(n8208), .A2(n8207), .ZN(n8214) );
  MUX2_X1 U9831 ( .A(n8209), .B(n8214), .S(n8213), .Z(n8220) );
  NAND2_X1 U9832 ( .A1(n9253), .A2(n9271), .ZN(n8219) );
  NAND2_X1 U9833 ( .A1(n8215), .A2(n9271), .ZN(n8216) );
  OR2_X1 U9834 ( .A1(n8224), .A2(n8223), .ZN(n8228) );
  OAI211_X1 U9835 ( .C1(n8226), .C2(n9350), .A(n8225), .B(n5698), .ZN(n8227)
         );
  AOI21_X1 U9836 ( .B1(n8229), .B2(n8228), .A(n8227), .ZN(n8230) );
  NOR2_X1 U9837 ( .A1(n8231), .A2(n8230), .ZN(n8233) );
  INV_X1 U9838 ( .A(n8238), .ZN(n8243) );
  OAI21_X1 U9839 ( .B1(n8238), .B2(n8237), .A(P1_B_REG_SCAN_IN), .ZN(n8239) );
  AOI21_X1 U9840 ( .B1(n8241), .B2(n8240), .A(n8239), .ZN(n8242) );
  XNOR2_X1 U9841 ( .A(n8829), .B(n8293), .ZN(n8292) );
  NAND2_X1 U9842 ( .A1(n8245), .A2(n8244), .ZN(n8247) );
  NAND2_X1 U9843 ( .A1(n8247), .A2(n8246), .ZN(n9738) );
  INV_X1 U9844 ( .A(n9738), .ZN(n8252) );
  XNOR2_X1 U9845 ( .A(n8248), .B(n8293), .ZN(n8250) );
  XNOR2_X1 U9846 ( .A(n8250), .B(n8249), .ZN(n9739) );
  INV_X1 U9847 ( .A(n9739), .ZN(n8251) );
  XNOR2_X1 U9848 ( .A(n8253), .B(n8293), .ZN(n8254) );
  XNOR2_X1 U9849 ( .A(n8254), .B(n8442), .ZN(n8429) );
  NAND2_X1 U9850 ( .A1(n8430), .A2(n8429), .ZN(n8428) );
  INV_X1 U9851 ( .A(n8254), .ZN(n8255) );
  NAND2_X1 U9852 ( .A1(n8255), .A2(n8442), .ZN(n8256) );
  XNOR2_X1 U9853 ( .A(n8809), .B(n6715), .ZN(n8354) );
  XNOR2_X1 U9854 ( .A(n9018), .B(n8293), .ZN(n8257) );
  NAND2_X1 U9855 ( .A1(n8257), .A2(n8755), .ZN(n8402) );
  INV_X1 U9856 ( .A(n8257), .ZN(n8258) );
  NAND2_X1 U9857 ( .A1(n8258), .A2(n8720), .ZN(n8259) );
  NAND2_X1 U9858 ( .A1(n8402), .A2(n8259), .ZN(n8365) );
  NAND2_X1 U9859 ( .A1(n8363), .A2(n8402), .ZN(n8260) );
  XNOR2_X1 U9860 ( .A(n9012), .B(n8293), .ZN(n8261) );
  XNOR2_X1 U9861 ( .A(n8261), .B(n8738), .ZN(n8403) );
  NAND2_X1 U9862 ( .A1(n8260), .A2(n8403), .ZN(n8406) );
  NAND2_X1 U9863 ( .A1(n8261), .A2(n8705), .ZN(n8262) );
  XNOR2_X1 U9864 ( .A(n8799), .B(n8293), .ZN(n8267) );
  XNOR2_X1 U9865 ( .A(n8267), .B(n8386), .ZN(n8321) );
  XNOR2_X1 U9866 ( .A(n9002), .B(n8293), .ZN(n8264) );
  NAND2_X1 U9867 ( .A1(n8264), .A2(n8706), .ZN(n8332) );
  INV_X1 U9868 ( .A(n8264), .ZN(n8265) );
  NAND2_X1 U9869 ( .A1(n8265), .A2(n8681), .ZN(n8266) );
  NAND2_X1 U9870 ( .A1(n8332), .A2(n8266), .ZN(n8380) );
  INV_X1 U9871 ( .A(n8267), .ZN(n8268) );
  AND2_X1 U9872 ( .A1(n8268), .A2(n8721), .ZN(n8379) );
  NOR2_X1 U9873 ( .A1(n8380), .A2(n8379), .ZN(n8331) );
  XNOR2_X1 U9874 ( .A(n8996), .B(n8293), .ZN(n8271) );
  XNOR2_X1 U9875 ( .A(n8271), .B(n8693), .ZN(n8333) );
  AND2_X1 U9876 ( .A1(n8331), .A2(n8333), .ZN(n8269) );
  NAND2_X1 U9877 ( .A1(n8271), .A2(n8270), .ZN(n8273) );
  INV_X1 U9878 ( .A(n8333), .ZN(n8272) );
  AND2_X1 U9879 ( .A1(n8273), .A2(n8335), .ZN(n8274) );
  XNOR2_X1 U9880 ( .A(n8788), .B(n8293), .ZN(n8275) );
  XNOR2_X1 U9881 ( .A(n8275), .B(n8316), .ZN(n8392) );
  INV_X1 U9882 ( .A(n8275), .ZN(n8276) );
  NAND2_X1 U9883 ( .A1(n8276), .A2(n8682), .ZN(n8277) );
  XNOR2_X1 U9884 ( .A(n8853), .B(n6715), .ZN(n8279) );
  XNOR2_X1 U9885 ( .A(n8847), .B(n8293), .ZN(n8283) );
  NAND2_X1 U9886 ( .A1(n8283), .A2(n8282), .ZN(n8286) );
  INV_X1 U9887 ( .A(n8283), .ZN(n8284) );
  NAND2_X1 U9888 ( .A1(n8284), .A2(n8653), .ZN(n8285) );
  NAND2_X1 U9889 ( .A1(n8286), .A2(n8285), .ZN(n8372) );
  AOI21_X1 U9890 ( .B1(n8373), .B2(n8281), .A(n8372), .ZN(n8343) );
  INV_X1 U9891 ( .A(n8286), .ZN(n8345) );
  XNOR2_X1 U9892 ( .A(n8841), .B(n8293), .ZN(n8288) );
  NAND2_X1 U9893 ( .A1(n8288), .A2(n8287), .ZN(n8417) );
  INV_X1 U9894 ( .A(n8288), .ZN(n8289) );
  NAND2_X1 U9895 ( .A1(n8289), .A2(n8639), .ZN(n8290) );
  XNOR2_X1 U9896 ( .A(n8835), .B(n8293), .ZN(n8291) );
  XNOR2_X1 U9897 ( .A(n8291), .B(n8349), .ZN(n8418) );
  XNOR2_X1 U9898 ( .A(n8292), .B(n8617), .ZN(n8305) );
  OAI21_X1 U9899 ( .B1(n8423), .B2(n8292), .A(n8304), .ZN(n8295) );
  XNOR2_X1 U9900 ( .A(n8588), .B(n8293), .ZN(n8294) );
  XNOR2_X1 U9901 ( .A(n8295), .B(n8294), .ZN(n8301) );
  OAI22_X1 U9902 ( .A1(n8423), .A2(n8412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8296), .ZN(n8299) );
  INV_X1 U9903 ( .A(n8598), .ZN(n8297) );
  OAI22_X1 U9904 ( .A1(n8441), .A2(n9734), .B1(n8297), .B2(n9746), .ZN(n8298)
         );
  AOI211_X1 U9905 ( .C1(n8823), .C2(n8369), .A(n8299), .B(n8298), .ZN(n8300)
         );
  OAI21_X1 U9906 ( .B1(n8301), .B2(n8391), .A(n8300), .ZN(P2_U3160) );
  OAI222_X1 U9907 ( .A1(n8303), .A2(n8956), .B1(n9694), .B2(n8302), .C1(
        P1_U3086), .C2(n9350), .ZN(P1_U3336) );
  INV_X1 U9908 ( .A(n8829), .ZN(n8312) );
  OAI211_X1 U9909 ( .C1(n8306), .C2(n8305), .A(n8304), .B(n9742), .ZN(n8311)
         );
  INV_X1 U9910 ( .A(n8611), .ZN(n8308) );
  AOI22_X1 U9911 ( .A1(n8629), .A2(n9737), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8307) );
  OAI21_X1 U9912 ( .B1(n8308), .B2(n9746), .A(n8307), .ZN(n8309) );
  AOI21_X1 U9913 ( .B1(n8410), .B2(n8607), .A(n8309), .ZN(n8310) );
  OAI211_X1 U9914 ( .C1(n8312), .C2(n8438), .A(n8311), .B(n8310), .ZN(P2_U3154) );
  OAI21_X1 U9915 ( .B1(n8397), .B2(n8313), .A(n8373), .ZN(n8314) );
  NAND2_X1 U9916 ( .A1(n8314), .A2(n9742), .ZN(n8319) );
  AOI22_X1 U9917 ( .A1(n8653), .A2(n8410), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8315) );
  OAI21_X1 U9918 ( .B1(n8316), .B2(n8412), .A(n8315), .ZN(n8317) );
  AOI21_X1 U9919 ( .B1(n8656), .B2(n8434), .A(n8317), .ZN(n8318) );
  OAI211_X1 U9920 ( .C1(n8320), .C2(n8438), .A(n8319), .B(n8318), .ZN(P2_U3156) );
  INV_X1 U9921 ( .A(n8799), .ZN(n8330) );
  AOI21_X1 U9922 ( .B1(n8322), .B2(n8321), .A(n8391), .ZN(n8324) );
  NAND2_X1 U9923 ( .A1(n8324), .A2(n8383), .ZN(n8329) );
  NOR2_X1 U9924 ( .A1(n8412), .A2(n8705), .ZN(n8327) );
  OAI21_X1 U9925 ( .B1(n8706), .B2(n9734), .A(n8325), .ZN(n8326) );
  AOI211_X1 U9926 ( .C1(n8711), .C2(n8434), .A(n8327), .B(n8326), .ZN(n8328)
         );
  OAI211_X1 U9927 ( .C1(n8330), .C2(n8438), .A(n8329), .B(n8328), .ZN(P2_U3159) );
  INV_X1 U9928 ( .A(n8996), .ZN(n8342) );
  INV_X1 U9929 ( .A(n8332), .ZN(n8334) );
  NOR3_X1 U9930 ( .A1(n4881), .A2(n8334), .A3(n8333), .ZN(n8337) );
  OAI21_X1 U9931 ( .B1(n8337), .B2(n4340), .A(n9742), .ZN(n8341) );
  AOI22_X1 U9932 ( .A1(n8682), .A2(n8410), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8338) );
  OAI21_X1 U9933 ( .B1(n8706), .B2(n8412), .A(n8338), .ZN(n8339) );
  AOI21_X1 U9934 ( .B1(n8685), .B2(n8434), .A(n8339), .ZN(n8340) );
  OAI211_X1 U9935 ( .C1(n8342), .C2(n8438), .A(n8341), .B(n8340), .ZN(P2_U3163) );
  INV_X1 U9936 ( .A(n8841), .ZN(n8353) );
  INV_X1 U9937 ( .A(n8419), .ZN(n8347) );
  NOR3_X1 U9938 ( .A1(n8343), .A2(n8345), .A3(n8344), .ZN(n8346) );
  OAI21_X1 U9939 ( .B1(n8347), .B2(n8346), .A(n9742), .ZN(n8352) );
  AOI22_X1 U9940 ( .A1(n8653), .A2(n9737), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8348) );
  OAI21_X1 U9941 ( .B1(n8349), .B2(n9734), .A(n8348), .ZN(n8350) );
  AOI21_X1 U9942 ( .B1(n8631), .B2(n8434), .A(n8350), .ZN(n8351) );
  OAI211_X1 U9943 ( .C1(n8353), .C2(n8438), .A(n8352), .B(n8351), .ZN(P2_U3165) );
  XNOR2_X1 U9944 ( .A(n8354), .B(n8432), .ZN(n8355) );
  XNOR2_X1 U9945 ( .A(n8356), .B(n8355), .ZN(n8362) );
  NAND2_X1 U9946 ( .A1(n8434), .A2(n8760), .ZN(n8359) );
  INV_X1 U9947 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8357) );
  NOR2_X1 U9948 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8357), .ZN(n8520) );
  AOI21_X1 U9949 ( .B1(n9737), .B2(n8442), .A(n8520), .ZN(n8358) );
  OAI211_X1 U9950 ( .C1(n8755), .C2(n9734), .A(n8359), .B(n8358), .ZN(n8360)
         );
  AOI21_X1 U9951 ( .B1(n8809), .B2(n8369), .A(n8360), .ZN(n8361) );
  OAI21_X1 U9952 ( .B1(n8362), .B2(n8391), .A(n8361), .ZN(P2_U3166) );
  INV_X1 U9953 ( .A(n8363), .ZN(n8405) );
  AOI21_X1 U9954 ( .B1(n8365), .B2(n8364), .A(n8405), .ZN(n8371) );
  NAND2_X1 U9955 ( .A1(n8434), .A2(n8732), .ZN(n8367) );
  AND2_X1 U9956 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8538) );
  AOI21_X1 U9957 ( .B1(n8410), .B2(n8738), .A(n8538), .ZN(n8366) );
  OAI211_X1 U9958 ( .C1(n8432), .C2(n8412), .A(n8367), .B(n8366), .ZN(n8368)
         );
  AOI21_X1 U9959 ( .B1(n9018), .B2(n8369), .A(n8368), .ZN(n8370) );
  OAI21_X1 U9960 ( .B1(n8371), .B2(n8391), .A(n8370), .ZN(P2_U3168) );
  INV_X1 U9961 ( .A(n8847), .ZN(n8645) );
  AND3_X1 U9962 ( .A1(n8373), .A2(n8281), .A3(n8372), .ZN(n8374) );
  OAI21_X1 U9963 ( .B1(n8343), .B2(n8374), .A(n9742), .ZN(n8378) );
  AOI22_X1 U9964 ( .A1(n8639), .A2(n8410), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8375) );
  OAI21_X1 U9965 ( .B1(n8397), .B2(n8412), .A(n8375), .ZN(n8376) );
  AOI21_X1 U9966 ( .B1(n8641), .B2(n8434), .A(n8376), .ZN(n8377) );
  OAI211_X1 U9967 ( .C1(n8645), .C2(n8438), .A(n8378), .B(n8377), .ZN(P2_U3169) );
  INV_X1 U9968 ( .A(n9002), .ZN(n8390) );
  INV_X1 U9969 ( .A(n8379), .ZN(n8382) );
  INV_X1 U9970 ( .A(n8380), .ZN(n8381) );
  AOI21_X1 U9971 ( .B1(n8383), .B2(n8382), .A(n8381), .ZN(n8384) );
  OAI21_X1 U9972 ( .B1(n4881), .B2(n8384), .A(n9742), .ZN(n8389) );
  AOI22_X1 U9973 ( .A1(n8693), .A2(n8410), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8385) );
  OAI21_X1 U9974 ( .B1(n8386), .B2(n8412), .A(n8385), .ZN(n8387) );
  AOI21_X1 U9975 ( .B1(n8696), .B2(n8434), .A(n8387), .ZN(n8388) );
  OAI211_X1 U9976 ( .C1(n8390), .C2(n8438), .A(n8389), .B(n8388), .ZN(P2_U3173) );
  INV_X1 U9977 ( .A(n8788), .ZN(n8401) );
  AOI21_X1 U9978 ( .B1(n8393), .B2(n8392), .A(n8391), .ZN(n8395) );
  NAND2_X1 U9979 ( .A1(n8395), .A2(n8394), .ZN(n8400) );
  AOI22_X1 U9980 ( .A1(n8693), .A2(n9737), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8396) );
  OAI21_X1 U9981 ( .B1(n8397), .B2(n9734), .A(n8396), .ZN(n8398) );
  AOI21_X1 U9982 ( .B1(n8667), .B2(n8434), .A(n8398), .ZN(n8399) );
  OAI211_X1 U9983 ( .C1(n8401), .C2(n8438), .A(n8400), .B(n8399), .ZN(P2_U3175) );
  INV_X1 U9984 ( .A(n9012), .ZN(n8416) );
  INV_X1 U9985 ( .A(n8402), .ZN(n8404) );
  NOR3_X1 U9986 ( .A1(n8405), .A2(n8404), .A3(n8403), .ZN(n8408) );
  INV_X1 U9987 ( .A(n8406), .ZN(n8407) );
  OAI21_X1 U9988 ( .B1(n8408), .B2(n8407), .A(n9742), .ZN(n8415) );
  NOR2_X1 U9989 ( .A1(n8409), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8567) );
  AOI21_X1 U9990 ( .B1(n8721), .B2(n8410), .A(n8567), .ZN(n8411) );
  OAI21_X1 U9991 ( .B1(n8755), .B2(n8412), .A(n8411), .ZN(n8413) );
  AOI21_X1 U9992 ( .B1(n8725), .B2(n8434), .A(n8413), .ZN(n8414) );
  OAI211_X1 U9993 ( .C1(n8416), .C2(n8438), .A(n8415), .B(n8414), .ZN(P2_U3178) );
  INV_X1 U9994 ( .A(n8835), .ZN(n8427) );
  AND3_X1 U9995 ( .A1(n8419), .A2(n8418), .A3(n8417), .ZN(n8420) );
  OAI21_X1 U9996 ( .B1(n8421), .B2(n8420), .A(n9742), .ZN(n8426) );
  AOI22_X1 U9997 ( .A1(n8639), .A2(n9737), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8422) );
  OAI21_X1 U9998 ( .B1(n8423), .B2(n9734), .A(n8422), .ZN(n8424) );
  AOI21_X1 U9999 ( .B1(n8620), .B2(n8434), .A(n8424), .ZN(n8425) );
  OAI211_X1 U10000 ( .C1(n8427), .C2(n8438), .A(n8426), .B(n8425), .ZN(
        P2_U3180) );
  OAI211_X1 U10001 ( .C1(n8430), .C2(n8429), .A(n8428), .B(n9742), .ZN(n8437)
         );
  AND2_X1 U10002 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8499) );
  AOI21_X1 U10003 ( .B1(n9737), .B2(n8443), .A(n8499), .ZN(n8431) );
  OAI21_X1 U10004 ( .B1(n8432), .B2(n9734), .A(n8431), .ZN(n8433) );
  AOI21_X1 U10005 ( .B1(n8435), .B2(n8434), .A(n8433), .ZN(n8436) );
  OAI211_X1 U10006 ( .C1(n8439), .C2(n8438), .A(n8437), .B(n8436), .ZN(
        P2_U3181) );
  MUX2_X1 U10007 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8572), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10008 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8440), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10009 ( .A(n8441), .ZN(n8592) );
  MUX2_X1 U10010 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8592), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10011 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8607), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10012 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8617), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10013 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8629), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10014 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8639), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10015 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8653), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10016 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8682), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10017 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8693), .S(n8455), .Z(
        P2_U3512) );
  MUX2_X1 U10018 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8681), .S(n8455), .Z(
        P2_U3511) );
  MUX2_X1 U10019 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8721), .S(n8455), .Z(
        P2_U3510) );
  MUX2_X1 U10020 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8738), .S(n8455), .Z(
        P2_U3509) );
  MUX2_X1 U10021 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8720), .S(n8455), .Z(
        P2_U3508) );
  MUX2_X1 U10022 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8740), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10023 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8442), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10024 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8443), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10025 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9736), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10026 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8444), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10027 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8445), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8446), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8447), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10030 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8448), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10031 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8449), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8450), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10033 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8451), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8452), .S(n8455), .Z(
        P2_U3495) );
  MUX2_X1 U10035 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8453), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10036 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8454), .S(n8455), .Z(
        P2_U3493) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8456), .S(n8455), .Z(
        P2_U3492) );
  AOI21_X1 U10038 ( .B1(n9752), .B2(n8458), .A(n8457), .ZN(n8474) );
  AOI21_X1 U10039 ( .B1(n8460), .B2(n8958), .A(n8459), .ZN(n8461) );
  OR2_X1 U10040 ( .A1(n8565), .A2(n8461), .ZN(n8464) );
  INV_X1 U10041 ( .A(n8462), .ZN(n8463) );
  OAI211_X1 U10042 ( .C1(n8465), .C2(n8561), .A(n8464), .B(n8463), .ZN(n8466)
         );
  AOI21_X1 U10043 ( .B1(n8467), .B2(n8553), .A(n8466), .ZN(n8473) );
  OAI21_X1 U10044 ( .B1(n8470), .B2(n8469), .A(n8468), .ZN(n8471) );
  NAND2_X1 U10045 ( .A1(n8471), .A2(n9981), .ZN(n8472) );
  OAI211_X1 U10046 ( .C1(n8474), .C2(n8559), .A(n8473), .B(n8472), .ZN(
        P2_U3195) );
  AOI21_X1 U10047 ( .B1(n8477), .B2(n8476), .A(n8475), .ZN(n8493) );
  OAI21_X1 U10048 ( .B1(n8480), .B2(n8479), .A(n8478), .ZN(n8491) );
  INV_X1 U10049 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U10050 ( .A1(n8553), .A2(n8481), .ZN(n8483) );
  NAND2_X1 U10051 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9732) );
  OAI211_X1 U10052 ( .C1(n8561), .C2(n8484), .A(n8483), .B(n9732), .ZN(n8490)
         );
  AOI21_X1 U10053 ( .B1(n8487), .B2(n8486), .A(n8485), .ZN(n8488) );
  NOR2_X1 U10054 ( .A1(n8488), .A2(n8565), .ZN(n8489) );
  AOI211_X1 U10055 ( .C1(n9981), .C2(n8491), .A(n8490), .B(n8489), .ZN(n8492)
         );
  OAI21_X1 U10056 ( .B1(n8493), .B2(n8559), .A(n8492), .ZN(P2_U3196) );
  AOI21_X1 U10057 ( .B1(n8495), .B2(n8917), .A(n8494), .ZN(n8512) );
  AOI21_X1 U10058 ( .B1(n8498), .B2(n8497), .A(n8496), .ZN(n8509) );
  INV_X1 U10059 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8968) );
  INV_X1 U10060 ( .A(n8499), .ZN(n8500) );
  OAI21_X1 U10061 ( .B1(n8561), .B2(n8968), .A(n8500), .ZN(n8501) );
  AOI21_X1 U10062 ( .B1(n8502), .B2(n8553), .A(n8501), .ZN(n8508) );
  OAI21_X1 U10063 ( .B1(n8505), .B2(n8504), .A(n8503), .ZN(n8506) );
  NAND2_X1 U10064 ( .A1(n8506), .A2(n9981), .ZN(n8507) );
  OAI211_X1 U10065 ( .C1(n8509), .C2(n8559), .A(n8508), .B(n8507), .ZN(n8510)
         );
  INV_X1 U10066 ( .A(n8510), .ZN(n8511) );
  OAI21_X1 U10067 ( .B1(n8512), .B2(n8565), .A(n8511), .ZN(P2_U3197) );
  AOI21_X1 U10068 ( .B1(n8515), .B2(n8514), .A(n8513), .ZN(n8531) );
  OAI21_X1 U10069 ( .B1(n8518), .B2(n8517), .A(n8516), .ZN(n8529) );
  INV_X1 U10070 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U10071 ( .A1(n8553), .A2(n8519), .ZN(n8522) );
  INV_X1 U10072 ( .A(n8520), .ZN(n8521) );
  OAI211_X1 U10073 ( .C1(n8523), .C2(n8561), .A(n8522), .B(n8521), .ZN(n8528)
         );
  AOI21_X1 U10074 ( .B1(n4330), .B2(n8525), .A(n8524), .ZN(n8526) );
  NOR2_X1 U10075 ( .A1(n8526), .A2(n8565), .ZN(n8527) );
  AOI211_X1 U10076 ( .C1(n9981), .C2(n8529), .A(n8528), .B(n8527), .ZN(n8530)
         );
  OAI21_X1 U10077 ( .B1(n8531), .B2(n8559), .A(n8530), .ZN(P2_U3198) );
  AOI21_X1 U10078 ( .B1(n8533), .B2(n8805), .A(n8532), .ZN(n8550) );
  NOR2_X1 U10079 ( .A1(n8561), .A2(n8534), .ZN(n8542) );
  AOI21_X1 U10080 ( .B1(n8537), .B2(n8536), .A(n8535), .ZN(n8540) );
  INV_X1 U10081 ( .A(n8538), .ZN(n8539) );
  OAI21_X1 U10082 ( .B1(n8540), .B2(n8565), .A(n8539), .ZN(n8541) );
  AOI211_X1 U10083 ( .C1(n8553), .C2(n8543), .A(n8542), .B(n8541), .ZN(n8549)
         );
  OAI21_X1 U10084 ( .B1(n8546), .B2(n8545), .A(n8544), .ZN(n8547) );
  NAND2_X1 U10085 ( .A1(n8547), .A2(n9981), .ZN(n8548) );
  OAI211_X1 U10086 ( .C1(n8550), .C2(n8559), .A(n8549), .B(n8548), .ZN(
        P2_U3199) );
  AOI21_X1 U10087 ( .B1(n8554), .B2(P2_U3893), .A(n8553), .ZN(n8570) );
  AOI21_X1 U10088 ( .B1(n4326), .B2(n8556), .A(n8555), .ZN(n8560) );
  NAND3_X1 U10089 ( .A1(n8557), .A2(n9981), .A3(n8569), .ZN(n8558) );
  OAI21_X1 U10090 ( .B1(n8560), .B2(n8559), .A(n8558), .ZN(n8568) );
  INV_X1 U10091 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10116) );
  NOR2_X1 U10092 ( .A1(n8561), .A2(n10116), .ZN(n8566) );
  AND2_X1 U10093 ( .A1(n8572), .A2(n8571), .ZN(n8815) );
  NOR2_X1 U10094 ( .A1(n8573), .A2(n8642), .ZN(n8581) );
  AOI21_X1 U10095 ( .B1(n8815), .B2(n8715), .A(n8581), .ZN(n8577) );
  NAND2_X1 U10096 ( .A1(n7496), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8574) );
  OAI211_X1 U10097 ( .C1(n8576), .C2(n8575), .A(n8577), .B(n8574), .ZN(
        P2_U3202) );
  NAND2_X1 U10098 ( .A1(n8818), .A2(n8762), .ZN(n8578) );
  OAI211_X1 U10099 ( .C1(n8723), .C2(n8986), .A(n8578), .B(n8577), .ZN(
        P2_U3203) );
  NAND2_X1 U10100 ( .A1(n8579), .A2(n8715), .ZN(n8585) );
  NOR2_X1 U10101 ( .A1(n8723), .A2(n8580), .ZN(n8582) );
  AOI211_X1 U10102 ( .C1(n8583), .C2(n8762), .A(n8582), .B(n8581), .ZN(n8584)
         );
  OAI211_X1 U10103 ( .C1(n8587), .C2(n8586), .A(n8585), .B(n8584), .ZN(
        P2_U3204) );
  XNOR2_X1 U10104 ( .A(n8589), .B(n8588), .ZN(n8826) );
  INV_X1 U10105 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8597) );
  XNOR2_X1 U10106 ( .A(n8591), .B(n8590), .ZN(n8596) );
  NAND2_X1 U10107 ( .A1(n8617), .A2(n8739), .ZN(n8593) );
  MUX2_X1 U10108 ( .A(n8597), .B(n8822), .S(n8723), .Z(n8600) );
  AOI22_X1 U10109 ( .A1(n8823), .A2(n8762), .B1(n8761), .B2(n8598), .ZN(n8599)
         );
  OAI211_X1 U10110 ( .C1(n8826), .C2(n8765), .A(n8600), .B(n8599), .ZN(
        P2_U3205) );
  XNOR2_X1 U10111 ( .A(n8602), .B(n8601), .ZN(n8832) );
  OAI21_X1 U10112 ( .B1(n8604), .B2(n8603), .A(n8752), .ZN(n8606) );
  OR2_X1 U10113 ( .A1(n8606), .A2(n8605), .ZN(n8609) );
  AOI22_X1 U10114 ( .A1(n8607), .A2(n8737), .B1(n8739), .B2(n8629), .ZN(n8608)
         );
  MUX2_X1 U10115 ( .A(n8610), .B(n8828), .S(n8723), .Z(n8613) );
  AOI22_X1 U10116 ( .A1(n8829), .A2(n8762), .B1(n8761), .B2(n8611), .ZN(n8612)
         );
  OAI211_X1 U10117 ( .C1(n8832), .C2(n8765), .A(n8613), .B(n8612), .ZN(
        P2_U3206) );
  XNOR2_X1 U10118 ( .A(n8614), .B(n8615), .ZN(n8838) );
  XOR2_X1 U10119 ( .A(n8616), .B(n8615), .Z(n8618) );
  AOI222_X1 U10120 ( .A1(n8752), .A2(n8618), .B1(n8617), .B2(n8737), .C1(n8639), .C2(n8739), .ZN(n8833) );
  MUX2_X1 U10121 ( .A(n8619), .B(n8833), .S(n8723), .Z(n8622) );
  AOI22_X1 U10122 ( .A1(n8835), .A2(n8762), .B1(n8761), .B2(n8620), .ZN(n8621)
         );
  OAI211_X1 U10123 ( .C1(n8838), .C2(n8765), .A(n8622), .B(n8621), .ZN(
        P2_U3207) );
  XNOR2_X1 U10124 ( .A(n8623), .B(n8625), .ZN(n8844) );
  INV_X1 U10125 ( .A(n8624), .ZN(n8628) );
  INV_X1 U10126 ( .A(n8625), .ZN(n8627) );
  OAI21_X1 U10127 ( .B1(n8628), .B2(n8627), .A(n8626), .ZN(n8630) );
  AOI222_X1 U10128 ( .A1(n8752), .A2(n8630), .B1(n8653), .B2(n8739), .C1(n8629), .C2(n8737), .ZN(n8839) );
  INV_X1 U10129 ( .A(n8644), .ZN(n8632) );
  AOI22_X1 U10130 ( .A1(n8841), .A2(n8632), .B1(n8761), .B2(n8631), .ZN(n8633)
         );
  AOI21_X1 U10131 ( .B1(n8839), .B2(n8633), .A(n7496), .ZN(n8634) );
  AOI21_X1 U10132 ( .B1(n7496), .B2(P2_REG2_REG_25__SCAN_IN), .A(n8634), .ZN(
        n8635) );
  OAI21_X1 U10133 ( .B1(n8844), .B2(n8765), .A(n8635), .ZN(P2_U3208) );
  XOR2_X1 U10134 ( .A(n8636), .B(n8638), .Z(n8850) );
  XOR2_X1 U10135 ( .A(n8638), .B(n8637), .Z(n8640) );
  AOI222_X1 U10136 ( .A1(n8752), .A2(n8640), .B1(n8639), .B2(n8737), .C1(n8665), .C2(n8739), .ZN(n8845) );
  INV_X1 U10137 ( .A(n8845), .ZN(n8647) );
  INV_X1 U10138 ( .A(n8641), .ZN(n8643) );
  OAI22_X1 U10139 ( .A1(n8645), .A2(n8644), .B1(n8643), .B2(n8642), .ZN(n8646)
         );
  OAI21_X1 U10140 ( .B1(n8647), .B2(n8646), .A(n8715), .ZN(n8649) );
  NAND2_X1 U10141 ( .A1(n7496), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8648) );
  OAI211_X1 U10142 ( .C1(n8850), .C2(n8765), .A(n8649), .B(n8648), .ZN(
        P2_U3209) );
  XOR2_X1 U10143 ( .A(n8650), .B(n8651), .Z(n8856) );
  XNOR2_X1 U10144 ( .A(n8652), .B(n8651), .ZN(n8654) );
  AOI222_X1 U10145 ( .A1(n8752), .A2(n8654), .B1(n8653), .B2(n8737), .C1(n8682), .C2(n8739), .ZN(n8851) );
  MUX2_X1 U10146 ( .A(n8655), .B(n8851), .S(n8723), .Z(n8658) );
  AOI22_X1 U10147 ( .A1(n8853), .A2(n8762), .B1(n8761), .B2(n8656), .ZN(n8657)
         );
  OAI211_X1 U10148 ( .C1(n8856), .C2(n8765), .A(n8658), .B(n8657), .ZN(
        P2_U3210) );
  OAI21_X1 U10149 ( .B1(n8661), .B2(n8660), .A(n8659), .ZN(n8791) );
  OAI21_X1 U10150 ( .B1(n8664), .B2(n8663), .A(n8662), .ZN(n8666) );
  AOI222_X1 U10151 ( .A1(n8752), .A2(n8666), .B1(n8693), .B2(n8739), .C1(n8665), .C2(n8737), .ZN(n8790) );
  OR2_X1 U10152 ( .A1(n8790), .A2(n7496), .ZN(n8672) );
  NAND2_X1 U10153 ( .A1(n8667), .A2(n8761), .ZN(n8668) );
  OAI21_X1 U10154 ( .B1(n8723), .B2(n8669), .A(n8668), .ZN(n8670) );
  AOI21_X1 U10155 ( .B1(n8788), .B2(n8762), .A(n8670), .ZN(n8671) );
  OAI211_X1 U10156 ( .C1(n8791), .C2(n8765), .A(n8672), .B(n8671), .ZN(
        P2_U3211) );
  NAND2_X1 U10157 ( .A1(n8674), .A2(n8673), .ZN(n8675) );
  XNOR2_X1 U10158 ( .A(n8675), .B(n8676), .ZN(n8999) );
  INV_X1 U10159 ( .A(n8676), .ZN(n8678) );
  NAND3_X1 U10160 ( .A1(n4303), .A2(n8678), .A3(n8677), .ZN(n8679) );
  NAND2_X1 U10161 ( .A1(n8680), .A2(n8679), .ZN(n8683) );
  AOI222_X1 U10162 ( .A1(n8752), .A2(n8683), .B1(n8682), .B2(n8737), .C1(n8681), .C2(n8739), .ZN(n8994) );
  MUX2_X1 U10163 ( .A(n8684), .B(n8994), .S(n8723), .Z(n8687) );
  AOI22_X1 U10164 ( .A1(n8996), .A2(n8762), .B1(n8685), .B2(n8761), .ZN(n8686)
         );
  OAI211_X1 U10165 ( .C1(n8999), .C2(n8765), .A(n8687), .B(n8686), .ZN(
        P2_U3212) );
  XNOR2_X1 U10166 ( .A(n8688), .B(n8690), .ZN(n9005) );
  INV_X1 U10167 ( .A(n8689), .ZN(n8692) );
  INV_X1 U10168 ( .A(n8690), .ZN(n8691) );
  OAI21_X1 U10169 ( .B1(n8692), .B2(n8691), .A(n4303), .ZN(n8694) );
  AOI222_X1 U10170 ( .A1(n8752), .A2(n8694), .B1(n8693), .B2(n8737), .C1(n8721), .C2(n8739), .ZN(n9000) );
  MUX2_X1 U10171 ( .A(n8695), .B(n9000), .S(n8723), .Z(n8698) );
  AOI22_X1 U10172 ( .A1(n9002), .A2(n8762), .B1(n8761), .B2(n8696), .ZN(n8697)
         );
  OAI211_X1 U10173 ( .C1(n9005), .C2(n8765), .A(n8698), .B(n8697), .ZN(
        P2_U3213) );
  NAND2_X1 U10174 ( .A1(n8719), .A2(n8699), .ZN(n8701) );
  NAND2_X1 U10175 ( .A1(n8701), .A2(n8700), .ZN(n8703) );
  XNOR2_X1 U10176 ( .A(n8703), .B(n8702), .ZN(n8704) );
  OAI222_X1 U10177 ( .A1(n8754), .A2(n8706), .B1(n8753), .B2(n8705), .C1(n8704), .C2(n10004), .ZN(n8798) );
  OR2_X1 U10178 ( .A1(n8708), .A2(n8707), .ZN(n8710) );
  NAND2_X1 U10179 ( .A1(n8710), .A2(n8709), .ZN(n9009) );
  AOI22_X1 U10180 ( .A1(n7496), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8761), .B2(
        n8711), .ZN(n8713) );
  NAND2_X1 U10181 ( .A1(n8799), .A2(n8762), .ZN(n8712) );
  OAI211_X1 U10182 ( .C1(n9009), .C2(n8765), .A(n8713), .B(n8712), .ZN(n8714)
         );
  AOI21_X1 U10183 ( .B1(n8798), .B2(n8715), .A(n8714), .ZN(n8716) );
  INV_X1 U10184 ( .A(n8716), .ZN(P2_U3214) );
  OAI21_X1 U10185 ( .B1(n4352), .B2(n8718), .A(n8717), .ZN(n9015) );
  XNOR2_X1 U10186 ( .A(n8719), .B(n8718), .ZN(n8722) );
  AOI222_X1 U10187 ( .A1(n8752), .A2(n8722), .B1(n8721), .B2(n8737), .C1(n8720), .C2(n8739), .ZN(n9010) );
  MUX2_X1 U10188 ( .A(n8724), .B(n9010), .S(n8723), .Z(n8727) );
  AOI22_X1 U10189 ( .A1(n9012), .A2(n8762), .B1(n8725), .B2(n8761), .ZN(n8726)
         );
  OAI211_X1 U10190 ( .C1(n9015), .C2(n8765), .A(n8727), .B(n8726), .ZN(
        P2_U3215) );
  INV_X1 U10191 ( .A(n8728), .ZN(n8729) );
  AOI21_X1 U10192 ( .B1(n8731), .B2(n8730), .A(n8729), .ZN(n9021) );
  AOI22_X1 U10193 ( .A1(n9018), .A2(n8762), .B1(n8761), .B2(n8732), .ZN(n8744)
         );
  NAND3_X1 U10194 ( .A1(n8733), .A2(n4838), .A3(n8734), .ZN(n8735) );
  NAND3_X1 U10195 ( .A1(n8736), .A2(n8752), .A3(n8735), .ZN(n8742) );
  AOI22_X1 U10196 ( .A1(n8740), .A2(n8739), .B1(n8738), .B2(n8737), .ZN(n8741)
         );
  AND2_X1 U10197 ( .A1(n8742), .A2(n8741), .ZN(n9017) );
  MUX2_X1 U10198 ( .A(n9017), .B(n8537), .S(n7496), .Z(n8743) );
  OAI211_X1 U10199 ( .C1(n9021), .C2(n8765), .A(n8744), .B(n8743), .ZN(
        P2_U3216) );
  OR2_X1 U10200 ( .A1(n8745), .A2(n8749), .ZN(n8746) );
  NAND2_X1 U10201 ( .A1(n8747), .A2(n8746), .ZN(n9026) );
  NAND3_X1 U10202 ( .A1(n8750), .A2(n8749), .A3(n8748), .ZN(n8751) );
  NAND3_X1 U10203 ( .A1(n8733), .A2(n8752), .A3(n8751), .ZN(n8758) );
  OAI22_X1 U10204 ( .A1(n8755), .A2(n8754), .B1(n9733), .B2(n8753), .ZN(n8756)
         );
  INV_X1 U10205 ( .A(n8756), .ZN(n8757) );
  NAND2_X1 U10206 ( .A1(n8758), .A2(n8757), .ZN(n9022) );
  MUX2_X1 U10207 ( .A(n9022), .B(P2_REG2_REG_16__SCAN_IN), .S(n7496), .Z(n8759) );
  INV_X1 U10208 ( .A(n8759), .ZN(n8764) );
  AOI22_X1 U10209 ( .A1(n8809), .A2(n8762), .B1(n8761), .B2(n8760), .ZN(n8763)
         );
  OAI211_X1 U10210 ( .C1(n9026), .C2(n8765), .A(n8764), .B(n8763), .ZN(
        P2_U3217) );
  INV_X1 U10211 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8767) );
  INV_X1 U10212 ( .A(n8810), .ZN(n8806) );
  NAND2_X1 U10213 ( .A1(n8814), .A2(n8806), .ZN(n8766) );
  NAND2_X1 U10214 ( .A1(n8815), .A2(n10107), .ZN(n8768) );
  OAI211_X1 U10215 ( .C1(n10107), .C2(n8767), .A(n8766), .B(n8768), .ZN(
        P2_U3490) );
  INV_X1 U10216 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8770) );
  NAND2_X1 U10217 ( .A1(n8818), .A2(n8806), .ZN(n8769) );
  OAI211_X1 U10218 ( .C1(n10107), .C2(n8770), .A(n8769), .B(n8768), .ZN(
        P2_U3489) );
  NAND2_X1 U10219 ( .A1(n8823), .A2(n8806), .ZN(n8772) );
  OAI211_X1 U10220 ( .C1(n8826), .C2(n8811), .A(n8773), .B(n8772), .ZN(
        P2_U3487) );
  INV_X1 U10221 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8774) );
  MUX2_X1 U10222 ( .A(n8774), .B(n8828), .S(n10107), .Z(n8776) );
  NAND2_X1 U10223 ( .A1(n8829), .A2(n8806), .ZN(n8775) );
  OAI211_X1 U10224 ( .C1(n8811), .C2(n8832), .A(n8776), .B(n8775), .ZN(
        P2_U3486) );
  INV_X1 U10225 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8777) );
  MUX2_X1 U10226 ( .A(n8777), .B(n8833), .S(n10107), .Z(n8779) );
  NAND2_X1 U10227 ( .A1(n8835), .A2(n8806), .ZN(n8778) );
  OAI211_X1 U10228 ( .C1(n8838), .C2(n8811), .A(n8779), .B(n8778), .ZN(
        P2_U3485) );
  INV_X1 U10229 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8780) );
  MUX2_X1 U10230 ( .A(n8780), .B(n8839), .S(n10107), .Z(n8782) );
  NAND2_X1 U10231 ( .A1(n8841), .A2(n8806), .ZN(n8781) );
  OAI211_X1 U10232 ( .C1(n8844), .C2(n8811), .A(n8782), .B(n8781), .ZN(
        P2_U3484) );
  MUX2_X1 U10233 ( .A(n8899), .B(n8845), .S(n10107), .Z(n8784) );
  NAND2_X1 U10234 ( .A1(n8847), .A2(n8806), .ZN(n8783) );
  OAI211_X1 U10235 ( .C1(n8811), .C2(n8850), .A(n8784), .B(n8783), .ZN(
        P2_U3483) );
  INV_X1 U10236 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8785) );
  MUX2_X1 U10237 ( .A(n8785), .B(n8851), .S(n10107), .Z(n8787) );
  NAND2_X1 U10238 ( .A1(n8853), .A2(n8806), .ZN(n8786) );
  OAI211_X1 U10239 ( .C1(n8856), .C2(n8811), .A(n8787), .B(n8786), .ZN(
        P2_U3482) );
  NAND2_X1 U10240 ( .A1(n8788), .A2(n10062), .ZN(n8789) );
  OAI211_X1 U10241 ( .C1(n10028), .C2(n8791), .A(n8790), .B(n8789), .ZN(n8857)
         );
  MUX2_X1 U10242 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8857), .S(n10107), .Z(
        P2_U3481) );
  INV_X1 U10243 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8792) );
  MUX2_X1 U10244 ( .A(n8792), .B(n8994), .S(n10107), .Z(n8794) );
  NAND2_X1 U10245 ( .A1(n8996), .A2(n8806), .ZN(n8793) );
  OAI211_X1 U10246 ( .C1(n8811), .C2(n8999), .A(n8794), .B(n8793), .ZN(
        P2_U3480) );
  INV_X1 U10247 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8795) );
  MUX2_X1 U10248 ( .A(n8795), .B(n9000), .S(n10107), .Z(n8797) );
  NAND2_X1 U10249 ( .A1(n9002), .A2(n8806), .ZN(n8796) );
  OAI211_X1 U10250 ( .C1(n9005), .C2(n8811), .A(n8797), .B(n8796), .ZN(
        P2_U3479) );
  INV_X1 U10251 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8800) );
  AOI21_X1 U10252 ( .B1(n10062), .B2(n8799), .A(n8798), .ZN(n9006) );
  MUX2_X1 U10253 ( .A(n8800), .B(n9006), .S(n10107), .Z(n8801) );
  OAI21_X1 U10254 ( .B1(n8811), .B2(n9009), .A(n8801), .ZN(P2_U3478) );
  MUX2_X1 U10255 ( .A(n8802), .B(n9010), .S(n10107), .Z(n8804) );
  NAND2_X1 U10256 ( .A1(n9012), .A2(n8806), .ZN(n8803) );
  OAI211_X1 U10257 ( .C1(n8811), .C2(n9015), .A(n8804), .B(n8803), .ZN(
        P2_U3477) );
  MUX2_X1 U10258 ( .A(n9017), .B(n8805), .S(n6337), .Z(n8808) );
  NAND2_X1 U10259 ( .A1(n9018), .A2(n8806), .ZN(n8807) );
  OAI211_X1 U10260 ( .C1(n9021), .C2(n8811), .A(n8808), .B(n8807), .ZN(
        P2_U3476) );
  MUX2_X1 U10261 ( .A(n9022), .B(P2_REG1_REG_16__SCAN_IN), .S(n6337), .Z(n8813) );
  INV_X1 U10262 ( .A(n8809), .ZN(n9024) );
  OAI22_X1 U10263 ( .A1(n9026), .A2(n8811), .B1(n9024), .B2(n8810), .ZN(n8812)
         );
  OR2_X1 U10264 ( .A1(n8813), .A2(n8812), .ZN(P2_U3475) );
  INV_X1 U10265 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U10266 ( .A1(n8814), .A2(n6352), .ZN(n8816) );
  NAND2_X1 U10267 ( .A1(n8815), .A2(n10080), .ZN(n8819) );
  OAI211_X1 U10268 ( .C1(n8817), .C2(n10080), .A(n8816), .B(n8819), .ZN(
        P2_U3458) );
  INV_X1 U10269 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U10270 ( .A1(n8818), .A2(n6352), .ZN(n8820) );
  OAI211_X1 U10271 ( .C1(n8821), .C2(n10080), .A(n8820), .B(n8819), .ZN(
        P2_U3457) );
  MUX2_X1 U10272 ( .A(n8970), .B(n8822), .S(n10080), .Z(n8825) );
  NAND2_X1 U10273 ( .A1(n8823), .A2(n6352), .ZN(n8824) );
  OAI211_X1 U10274 ( .C1(n8826), .C2(n9025), .A(n8825), .B(n8824), .ZN(
        P2_U3455) );
  INV_X1 U10275 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8827) );
  MUX2_X1 U10276 ( .A(n8828), .B(n8827), .S(n10078), .Z(n8831) );
  NAND2_X1 U10277 ( .A1(n8829), .A2(n6352), .ZN(n8830) );
  OAI211_X1 U10278 ( .C1(n8832), .C2(n9025), .A(n8831), .B(n8830), .ZN(
        P2_U3454) );
  INV_X1 U10279 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8834) );
  MUX2_X1 U10280 ( .A(n8834), .B(n8833), .S(n10080), .Z(n8837) );
  NAND2_X1 U10281 ( .A1(n8835), .A2(n6352), .ZN(n8836) );
  OAI211_X1 U10282 ( .C1(n8838), .C2(n9025), .A(n8837), .B(n8836), .ZN(
        P2_U3453) );
  INV_X1 U10283 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8840) );
  MUX2_X1 U10284 ( .A(n8840), .B(n8839), .S(n10080), .Z(n8843) );
  NAND2_X1 U10285 ( .A1(n8841), .A2(n6352), .ZN(n8842) );
  OAI211_X1 U10286 ( .C1(n8844), .C2(n9025), .A(n8843), .B(n8842), .ZN(
        P2_U3452) );
  INV_X1 U10287 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8846) );
  MUX2_X1 U10288 ( .A(n8846), .B(n8845), .S(n10080), .Z(n8849) );
  NAND2_X1 U10289 ( .A1(n8847), .A2(n6352), .ZN(n8848) );
  OAI211_X1 U10290 ( .C1(n8850), .C2(n9025), .A(n8849), .B(n8848), .ZN(
        P2_U3451) );
  INV_X1 U10291 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8852) );
  MUX2_X1 U10292 ( .A(n8852), .B(n8851), .S(n10080), .Z(n8855) );
  NAND2_X1 U10293 ( .A1(n8853), .A2(n6352), .ZN(n8854) );
  OAI211_X1 U10294 ( .C1(n8856), .C2(n9025), .A(n8855), .B(n8854), .ZN(
        P2_U3450) );
  MUX2_X1 U10295 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8857), .S(n10080), .Z(
        n8993) );
  AOI22_X1 U10296 ( .A1(n7214), .A2(keyinput16), .B1(n8859), .B2(keyinput25), 
        .ZN(n8858) );
  OAI221_X1 U10297 ( .B1(n7214), .B2(keyinput16), .C1(n8859), .C2(keyinput25), 
        .A(n8858), .ZN(n8870) );
  AOI22_X1 U10298 ( .A1(n8958), .A2(keyinput4), .B1(n6004), .B2(keyinput31), 
        .ZN(n8860) );
  OAI221_X1 U10299 ( .B1(n8958), .B2(keyinput4), .C1(n6004), .C2(keyinput31), 
        .A(n8860), .ZN(n8869) );
  AOI22_X1 U10300 ( .A1(n7108), .A2(keyinput46), .B1(n8862), .B2(keyinput62), 
        .ZN(n8861) );
  OAI221_X1 U10301 ( .B1(n7108), .B2(keyinput46), .C1(n8862), .C2(keyinput62), 
        .A(n8861), .ZN(n8868) );
  XNOR2_X1 U10302 ( .A(keyinput37), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(n8866) );
  XNOR2_X1 U10303 ( .A(P2_D_REG_6__SCAN_IN), .B(keyinput49), .ZN(n8865) );
  XOR2_X1 U10304 ( .A(n7380), .B(keyinput11), .Z(n8864) );
  XOR2_X1 U10305 ( .A(n5486), .B(keyinput9), .Z(n8863) );
  NAND4_X1 U10306 ( .A1(n8866), .A2(n8865), .A3(n8864), .A4(n8863), .ZN(n8867)
         );
  NOR4_X1 U10307 ( .A1(n8870), .A2(n8869), .A3(n8868), .A4(n8867), .ZN(n8891)
         );
  OAI22_X1 U10308 ( .A1(n5826), .A2(keyinput39), .B1(n9664), .B2(keyinput33), 
        .ZN(n8871) );
  AOI221_X1 U10309 ( .B1(n5826), .B2(keyinput39), .C1(keyinput33), .C2(n9664), 
        .A(n8871), .ZN(n8890) );
  INV_X1 U10310 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9055) );
  AOI22_X1 U10311 ( .A1(n9586), .A2(keyinput15), .B1(n9055), .B2(keyinput32), 
        .ZN(n8872) );
  OAI221_X1 U10312 ( .B1(n9586), .B2(keyinput15), .C1(n9055), .C2(keyinput32), 
        .A(n8872), .ZN(n8888) );
  XNOR2_X1 U10313 ( .A(SI_0_), .B(keyinput3), .ZN(n8876) );
  XNOR2_X1 U10314 ( .A(SI_23_), .B(keyinput63), .ZN(n8875) );
  XNOR2_X1 U10315 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput59), .ZN(n8874) );
  XNOR2_X1 U10316 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput56), .ZN(n8873)
         );
  NAND4_X1 U10317 ( .A1(n8876), .A2(n8875), .A3(n8874), .A4(n8873), .ZN(n8887)
         );
  XNOR2_X1 U10318 ( .A(P1_REG0_REG_29__SCAN_IN), .B(keyinput24), .ZN(n8880) );
  XNOR2_X1 U10319 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput61), .ZN(n8879) );
  XNOR2_X1 U10320 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput14), .ZN(n8878) );
  XNOR2_X1 U10321 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput22), .ZN(n8877) );
  NAND4_X1 U10322 ( .A1(n8880), .A2(n8879), .A3(n8878), .A4(n8877), .ZN(n8886)
         );
  XNOR2_X1 U10323 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput40), .ZN(n8884) );
  XNOR2_X1 U10324 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput26), .ZN(n8883) );
  XNOR2_X1 U10325 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput13), .ZN(n8882) );
  XNOR2_X1 U10326 ( .A(P2_REG2_REG_30__SCAN_IN), .B(keyinput6), .ZN(n8881) );
  NAND4_X1 U10327 ( .A1(n8884), .A2(n8883), .A3(n8882), .A4(n8881), .ZN(n8885)
         );
  NOR4_X1 U10328 ( .A1(n8888), .A2(n8887), .A3(n8886), .A4(n8885), .ZN(n8889)
         );
  AND3_X1 U10329 ( .A1(n8891), .A2(n8890), .A3(n8889), .ZN(n8930) );
  AOI22_X1 U10330 ( .A1(n5748), .A2(keyinput52), .B1(keyinput44), .B2(n8597), 
        .ZN(n8892) );
  OAI221_X1 U10331 ( .B1(n5748), .B2(keyinput52), .C1(n8597), .C2(keyinput44), 
        .A(n8892), .ZN(n8903) );
  AOI22_X1 U10332 ( .A1(n8894), .A2(keyinput53), .B1(keyinput42), .B2(n9834), 
        .ZN(n8893) );
  OAI221_X1 U10333 ( .B1(n8894), .B2(keyinput53), .C1(n9834), .C2(keyinput42), 
        .A(n8893), .ZN(n8902) );
  INV_X1 U10334 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8896) );
  AOI22_X1 U10335 ( .A1(n4738), .A2(keyinput20), .B1(n8896), .B2(keyinput8), 
        .ZN(n8895) );
  OAI221_X1 U10336 ( .B1(n4738), .B2(keyinput20), .C1(n8896), .C2(keyinput8), 
        .A(n8895), .ZN(n8901) );
  INV_X1 U10337 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8898) );
  AOI22_X1 U10338 ( .A1(n8899), .A2(keyinput45), .B1(n8898), .B2(keyinput30), 
        .ZN(n8897) );
  OAI221_X1 U10339 ( .B1(n8899), .B2(keyinput45), .C1(n8898), .C2(keyinput30), 
        .A(n8897), .ZN(n8900) );
  NOR4_X1 U10340 ( .A1(n8903), .A2(n8902), .A3(n8901), .A4(n8900), .ZN(n8929)
         );
  INV_X1 U10341 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10030) );
  AOI22_X1 U10342 ( .A1(n8905), .A2(keyinput28), .B1(keyinput47), .B2(n10030), 
        .ZN(n8904) );
  OAI221_X1 U10343 ( .B1(n8905), .B2(keyinput28), .C1(n10030), .C2(keyinput47), 
        .A(n8904), .ZN(n8915) );
  AOI22_X1 U10344 ( .A1(n9533), .A2(keyinput48), .B1(keyinput1), .B2(n8907), 
        .ZN(n8906) );
  OAI221_X1 U10345 ( .B1(n9533), .B2(keyinput48), .C1(n8907), .C2(keyinput1), 
        .A(n8906), .ZN(n8914) );
  INV_X1 U10346 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9199) );
  AOI22_X1 U10347 ( .A1(n8909), .A2(keyinput54), .B1(keyinput36), .B2(n9199), 
        .ZN(n8908) );
  OAI221_X1 U10348 ( .B1(n8909), .B2(keyinput54), .C1(n9199), .C2(keyinput36), 
        .A(n8908), .ZN(n8913) );
  INV_X1 U10349 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8985) );
  INV_X1 U10350 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8911) );
  AOI22_X1 U10351 ( .A1(n8985), .A2(keyinput17), .B1(keyinput12), .B2(n8911), 
        .ZN(n8910) );
  OAI221_X1 U10352 ( .B1(n8985), .B2(keyinput17), .C1(n8911), .C2(keyinput12), 
        .A(n8910), .ZN(n8912) );
  NOR4_X1 U10353 ( .A1(n8915), .A2(n8914), .A3(n8913), .A4(n8912), .ZN(n8928)
         );
  AOI22_X1 U10354 ( .A1(n8918), .A2(keyinput7), .B1(keyinput50), .B2(n8917), 
        .ZN(n8916) );
  OAI221_X1 U10355 ( .B1(n8918), .B2(keyinput7), .C1(n8917), .C2(keyinput50), 
        .A(n8916), .ZN(n8926) );
  AOI22_X1 U10356 ( .A1(n8920), .A2(keyinput43), .B1(n10095), .B2(keyinput51), 
        .ZN(n8919) );
  OAI221_X1 U10357 ( .B1(n8920), .B2(keyinput43), .C1(n10095), .C2(keyinput51), 
        .A(n8919), .ZN(n8925) );
  INV_X1 U10358 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8921) );
  XNOR2_X1 U10359 ( .A(n8921), .B(keyinput60), .ZN(n8924) );
  XNOR2_X1 U10360 ( .A(n8922), .B(keyinput58), .ZN(n8923) );
  NOR4_X1 U10361 ( .A1(n8926), .A2(n8925), .A3(n8924), .A4(n8923), .ZN(n8927)
         );
  AND4_X1 U10362 ( .A1(n8930), .A2(n8929), .A3(n8928), .A4(n8927), .ZN(n8955)
         );
  AOI22_X1 U10363 ( .A1(n8933), .A2(keyinput35), .B1(keyinput2), .B2(n8932), 
        .ZN(n8931) );
  OAI221_X1 U10364 ( .B1(n8933), .B2(keyinput35), .C1(n8932), .C2(keyinput2), 
        .A(n8931), .ZN(n8942) );
  AOI22_X1 U10365 ( .A1(n8935), .A2(keyinput21), .B1(n10103), .B2(keyinput10), 
        .ZN(n8934) );
  OAI221_X1 U10366 ( .B1(n8935), .B2(keyinput21), .C1(n10103), .C2(keyinput10), 
        .A(n8934), .ZN(n8941) );
  AOI22_X1 U10367 ( .A1(n8937), .A2(keyinput38), .B1(keyinput27), .B2(n8981), 
        .ZN(n8936) );
  OAI221_X1 U10368 ( .B1(n8937), .B2(keyinput38), .C1(n8981), .C2(keyinput27), 
        .A(n8936), .ZN(n8940) );
  INV_X1 U10369 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9216) );
  AOI22_X1 U10370 ( .A1(n9857), .A2(keyinput19), .B1(keyinput5), .B2(n9216), 
        .ZN(n8938) );
  OAI221_X1 U10371 ( .B1(n9857), .B2(keyinput19), .C1(n9216), .C2(keyinput5), 
        .A(n8938), .ZN(n8939) );
  NOR4_X1 U10372 ( .A1(n8942), .A2(n8941), .A3(n8940), .A4(n8939), .ZN(n8954)
         );
  AOI22_X1 U10373 ( .A1(n8970), .A2(keyinput55), .B1(keyinput34), .B2(n9094), 
        .ZN(n8943) );
  OAI221_X1 U10374 ( .B1(n8970), .B2(keyinput55), .C1(n9094), .C2(keyinput34), 
        .A(n8943), .ZN(n8952) );
  INV_X1 U10375 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8945) );
  INV_X1 U10376 ( .A(SI_30_), .ZN(n8969) );
  AOI22_X1 U10377 ( .A1(n8945), .A2(keyinput41), .B1(keyinput23), .B2(n8969), 
        .ZN(n8944) );
  OAI221_X1 U10378 ( .B1(n8945), .B2(keyinput41), .C1(n8969), .C2(keyinput23), 
        .A(n8944), .ZN(n8951) );
  AOI22_X1 U10379 ( .A1(n8963), .A2(keyinput29), .B1(n8947), .B2(keyinput18), 
        .ZN(n8946) );
  OAI221_X1 U10380 ( .B1(n8963), .B2(keyinput29), .C1(n8947), .C2(keyinput18), 
        .A(n8946), .ZN(n8950) );
  INV_X1 U10381 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9939) );
  AOI22_X1 U10382 ( .A1(n9939), .A2(keyinput57), .B1(n8957), .B2(keyinput0), 
        .ZN(n8948) );
  OAI221_X1 U10383 ( .B1(n9939), .B2(keyinput57), .C1(n8957), .C2(keyinput0), 
        .A(n8948), .ZN(n8949) );
  NOR4_X1 U10384 ( .A1(n8952), .A2(n8951), .A3(n8950), .A4(n8949), .ZN(n8953)
         );
  NAND3_X1 U10385 ( .A1(n8955), .A2(n8954), .A3(n8953), .ZN(n8991) );
  NOR4_X1 U10386 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .A3(P2_ADDR_REG_19__SCAN_IN), .A4(SI_20_), .ZN(n8962) );
  NOR4_X1 U10387 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(SI_0_), .A3(n8957), .A4(
        n8956), .ZN(n8961) );
  NOR4_X1 U10388 ( .A1(P2_REG0_REG_16__SCAN_IN), .A2(P2_REG2_REG_16__SCAN_IN), 
        .A3(P2_REG2_REG_15__SCAN_IN), .A4(n8958), .ZN(n8960) );
  NOR4_X1 U10389 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(P2_REG1_REG_11__SCAN_IN), 
        .A3(P2_REG2_REG_10__SCAN_IN), .A4(P2_REG1_REG_7__SCAN_IN), .ZN(n8959)
         );
  NAND4_X1 U10390 ( .A1(n8962), .A2(n8961), .A3(n8960), .A4(n8959), .ZN(n8980)
         );
  NOR3_X1 U10391 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_15__SCAN_IN), .ZN(n8965) );
  NOR3_X1 U10392 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .A3(n8963), .ZN(n8964) );
  NAND4_X1 U10393 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        n8965), .A4(n8964), .ZN(n8979) );
  NOR4_X1 U10394 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .A3(P2_IR_REG_26__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8966) );
  NAND4_X1 U10395 ( .A1(n8967), .A2(P1_ADDR_REG_3__SCAN_IN), .A3(n8966), .A4(
        n9216), .ZN(n8978) );
  NAND4_X1 U10396 ( .A1(P1_REG0_REG_19__SCAN_IN), .A2(P1_DATAO_REG_25__SCAN_IN), .A3(P2_ADDR_REG_11__SCAN_IN), .A4(n8968), .ZN(n8976) );
  INV_X1 U10397 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n8972) );
  NOR4_X1 U10398 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .A3(n8970), .A4(n8969), .ZN(n8971) );
  NAND4_X1 U10399 ( .A1(n4975), .A2(n8911), .A3(n8972), .A4(n8971), .ZN(n8975)
         );
  NAND3_X1 U10400 ( .A1(SI_23_), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_REG3_REG_16__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U10401 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(P1_REG1_REG_22__SCAN_IN), 
        .ZN(n8973) );
  OR4_X1 U10402 ( .A1(n8976), .A2(n8975), .A3(n8974), .A4(n8973), .ZN(n8977)
         );
  NOR4_X1 U10403 ( .A1(n8980), .A2(n8979), .A3(n8978), .A4(n8977), .ZN(n8989)
         );
  NAND4_X1 U10404 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG1_REG_11__SCAN_IN), .A4(n8981), .ZN(n8984) );
  NAND3_X1 U10405 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(P2_REG1_REG_24__SCAN_IN), 
        .A3(P1_DATAO_REG_31__SCAN_IN), .ZN(n8983) );
  NAND4_X1 U10406 ( .A1(P1_REG0_REG_5__SCAN_IN), .A2(P1_REG3_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_12__SCAN_IN), .A4(n9533), .ZN(n8982) );
  NOR4_X1 U10407 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n8984), .A3(n8983), .A4(
        n8982), .ZN(n8988) );
  NOR4_X1 U10408 ( .A1(P2_REG0_REG_4__SCAN_IN), .A2(n8986), .A3(n8985), .A4(
        n7108), .ZN(n8987) );
  NAND3_X1 U10409 ( .A1(n8989), .A2(n8988), .A3(n8987), .ZN(n8990) );
  XNOR2_X1 U10410 ( .A(n8991), .B(n8990), .ZN(n8992) );
  XNOR2_X1 U10411 ( .A(n8993), .B(n8992), .ZN(P2_U3449) );
  INV_X1 U10412 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8995) );
  MUX2_X1 U10413 ( .A(n8995), .B(n8994), .S(n10080), .Z(n8998) );
  NAND2_X1 U10414 ( .A1(n8996), .A2(n6352), .ZN(n8997) );
  OAI211_X1 U10415 ( .C1(n8999), .C2(n9025), .A(n8998), .B(n8997), .ZN(
        P2_U3448) );
  INV_X1 U10416 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9001) );
  MUX2_X1 U10417 ( .A(n9001), .B(n9000), .S(n10080), .Z(n9004) );
  NAND2_X1 U10418 ( .A1(n9002), .A2(n6352), .ZN(n9003) );
  OAI211_X1 U10419 ( .C1(n9005), .C2(n9025), .A(n9004), .B(n9003), .ZN(
        P2_U3447) );
  INV_X1 U10420 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9007) );
  MUX2_X1 U10421 ( .A(n9007), .B(n9006), .S(n10080), .Z(n9008) );
  OAI21_X1 U10422 ( .B1(n9009), .B2(n9025), .A(n9008), .ZN(P2_U3446) );
  INV_X1 U10423 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9011) );
  MUX2_X1 U10424 ( .A(n9011), .B(n9010), .S(n10080), .Z(n9014) );
  NAND2_X1 U10425 ( .A1(n9012), .A2(n6352), .ZN(n9013) );
  OAI211_X1 U10426 ( .C1(n9015), .C2(n9025), .A(n9014), .B(n9013), .ZN(
        P2_U3444) );
  INV_X1 U10427 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9016) );
  MUX2_X1 U10428 ( .A(n9017), .B(n9016), .S(n10078), .Z(n9020) );
  NAND2_X1 U10429 ( .A1(n9018), .A2(n6352), .ZN(n9019) );
  OAI211_X1 U10430 ( .C1(n9021), .C2(n9025), .A(n9020), .B(n9019), .ZN(
        P2_U3441) );
  MUX2_X1 U10431 ( .A(n9022), .B(P2_REG0_REG_16__SCAN_IN), .S(n10078), .Z(
        n9028) );
  OAI22_X1 U10432 ( .A1(n9026), .A2(n9025), .B1(n9024), .B2(n9023), .ZN(n9027)
         );
  OR2_X1 U10433 ( .A1(n9028), .A2(n9027), .ZN(P2_U3438) );
  INV_X1 U10434 ( .A(n9029), .ZN(n9695) );
  NAND3_X1 U10435 ( .A1(n5957), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9031) );
  OAI22_X1 U10436 ( .A1(n9032), .A2(n9031), .B1(n8894), .B2(n9030), .ZN(n9033)
         );
  INV_X1 U10437 ( .A(n9033), .ZN(n9034) );
  OAI21_X1 U10438 ( .B1(n9695), .B2(n9035), .A(n9034), .ZN(P2_U3264) );
  MUX2_X1 U10439 ( .A(n9036), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10440 ( .A1(n4780), .A2(n9037), .ZN(n9039) );
  XNOR2_X1 U10441 ( .A(n9039), .B(n9038), .ZN(n9046) );
  OAI22_X1 U10442 ( .A1(n9787), .A2(n9041), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9040), .ZN(n9043) );
  NOR2_X1 U10443 ( .A1(n9686), .A2(n9143), .ZN(n9042) );
  AOI211_X1 U10444 ( .C1(n9044), .C2(n9140), .A(n9043), .B(n9042), .ZN(n9045)
         );
  OAI21_X1 U10445 ( .B1(n9046), .B2(n9792), .A(n9045), .ZN(P1_U3215) );
  INV_X1 U10446 ( .A(n9047), .ZN(n9052) );
  NOR3_X1 U10447 ( .A1(n9048), .A2(n9050), .A3(n9049), .ZN(n9051) );
  OAI21_X1 U10448 ( .B1(n9052), .B2(n9051), .A(n9158), .ZN(n9058) );
  OR2_X1 U10449 ( .A1(n9172), .A2(n9161), .ZN(n9054) );
  INV_X1 U10450 ( .A(n9299), .ZN(n9298) );
  NAND2_X1 U10451 ( .A1(n9298), .A2(n9761), .ZN(n9053) );
  AND2_X1 U10452 ( .A1(n9054), .A2(n9053), .ZN(n9410) );
  OAI22_X1 U10453 ( .A1(n9410), .A2(n9787), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9055), .ZN(n9056) );
  AOI21_X1 U10454 ( .B1(n4888), .B2(n9140), .A(n9056), .ZN(n9057) );
  OAI211_X1 U10455 ( .C1(n9407), .C2(n9143), .A(n9058), .B(n9057), .ZN(
        P1_U3216) );
  NAND2_X1 U10456 ( .A1(n9135), .A2(n9059), .ZN(n9065) );
  XNOR2_X1 U10457 ( .A(n9060), .B(n9062), .ZN(n9152) );
  AOI22_X1 U10458 ( .A1(n9152), .A2(n9063), .B1(n9062), .B2(n9061), .ZN(n9064)
         );
  XOR2_X1 U10459 ( .A(n9065), .B(n9064), .Z(n9071) );
  OR2_X1 U10460 ( .A1(n9173), .A2(n9161), .ZN(n9067) );
  INV_X1 U10461 ( .A(n9287), .ZN(n9286) );
  NAND2_X1 U10462 ( .A1(n9286), .A2(n9761), .ZN(n9066) );
  NAND2_X1 U10463 ( .A1(n9067), .A2(n9066), .ZN(n9467) );
  AOI22_X1 U10464 ( .A1(n9467), .A2(n9164), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9068) );
  OAI21_X1 U10465 ( .B1(n9797), .B2(n9475), .A(n9068), .ZN(n9069) );
  AOI21_X1 U10466 ( .B1(n9474), .B2(n4282), .A(n9069), .ZN(n9070) );
  OAI21_X1 U10467 ( .B1(n9071), .B2(n9792), .A(n9070), .ZN(P1_U3219) );
  OAI21_X1 U10468 ( .B1(n9075), .B2(n9072), .A(n9074), .ZN(n9076) );
  NAND2_X1 U10469 ( .A1(n9076), .A2(n9158), .ZN(n9081) );
  NOR2_X1 U10470 ( .A1(n9173), .A2(n9163), .ZN(n9077) );
  AOI21_X1 U10471 ( .B1(n9298), .B2(n9758), .A(n9077), .ZN(n9441) );
  OAI22_X1 U10472 ( .A1(n9441), .A2(n9787), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9078), .ZN(n9079) );
  AOI21_X1 U10473 ( .B1(n9445), .B2(n9140), .A(n9079), .ZN(n9080) );
  OAI211_X1 U10474 ( .C1(n9295), .C2(n9143), .A(n9081), .B(n9080), .ZN(
        P1_U3223) );
  OAI21_X1 U10475 ( .B1(n9084), .B2(n9082), .A(n9083), .ZN(n9085) );
  NAND2_X1 U10476 ( .A1(n9085), .A2(n9158), .ZN(n9091) );
  OR2_X1 U10477 ( .A1(n9172), .A2(n9163), .ZN(n9087) );
  NAND2_X1 U10478 ( .A1(n9171), .A2(n9758), .ZN(n9086) );
  AND2_X1 U10479 ( .A1(n9087), .A2(n9086), .ZN(n9376) );
  INV_X1 U10480 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9088) );
  OAI22_X1 U10481 ( .A1(n9376), .A2(n9787), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9088), .ZN(n9089) );
  AOI21_X1 U10482 ( .B1(n9382), .B2(n9140), .A(n9089), .ZN(n9090) );
  OAI211_X1 U10483 ( .C1(n9649), .C2(n9143), .A(n9091), .B(n9090), .ZN(
        P1_U3225) );
  AOI21_X1 U10484 ( .B1(n9093), .B2(n9092), .A(n9101), .ZN(n9098) );
  OAI22_X1 U10485 ( .A1(n9284), .A2(n9161), .B1(n9279), .B2(n9163), .ZN(n9522)
         );
  NOR2_X1 U10486 ( .A1(n9094), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9868) );
  AOI21_X1 U10487 ( .B1(n9164), .B2(n9522), .A(n9868), .ZN(n9095) );
  OAI21_X1 U10488 ( .B1(n9797), .B2(n9532), .A(n9095), .ZN(n9096) );
  AOI21_X1 U10489 ( .B1(n9529), .B2(n4282), .A(n9096), .ZN(n9097) );
  OAI21_X1 U10490 ( .B1(n9098), .B2(n9792), .A(n9097), .ZN(P1_U3226) );
  OAI21_X1 U10491 ( .B1(n9101), .B2(n9100), .A(n9099), .ZN(n9102) );
  NAND3_X1 U10492 ( .A1(n4811), .A2(n9158), .A3(n9102), .ZN(n9107) );
  OAI22_X1 U10493 ( .A1(n9287), .A2(n9161), .B1(n9103), .B2(n9163), .ZN(n9104)
         );
  INV_X1 U10494 ( .A(n9104), .ZN(n9507) );
  NAND2_X1 U10495 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9886) );
  OAI21_X1 U10496 ( .B1(n9787), .B2(n9507), .A(n9886), .ZN(n9105) );
  AOI21_X1 U10497 ( .B1(n9140), .B2(n9513), .A(n9105), .ZN(n9106) );
  OAI211_X1 U10498 ( .C1(n9674), .C2(n9143), .A(n9107), .B(n9106), .ZN(
        P1_U3228) );
  OAI22_X1 U10499 ( .A1(n9307), .A2(n9161), .B1(n9301), .B2(n9163), .ZN(n9392)
         );
  AOI22_X1 U10500 ( .A1(n9392), .A2(n9164), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9108) );
  OAI21_X1 U10501 ( .B1(n9797), .B2(n9109), .A(n9108), .ZN(n9114) );
  INV_X1 U10502 ( .A(n9111), .ZN(n9112) );
  INV_X1 U10503 ( .A(n6874), .ZN(n9116) );
  NAND2_X1 U10504 ( .A1(n9116), .A2(n9115), .ZN(n9117) );
  XNOR2_X1 U10505 ( .A(n9117), .B(n9118), .ZN(n9784) );
  NOR2_X1 U10506 ( .A1(n9784), .A2(n9783), .ZN(n9782) );
  AOI21_X1 U10507 ( .B1(n9118), .B2(n9117), .A(n9782), .ZN(n9121) );
  OAI211_X1 U10508 ( .C1(n9121), .C2(n9120), .A(n9158), .B(n9119), .ZN(n9131)
         );
  NAND2_X1 U10509 ( .A1(n9123), .A2(n9122), .ZN(n9125) );
  NOR2_X1 U10510 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9124), .ZN(n9243) );
  AOI21_X1 U10511 ( .B1(n9164), .B2(n9125), .A(n9243), .ZN(n9130) );
  NAND2_X1 U10512 ( .A1(n4282), .A2(n5265), .ZN(n9129) );
  NAND2_X1 U10513 ( .A1(n9140), .A2(n9127), .ZN(n9128) );
  NAND4_X1 U10514 ( .A1(n9131), .A2(n9130), .A3(n9129), .A4(n9128), .ZN(
        P1_U3231) );
  INV_X1 U10515 ( .A(n9132), .ZN(n9137) );
  AOI21_X1 U10516 ( .B1(n9133), .B2(n9135), .A(n9134), .ZN(n9136) );
  OAI21_X1 U10517 ( .B1(n9137), .B2(n9136), .A(n9158), .ZN(n9142) );
  AOI22_X1 U10518 ( .A1(n9294), .A2(n9758), .B1(n9761), .B2(n9288), .ZN(n9452)
         );
  OAI22_X1 U10519 ( .A1(n9452), .A2(n9787), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9138), .ZN(n9139) );
  AOI21_X1 U10520 ( .B1(n9454), .B2(n9140), .A(n9139), .ZN(n9141) );
  OAI211_X1 U10521 ( .C1(n9662), .C2(n9143), .A(n9142), .B(n9141), .ZN(
        P1_U3233) );
  AOI21_X1 U10522 ( .B1(n9145), .B2(n9144), .A(n9048), .ZN(n9151) );
  OR2_X1 U10523 ( .A1(n9301), .A2(n9161), .ZN(n9147) );
  NAND2_X1 U10524 ( .A1(n9294), .A2(n9761), .ZN(n9146) );
  NAND2_X1 U10525 ( .A1(n9147), .A2(n9146), .ZN(n9420) );
  AOI22_X1 U10526 ( .A1(n9420), .A2(n9164), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9148) );
  OAI21_X1 U10527 ( .B1(n9797), .B2(n9425), .A(n9148), .ZN(n9149) );
  AOI21_X1 U10528 ( .B1(n9424), .B2(n4282), .A(n9149), .ZN(n9150) );
  OAI21_X1 U10529 ( .B1(n9151), .B2(n9792), .A(n9150), .ZN(P1_U3235) );
  XNOR2_X1 U10530 ( .A(n9152), .B(n4809), .ZN(n9156) );
  OAI22_X1 U10531 ( .A1(n9290), .A2(n9161), .B1(n9284), .B2(n9163), .ZN(n9488)
         );
  AOI22_X1 U10532 ( .A1(n9164), .A2(n9488), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9153) );
  OAI21_X1 U10533 ( .B1(n9797), .B2(n9494), .A(n9153), .ZN(n9154) );
  AOI21_X1 U10534 ( .B1(n9493), .B2(n4282), .A(n9154), .ZN(n9155) );
  OAI21_X1 U10535 ( .B1(n9156), .B2(n9792), .A(n9155), .ZN(P1_U3238) );
  NAND2_X1 U10536 ( .A1(n9157), .A2(n9158), .ZN(n9170) );
  AOI21_X1 U10537 ( .B1(n9083), .B2(n9160), .A(n9159), .ZN(n9169) );
  INV_X1 U10538 ( .A(n9361), .ZN(n9166) );
  OAI22_X1 U10539 ( .A1(n9307), .A2(n9163), .B1(n9162), .B2(n9161), .ZN(n9367)
         );
  AOI22_X1 U10540 ( .A1(n9367), .A2(n9164), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9165) );
  OAI21_X1 U10541 ( .B1(n9797), .B2(n9166), .A(n9165), .ZN(n9167) );
  AOI21_X1 U10542 ( .B1(n9563), .B2(n4282), .A(n9167), .ZN(n9168) );
  OAI21_X1 U10543 ( .B1(n9170), .B2(n9169), .A(n9168), .ZN(P1_U3240) );
  MUX2_X1 U10544 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9271), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10545 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9317), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10546 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9315), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10547 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9171), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10548 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9309), .S(P1_U3973), .Z(
        P1_U3579) );
  INV_X1 U10549 ( .A(n9172), .ZN(n9304) );
  MUX2_X1 U10550 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9304), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10551 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9298), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10552 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9294), .S(P1_U3973), .Z(
        P1_U3575) );
  INV_X1 U10553 ( .A(n9173), .ZN(n9291) );
  MUX2_X1 U10554 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9291), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10555 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9288), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10556 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9286), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10557 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9281), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10558 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9275), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10559 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9174), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10560 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9175), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10561 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9176), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10562 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9759), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10563 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9177), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10564 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9760), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10565 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9178), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10566 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9179), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10567 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9180), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10568 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9181), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10569 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9182), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10570 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9183), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10571 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9184), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10572 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9185), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10573 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9186), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10574 ( .C1(n9189), .C2(n9188), .A(n9884), .B(n9187), .ZN(n9197)
         );
  AND2_X1 U10575 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9191) );
  OAI211_X1 U10576 ( .C1(n9192), .C2(n9191), .A(n9892), .B(n9190), .ZN(n9196)
         );
  AOI22_X1 U10577 ( .A1(n9869), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9195) );
  NAND2_X1 U10578 ( .A1(n9881), .A2(n9193), .ZN(n9194) );
  NAND4_X1 U10579 ( .A1(n9197), .A2(n9196), .A3(n9195), .A4(n9194), .ZN(
        P1_U3244) );
  NAND2_X1 U10580 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9198) );
  OAI21_X1 U10581 ( .B1(n9904), .B2(n9199), .A(n9198), .ZN(n9200) );
  AOI21_X1 U10582 ( .B1(n9201), .B2(n9881), .A(n9200), .ZN(n9210) );
  OAI211_X1 U10583 ( .C1(n9204), .C2(n9203), .A(n9884), .B(n9202), .ZN(n9209)
         );
  OAI211_X1 U10584 ( .C1(n9207), .C2(n9206), .A(n9892), .B(n9205), .ZN(n9208)
         );
  NAND3_X1 U10585 ( .A1(n9210), .A2(n9209), .A3(n9208), .ZN(P1_U3246) );
  AOI211_X1 U10586 ( .C1(n9213), .C2(n9212), .A(n9211), .B(n9851), .ZN(n9214)
         );
  INV_X1 U10587 ( .A(n9214), .ZN(n9224) );
  NAND2_X1 U10588 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9215) );
  OAI21_X1 U10589 ( .B1(n9904), .B2(n9216), .A(n9215), .ZN(n9217) );
  AOI21_X1 U10590 ( .B1(n9218), .B2(n9881), .A(n9217), .ZN(n9223) );
  OAI211_X1 U10591 ( .C1(n9221), .C2(n9220), .A(n9884), .B(n9219), .ZN(n9222)
         );
  NAND3_X1 U10592 ( .A1(n9224), .A2(n9223), .A3(n9222), .ZN(P1_U3248) );
  AOI211_X1 U10593 ( .C1(n9227), .C2(n9226), .A(n9851), .B(n9225), .ZN(n9228)
         );
  INV_X1 U10594 ( .A(n9228), .ZN(n9238) );
  INV_X1 U10595 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U10596 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9229) );
  OAI21_X1 U10597 ( .B1(n9904), .B2(n9230), .A(n9229), .ZN(n9231) );
  AOI21_X1 U10598 ( .B1(n9232), .B2(n9881), .A(n9231), .ZN(n9237) );
  OAI211_X1 U10599 ( .C1(n9235), .C2(n9234), .A(n9884), .B(n9233), .ZN(n9236)
         );
  NAND3_X1 U10600 ( .A1(n9238), .A2(n9237), .A3(n9236), .ZN(P1_U3249) );
  OAI21_X1 U10601 ( .B1(n9241), .B2(n9240), .A(n9239), .ZN(n9242) );
  NAND2_X1 U10602 ( .A1(n9242), .A2(n9884), .ZN(n9252) );
  AOI21_X1 U10603 ( .B1(n9869), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9243), .ZN(
        n9251) );
  OAI21_X1 U10604 ( .B1(n9246), .B2(n9245), .A(n9244), .ZN(n9247) );
  NAND2_X1 U10605 ( .A1(n9247), .A2(n9892), .ZN(n9250) );
  NAND2_X1 U10606 ( .A1(n9881), .A2(n9248), .ZN(n9249) );
  NAND4_X1 U10607 ( .A1(n9252), .A2(n9251), .A3(n9250), .A4(n9249), .ZN(
        P1_U3252) );
  INV_X1 U10608 ( .A(n9253), .ZN(n9632) );
  XNOR2_X1 U10609 ( .A(n9254), .B(n9253), .ZN(n9255) );
  NAND2_X1 U10610 ( .A1(n9540), .A2(n9921), .ZN(n9258) );
  AOI21_X1 U10611 ( .B1(n9928), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9256), .ZN(
        n9257) );
  OAI211_X1 U10612 ( .C1(n9632), .C2(n9530), .A(n9258), .B(n9257), .ZN(
        P1_U3263) );
  NAND3_X1 U10613 ( .A1(n9434), .A2(n9435), .A3(n9433), .ZN(n9438) );
  INV_X1 U10614 ( .A(n9261), .ZN(n9263) );
  NAND3_X1 U10615 ( .A1(n9389), .A2(n9379), .A3(n9373), .ZN(n9372) );
  NAND2_X1 U10616 ( .A1(n9372), .A2(n9265), .ZN(n9365) );
  INV_X1 U10617 ( .A(n9356), .ZN(n9366) );
  NAND2_X1 U10618 ( .A1(n9365), .A2(n9366), .ZN(n9364) );
  NAND2_X1 U10619 ( .A1(n9364), .A2(n9266), .ZN(n9345) );
  NAND2_X1 U10620 ( .A1(n9345), .A2(n4676), .ZN(n9344) );
  INV_X1 U10621 ( .A(n9267), .ZN(n9269) );
  AOI22_X1 U10622 ( .A1(n9344), .A2(n9269), .B1(n9268), .B2(n9316), .ZN(n9270)
         );
  AOI22_X1 U10623 ( .A1(n9317), .A2(n9761), .B1(n9272), .B2(n9271), .ZN(n9273)
         );
  INV_X1 U10624 ( .A(n9474), .ZN(n9666) );
  NAND2_X1 U10625 ( .A1(n9276), .A2(n9279), .ZN(n9277) );
  NAND2_X1 U10626 ( .A1(n9280), .A2(n4874), .ZN(n9525) );
  AOI21_X2 U10627 ( .B1(n9525), .B2(n9283), .A(n9282), .ZN(n9501) );
  AOI21_X2 U10628 ( .B1(n9456), .B2(n9455), .A(n9292), .ZN(n9432) );
  NAND2_X1 U10629 ( .A1(n9432), .A2(n4872), .ZN(n9297) );
  NAND2_X1 U10630 ( .A1(n9297), .A2(n9296), .ZN(n9417) );
  NAND2_X1 U10631 ( .A1(n9424), .A2(n9298), .ZN(n9300) );
  AOI22_X2 U10632 ( .A1(n9417), .A2(n9300), .B1(n9299), .B2(n9655), .ZN(n9402)
         );
  NAND2_X1 U10633 ( .A1(n9407), .A2(n9301), .ZN(n9303) );
  NOR2_X1 U10634 ( .A1(n9407), .A2(n9301), .ZN(n9302) );
  AOI21_X2 U10635 ( .B1(n9402), .B2(n9303), .A(n9302), .ZN(n9388) );
  NAND2_X1 U10636 ( .A1(n9574), .A2(n9304), .ZN(n9306) );
  NOR2_X1 U10637 ( .A1(n9574), .A2(n9304), .ZN(n9305) );
  AOI21_X2 U10638 ( .B1(n9388), .B2(n9306), .A(n9305), .ZN(n9378) );
  NAND2_X1 U10639 ( .A1(n9649), .A2(n9307), .ZN(n9308) );
  NAND2_X1 U10640 ( .A1(n9378), .A2(n9308), .ZN(n9311) );
  NAND2_X1 U10641 ( .A1(n9381), .A2(n9309), .ZN(n9310) );
  NOR2_X1 U10642 ( .A1(n9363), .A2(n9312), .ZN(n9314) );
  NAND2_X1 U10643 ( .A1(n9363), .A2(n9312), .ZN(n9313) );
  XNOR2_X1 U10644 ( .A(n9319), .B(n9318), .ZN(n9547) );
  NAND2_X1 U10645 ( .A1(n9547), .A2(n9935), .ZN(n9327) );
  AOI21_X1 U10646 ( .B1(n9321), .B2(n9335), .A(n9320), .ZN(n9549) );
  AOI22_X1 U10647 ( .A1(n9928), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9322), .B2(
        n9927), .ZN(n9323) );
  OAI21_X1 U10648 ( .B1(n4461), .B2(n9530), .A(n9323), .ZN(n9324) );
  AOI21_X1 U10649 ( .B1(n9549), .B2(n9325), .A(n9324), .ZN(n9326) );
  OAI211_X1 U10650 ( .C1(n4338), .C2(n9938), .A(n9327), .B(n9326), .ZN(
        P1_U3356) );
  NAND2_X1 U10651 ( .A1(n9344), .A2(n9328), .ZN(n9329) );
  XNOR2_X1 U10652 ( .A(n9329), .B(n9332), .ZN(n9331) );
  AOI21_X1 U10653 ( .B1(n9331), .B2(n9910), .A(n9330), .ZN(n9551) );
  NAND2_X1 U10654 ( .A1(n9553), .A2(n9935), .ZN(n9341) );
  OAI211_X1 U10655 ( .C1(n7725), .C2(n4316), .A(n9917), .B(n9335), .ZN(n9550)
         );
  INV_X1 U10656 ( .A(n9550), .ZN(n9339) );
  AOI22_X1 U10657 ( .A1(n9928), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9336), .B2(
        n9927), .ZN(n9337) );
  OAI21_X1 U10658 ( .B1(n7725), .B2(n9530), .A(n9337), .ZN(n9338) );
  AOI21_X1 U10659 ( .B1(n9339), .B2(n9921), .A(n9338), .ZN(n9340) );
  OAI211_X1 U10660 ( .C1(n9551), .C2(n9928), .A(n9341), .B(n9340), .ZN(
        P1_U3265) );
  INV_X1 U10661 ( .A(n9342), .ZN(n9343) );
  NOR2_X1 U10662 ( .A1(n9531), .A2(n9343), .ZN(n9349) );
  OAI21_X1 U10663 ( .B1(n4676), .B2(n9345), .A(n9344), .ZN(n9347) );
  AOI21_X1 U10664 ( .B1(n9347), .B2(n9910), .A(n9346), .ZN(n9348) );
  INV_X1 U10665 ( .A(n9348), .ZN(n9557) );
  AOI211_X1 U10666 ( .C1(n9558), .C2(n9350), .A(n9349), .B(n9557), .ZN(n9355)
         );
  NAND2_X1 U10667 ( .A1(n9559), .A2(n9935), .ZN(n9354) );
  AOI22_X1 U10668 ( .A1(n9556), .A2(n9925), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9928), .ZN(n9353) );
  OAI211_X1 U10669 ( .C1(n9938), .C2(n9355), .A(n9354), .B(n9353), .ZN(
        P1_U3266) );
  XNOR2_X1 U10670 ( .A(n9357), .B(n9356), .ZN(n9566) );
  INV_X1 U10671 ( .A(n9380), .ZN(n9360) );
  INV_X1 U10672 ( .A(n9358), .ZN(n9359) );
  AOI211_X1 U10673 ( .C1(n9563), .C2(n9360), .A(n9527), .B(n9359), .ZN(n9562)
         );
  AOI22_X1 U10674 ( .A1(n9938), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9361), .B2(
        n9927), .ZN(n9362) );
  OAI21_X1 U10675 ( .B1(n9363), .B2(n9530), .A(n9362), .ZN(n9370) );
  OAI21_X1 U10676 ( .B1(n9366), .B2(n9365), .A(n9364), .ZN(n9368) );
  AOI21_X1 U10677 ( .B1(n9368), .B2(n9910), .A(n9367), .ZN(n9565) );
  NOR2_X1 U10678 ( .A1(n9565), .A2(n9928), .ZN(n9369) );
  AOI211_X1 U10679 ( .C1(n9562), .C2(n9921), .A(n9370), .B(n9369), .ZN(n9371)
         );
  OAI21_X1 U10680 ( .B1(n9566), .B2(n9518), .A(n9371), .ZN(P1_U3267) );
  INV_X1 U10681 ( .A(n9372), .ZN(n9375) );
  AOI21_X1 U10682 ( .B1(n9389), .B2(n9373), .A(n9379), .ZN(n9374) );
  OAI21_X1 U10683 ( .B1(n9375), .B2(n9374), .A(n9910), .ZN(n9377) );
  NAND2_X1 U10684 ( .A1(n9377), .A2(n9376), .ZN(n9567) );
  INV_X1 U10685 ( .A(n9567), .ZN(n9387) );
  XNOR2_X1 U10686 ( .A(n9378), .B(n9379), .ZN(n9569) );
  NAND2_X1 U10687 ( .A1(n9569), .A2(n9935), .ZN(n9386) );
  AOI211_X1 U10688 ( .C1(n9381), .C2(n9395), .A(n9527), .B(n9380), .ZN(n9568)
         );
  AOI22_X1 U10689 ( .A1(n9382), .A2(n9927), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9938), .ZN(n9383) );
  OAI21_X1 U10690 ( .B1(n9649), .B2(n9530), .A(n9383), .ZN(n9384) );
  AOI21_X1 U10691 ( .B1(n9568), .B2(n9921), .A(n9384), .ZN(n9385) );
  OAI211_X1 U10692 ( .C1(n9938), .C2(n9387), .A(n9386), .B(n9385), .ZN(
        P1_U3268) );
  XNOR2_X1 U10693 ( .A(n9388), .B(n9390), .ZN(n9576) );
  OAI211_X1 U10694 ( .C1(n9391), .C2(n9390), .A(n9389), .B(n9910), .ZN(n9394)
         );
  INV_X1 U10695 ( .A(n9392), .ZN(n9393) );
  NAND2_X1 U10696 ( .A1(n9394), .A2(n9393), .ZN(n9572) );
  INV_X1 U10697 ( .A(n9574), .ZN(n9399) );
  AOI211_X1 U10698 ( .C1(n9574), .C2(n9403), .A(n9527), .B(n7724), .ZN(n9573)
         );
  NAND2_X1 U10699 ( .A1(n9573), .A2(n9921), .ZN(n9398) );
  AOI22_X1 U10700 ( .A1(n9396), .A2(n9927), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9938), .ZN(n9397) );
  OAI211_X1 U10701 ( .C1(n9399), .C2(n9530), .A(n9398), .B(n9397), .ZN(n9400)
         );
  AOI21_X1 U10702 ( .B1(n9534), .B2(n9572), .A(n9400), .ZN(n9401) );
  OAI21_X1 U10703 ( .B1(n9576), .B2(n9518), .A(n9401), .ZN(P1_U3269) );
  XOR2_X1 U10704 ( .A(n9409), .B(n9402), .Z(n9582) );
  INV_X1 U10705 ( .A(n9423), .ZN(n9405) );
  INV_X1 U10706 ( .A(n9403), .ZN(n9404) );
  AOI211_X1 U10707 ( .C1(n9579), .C2(n9405), .A(n9527), .B(n9404), .ZN(n9578)
         );
  OAI22_X1 U10708 ( .A1(n9407), .A2(n9530), .B1(n9406), .B2(n9534), .ZN(n9414)
         );
  XOR2_X1 U10709 ( .A(n9409), .B(n9408), .Z(n9411) );
  OAI21_X1 U10710 ( .B1(n9411), .B2(n9469), .A(n9410), .ZN(n9577) );
  AOI21_X1 U10711 ( .B1(n4888), .B2(n9927), .A(n9577), .ZN(n9412) );
  NOR2_X1 U10712 ( .A1(n9412), .A2(n9928), .ZN(n9413) );
  AOI211_X1 U10713 ( .C1(n9578), .C2(n9921), .A(n9414), .B(n9413), .ZN(n9415)
         );
  OAI21_X1 U10714 ( .B1(n9582), .B2(n9518), .A(n9415), .ZN(P1_U3270) );
  XNOR2_X1 U10715 ( .A(n9417), .B(n9416), .ZN(n9585) );
  INV_X1 U10716 ( .A(n9585), .ZN(n9431) );
  XNOR2_X1 U10717 ( .A(n9419), .B(n9418), .ZN(n9422) );
  INV_X1 U10718 ( .A(n9420), .ZN(n9421) );
  OAI21_X1 U10719 ( .B1(n9422), .B2(n9469), .A(n9421), .ZN(n9583) );
  AOI211_X1 U10720 ( .C1(n9424), .C2(n9443), .A(n9527), .B(n9423), .ZN(n9584)
         );
  NAND2_X1 U10721 ( .A1(n9584), .A2(n9921), .ZN(n9428) );
  INV_X1 U10722 ( .A(n9425), .ZN(n9426) );
  AOI22_X1 U10723 ( .A1(n9426), .A2(n9927), .B1(n9928), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9427) );
  OAI211_X1 U10724 ( .C1(n9655), .C2(n9530), .A(n9428), .B(n9427), .ZN(n9429)
         );
  AOI21_X1 U10725 ( .B1(n9534), .B2(n9583), .A(n9429), .ZN(n9430) );
  OAI21_X1 U10726 ( .B1(n9431), .B2(n9518), .A(n9430), .ZN(P1_U3271) );
  XOR2_X1 U10727 ( .A(n9432), .B(n9435), .Z(n9590) );
  INV_X1 U10728 ( .A(n9590), .ZN(n9450) );
  NAND2_X1 U10729 ( .A1(n9434), .A2(n9433), .ZN(n9437) );
  INV_X1 U10730 ( .A(n9435), .ZN(n9436) );
  NAND2_X1 U10731 ( .A1(n9437), .A2(n9436), .ZN(n9439) );
  NAND2_X1 U10732 ( .A1(n9439), .A2(n9438), .ZN(n9440) );
  NAND2_X1 U10733 ( .A1(n9440), .A2(n9910), .ZN(n9442) );
  NAND2_X1 U10734 ( .A1(n9442), .A2(n9441), .ZN(n9588) );
  AOI211_X1 U10735 ( .C1(n9444), .C2(n9457), .A(n9527), .B(n7723), .ZN(n9589)
         );
  NAND2_X1 U10736 ( .A1(n9589), .A2(n9921), .ZN(n9447) );
  AOI22_X1 U10737 ( .A1(n9928), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9445), .B2(
        n9927), .ZN(n9446) );
  OAI211_X1 U10738 ( .C1(n9295), .C2(n9530), .A(n9447), .B(n9446), .ZN(n9448)
         );
  AOI21_X1 U10739 ( .B1(n9534), .B2(n9588), .A(n9448), .ZN(n9449) );
  OAI21_X1 U10740 ( .B1(n9450), .B2(n9518), .A(n9449), .ZN(P1_U3272) );
  XOR2_X1 U10741 ( .A(n9455), .B(n9451), .Z(n9453) );
  OAI21_X1 U10742 ( .B1(n9453), .B2(n9469), .A(n9452), .ZN(n9593) );
  AOI21_X1 U10743 ( .B1(n9454), .B2(n9927), .A(n9593), .ZN(n9465) );
  XOR2_X1 U10744 ( .A(n9456), .B(n9455), .Z(n9595) );
  NAND2_X1 U10745 ( .A1(n9595), .A2(n9935), .ZN(n9464) );
  INV_X1 U10746 ( .A(n9473), .ZN(n9459) );
  INV_X1 U10747 ( .A(n9457), .ZN(n9458) );
  AOI211_X1 U10748 ( .C1(n9460), .C2(n9459), .A(n9527), .B(n9458), .ZN(n9594)
         );
  OAI22_X1 U10749 ( .A1(n9662), .A2(n9530), .B1(n9461), .B2(n9534), .ZN(n9462)
         );
  AOI21_X1 U10750 ( .B1(n9594), .B2(n9921), .A(n9462), .ZN(n9463) );
  OAI211_X1 U10751 ( .C1(n9938), .C2(n9465), .A(n9464), .B(n9463), .ZN(
        P1_U3273) );
  XOR2_X1 U10752 ( .A(n9471), .B(n9466), .Z(n9470) );
  INV_X1 U10753 ( .A(n9467), .ZN(n9468) );
  OAI21_X1 U10754 ( .B1(n9470), .B2(n9469), .A(n9468), .ZN(n9598) );
  INV_X1 U10755 ( .A(n9598), .ZN(n9481) );
  XNOR2_X1 U10756 ( .A(n9472), .B(n9471), .ZN(n9600) );
  NAND2_X1 U10757 ( .A1(n9600), .A2(n9935), .ZN(n9480) );
  AOI211_X1 U10758 ( .C1(n9474), .C2(n9491), .A(n9527), .B(n9473), .ZN(n9599)
         );
  NOR2_X1 U10759 ( .A1(n9666), .A2(n9530), .ZN(n9478) );
  OAI22_X1 U10760 ( .A1(n9534), .A2(n9476), .B1(n9475), .B2(n9531), .ZN(n9477)
         );
  AOI211_X1 U10761 ( .C1(n9599), .C2(n9921), .A(n9478), .B(n9477), .ZN(n9479)
         );
  OAI211_X1 U10762 ( .C1(n9938), .C2(n9481), .A(n9480), .B(n9479), .ZN(
        P1_U3274) );
  XNOR2_X1 U10763 ( .A(n9482), .B(n9486), .ZN(n9604) );
  INV_X1 U10764 ( .A(n9604), .ZN(n9500) );
  AND2_X1 U10765 ( .A1(n9506), .A2(n9483), .ZN(n9485) );
  OAI21_X1 U10766 ( .B1(n9486), .B2(n9485), .A(n9484), .ZN(n9487) );
  NAND2_X1 U10767 ( .A1(n9487), .A2(n9910), .ZN(n9490) );
  INV_X1 U10768 ( .A(n9488), .ZN(n9489) );
  NAND2_X1 U10769 ( .A1(n9490), .A2(n9489), .ZN(n9602) );
  INV_X1 U10770 ( .A(n9491), .ZN(n9492) );
  AOI211_X1 U10771 ( .C1(n9493), .C2(n9509), .A(n9527), .B(n9492), .ZN(n9603)
         );
  NAND2_X1 U10772 ( .A1(n9603), .A2(n9921), .ZN(n9497) );
  INV_X1 U10773 ( .A(n9494), .ZN(n9495) );
  AOI22_X1 U10774 ( .A1(n9928), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9495), .B2(
        n9927), .ZN(n9496) );
  OAI211_X1 U10775 ( .C1(n9670), .C2(n9530), .A(n9497), .B(n9496), .ZN(n9498)
         );
  AOI21_X1 U10776 ( .B1(n9534), .B2(n9602), .A(n9498), .ZN(n9499) );
  OAI21_X1 U10777 ( .B1(n9500), .B2(n9518), .A(n9499), .ZN(P1_U3275) );
  XNOR2_X1 U10778 ( .A(n9501), .B(n9503), .ZN(n9609) );
  INV_X1 U10779 ( .A(n9609), .ZN(n9519) );
  NAND2_X1 U10780 ( .A1(n9520), .A2(n9502), .ZN(n9504) );
  NAND2_X1 U10781 ( .A1(n9504), .A2(n9503), .ZN(n9505) );
  NAND3_X1 U10782 ( .A1(n9506), .A2(n9505), .A3(n9910), .ZN(n9508) );
  NAND2_X1 U10783 ( .A1(n9508), .A2(n9507), .ZN(n9607) );
  INV_X1 U10784 ( .A(n9526), .ZN(n9511) );
  INV_X1 U10785 ( .A(n9509), .ZN(n9510) );
  AOI211_X1 U10786 ( .C1(n9512), .C2(n9511), .A(n9527), .B(n9510), .ZN(n9608)
         );
  NAND2_X1 U10787 ( .A1(n9608), .A2(n9921), .ZN(n9515) );
  AOI22_X1 U10788 ( .A1(n9928), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9513), .B2(
        n9927), .ZN(n9514) );
  OAI211_X1 U10789 ( .C1(n9674), .C2(n9530), .A(n9515), .B(n9514), .ZN(n9516)
         );
  AOI21_X1 U10790 ( .B1(n9534), .B2(n9607), .A(n9516), .ZN(n9517) );
  OAI21_X1 U10791 ( .B1(n9519), .B2(n9518), .A(n9517), .ZN(P1_U3276) );
  OAI21_X1 U10792 ( .B1(n9524), .B2(n9521), .A(n9520), .ZN(n9523) );
  AOI21_X1 U10793 ( .B1(n9523), .B2(n9910), .A(n9522), .ZN(n9612) );
  XNOR2_X1 U10794 ( .A(n9525), .B(n9524), .ZN(n9615) );
  NAND2_X1 U10795 ( .A1(n9615), .A2(n9935), .ZN(n9538) );
  AOI211_X1 U10796 ( .C1(n9529), .C2(n9528), .A(n9527), .B(n9526), .ZN(n9614)
         );
  INV_X1 U10797 ( .A(n9529), .ZN(n9678) );
  NOR2_X1 U10798 ( .A1(n9678), .A2(n9530), .ZN(n9536) );
  OAI22_X1 U10799 ( .A1(n9534), .A2(n9533), .B1(n9532), .B2(n9531), .ZN(n9535)
         );
  AOI211_X1 U10800 ( .C1(n9614), .C2(n9921), .A(n9536), .B(n9535), .ZN(n9537)
         );
  OAI211_X1 U10801 ( .C1(n9938), .C2(n9612), .A(n9538), .B(n9537), .ZN(
        P1_U3277) );
  INV_X1 U10802 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9541) );
  NOR2_X1 U10803 ( .A1(n9540), .A2(n9539), .ZN(n9629) );
  MUX2_X1 U10804 ( .A(n9541), .B(n9629), .S(n9978), .Z(n9542) );
  OAI21_X1 U10805 ( .B1(n9632), .B2(n9627), .A(n9542), .ZN(P1_U3553) );
  AND2_X1 U10806 ( .A1(n9544), .A2(n9543), .ZN(n9633) );
  MUX2_X1 U10807 ( .A(n9545), .B(n9633), .S(n9978), .Z(n9546) );
  OAI21_X1 U10808 ( .B1(n9636), .B2(n9627), .A(n9546), .ZN(P1_U3552) );
  NOR2_X1 U10809 ( .A1(n4461), .A2(n9965), .ZN(n9548) );
  MUX2_X1 U10810 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9637), .S(n9978), .Z(
        P1_U3551) );
  INV_X1 U10811 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9554) );
  NAND2_X1 U10812 ( .A1(n9551), .A2(n9550), .ZN(n9552) );
  MUX2_X1 U10813 ( .A(n9554), .B(n9638), .S(n9978), .Z(n9555) );
  OAI21_X1 U10814 ( .B1(n7725), .B2(n9627), .A(n9555), .ZN(P1_U3550) );
  INV_X1 U10815 ( .A(n9556), .ZN(n9644) );
  INV_X1 U10816 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9560) );
  MUX2_X1 U10817 ( .A(n9560), .B(n9641), .S(n9978), .Z(n9561) );
  OAI21_X1 U10818 ( .B1(n9644), .B2(n9627), .A(n9561), .ZN(P1_U3549) );
  AOI21_X1 U10819 ( .B1(n9580), .B2(n9563), .A(n9562), .ZN(n9564) );
  OAI211_X1 U10820 ( .C1(n9566), .C2(n9962), .A(n9565), .B(n9564), .ZN(n9645)
         );
  MUX2_X1 U10821 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9645), .S(n9978), .Z(
        P1_U3548) );
  INV_X1 U10822 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9570) );
  AOI211_X1 U10823 ( .C1(n9569), .C2(n9958), .A(n9568), .B(n9567), .ZN(n9646)
         );
  MUX2_X1 U10824 ( .A(n9570), .B(n9646), .S(n9978), .Z(n9571) );
  OAI21_X1 U10825 ( .B1(n9649), .B2(n9627), .A(n9571), .ZN(P1_U3547) );
  AOI211_X1 U10826 ( .C1(n9580), .C2(n9574), .A(n9573), .B(n9572), .ZN(n9575)
         );
  OAI21_X1 U10827 ( .B1(n9576), .B2(n9962), .A(n9575), .ZN(n9650) );
  MUX2_X1 U10828 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9650), .S(n9978), .Z(
        P1_U3546) );
  AOI211_X1 U10829 ( .C1(n9580), .C2(n9579), .A(n9578), .B(n9577), .ZN(n9581)
         );
  OAI21_X1 U10830 ( .B1(n9582), .B2(n9962), .A(n9581), .ZN(n9651) );
  MUX2_X1 U10831 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9651), .S(n9978), .Z(
        P1_U3545) );
  AOI211_X1 U10832 ( .C1(n9585), .C2(n9958), .A(n9584), .B(n9583), .ZN(n9652)
         );
  MUX2_X1 U10833 ( .A(n9586), .B(n9652), .S(n9978), .Z(n9587) );
  OAI21_X1 U10834 ( .B1(n9655), .B2(n9627), .A(n9587), .ZN(P1_U3544) );
  INV_X1 U10835 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9591) );
  AOI211_X1 U10836 ( .C1(n9590), .C2(n9958), .A(n9589), .B(n9588), .ZN(n9656)
         );
  MUX2_X1 U10837 ( .A(n9591), .B(n9656), .S(n9978), .Z(n9592) );
  OAI21_X1 U10838 ( .B1(n9295), .B2(n9627), .A(n9592), .ZN(P1_U3543) );
  INV_X1 U10839 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9596) );
  AOI211_X1 U10840 ( .C1(n9595), .C2(n9958), .A(n9594), .B(n9593), .ZN(n9659)
         );
  MUX2_X1 U10841 ( .A(n9596), .B(n9659), .S(n9978), .Z(n9597) );
  OAI21_X1 U10842 ( .B1(n9662), .B2(n9627), .A(n9597), .ZN(P1_U3542) );
  AOI211_X1 U10843 ( .C1(n9600), .C2(n9958), .A(n9599), .B(n9598), .ZN(n9663)
         );
  MUX2_X1 U10844 ( .A(n4379), .B(n9663), .S(n9978), .Z(n9601) );
  OAI21_X1 U10845 ( .B1(n9666), .B2(n9627), .A(n9601), .ZN(P1_U3541) );
  AOI211_X1 U10846 ( .C1(n9604), .C2(n9958), .A(n9603), .B(n9602), .ZN(n9667)
         );
  MUX2_X1 U10847 ( .A(n9605), .B(n9667), .S(n9978), .Z(n9606) );
  OAI21_X1 U10848 ( .B1(n9670), .B2(n9627), .A(n9606), .ZN(P1_U3540) );
  AOI211_X1 U10849 ( .C1(n9609), .C2(n9958), .A(n9608), .B(n9607), .ZN(n9671)
         );
  MUX2_X1 U10850 ( .A(n9610), .B(n9671), .S(n9978), .Z(n9611) );
  OAI21_X1 U10851 ( .B1(n9674), .B2(n9627), .A(n9611), .ZN(P1_U3539) );
  INV_X1 U10852 ( .A(n9612), .ZN(n9613) );
  AOI211_X1 U10853 ( .C1(n9615), .C2(n9958), .A(n9614), .B(n9613), .ZN(n9675)
         );
  MUX2_X1 U10854 ( .A(n9616), .B(n9675), .S(n9978), .Z(n9617) );
  OAI21_X1 U10855 ( .B1(n9678), .B2(n9627), .A(n9617), .ZN(P1_U3538) );
  INV_X1 U10856 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9854) );
  AOI211_X1 U10857 ( .C1(n9620), .C2(n9958), .A(n9619), .B(n9618), .ZN(n9679)
         );
  MUX2_X1 U10858 ( .A(n9854), .B(n9679), .S(n9978), .Z(n9621) );
  OAI21_X1 U10859 ( .B1(n9276), .B2(n9627), .A(n9621), .ZN(P1_U3537) );
  INV_X1 U10860 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9625) );
  AOI211_X1 U10861 ( .C1(n9624), .C2(n9958), .A(n9623), .B(n9622), .ZN(n9682)
         );
  MUX2_X1 U10862 ( .A(n9625), .B(n9682), .S(n9978), .Z(n9626) );
  OAI21_X1 U10863 ( .B1(n9686), .B2(n9627), .A(n9626), .ZN(P1_U3536) );
  MUX2_X1 U10864 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9628), .S(n9978), .Z(
        P1_U3522) );
  INV_X1 U10865 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9630) );
  MUX2_X1 U10866 ( .A(n9630), .B(n9629), .S(n9971), .Z(n9631) );
  OAI21_X1 U10867 ( .B1(n9632), .B2(n9685), .A(n9631), .ZN(P1_U3521) );
  INV_X1 U10868 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9634) );
  MUX2_X1 U10869 ( .A(n9634), .B(n9633), .S(n9971), .Z(n9635) );
  OAI21_X1 U10870 ( .B1(n9636), .B2(n9685), .A(n9635), .ZN(P1_U3520) );
  MUX2_X1 U10871 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9637), .S(n9961), .Z(
        P1_U3519) );
  INV_X1 U10872 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9639) );
  MUX2_X1 U10873 ( .A(n9639), .B(n9638), .S(n9971), .Z(n9640) );
  OAI21_X1 U10874 ( .B1(n7725), .B2(n9685), .A(n9640), .ZN(P1_U3518) );
  INV_X1 U10875 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9642) );
  MUX2_X1 U10876 ( .A(n9642), .B(n9641), .S(n9971), .Z(n9643) );
  OAI21_X1 U10877 ( .B1(n9644), .B2(n9685), .A(n9643), .ZN(P1_U3517) );
  MUX2_X1 U10878 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9645), .S(n9961), .Z(
        P1_U3516) );
  INV_X1 U10879 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9647) );
  MUX2_X1 U10880 ( .A(n9647), .B(n9646), .S(n9971), .Z(n9648) );
  OAI21_X1 U10881 ( .B1(n9649), .B2(n9685), .A(n9648), .ZN(P1_U3515) );
  MUX2_X1 U10882 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9650), .S(n9961), .Z(
        P1_U3514) );
  MUX2_X1 U10883 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9651), .S(n9961), .Z(
        P1_U3513) );
  INV_X1 U10884 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9653) );
  MUX2_X1 U10885 ( .A(n9653), .B(n9652), .S(n9971), .Z(n9654) );
  OAI21_X1 U10886 ( .B1(n9655), .B2(n9685), .A(n9654), .ZN(P1_U3512) );
  INV_X1 U10887 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9657) );
  MUX2_X1 U10888 ( .A(n9657), .B(n9656), .S(n9971), .Z(n9658) );
  OAI21_X1 U10889 ( .B1(n9295), .B2(n9685), .A(n9658), .ZN(P1_U3511) );
  INV_X1 U10890 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9660) );
  MUX2_X1 U10891 ( .A(n9660), .B(n9659), .S(n9971), .Z(n9661) );
  OAI21_X1 U10892 ( .B1(n9662), .B2(n9685), .A(n9661), .ZN(P1_U3510) );
  MUX2_X1 U10893 ( .A(n9664), .B(n9663), .S(n9961), .Z(n9665) );
  OAI21_X1 U10894 ( .B1(n9666), .B2(n9685), .A(n9665), .ZN(P1_U3509) );
  INV_X1 U10895 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9668) );
  MUX2_X1 U10896 ( .A(n9668), .B(n9667), .S(n9971), .Z(n9669) );
  OAI21_X1 U10897 ( .B1(n9670), .B2(n9685), .A(n9669), .ZN(P1_U3507) );
  INV_X1 U10898 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9672) );
  MUX2_X1 U10899 ( .A(n9672), .B(n9671), .S(n9971), .Z(n9673) );
  OAI21_X1 U10900 ( .B1(n9674), .B2(n9685), .A(n9673), .ZN(P1_U3504) );
  MUX2_X1 U10901 ( .A(n9676), .B(n9675), .S(n9971), .Z(n9677) );
  OAI21_X1 U10902 ( .B1(n9678), .B2(n9685), .A(n9677), .ZN(P1_U3501) );
  INV_X1 U10903 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9680) );
  MUX2_X1 U10904 ( .A(n9680), .B(n9679), .S(n9971), .Z(n9681) );
  OAI21_X1 U10905 ( .B1(n9276), .B2(n9685), .A(n9681), .ZN(P1_U3498) );
  INV_X1 U10906 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9683) );
  MUX2_X1 U10907 ( .A(n9683), .B(n9682), .S(n9971), .Z(n9684) );
  OAI21_X1 U10908 ( .B1(n9686), .B2(n9685), .A(n9684), .ZN(P1_U3495) );
  INV_X1 U10909 ( .A(n9687), .ZN(n9692) );
  NOR4_X1 U10910 ( .A1(n9689), .A2(P1_U3086), .A3(n9688), .A4(
        P1_IR_REG_30__SCAN_IN), .ZN(n9691) );
  AOI22_X1 U10911 ( .A1(n9692), .A2(n9691), .B1(P2_DATAO_REG_31__SCAN_IN), 
        .B2(n9690), .ZN(n9693) );
  OAI21_X1 U10912 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(P1_U3324) );
  MUX2_X1 U10913 ( .A(n9696), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10914 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9707) );
  AOI211_X1 U10915 ( .C1(n9699), .C2(n9698), .A(n9697), .B(n9851), .ZN(n9704)
         );
  AOI211_X1 U10916 ( .C1(n9702), .C2(n9701), .A(n9700), .B(n9889), .ZN(n9703)
         );
  AOI211_X1 U10917 ( .C1(n9881), .C2(n9705), .A(n9704), .B(n9703), .ZN(n9706)
         );
  NAND2_X1 U10918 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9757) );
  OAI211_X1 U10919 ( .C1(n9904), .C2(n9707), .A(n9706), .B(n9757), .ZN(
        P1_U3253) );
  INV_X1 U10920 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9720) );
  OAI21_X1 U10921 ( .B1(n9709), .B2(n9708), .A(n9884), .ZN(n9711) );
  NOR2_X1 U10922 ( .A1(n9711), .A2(n9710), .ZN(n9716) );
  AOI211_X1 U10923 ( .C1(n9714), .C2(n9713), .A(n9851), .B(n9712), .ZN(n9715)
         );
  AOI211_X1 U10924 ( .C1(n9881), .C2(n9717), .A(n9716), .B(n9715), .ZN(n9719)
         );
  OAI211_X1 U10925 ( .C1(n9904), .C2(n9720), .A(n9719), .B(n9718), .ZN(
        P1_U3250) );
  INV_X1 U10926 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9731) );
  AOI211_X1 U10927 ( .C1(n9723), .C2(n9722), .A(n9721), .B(n9889), .ZN(n9728)
         );
  AOI211_X1 U10928 ( .C1(n9726), .C2(n9725), .A(n9724), .B(n9851), .ZN(n9727)
         );
  AOI211_X1 U10929 ( .C1(n9881), .C2(n9729), .A(n9728), .B(n9727), .ZN(n9730)
         );
  NAND2_X1 U10930 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9785) );
  OAI211_X1 U10931 ( .C1(n9904), .C2(n9731), .A(n9730), .B(n9785), .ZN(
        P1_U3251) );
  OAI21_X1 U10932 ( .B1(n9734), .B2(n9733), .A(n9732), .ZN(n9735) );
  AOI21_X1 U10933 ( .B1(n9737), .B2(n9736), .A(n9735), .ZN(n9745) );
  XNOR2_X1 U10934 ( .A(n9738), .B(n9739), .ZN(n9743) );
  AOI22_X1 U10935 ( .A1(n9743), .A2(n9742), .B1(n9741), .B2(n9740), .ZN(n9744)
         );
  OAI211_X1 U10936 ( .C1(n9747), .C2(n9746), .A(n9745), .B(n9744), .ZN(
        P2_U3155) );
  NOR2_X1 U10937 ( .A1(n9748), .A2(n10072), .ZN(n9750) );
  AOI211_X1 U10938 ( .C1(n10070), .C2(n9751), .A(n9750), .B(n9749), .ZN(n9754)
         );
  AOI22_X1 U10939 ( .A1(n10107), .A2(n9754), .B1(n9752), .B2(n6337), .ZN(
        P2_U3472) );
  INV_X1 U10940 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9753) );
  AOI22_X1 U10941 ( .A1(n10080), .A2(n9754), .B1(n9753), .B2(n10078), .ZN(
        P2_U3429) );
  AOI21_X1 U10942 ( .B1(n9756), .B2(n9755), .A(n4349), .ZN(n9765) );
  INV_X1 U10943 ( .A(n9757), .ZN(n9763) );
  AOI22_X1 U10944 ( .A1(n9761), .A2(n9760), .B1(n9759), .B2(n9758), .ZN(n9908)
         );
  NOR2_X1 U10945 ( .A1(n9787), .A2(n9908), .ZN(n9762) );
  AOI211_X1 U10946 ( .C1(n9913), .C2(n4282), .A(n9763), .B(n9762), .ZN(n9764)
         );
  OAI21_X1 U10947 ( .B1(n9765), .B2(n9792), .A(n9764), .ZN(n9766) );
  INV_X1 U10948 ( .A(n9766), .ZN(n9767) );
  OAI21_X1 U10949 ( .B1(n9797), .B2(n9768), .A(n9767), .ZN(P1_U3217) );
  INV_X1 U10950 ( .A(n9769), .ZN(n9770) );
  OAI21_X1 U10951 ( .B1(n9787), .B2(n9771), .A(n9770), .ZN(n9778) );
  INV_X1 U10952 ( .A(n9772), .ZN(n9776) );
  NAND3_X1 U10953 ( .A1(n7399), .A2(n9774), .A3(n9773), .ZN(n9775) );
  AOI21_X1 U10954 ( .B1(n9776), .B2(n9775), .A(n9792), .ZN(n9777) );
  AOI211_X1 U10955 ( .C1(n9779), .C2(n4282), .A(n9778), .B(n9777), .ZN(n9780)
         );
  OAI21_X1 U10956 ( .B1(n9797), .B2(n9781), .A(n9780), .ZN(P1_U3224) );
  XNOR2_X1 U10957 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10958 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U10959 ( .B1(n9784), .B2(n9783), .A(n9782), .ZN(n9793) );
  INV_X1 U10960 ( .A(n9785), .ZN(n9789) );
  NOR2_X1 U10961 ( .A1(n9787), .A2(n9786), .ZN(n9788) );
  AOI211_X1 U10962 ( .C1(n9790), .C2(n4282), .A(n9789), .B(n9788), .ZN(n9791)
         );
  OAI21_X1 U10963 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(n9794) );
  INV_X1 U10964 ( .A(n9794), .ZN(n9795) );
  OAI21_X1 U10965 ( .B1(n9797), .B2(n9796), .A(n9795), .ZN(P1_U3221) );
  NAND2_X1 U10966 ( .A1(n6469), .A2(n9798), .ZN(n9802) );
  INV_X1 U10967 ( .A(n9799), .ZN(n9800) );
  NAND2_X1 U10968 ( .A1(n9800), .A2(n9802), .ZN(n9801) );
  MUX2_X1 U10969 ( .A(n9802), .B(n9801), .S(P1_IR_REG_0__SCAN_IN), .Z(n9804)
         );
  NAND2_X1 U10970 ( .A1(n9804), .A2(n9803), .ZN(n9806) );
  AOI22_X1 U10971 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9869), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9805) );
  OAI21_X1 U10972 ( .B1(n9807), .B2(n9806), .A(n9805), .ZN(P1_U3243) );
  INV_X1 U10973 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9822) );
  AOI21_X1 U10974 ( .B1(n9810), .B2(n9809), .A(n9808), .ZN(n9811) );
  NAND2_X1 U10975 ( .A1(n9884), .A2(n9811), .ZN(n9817) );
  AOI21_X1 U10976 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n9815) );
  NAND2_X1 U10977 ( .A1(n9892), .A2(n9815), .ZN(n9816) );
  OAI211_X1 U10978 ( .C1(n9898), .C2(n9818), .A(n9817), .B(n9816), .ZN(n9819)
         );
  INV_X1 U10979 ( .A(n9819), .ZN(n9821) );
  OAI211_X1 U10980 ( .C1(n9904), .C2(n9822), .A(n9821), .B(n9820), .ZN(
        P1_U3254) );
  AOI211_X1 U10981 ( .C1(n9825), .C2(n9824), .A(n9823), .B(n9851), .ZN(n9830)
         );
  AOI211_X1 U10982 ( .C1(n9828), .C2(n9827), .A(n9826), .B(n9889), .ZN(n9829)
         );
  AOI211_X1 U10983 ( .C1(n9881), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9833)
         );
  OAI211_X1 U10984 ( .C1(n9834), .C2(n9904), .A(n9833), .B(n9832), .ZN(
        P1_U3256) );
  INV_X1 U10985 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9849) );
  AOI21_X1 U10986 ( .B1(n9837), .B2(n9836), .A(n9835), .ZN(n9838) );
  NAND2_X1 U10987 ( .A1(n9884), .A2(n9838), .ZN(n9844) );
  AOI21_X1 U10988 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(n9842) );
  NAND2_X1 U10989 ( .A1(n9892), .A2(n9842), .ZN(n9843) );
  OAI211_X1 U10990 ( .C1(n9898), .C2(n9845), .A(n9844), .B(n9843), .ZN(n9846)
         );
  INV_X1 U10991 ( .A(n9846), .ZN(n9848) );
  NAND2_X1 U10992 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9847) );
  OAI211_X1 U10993 ( .C1(n9904), .C2(n9849), .A(n9848), .B(n9847), .ZN(
        P1_U3257) );
  INV_X1 U10994 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9863) );
  INV_X1 U10995 ( .A(n9850), .ZN(n9853) );
  AOI211_X1 U10996 ( .C1(n9854), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9859)
         );
  AOI211_X1 U10997 ( .C1(n9857), .C2(n9856), .A(n9855), .B(n9889), .ZN(n9858)
         );
  AOI211_X1 U10998 ( .C1(n9881), .C2(n9860), .A(n9859), .B(n9858), .ZN(n9862)
         );
  OAI211_X1 U10999 ( .C1(n9904), .C2(n9863), .A(n9862), .B(n9861), .ZN(
        P1_U3258) );
  AOI211_X1 U11000 ( .C1(n9866), .C2(n9865), .A(n9864), .B(n9889), .ZN(n9867)
         );
  AOI211_X1 U11001 ( .C1(n9869), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9868), .B(
        n9867), .ZN(n9876) );
  OAI21_X1 U11002 ( .B1(n9872), .B2(n9871), .A(n9870), .ZN(n9874) );
  AOI22_X1 U11003 ( .A1(n9874), .A2(n9892), .B1(n9873), .B2(n9881), .ZN(n9875)
         );
  NAND2_X1 U11004 ( .A1(n9876), .A2(n9875), .ZN(P1_U3259) );
  XNOR2_X1 U11005 ( .A(n9878), .B(n9877), .ZN(n9885) );
  XNOR2_X1 U11006 ( .A(n9880), .B(n9879), .ZN(n9883) );
  AOI222_X1 U11007 ( .A1(n9885), .A2(n9884), .B1(n9892), .B2(n9883), .C1(n9882), .C2(n9881), .ZN(n9887) );
  OAI211_X1 U11008 ( .C1(n9904), .C2(n9888), .A(n9887), .B(n9886), .ZN(
        P1_U3260) );
  AOI21_X1 U11009 ( .B1(n9891), .B2(n9890), .A(n9889), .ZN(n9901) );
  OAI211_X1 U11010 ( .C1(n9895), .C2(n9894), .A(n9893), .B(n9892), .ZN(n9896)
         );
  OAI21_X1 U11011 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(n9899) );
  AOI21_X1 U11012 ( .B1(n9901), .B2(n9900), .A(n9899), .ZN(n9903) );
  NAND2_X1 U11013 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9902) );
  OAI211_X1 U11014 ( .C1(n9904), .C2(n10114), .A(n9903), .B(n9902), .ZN(
        P1_U3261) );
  INV_X1 U11015 ( .A(n9905), .ZN(n9907) );
  OAI21_X1 U11016 ( .B1(n9907), .B2(n4643), .A(n9906), .ZN(n9911) );
  INV_X1 U11017 ( .A(n9908), .ZN(n9909) );
  AOI21_X1 U11018 ( .B1(n9911), .B2(n9910), .A(n9909), .ZN(n9955) );
  AOI222_X1 U11019 ( .A1(n9913), .A2(n9925), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n9938), .C1(n9912), .C2(n9927), .ZN(n9923) );
  XNOR2_X1 U11020 ( .A(n9915), .B(n9914), .ZN(n9959) );
  INV_X1 U11021 ( .A(n9916), .ZN(n9918) );
  OAI211_X1 U11022 ( .C1(n9956), .C2(n9919), .A(n9918), .B(n9917), .ZN(n9954)
         );
  INV_X1 U11023 ( .A(n9954), .ZN(n9920) );
  AOI22_X1 U11024 ( .A1(n9959), .A2(n9935), .B1(n9921), .B2(n9920), .ZN(n9922)
         );
  OAI211_X1 U11025 ( .C1(n9938), .C2(n9955), .A(n9923), .B(n9922), .ZN(
        P1_U3283) );
  NAND2_X1 U11026 ( .A1(n9925), .A2(n9924), .ZN(n9930) );
  AOI22_X1 U11027 ( .A1(n9928), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9927), .B2(
        n9926), .ZN(n9929) );
  OAI211_X1 U11028 ( .C1(n9932), .C2(n9931), .A(n9930), .B(n9929), .ZN(n9933)
         );
  AOI21_X1 U11029 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(n9936) );
  OAI21_X1 U11030 ( .B1(n9938), .B2(n9937), .A(n9936), .ZN(P1_U3290) );
  AND2_X1 U11031 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9941), .ZN(P1_U3294) );
  AND2_X1 U11032 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9941), .ZN(P1_U3295) );
  AND2_X1 U11033 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9941), .ZN(P1_U3296) );
  AND2_X1 U11034 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9941), .ZN(P1_U3297) );
  AND2_X1 U11035 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9941), .ZN(P1_U3298) );
  AND2_X1 U11036 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9941), .ZN(P1_U3299) );
  AND2_X1 U11037 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9941), .ZN(P1_U3300) );
  AND2_X1 U11038 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9941), .ZN(P1_U3301) );
  AND2_X1 U11039 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9941), .ZN(P1_U3302) );
  AND2_X1 U11040 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9941), .ZN(P1_U3303) );
  NOR2_X1 U11041 ( .A1(n9940), .A2(n9939), .ZN(P1_U3304) );
  AND2_X1 U11042 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9941), .ZN(P1_U3305) );
  AND2_X1 U11043 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9941), .ZN(P1_U3306) );
  AND2_X1 U11044 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9941), .ZN(P1_U3307) );
  AND2_X1 U11045 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9941), .ZN(P1_U3308) );
  AND2_X1 U11046 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9941), .ZN(P1_U3309) );
  AND2_X1 U11047 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9941), .ZN(P1_U3310) );
  AND2_X1 U11048 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9941), .ZN(P1_U3311) );
  AND2_X1 U11049 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9941), .ZN(P1_U3312) );
  AND2_X1 U11050 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9941), .ZN(P1_U3313) );
  AND2_X1 U11051 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9941), .ZN(P1_U3314) );
  AND2_X1 U11052 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9941), .ZN(P1_U3315) );
  AND2_X1 U11053 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9941), .ZN(P1_U3316) );
  AND2_X1 U11054 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9941), .ZN(P1_U3317) );
  AND2_X1 U11055 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9941), .ZN(P1_U3318) );
  AND2_X1 U11056 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9941), .ZN(P1_U3319) );
  AND2_X1 U11057 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9941), .ZN(P1_U3320) );
  AND2_X1 U11058 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9941), .ZN(P1_U3321) );
  AND2_X1 U11059 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9941), .ZN(P1_U3322) );
  AND2_X1 U11060 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9941), .ZN(P1_U3323) );
  OAI21_X1 U11061 ( .B1(n9943), .B2(n9965), .A(n9942), .ZN(n9945) );
  AOI211_X1 U11062 ( .C1(n9958), .C2(n9946), .A(n9945), .B(n9944), .ZN(n9973)
         );
  INV_X1 U11063 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U11064 ( .A1(n9961), .A2(n9973), .B1(n9947), .B2(n6560), .ZN(
        P1_U3465) );
  INV_X1 U11065 ( .A(n5265), .ZN(n9949) );
  OAI21_X1 U11066 ( .B1(n9949), .B2(n9965), .A(n9948), .ZN(n9951) );
  AOI211_X1 U11067 ( .C1(n9958), .C2(n9952), .A(n9951), .B(n9950), .ZN(n9975)
         );
  INV_X1 U11068 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9953) );
  AOI22_X1 U11069 ( .A1(n9971), .A2(n9975), .B1(n9953), .B2(n6560), .ZN(
        P1_U3480) );
  OAI211_X1 U11070 ( .C1(n9956), .C2(n9965), .A(n9955), .B(n9954), .ZN(n9957)
         );
  AOI21_X1 U11071 ( .B1(n9959), .B2(n9958), .A(n9957), .ZN(n9977) );
  INV_X1 U11072 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U11073 ( .A1(n9961), .A2(n9977), .B1(n9960), .B2(n6560), .ZN(
        P1_U3483) );
  NOR3_X1 U11074 ( .A1(n7596), .A2(n9963), .A3(n9962), .ZN(n9969) );
  OAI21_X1 U11075 ( .B1(n9966), .B2(n9965), .A(n9964), .ZN(n9967) );
  NOR3_X1 U11076 ( .A1(n9969), .A2(n9968), .A3(n9967), .ZN(n9980) );
  INV_X1 U11077 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9970) );
  AOI22_X1 U11078 ( .A1(n9971), .A2(n9980), .B1(n9970), .B2(n6560), .ZN(
        P1_U3492) );
  AOI22_X1 U11079 ( .A1(n9978), .A2(n9973), .B1(n9972), .B2(n9979), .ZN(
        P1_U3526) );
  INV_X1 U11080 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11081 ( .A1(n9978), .A2(n9975), .B1(n9974), .B2(n9979), .ZN(
        P1_U3531) );
  INV_X1 U11082 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9976) );
  AOI22_X1 U11083 ( .A1(n9978), .A2(n9977), .B1(n9976), .B2(n9979), .ZN(
        P1_U3532) );
  AOI22_X1 U11084 ( .A1(n9978), .A2(n9980), .B1(n7698), .B2(n9979), .ZN(
        P1_U3535) );
  OAI211_X1 U11085 ( .C1(n9984), .C2(n9983), .A(n9982), .B(n9981), .ZN(n9985)
         );
  INV_X1 U11086 ( .A(n9985), .ZN(n9995) );
  OAI21_X1 U11087 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(n9989) );
  AOI22_X1 U11088 ( .A1(n9991), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n9990), .B2(
        n9989), .ZN(n9992) );
  OAI21_X1 U11089 ( .B1(n9993), .B2(n4286), .A(n9992), .ZN(n9994) );
  NOR2_X1 U11090 ( .A1(n9995), .A2(n9994), .ZN(n10002) );
  OAI21_X1 U11091 ( .B1(n9998), .B2(n9997), .A(n9996), .ZN(n9999) );
  NAND2_X1 U11092 ( .A1(n10000), .A2(n9999), .ZN(n10001) );
  OAI211_X1 U11093 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6525), .A(n10002), .B(
        n10001), .ZN(P2_U3184) );
  AOI21_X1 U11094 ( .B1(n10004), .B2(n10028), .A(n10003), .ZN(n10005) );
  AOI211_X1 U11095 ( .C1(n10007), .C2(n10062), .A(n10006), .B(n10005), .ZN(
        n10082) );
  INV_X1 U11096 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10008) );
  AOI22_X1 U11097 ( .A1(n10080), .A2(n10082), .B1(n10008), .B2(n10078), .ZN(
        P2_U3390) );
  OAI211_X1 U11098 ( .C1(n10028), .C2(n10011), .A(n10010), .B(n10009), .ZN(
        n10012) );
  INV_X1 U11099 ( .A(n10012), .ZN(n10084) );
  INV_X1 U11100 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10013) );
  AOI22_X1 U11101 ( .A1(n10080), .A2(n10084), .B1(n10013), .B2(n10078), .ZN(
        P2_U3393) );
  INV_X1 U11102 ( .A(n10014), .ZN(n10017) );
  INV_X1 U11103 ( .A(n10015), .ZN(n10016) );
  AOI211_X1 U11104 ( .C1(n10032), .C2(n10018), .A(n10017), .B(n10016), .ZN(
        n10086) );
  INV_X1 U11105 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10019) );
  AOI22_X1 U11106 ( .A1(n10080), .A2(n10086), .B1(n10019), .B2(n10078), .ZN(
        P2_U3396) );
  NOR2_X1 U11107 ( .A1(n10020), .A2(n10072), .ZN(n10022) );
  AOI211_X1 U11108 ( .C1(n10070), .C2(n10023), .A(n10022), .B(n10021), .ZN(
        n10088) );
  INV_X1 U11109 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10024) );
  AOI22_X1 U11110 ( .A1(n10080), .A2(n10088), .B1(n10024), .B2(n10078), .ZN(
        P2_U3399) );
  OAI211_X1 U11111 ( .C1(n10028), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10029) );
  INV_X1 U11112 ( .A(n10029), .ZN(n10090) );
  AOI22_X1 U11113 ( .A1(n10080), .A2(n10090), .B1(n10030), .B2(n10078), .ZN(
        P2_U3402) );
  AOI21_X1 U11114 ( .B1(n10033), .B2(n10032), .A(n10031), .ZN(n10034) );
  AND2_X1 U11115 ( .A1(n10035), .A2(n10034), .ZN(n10092) );
  INV_X1 U11116 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U11117 ( .A1(n10080), .A2(n10092), .B1(n10036), .B2(n10078), .ZN(
        P2_U3405) );
  INV_X1 U11118 ( .A(n10037), .ZN(n10041) );
  OAI21_X1 U11119 ( .B1(n10039), .B2(n10072), .A(n10038), .ZN(n10040) );
  AOI21_X1 U11120 ( .B1(n10070), .B2(n10041), .A(n10040), .ZN(n10094) );
  INV_X1 U11121 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10042) );
  AOI22_X1 U11122 ( .A1(n10080), .A2(n10094), .B1(n10042), .B2(n10078), .ZN(
        P2_U3408) );
  OAI22_X1 U11123 ( .A1(n10044), .A2(n10057), .B1(n10043), .B2(n10072), .ZN(
        n10045) );
  NOR2_X1 U11124 ( .A1(n10046), .A2(n10045), .ZN(n10096) );
  INV_X1 U11125 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10047) );
  AOI22_X1 U11126 ( .A1(n10080), .A2(n10096), .B1(n10047), .B2(n10078), .ZN(
        P2_U3411) );
  AOI211_X1 U11127 ( .C1(n10070), .C2(n10050), .A(n10049), .B(n10048), .ZN(
        n10098) );
  INV_X1 U11128 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10051) );
  AOI22_X1 U11129 ( .A1(n10080), .A2(n10098), .B1(n10051), .B2(n10078), .ZN(
        P2_U3414) );
  NOR2_X1 U11130 ( .A1(n10052), .A2(n10057), .ZN(n10054) );
  AOI211_X1 U11131 ( .C1(n10062), .C2(n10055), .A(n10054), .B(n10053), .ZN(
        n10100) );
  INV_X1 U11132 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10056) );
  AOI22_X1 U11133 ( .A1(n10080), .A2(n10100), .B1(n10056), .B2(n10078), .ZN(
        P2_U3417) );
  NOR2_X1 U11134 ( .A1(n10058), .A2(n10057), .ZN(n10060) );
  AOI211_X1 U11135 ( .C1(n10062), .C2(n10061), .A(n10060), .B(n10059), .ZN(
        n10102) );
  INV_X1 U11136 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10063) );
  AOI22_X1 U11137 ( .A1(n10080), .A2(n10102), .B1(n10063), .B2(n10078), .ZN(
        P2_U3420) );
  AND2_X1 U11138 ( .A1(n10064), .A2(n10070), .ZN(n10065) );
  NOR3_X1 U11139 ( .A1(n10067), .A2(n10066), .A3(n10065), .ZN(n10104) );
  INV_X1 U11140 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10068) );
  AOI22_X1 U11141 ( .A1(n10080), .A2(n10104), .B1(n10068), .B2(n10078), .ZN(
        P2_U3423) );
  AND3_X1 U11142 ( .A1(n7492), .A2(n10070), .A3(n10069), .ZN(n10076) );
  INV_X1 U11143 ( .A(n10071), .ZN(n10073) );
  NOR2_X1 U11144 ( .A1(n10073), .A2(n10072), .ZN(n10074) );
  NOR4_X1 U11145 ( .A1(n10077), .A2(n10076), .A3(n10075), .A4(n10074), .ZN(
        n10106) );
  INV_X1 U11146 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10079) );
  AOI22_X1 U11147 ( .A1(n10080), .A2(n10106), .B1(n10079), .B2(n10078), .ZN(
        P2_U3426) );
  AOI22_X1 U11148 ( .A1(n10107), .A2(n10082), .B1(n10081), .B2(n6337), .ZN(
        P2_U3459) );
  AOI22_X1 U11149 ( .A1(n10107), .A2(n10084), .B1(n10083), .B2(n6337), .ZN(
        P2_U3460) );
  AOI22_X1 U11150 ( .A1(n10107), .A2(n10086), .B1(n10085), .B2(n6337), .ZN(
        P2_U3461) );
  AOI22_X1 U11151 ( .A1(n10107), .A2(n10088), .B1(n10087), .B2(n6337), .ZN(
        P2_U3462) );
  INV_X1 U11152 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10089) );
  AOI22_X1 U11153 ( .A1(n10107), .A2(n10090), .B1(n10089), .B2(n6337), .ZN(
        P2_U3463) );
  AOI22_X1 U11154 ( .A1(n10107), .A2(n10092), .B1(n10091), .B2(n6337), .ZN(
        P2_U3464) );
  AOI22_X1 U11155 ( .A1(n10107), .A2(n10094), .B1(n10093), .B2(n6337), .ZN(
        P2_U3465) );
  AOI22_X1 U11156 ( .A1(n10107), .A2(n10096), .B1(n10095), .B2(n6337), .ZN(
        P2_U3466) );
  AOI22_X1 U11157 ( .A1(n10107), .A2(n10098), .B1(n10097), .B2(n6337), .ZN(
        P2_U3467) );
  AOI22_X1 U11158 ( .A1(n10107), .A2(n10100), .B1(n10099), .B2(n6337), .ZN(
        P2_U3468) );
  AOI22_X1 U11159 ( .A1(n10107), .A2(n10102), .B1(n10101), .B2(n6337), .ZN(
        P2_U3469) );
  AOI22_X1 U11160 ( .A1(n10107), .A2(n10104), .B1(n10103), .B2(n6337), .ZN(
        P2_U3470) );
  INV_X1 U11161 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U11162 ( .A1(n10107), .A2(n10106), .B1(n10105), .B2(n6337), .ZN(
        P2_U3471) );
  OAI222_X1 U11163 ( .A1(n10112), .A2(n10111), .B1(n10112), .B2(n10110), .C1(
        n10109), .C2(n10108), .ZN(ADD_1068_U5) );
  XOR2_X1 U11164 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11165 ( .B1(n10115), .B2(n10114), .A(n10113), .ZN(n10117) );
  XNOR2_X1 U11166 ( .A(n10117), .B(n10116), .ZN(ADD_1068_U55) );
  OAI21_X1 U11167 ( .B1(n10120), .B2(n10119), .A(n10118), .ZN(ADD_1068_U56) );
  OAI21_X1 U11168 ( .B1(n10123), .B2(n10122), .A(n10121), .ZN(ADD_1068_U57) );
  OAI21_X1 U11169 ( .B1(n10126), .B2(n10125), .A(n10124), .ZN(ADD_1068_U58) );
  OAI21_X1 U11170 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(ADD_1068_U59) );
  OAI21_X1 U11171 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(ADD_1068_U60) );
  OAI21_X1 U11172 ( .B1(n10135), .B2(n10134), .A(n10133), .ZN(ADD_1068_U61) );
  OAI21_X1 U11173 ( .B1(n10138), .B2(n10137), .A(n10136), .ZN(ADD_1068_U62) );
  OAI21_X1 U11174 ( .B1(n10141), .B2(n10140), .A(n10139), .ZN(ADD_1068_U63) );
  OAI21_X1 U11175 ( .B1(n10144), .B2(n10143), .A(n10142), .ZN(ADD_1068_U50) );
  OAI21_X1 U11176 ( .B1(n10147), .B2(n10146), .A(n10145), .ZN(ADD_1068_U51) );
  OAI21_X1 U11177 ( .B1(n10150), .B2(n10149), .A(n10148), .ZN(ADD_1068_U47) );
  OAI21_X1 U11178 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(ADD_1068_U49) );
  OAI21_X1 U11179 ( .B1(n10156), .B2(n10155), .A(n10154), .ZN(ADD_1068_U48) );
  AOI21_X1 U11180 ( .B1(n10159), .B2(n10158), .A(n10157), .ZN(ADD_1068_U54) );
  AOI21_X1 U11181 ( .B1(n10162), .B2(n10161), .A(n10160), .ZN(ADD_1068_U53) );
  OAI21_X1 U11182 ( .B1(n10165), .B2(n10164), .A(n10163), .ZN(ADD_1068_U52) );
  CLKBUF_X2 U4795 ( .A(n6028), .Z(n7755) );
  CLKBUF_X1 U4801 ( .A(n5105), .Z(n7985) );
  AND3_X1 U4815 ( .A1(n5970), .A2(n5969), .A3(n5968), .ZN(n6459) );
  CLKBUF_X1 U4859 ( .A(n5833), .Z(n4286) );
endmodule

