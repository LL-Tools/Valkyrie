

module b14_C_gen_AntiSAT_k_128_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, 
        U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, 
        U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, 
        U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, 
        U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, 
        U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, 
        U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, 
        U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, 
        U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, 
        U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, 
        U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, 
        U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, 
        U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, 
        U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, 
        U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, 
        U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, 
        U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, 
        U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, 
        U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, 
        U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, 
        U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, 
        U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, 
        U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, 
        U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, 
        U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4728, n4729;

  CLKBUF_X2 U2286 ( .A(n2341), .Z(n3230) );
  INV_X1 U2287 ( .A(n3682), .ZN(n2968) );
  INV_X1 U2288 ( .A(n3529), .ZN(n3657) );
  INV_X2 U2289 ( .A(n3579), .ZN(n3529) );
  CLKBUF_X2 U2290 ( .A(n2344), .Z(n3229) );
  INV_X1 U2291 ( .A(n3959), .ZN(n2999) );
  CLKBUF_X3 U2292 ( .A(n2343), .Z(n3234) );
  NAND3_X2 U2293 ( .A1(n4371), .A2(n2678), .A3(n2736), .ZN(n2800) );
  AOI21_X2 U2294 ( .B1(n4377), .B2(n2824), .A(n2823), .ZN(n2914) );
  OAI21_X2 U2295 ( .B1(n4098), .B2(n2578), .A(n2577), .ZN(n4073) );
  OAI21_X2 U2296 ( .B1(n2950), .B2(n2215), .A(n2212), .ZN(n3096) );
  NAND2_X2 U2297 ( .A1(n2942), .A2(n2373), .ZN(n2950) );
  NAND2_X1 U2298 ( .A1(n3332), .A2(n2632), .ZN(n2631) );
  NAND2_X1 U2299 ( .A1(n3726), .A2(n3654), .ZN(n3729) );
  NAND2_X1 U2300 ( .A1(n2109), .A2(n2075), .ZN(n2282) );
  NAND2_X1 U2301 ( .A1(n3846), .A2(n3850), .ZN(n3771) );
  NAND2_X1 U2302 ( .A1(n3630), .A2(n3629), .ZN(n3631) );
  INV_X1 U2303 ( .A(n3628), .ZN(n3629) );
  OAI211_X1 U2304 ( .C1(n3234), .C2(n4300), .A(n2532), .B(n2531), .ZN(n4288)
         );
  INV_X2 U2305 ( .A(n4493), .ZN(n4229) );
  INV_X2 U2306 ( .A(n3540), .ZN(n3684) );
  AND2_X2 U2307 ( .A1(n2968), .A2(n2985), .ZN(n3540) );
  INV_X1 U2308 ( .A(n3065), .ZN(n3958) );
  NAND4_X2 U2309 ( .A1(n2358), .A2(n2357), .A3(n2356), .A4(n2355), .ZN(n3959)
         );
  NAND2_X2 U2310 ( .A1(n2800), .A2(n2799), .ZN(n3682) );
  INV_X2 U2311 ( .A(n2044), .ZN(n2046) );
  NAND4_X1 U2312 ( .A1(n2337), .A2(n2336), .A3(n2335), .A4(n2334), .ZN(n3962)
         );
  INV_X2 U2313 ( .A(n3234), .ZN(n2536) );
  BUF_X2 U2314 ( .A(n2340), .Z(n2601) );
  INV_X1 U2315 ( .A(n2351), .ZN(n2044) );
  INV_X1 U2316 ( .A(n2932), .ZN(n2987) );
  INV_X1 U2317 ( .A(n2677), .ZN(n4371) );
  AND2_X1 U2318 ( .A1(n2309), .A2(n2310), .ZN(n2341) );
  NAND2_X1 U2319 ( .A1(n4370), .A2(n2309), .ZN(n2343) );
  AND2_X1 U2320 ( .A1(n2674), .A2(n2673), .ZN(n2736) );
  INV_X1 U2321 ( .A(n2310), .ZN(n4370) );
  XNOR2_X1 U2322 ( .A(n2302), .B(IR_REG_30__SCAN_IN), .ZN(n2305) );
  NAND2_X1 U2323 ( .A1(n2304), .A2(IR_REG_31__SCAN_IN), .ZN(n2302) );
  XNOR2_X1 U2324 ( .A(n2350), .B(IR_REG_2__SCAN_IN), .ZN(n4381) );
  OR2_X1 U2325 ( .A1(IR_REG_21__SCAN_IN), .A2(n2298), .ZN(n2299) );
  AND2_X1 U2326 ( .A1(n2296), .A2(n2667), .ZN(n2297) );
  XNOR2_X1 U2327 ( .A(n2331), .B(IR_REG_1__SCAN_IN), .ZN(n4382) );
  AND4_X1 U2328 ( .A1(n2421), .A2(n4614), .A3(n2434), .A4(n2437), .ZN(n2290)
         );
  AND4_X1 U2329 ( .A1(n2288), .A2(n2287), .A3(n4696), .A4(n2317), .ZN(n2291)
         );
  NOR2_X1 U2330 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2287)
         );
  NOR2_X1 U2331 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2288)
         );
  INV_X1 U2332 ( .A(IR_REG_22__SCAN_IN), .ZN(n2667) );
  INV_X1 U2333 ( .A(IR_REG_3__SCAN_IN), .ZN(n4696) );
  NOR2_X1 U2334 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2502)
         );
  INV_X2 U2335 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2336 ( .A(n2044), .ZN(n2045) );
  NAND2_X1 U2337 ( .A1(n3548), .A2(n3549), .ZN(n2266) );
  AND2_X1 U2338 ( .A1(n2323), .A2(n2322), .ZN(n2619) );
  NAND2_X1 U2339 ( .A1(n2586), .A2(n2070), .ZN(n2273) );
  AND2_X1 U2340 ( .A1(n2134), .A2(n3903), .ZN(n2141) );
  INV_X1 U2341 ( .A(n2158), .ZN(n2153) );
  NAND2_X1 U2342 ( .A1(n3982), .A2(n2195), .ZN(n2194) );
  NAND2_X1 U2343 ( .A1(n4381), .A2(REG2_REG_2__SCAN_IN), .ZN(n2195) );
  INV_X1 U2344 ( .A(n2255), .ZN(n2254) );
  INV_X1 U2345 ( .A(IR_REG_28__SCAN_IN), .ZN(n2325) );
  AOI21_X1 U2346 ( .B1(n2131), .B2(n2129), .A(n2074), .ZN(n2128) );
  INV_X1 U2347 ( .A(n3788), .ZN(n2129) );
  NAND2_X1 U2348 ( .A1(n2548), .A2(n2547), .ZN(n2560) );
  INV_X1 U2349 ( .A(n2601), .ZN(n2628) );
  AND2_X1 U2350 ( .A1(n2305), .A2(n4370), .ZN(n2340) );
  XNOR2_X1 U2351 ( .A(n2822), .B(n2104), .ZN(n2778) );
  INV_X1 U2352 ( .A(n4377), .ZN(n2104) );
  NAND2_X1 U2353 ( .A1(n4387), .A2(n4388), .ZN(n4386) );
  NAND2_X1 U2354 ( .A1(n4454), .A2(n4040), .ZN(n4042) );
  NAND2_X1 U2355 ( .A1(n2516), .A2(n2147), .ZN(n2146) );
  INV_X1 U2356 ( .A(IR_REG_18__SCAN_IN), .ZN(n2147) );
  OR2_X1 U2357 ( .A1(n2454), .A2(IR_REG_13__SCAN_IN), .ZN(n2504) );
  OR3_X1 U2358 ( .A1(n4113), .A2(n3274), .A3(n3372), .ZN(n2178) );
  OAI21_X1 U2359 ( .B1(n4115), .B2(n2567), .A(n2568), .ZN(n4098) );
  NOR2_X1 U2360 ( .A1(n4312), .A2(n3813), .ZN(n2506) );
  NOR2_X1 U2361 ( .A1(n2464), .A2(n2209), .ZN(n2208) );
  INV_X1 U2362 ( .A(n2452), .ZN(n2209) );
  NOR2_X1 U2363 ( .A1(n3863), .A2(n3949), .ZN(n2464) );
  NAND2_X1 U2364 ( .A1(n2207), .A2(n2205), .ZN(n3398) );
  NOR2_X1 U2365 ( .A1(n2206), .A2(n2283), .ZN(n2205) );
  INV_X1 U2366 ( .A(n2256), .ZN(n3164) );
  INV_X1 U2367 ( .A(n2259), .ZN(n2257) );
  AND2_X1 U2368 ( .A1(n2072), .A2(n2587), .ZN(n2272) );
  AOI22_X1 U2369 ( .A1(n2710), .A2(n4197), .B1(n4056), .B2(n3941), .ZN(n4065)
         );
  NOR2_X2 U2370 ( .A1(n2613), .A2(n2299), .ZN(n2323) );
  AND2_X1 U2371 ( .A1(n2325), .A2(n2322), .ZN(n2303) );
  NOR3_X1 U2372 ( .A1(n2712), .A2(n4540), .A3(n4527), .ZN(n2217) );
  NAND2_X1 U2373 ( .A1(n3524), .A2(n2140), .ZN(n2143) );
  OR2_X1 U2374 ( .A1(n2141), .A2(n2059), .ZN(n2139) );
  AND2_X1 U2375 ( .A1(n2141), .A2(n2142), .ZN(n2137) );
  INV_X1 U2376 ( .A(n3524), .ZN(n2142) );
  NAND2_X1 U2377 ( .A1(n2234), .A2(n3858), .ZN(n2233) );
  NAND2_X1 U2378 ( .A1(n2121), .A2(n2120), .ZN(n2119) );
  INV_X1 U2379 ( .A(n3881), .ZN(n2121) );
  NOR2_X1 U2380 ( .A1(n2154), .A2(n2150), .ZN(n2149) );
  INV_X1 U2381 ( .A(n2155), .ZN(n2154) );
  INV_X1 U2382 ( .A(n3800), .ZN(n2150) );
  NOR2_X1 U2383 ( .A1(n3891), .A2(n2156), .ZN(n2155) );
  INV_X1 U2384 ( .A(n3616), .ZN(n2156) );
  INV_X1 U2385 ( .A(n2279), .ZN(n2277) );
  INV_X1 U2386 ( .A(n3660), .ZN(n2276) );
  INV_X1 U2387 ( .A(n2075), .ZN(n2274) );
  INV_X1 U2388 ( .A(n3654), .ZN(n2278) );
  AND2_X1 U2389 ( .A1(n3576), .A2(n3575), .ZN(n3577) );
  NOR2_X1 U2390 ( .A1(n3871), .A2(n2280), .ZN(n2279) );
  INV_X1 U2391 ( .A(n2281), .ZN(n2280) );
  NOR2_X1 U2392 ( .A1(n3615), .A2(n2159), .ZN(n2158) );
  INV_X1 U2393 ( .A(n3609), .ZN(n2159) );
  AOI21_X1 U2394 ( .B1(n3479), .B2(n2519), .A(n2058), .ZN(n2255) );
  NAND2_X1 U2395 ( .A1(n4288), .A2(n4192), .ZN(n3304) );
  INV_X1 U2396 ( .A(n2385), .ZN(n2214) );
  NAND2_X1 U2397 ( .A1(n4117), .A2(n2088), .ZN(n2093) );
  NOR2_X1 U2398 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2322)
         );
  NOR2_X1 U2399 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2294)
         );
  AOI21_X1 U2400 ( .B1(n2050), .B2(IR_REG_31__SCAN_IN), .A(IR_REG_19__SCAN_IN), 
        .ZN(n2145) );
  INV_X1 U2401 ( .A(n3707), .ZN(n2126) );
  INV_X1 U2402 ( .A(n3789), .ZN(n2132) );
  NAND2_X1 U2403 ( .A1(n2233), .A2(n2231), .ZN(n2230) );
  INV_X1 U2404 ( .A(n3778), .ZN(n2231) );
  AND2_X1 U2405 ( .A1(n2227), .A2(n2115), .ZN(n2114) );
  NOR2_X1 U2406 ( .A1(n2232), .A2(n2228), .ZN(n2227) );
  AOI21_X1 U2407 ( .B1(n2119), .B2(n2117), .A(n2116), .ZN(n2115) );
  INV_X1 U2408 ( .A(n2087), .ZN(n2228) );
  INV_X1 U2409 ( .A(n2119), .ZN(n2118) );
  NOR2_X1 U2410 ( .A1(n3735), .A2(n2271), .ZN(n2270) );
  INV_X1 U2411 ( .A(n3557), .ZN(n2271) );
  INV_X1 U2412 ( .A(n3689), .ZN(n2246) );
  AOI21_X1 U2413 ( .B1(n2249), .B2(n3915), .A(n2248), .ZN(n2247) );
  NOR2_X1 U2414 ( .A1(n3680), .A2(n3681), .ZN(n2248) );
  OR2_X1 U2415 ( .A1(n2441), .A2(n4662), .ZN(n2458) );
  OR2_X1 U2416 ( .A1(n2236), .A2(n2235), .ZN(n2229) );
  NAND2_X1 U2417 ( .A1(n3570), .A2(n2087), .ZN(n2235) );
  INV_X1 U2418 ( .A(n3571), .ZN(n2236) );
  NAND2_X1 U2419 ( .A1(n2282), .A2(n2279), .ZN(n3726) );
  NAND2_X1 U2420 ( .A1(n2160), .A2(n2158), .ZN(n2157) );
  AND4_X1 U2421 ( .A1(n2515), .A2(n2514), .A3(n2513), .A4(n2512), .ZN(n3619)
         );
  AND4_X1 U2422 ( .A1(n2400), .A2(n2399), .A3(n2398), .A4(n2397), .ZN(n3533)
         );
  XNOR2_X1 U2423 ( .A(n2194), .B(n2193), .ZN(n3994) );
  NOR2_X1 U2424 ( .A1(n2777), .A2(n2076), .ZN(n2822) );
  NAND2_X1 U2425 ( .A1(n2185), .A2(n2190), .ZN(n2183) );
  OAI21_X1 U2426 ( .B1(n4028), .B2(n3137), .A(n2096), .ZN(n4387) );
  NAND2_X1 U2427 ( .A1(n4398), .A2(REG2_REG_10__SCAN_IN), .ZN(n4397) );
  NAND2_X1 U2428 ( .A1(n4402), .A2(n4031), .ZN(n4408) );
  NAND2_X1 U2429 ( .A1(n4408), .A2(n4409), .ZN(n4407) );
  NAND2_X1 U2430 ( .A1(n4410), .A2(n4010), .ZN(n4011) );
  NAND2_X1 U2431 ( .A1(n4419), .A2(REG2_REG_12__SCAN_IN), .ZN(n4418) );
  NAND2_X1 U2432 ( .A1(n2182), .A2(n2181), .ZN(n4013) );
  OR2_X1 U2433 ( .A1(n4022), .A2(REG2_REG_13__SCAN_IN), .ZN(n2181) );
  OR2_X1 U2434 ( .A1(n4431), .A2(n4427), .ZN(n2182) );
  NOR2_X1 U2435 ( .A1(n4449), .A2(n2179), .ZN(n4016) );
  AND2_X1 U2436 ( .A1(n4021), .A2(REG2_REG_15__SCAN_IN), .ZN(n2179) );
  NOR2_X1 U2437 ( .A1(n2203), .A2(n4480), .ZN(n4479) );
  AND2_X1 U2438 ( .A1(n3376), .A2(n3508), .ZN(n2177) );
  AND2_X1 U2439 ( .A1(n4066), .A2(n2600), .ZN(n3691) );
  INV_X1 U2440 ( .A(n2570), .ZN(n2569) );
  OR2_X1 U2441 ( .A1(n2560), .A2(n4648), .ZN(n2570) );
  AOI21_X1 U2442 ( .B1(n2164), .B2(n2168), .A(n2163), .ZN(n2162) );
  NAND2_X1 U2443 ( .A1(n4127), .A2(n2557), .ZN(n2237) );
  NAND2_X1 U2444 ( .A1(n4169), .A2(n2539), .ZN(n2268) );
  AND2_X1 U2445 ( .A1(n4212), .A2(n4213), .ZN(n3479) );
  OR2_X1 U2446 ( .A1(n3476), .A2(n3479), .ZN(n3474) );
  NAND2_X1 U2447 ( .A1(n3950), .A2(n2450), .ZN(n2451) );
  NAND2_X1 U2448 ( .A1(n2065), .A2(n2266), .ZN(n2261) );
  NOR2_X1 U2449 ( .A1(n3548), .A2(n3549), .ZN(n2267) );
  NAND2_X1 U2450 ( .A1(n2176), .A2(n3350), .ZN(n3101) );
  NAND2_X1 U2451 ( .A1(n3123), .A2(n3353), .ZN(n2176) );
  NOR2_X1 U2452 ( .A1(n3124), .A2(n3115), .ZN(n2263) );
  OAI21_X1 U2453 ( .B1(n2952), .B2(n2951), .A(n3321), .ZN(n3012) );
  INV_X1 U2454 ( .A(n3956), .ZN(n3527) );
  INV_X1 U2455 ( .A(DATAI_0_), .ZN(n2094) );
  INV_X1 U2456 ( .A(IR_REG_0__SCAN_IN), .ZN(n2095) );
  NAND2_X1 U2457 ( .A1(n2714), .A2(n4063), .ZN(n4239) );
  NOR2_X2 U2458 ( .A1(n2093), .A2(n3690), .ZN(n2714) );
  AND2_X1 U2459 ( .A1(n2585), .A2(n2584), .ZN(n4262) );
  OR2_X1 U2460 ( .A1(n4088), .A2(n2628), .ZN(n2585) );
  INV_X1 U2461 ( .A(n3909), .ZN(n3526) );
  AND4_X1 U2462 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n3053)
         );
  NAND2_X1 U2463 ( .A1(n3269), .A2(n2657), .ZN(n4197) );
  INV_X1 U2464 ( .A(n3057), .ZN(n3068) );
  AND2_X1 U2465 ( .A1(n2618), .A2(n2865), .ZN(n4317) );
  NAND2_X1 U2466 ( .A1(n2675), .A2(n2736), .ZN(n2732) );
  NAND2_X1 U2467 ( .A1(n2304), .A2(n2169), .ZN(n2310) );
  AOI21_X1 U2468 ( .B1(n2622), .B2(n2061), .A(n2170), .ZN(n2169) );
  NOR2_X1 U2469 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2170)
         );
  NAND2_X1 U2470 ( .A1(n2673), .A2(n2321), .ZN(n2705) );
  AND2_X1 U2471 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2321)
         );
  NAND2_X1 U2472 ( .A1(n2269), .A2(IR_REG_31__SCAN_IN), .ZN(n2680) );
  NOR2_X1 U2473 ( .A1(n2613), .A2(IR_REG_21__SCAN_IN), .ZN(n2668) );
  NOR2_X1 U2474 ( .A1(n2504), .A2(n2503), .ZN(n2517) );
  INV_X1 U2475 ( .A(IR_REG_7__SCAN_IN), .ZN(n2402) );
  OR2_X1 U2476 ( .A1(n2382), .A2(IR_REG_5__SCAN_IN), .ZN(n2401) );
  AND2_X1 U2477 ( .A1(n2241), .A2(n2083), .ZN(n2239) );
  AND2_X1 U2478 ( .A1(n2242), .A2(n3929), .ZN(n2241) );
  OAI21_X1 U2479 ( .B1(n2247), .B2(n3689), .A(n2243), .ZN(n2242) );
  NAND2_X1 U2480 ( .A1(n2247), .A2(n2244), .ZN(n2243) );
  NAND2_X1 U2481 ( .A1(n2250), .A2(n2246), .ZN(n2244) );
  NAND2_X1 U2482 ( .A1(n2247), .A2(n2246), .ZN(n2245) );
  NAND2_X1 U2483 ( .A1(n3056), .A2(n3055), .ZN(n3525) );
  AND2_X1 U2484 ( .A1(n2510), .A2(n2496), .ZN(n3814) );
  NAND2_X1 U2485 ( .A1(n2133), .A2(n3789), .ZN(n3917) );
  AND2_X1 U2486 ( .A1(n2861), .A2(n2860), .ZN(n3934) );
  AND2_X1 U2487 ( .A1(n2861), .A2(n2809), .ZN(n3931) );
  NAND2_X1 U2488 ( .A1(n2593), .A2(n2592), .ZN(n3943) );
  NAND2_X1 U2489 ( .A1(n2761), .A2(n2762), .ZN(n3982) );
  AND2_X1 U2490 ( .A1(n2106), .A2(n2105), .ZN(n2777) );
  INV_X1 U2491 ( .A(n2758), .ZN(n2105) );
  NAND2_X1 U2492 ( .A1(n4411), .A2(n4412), .ZN(n4410) );
  XNOR2_X1 U2493 ( .A(n4016), .B(n4041), .ZN(n4461) );
  NAND2_X1 U2494 ( .A1(n4461), .A2(n4459), .ZN(n4460) );
  NOR2_X1 U2495 ( .A1(n4465), .A2(n4043), .ZN(n4474) );
  OAI21_X1 U2496 ( .B1(n4479), .B2(n2201), .A(n2200), .ZN(n2199) );
  AOI21_X1 U2497 ( .B1(n4482), .B2(ADDR_REG_18__SCAN_IN), .A(n4481), .ZN(n2200) );
  NAND2_X1 U2498 ( .A1(n2202), .A2(n4429), .ZN(n2201) );
  NAND2_X1 U2499 ( .A1(n2203), .A2(n4480), .ZN(n2202) );
  XNOR2_X1 U2500 ( .A(n2609), .B(n2608), .ZN(n4051) );
  AND2_X1 U2501 ( .A1(n2768), .A2(n2765), .ZN(n4484) );
  OAI211_X1 U2502 ( .C1(n2701), .C2(n2223), .A(n2220), .B(n2218), .ZN(n4061)
         );
  INV_X1 U2503 ( .A(n2224), .ZN(n2223) );
  AND2_X1 U2504 ( .A1(n2221), .A2(n2225), .ZN(n2220) );
  AND2_X1 U2505 ( .A1(n4061), .A2(n4527), .ZN(n2173) );
  NAND2_X1 U2506 ( .A1(n4065), .A2(n2174), .ZN(n2712) );
  AND2_X1 U2507 ( .A1(n2711), .A2(n2175), .ZN(n2174) );
  NAND2_X1 U2508 ( .A1(n4310), .A2(n3258), .ZN(n2175) );
  NOR2_X1 U2509 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2292)
         );
  NOR2_X1 U2510 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2293)
         );
  INV_X1 U2511 ( .A(IR_REG_10__SCAN_IN), .ZN(n2434) );
  INV_X1 U2512 ( .A(IR_REG_8__SCAN_IN), .ZN(n4613) );
  AND2_X1 U2513 ( .A1(n3881), .A2(n3880), .ZN(n2116) );
  INV_X1 U2514 ( .A(n3566), .ZN(n2117) );
  INV_X1 U2515 ( .A(n2233), .ZN(n2232) );
  INV_X1 U2516 ( .A(n3880), .ZN(n2120) );
  INV_X1 U2517 ( .A(n3627), .ZN(n3630) );
  AND2_X1 U2518 ( .A1(n2414), .A2(REG3_REG_10__SCAN_IN), .ZN(n2426) );
  INV_X1 U2519 ( .A(n2415), .ZN(n2414) );
  INV_X1 U2520 ( .A(n2187), .ZN(n2185) );
  INV_X1 U2521 ( .A(n3248), .ZN(n2163) );
  OAI21_X1 U2522 ( .B1(n2261), .B2(n2260), .A(n2062), .ZN(n2259) );
  INV_X1 U2523 ( .A(n2425), .ZN(n2260) );
  NAND2_X1 U2524 ( .A1(n3345), .A2(n3341), .ZN(n2938) );
  INV_X1 U2525 ( .A(n2732), .ZN(n2689) );
  INV_X1 U2526 ( .A(n3317), .ZN(n2222) );
  NOR2_X1 U2527 ( .A1(n4080), .A2(n4258), .ZN(n2092) );
  AND2_X1 U2528 ( .A1(n2046), .A2(DATAI_20_), .ZN(n4192) );
  NOR2_X1 U2529 ( .A1(n3131), .A2(n3762), .ZN(n2091) );
  NOR2_X1 U2530 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2660)
         );
  INV_X1 U2531 ( .A(IR_REG_16__SCAN_IN), .ZN(n2501) );
  INV_X1 U2532 ( .A(IR_REG_9__SCAN_IN), .ZN(n2421) );
  INV_X1 U2533 ( .A(IR_REG_2__SCAN_IN), .ZN(n2289) );
  XNOR2_X1 U2534 ( .A(n4603), .B(keyinput_g27), .ZN(n2198) );
  XNOR2_X1 U2535 ( .A(n2197), .B(IR_REG_1__SCAN_IN), .ZN(n2196) );
  INV_X1 U2536 ( .A(keyinput_g56), .ZN(n2197) );
  INV_X1 U2537 ( .A(IR_REG_4__SCAN_IN), .ZN(n4614) );
  XNOR2_X1 U2538 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_f56), .ZN(n4585) );
  NAND2_X1 U2539 ( .A1(n2138), .A2(n2136), .ZN(n3698) );
  NOR2_X1 U2540 ( .A1(n2137), .A2(n2060), .ZN(n2136) );
  NAND2_X1 U2541 ( .A1(n3056), .A2(n2139), .ZN(n2138) );
  AOI21_X1 U2542 ( .B1(n2153), .B2(n2155), .A(n2152), .ZN(n2151) );
  INV_X1 U2543 ( .A(n3892), .ZN(n2152) );
  AND2_X1 U2544 ( .A1(n2799), .A2(n2849), .ZN(n3667) );
  INV_X1 U2545 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4662) );
  OAI21_X1 U2546 ( .B1(n2110), .B2(n2113), .A(n3881), .ZN(n3571) );
  NAND2_X1 U2547 ( .A1(n3566), .A2(n2120), .ZN(n2113) );
  NAND2_X1 U2548 ( .A1(n3883), .A2(n3880), .ZN(n3570) );
  INV_X1 U2549 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U2550 ( .A1(n3729), .A2(n2286), .ZN(n3819) );
  AOI21_X1 U2551 ( .B1(n3654), .B2(n2277), .A(n2276), .ZN(n2275) );
  AOI21_X1 U2552 ( .B1(n3540), .B2(n3962), .A(n2802), .ZN(n2804) );
  OAI21_X1 U2553 ( .B1(n3579), .B2(n2867), .A(n2801), .ZN(n2802) );
  NAND2_X1 U2554 ( .A1(n2973), .A2(IR_REG_0__SCAN_IN), .ZN(n2801) );
  NAND2_X1 U2555 ( .A1(n3769), .A2(n3768), .ZN(n2281) );
  INV_X1 U2556 ( .A(n3771), .ZN(n2109) );
  NAND2_X1 U2557 ( .A1(n3737), .A2(n3566), .ZN(n3883) );
  NAND2_X1 U2558 ( .A1(n2808), .A2(n3540), .ZN(n2853) );
  NOR2_X1 U2559 ( .A1(n2387), .A2(n2775), .ZN(n2395) );
  INV_X1 U2560 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2775) );
  AOI21_X1 U2561 ( .B1(n3994), .B2(REG2_REG_3__SCAN_IN), .A(n2064), .ZN(n2763)
         );
  OR2_X1 U2562 ( .A1(n2756), .A2(n2107), .ZN(n2106) );
  AND2_X1 U2563 ( .A1(n2757), .A2(n4379), .ZN(n2107) );
  AOI21_X1 U2564 ( .B1(n2192), .B2(n2188), .A(n2820), .ZN(n2187) );
  INV_X1 U2565 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2188) );
  XNOR2_X1 U2566 ( .A(n4005), .B(n4027), .ZN(n4006) );
  NAND2_X1 U2567 ( .A1(n4386), .A2(n4029), .ZN(n4030) );
  NAND2_X1 U2568 ( .A1(n4407), .A2(n4032), .ZN(n4034) );
  NAND2_X1 U2569 ( .A1(n4469), .A2(n2204), .ZN(n2203) );
  OR2_X1 U2570 ( .A1(n4044), .A2(REG2_REG_17__SCAN_IN), .ZN(n2204) );
  INV_X1 U2571 ( .A(n4048), .ZN(n2100) );
  NOR2_X1 U2572 ( .A1(n2103), .A2(n4048), .ZN(n2099) );
  OR2_X1 U2573 ( .A1(n4113), .A2(n3274), .ZN(n4094) );
  AND2_X1 U2574 ( .A1(n2566), .A2(n2565), .ZN(n4134) );
  NAND2_X1 U2575 ( .A1(n2165), .A2(n3369), .ZN(n4167) );
  NAND2_X1 U2576 ( .A1(n2167), .A2(n2166), .ZN(n2165) );
  AOI21_X1 U2577 ( .B1(n2255), .B2(n2253), .A(n2078), .ZN(n2252) );
  INV_X1 U2578 ( .A(n2519), .ZN(n2253) );
  NAND2_X1 U2579 ( .A1(n2167), .A2(n2054), .ZN(n4189) );
  INV_X1 U2580 ( .A(n3945), .ZN(n4195) );
  NAND2_X1 U2581 ( .A1(n2167), .A2(n2053), .ZN(n3478) );
  OR2_X1 U2582 ( .A1(n3429), .A2(n3432), .ZN(n3430) );
  NAND2_X1 U2583 ( .A1(n3572), .A2(n3574), .ZN(n2452) );
  OAI21_X1 U2584 ( .B1(n3101), .B2(n3100), .A(n3354), .ZN(n3142) );
  AND2_X1 U2585 ( .A1(n2395), .A2(REG3_REG_7__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U2586 ( .A1(n2637), .A2(n3351), .ZN(n3123) );
  OR2_X1 U2587 ( .A1(n3084), .A2(n2636), .ZN(n2637) );
  NAND2_X1 U2588 ( .A1(n2057), .A2(n2386), .ZN(n2215) );
  AND2_X1 U2589 ( .A1(n2213), .A2(n2394), .ZN(n2212) );
  AND2_X1 U2590 ( .A1(n2635), .A2(n3351), .ZN(n3348) );
  INV_X1 U2591 ( .A(n3701), .ZN(n3532) );
  OAI21_X1 U2592 ( .B1(n2939), .B2(n2633), .A(n3345), .ZN(n2952) );
  NAND2_X1 U2593 ( .A1(n2904), .A2(n3340), .ZN(n2939) );
  INV_X1 U2594 ( .A(n2938), .ZN(n3296) );
  AND2_X1 U2595 ( .A1(n4493), .A2(n4311), .ZN(n4175) );
  AND2_X1 U2596 ( .A1(n3340), .A2(n3337), .ZN(n3300) );
  NAND2_X1 U2597 ( .A1(n3338), .A2(n3335), .ZN(n2882) );
  INV_X1 U2598 ( .A(n2631), .ZN(n3297) );
  NAND2_X1 U2599 ( .A1(n3297), .A2(n2171), .ZN(n2926) );
  NOR2_X1 U2600 ( .A1(n3318), .A2(n2222), .ZN(n2219) );
  NAND2_X1 U2601 ( .A1(n2226), .A2(n2069), .ZN(n2225) );
  NOR2_X1 U2602 ( .A1(n2226), .A2(n2069), .ZN(n2224) );
  NOR2_X1 U2603 ( .A1(n4239), .A2(n4242), .ZN(n4238) );
  NAND2_X1 U2604 ( .A1(n4117), .A2(n2092), .ZN(n4084) );
  NAND2_X1 U2605 ( .A1(n4117), .A2(n4100), .ZN(n4099) );
  AND2_X1 U2606 ( .A1(n4140), .A2(n4267), .ZN(n4117) );
  AND2_X1 U2607 ( .A1(n4158), .A2(n4138), .ZN(n4140) );
  NOR2_X1 U2608 ( .A1(n4172), .A2(n3648), .ZN(n4158) );
  OR2_X1 U2609 ( .A1(n4201), .A2(n4286), .ZN(n4172) );
  INV_X1 U2610 ( .A(n4192), .ZN(n4202) );
  OR2_X1 U2611 ( .A1(n4224), .A2(n4192), .ZN(n4201) );
  NOR2_X1 U2612 ( .A1(n2090), .A2(n3897), .ZN(n4226) );
  NAND2_X1 U2613 ( .A1(n4226), .A2(n4225), .ZN(n4224) );
  AND4_X1 U2614 ( .A1(n2490), .A2(n2489), .A3(n2488), .A4(n2487), .ZN(n3602)
         );
  NAND2_X1 U2615 ( .A1(n3435), .A2(n3593), .ZN(n3434) );
  AND4_X1 U2616 ( .A1(n2470), .A2(n2469), .A3(n2468), .A4(n2467), .ZN(n3585)
         );
  AND2_X1 U2617 ( .A1(n3402), .A2(n3583), .ZN(n3435) );
  INV_X1 U2618 ( .A(n3719), .ZN(n3583) );
  NOR2_X1 U2619 ( .A1(n3221), .A2(n3863), .ZN(n3402) );
  OR2_X1 U2620 ( .A1(n3182), .A2(n2450), .ZN(n3221) );
  NAND2_X1 U2621 ( .A1(n3169), .A2(n3567), .ZN(n3182) );
  AND4_X1 U2622 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2417), .ZN(n3561)
         );
  NOR2_X1 U2623 ( .A1(n3146), .A2(n3740), .ZN(n3169) );
  NAND2_X1 U2624 ( .A1(n2091), .A2(n3548), .ZN(n3146) );
  NAND2_X1 U2625 ( .A1(n3089), .A2(n3532), .ZN(n3131) );
  INV_X1 U2626 ( .A(n2091), .ZN(n3133) );
  AND2_X1 U2627 ( .A1(n3016), .A2(n3526), .ZN(n3089) );
  NAND2_X1 U2628 ( .A1(n2937), .A2(n3046), .ZN(n2956) );
  NOR2_X1 U2629 ( .A1(n2956), .A2(n3068), .ZN(n3016) );
  AND2_X1 U2630 ( .A1(n2909), .A2(n3077), .ZN(n2937) );
  NAND2_X1 U2631 ( .A1(n2987), .A2(n2867), .ZN(n2934) );
  AND2_X1 U2632 ( .A1(n2728), .A2(n2790), .ZN(n4287) );
  INV_X1 U2633 ( .A(IR_REG_27__SCAN_IN), .ZN(n2324) );
  INV_X1 U2634 ( .A(IR_REG_26__SCAN_IN), .ZN(n2320) );
  INV_X1 U2635 ( .A(IR_REG_20__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U2636 ( .A1(n2610), .A2(IR_REG_31__SCAN_IN), .ZN(n2612) );
  AND2_X1 U2637 ( .A1(n2491), .A2(n2482), .ZN(n4021) );
  AND2_X1 U2638 ( .A1(n2198), .A2(n2196), .ZN(n4679) );
  OAI21_X1 U2639 ( .B1(n2128), .B2(n3707), .A(n2124), .ZN(n2123) );
  NAND2_X1 U2640 ( .A1(n2128), .A2(n2125), .ZN(n2124) );
  NAND2_X1 U2641 ( .A1(n2130), .A2(n2126), .ZN(n2125) );
  NAND2_X1 U2642 ( .A1(n2131), .A2(n3707), .ZN(n2127) );
  AOI21_X1 U2643 ( .B1(n2114), .B2(n2118), .A(n2080), .ZN(n2111) );
  INV_X1 U2644 ( .A(n2114), .ZN(n2112) );
  AND2_X1 U2645 ( .A1(n2474), .A2(n2466), .ZN(n3723) );
  INV_X1 U2646 ( .A(n3559), .ZN(n3740) );
  NAND2_X1 U2647 ( .A1(n3558), .A2(n3557), .ZN(n3736) );
  NAND2_X1 U2648 ( .A1(n2967), .A2(n2966), .ZN(n3043) );
  OR2_X1 U2649 ( .A1(n2965), .A2(n2964), .ZN(n2966) );
  AND2_X1 U2650 ( .A1(n2556), .A2(n2555), .ZN(n4151) );
  OR2_X1 U2651 ( .A1(n4141), .A2(n2628), .ZN(n2556) );
  NAND2_X1 U2652 ( .A1(n2229), .A2(n3778), .ZN(n3861) );
  INV_X1 U2653 ( .A(n3934), .ZN(n3919) );
  NAND2_X1 U2654 ( .A1(n2282), .A2(n2281), .ZN(n3870) );
  NAND2_X1 U2655 ( .A1(n2895), .A2(n2896), .ZN(n2967) );
  NAND2_X1 U2656 ( .A1(n2157), .A2(n3616), .ZN(n3895) );
  NAND2_X1 U2657 ( .A1(n3525), .A2(n3524), .ZN(n3906) );
  NAND2_X1 U2658 ( .A1(n2977), .A2(n2976), .ZN(n3936) );
  NAND2_X1 U2659 ( .A1(n2813), .A2(n4490), .ZN(n3933) );
  AND2_X1 U2660 ( .A1(n3529), .A2(n2788), .ZN(n3391) );
  NAND2_X1 U2661 ( .A1(n2576), .A2(n2575), .ZN(n4119) );
  OR2_X1 U2662 ( .A1(n4104), .A2(n2628), .ZN(n2576) );
  INV_X1 U2663 ( .A(n4134), .ZN(n4259) );
  NAND2_X1 U2664 ( .A1(n2545), .A2(n2544), .ZN(n4176) );
  OAI211_X1 U2665 ( .C1(n3772), .C2(n2628), .A(n2538), .B(n2537), .ZN(n4193)
         );
  OR2_X1 U2666 ( .A1(n4204), .A2(n2628), .ZN(n2532) );
  INV_X1 U2667 ( .A(n3619), .ZN(n4220) );
  NAND4_X1 U2668 ( .A1(n2500), .A2(n2499), .A3(n2498), .A4(n2497), .ZN(n4312)
         );
  INV_X1 U2669 ( .A(n3602), .ZN(n3946) );
  INV_X1 U2670 ( .A(n3561), .ZN(n3952) );
  CLKBUF_X2 U2671 ( .A(U4043), .Z(n3961) );
  INV_X1 U2672 ( .A(n2106), .ZN(n2759) );
  AOI21_X1 U2673 ( .B1(n2819), .B2(REG2_REG_6__SCAN_IN), .A(n2189), .ZN(n2821)
         );
  NAND2_X1 U2674 ( .A1(n4397), .A2(n4009), .ZN(n4411) );
  XNOR2_X1 U2675 ( .A(n4034), .B(n4510), .ZN(n4424) );
  NAND2_X1 U2676 ( .A1(n4418), .A2(n4012), .ZN(n4431) );
  XNOR2_X1 U2677 ( .A(n4013), .B(n2180), .ZN(n4441) );
  XNOR2_X1 U2678 ( .A(n4042), .B(n4041), .ZN(n4464) );
  NOR2_X1 U2679 ( .A1(n4464), .A2(REG1_REG_16__SCAN_IN), .ZN(n4465) );
  NAND2_X1 U2680 ( .A1(n4460), .A2(n4017), .ZN(n4468) );
  AND2_X1 U2681 ( .A1(n2747), .A2(n2746), .ZN(n4482) );
  NAND2_X1 U2682 ( .A1(n4486), .A2(n2102), .ZN(n2101) );
  AOI22_X1 U2683 ( .A1(n2101), .A2(n2099), .B1(n4048), .B2(n2103), .ZN(n2098)
         );
  AND2_X1 U2684 ( .A1(n4493), .A2(n4287), .ZN(n4174) );
  NAND2_X1 U2685 ( .A1(n2273), .A2(n2587), .ZN(n3501) );
  AND2_X1 U2686 ( .A1(n2178), .A2(n3376), .ZN(n3507) );
  AND2_X1 U2687 ( .A1(n2607), .A2(n2606), .ZN(n3685) );
  CLKBUF_X1 U2688 ( .A(n4154), .Z(n4155) );
  NAND2_X1 U2689 ( .A1(n3474), .A2(n2519), .ZN(n4211) );
  AND2_X1 U2690 ( .A1(n2207), .A2(n2210), .ZN(n3400) );
  NAND2_X1 U2691 ( .A1(n2258), .A2(n2261), .ZN(n3141) );
  NAND2_X1 U2692 ( .A1(n2265), .A2(n2049), .ZN(n2258) );
  INV_X1 U2693 ( .A(n2263), .ZN(n2262) );
  NAND2_X1 U2694 ( .A1(n2265), .A2(n2048), .ZN(n2264) );
  NAND2_X1 U2695 ( .A1(n2812), .A2(n2811), .ZN(n4490) );
  NAND2_X1 U2696 ( .A1(n2211), .A2(n2386), .ZN(n3011) );
  NAND2_X1 U2697 ( .A1(n2950), .A2(n2385), .ZN(n2211) );
  INV_X1 U2698 ( .A(n2980), .ZN(n3077) );
  INV_X1 U2699 ( .A(n4234), .ZN(n4171) );
  OAI21_X1 U2700 ( .B1(n2631), .B2(n2924), .A(n2923), .ZN(n2994) );
  INV_X1 U2701 ( .A(n4231), .ZN(n4497) );
  OR2_X1 U2702 ( .A1(n2714), .A2(n2695), .ZN(n3513) );
  INV_X2 U2703 ( .A(n4534), .ZN(n4536) );
  NAND2_X1 U2704 ( .A1(n2732), .A2(n2811), .ZN(n4503) );
  AND2_X1 U2705 ( .A1(n2300), .A2(n2303), .ZN(n2301) );
  INV_X1 U2706 ( .A(IR_REG_29__SCAN_IN), .ZN(n2300) );
  NAND2_X1 U2707 ( .A1(n2669), .A2(IR_REG_31__SCAN_IN), .ZN(n2670) );
  AND2_X1 U2708 ( .A1(n2743), .A2(STATE_REG_SCAN_IN), .ZN(n4504) );
  XNOR2_X1 U2709 ( .A(n2616), .B(IR_REG_22__SCAN_IN), .ZN(n4372) );
  XNOR2_X1 U2710 ( .A(n2614), .B(IR_REG_21__SCAN_IN), .ZN(n4373) );
  INV_X1 U2711 ( .A(n4051), .ZN(n4374) );
  INV_X1 U2712 ( .A(n4033), .ZN(n4510) );
  AND2_X1 U2713 ( .A1(n2412), .A2(n2404), .ZN(n4376) );
  NAND2_X1 U2714 ( .A1(n2108), .A2(IR_REG_31__SCAN_IN), .ZN(n2350) );
  INV_X1 U2715 ( .A(n2349), .ZN(n2108) );
  NAND2_X1 U2716 ( .A1(n2241), .A2(n2245), .ZN(n2240) );
  INV_X1 U2717 ( .A(n2199), .ZN(n4488) );
  OR2_X1 U2718 ( .A1(n4475), .A2(n2101), .ZN(n4483) );
  OR2_X1 U2719 ( .A1(n4067), .A2(n4305), .ZN(n2715) );
  OAI21_X1 U2720 ( .B1(n2712), .B2(n2173), .A(n4536), .ZN(n2172) );
  AND2_X1 U2721 ( .A1(n3435), .A2(n2055), .ZN(n2047) );
  OR2_X1 U2722 ( .A1(n3954), .A2(n3762), .ZN(n2048) );
  AND2_X1 U2723 ( .A1(n2266), .A2(n2048), .ZN(n2049) );
  OR2_X1 U2724 ( .A1(n2503), .A2(n2146), .ZN(n2050) );
  AND4_X1 U2725 ( .A1(n2502), .A2(n2294), .A3(n2293), .A4(n2292), .ZN(n2051)
         );
  AND2_X1 U2726 ( .A1(n3701), .A2(n3955), .ZN(n2052) );
  INV_X1 U2727 ( .A(n3582), .ZN(n3949) );
  NAND2_X1 U2728 ( .A1(n4312), .A2(n3469), .ZN(n2053) );
  INV_X1 U2729 ( .A(n3572), .ZN(n2450) );
  AND2_X1 U2730 ( .A1(n2648), .A2(n2053), .ZN(n2054) );
  AND2_X1 U2731 ( .A1(n3593), .A2(n3601), .ZN(n2055) );
  OR3_X1 U2732 ( .A1(n2504), .A2(n2503), .A3(IR_REG_17__SCAN_IN), .ZN(n2056)
         );
  INV_X1 U2733 ( .A(n4244), .ZN(n4310) );
  OAI21_X1 U2734 ( .B1(n2504), .B2(n2050), .A(IR_REG_31__SCAN_IN), .ZN(n2609)
         );
  XNOR2_X1 U2735 ( .A(n2612), .B(n2611), .ZN(n2618) );
  INV_X1 U2736 ( .A(n2867), .ZN(n2931) );
  NAND2_X1 U2737 ( .A1(n3956), .A2(n3909), .ZN(n2057) );
  AND2_X1 U2738 ( .A1(n2361), .A2(n2370), .ZN(n4380) );
  INV_X1 U2739 ( .A(n4380), .ZN(n2193) );
  NAND2_X1 U2740 ( .A1(n2618), .A2(n4373), .ZN(n2799) );
  INV_X1 U2741 ( .A(n3463), .ZN(n2167) );
  AND2_X1 U2742 ( .A1(n3945), .A2(n3750), .ZN(n2058) );
  AND2_X1 U2743 ( .A1(n2310), .A2(n2305), .ZN(n2344) );
  AND2_X1 U2744 ( .A1(n3055), .A2(n3904), .ZN(n2059) );
  AND2_X1 U2745 ( .A1(n2143), .A2(n3904), .ZN(n2060) );
  NAND2_X1 U2746 ( .A1(n2268), .A2(n2540), .ZN(n4156) );
  AND2_X1 U2747 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2061)
         );
  NAND2_X1 U2748 ( .A1(n3740), .A2(n3952), .ZN(n2062) );
  OR2_X1 U2749 ( .A1(n2712), .A2(n4540), .ZN(n2063) );
  AND2_X1 U2750 ( .A1(n2194), .A2(n4380), .ZN(n2064) );
  OR2_X1 U2751 ( .A1(n2267), .A2(n2263), .ZN(n2065) );
  AND2_X1 U2752 ( .A1(n2349), .A2(n2289), .ZN(n2315) );
  INV_X1 U2753 ( .A(n2250), .ZN(n2249) );
  OR2_X1 U2754 ( .A1(n3707), .A2(n2074), .ZN(n2250) );
  NAND2_X1 U2755 ( .A1(n2237), .A2(n2559), .ZN(n4115) );
  AND2_X1 U2756 ( .A1(n2324), .A2(n2723), .ZN(n2066) );
  AND2_X1 U2757 ( .A1(n2851), .A2(n3667), .ZN(n2067) );
  INV_X1 U2758 ( .A(n2192), .ZN(n2189) );
  NAND2_X1 U2759 ( .A1(n2818), .A2(n4377), .ZN(n2192) );
  INV_X1 U2760 ( .A(n3903), .ZN(n2140) );
  AND2_X1 U2761 ( .A1(n3369), .A2(n3370), .ZN(n2164) );
  NAND2_X1 U2762 ( .A1(n2049), .A2(n2425), .ZN(n2068) );
  XNOR2_X1 U2763 ( .A(n2670), .B(IR_REG_24__SCAN_IN), .ZN(n2678) );
  INV_X1 U2764 ( .A(n3399), .ZN(n2206) );
  INV_X1 U2765 ( .A(n3859), .ZN(n2234) );
  NOR2_X1 U2766 ( .A1(n3685), .A2(n3683), .ZN(n2069) );
  OR2_X1 U2767 ( .A1(n4262), .A2(n4085), .ZN(n2070) );
  INV_X1 U2768 ( .A(n2925), .ZN(n2171) );
  AND2_X1 U2769 ( .A1(n3536), .A2(n3535), .ZN(n2071) );
  AND2_X1 U2770 ( .A1(n4131), .A2(n2652), .ZN(n4157) );
  NAND2_X1 U2771 ( .A1(n2160), .A2(n3609), .ZN(n3808) );
  INV_X1 U2772 ( .A(n3318), .ZN(n2226) );
  OR2_X1 U2773 ( .A1(n3943), .A2(n3708), .ZN(n2072) );
  OR2_X1 U2774 ( .A1(n3948), .A2(n3719), .ZN(n2073) );
  AND2_X1 U2775 ( .A1(n3678), .A2(n3677), .ZN(n2074) );
  NAND2_X1 U2776 ( .A1(n3435), .A2(n2077), .ZN(n2090) );
  OR2_X1 U2777 ( .A1(n3769), .A2(n3768), .ZN(n2075) );
  AND2_X1 U2778 ( .A1(n4378), .A2(REG1_REG_5__SCAN_IN), .ZN(n2076) );
  INV_X1 U2779 ( .A(n2168), .ZN(n2166) );
  NAND2_X1 U2780 ( .A1(n2054), .A2(n3237), .ZN(n2168) );
  AND2_X1 U2781 ( .A1(n2055), .A2(n3469), .ZN(n2077) );
  AND2_X1 U2782 ( .A1(n4195), .A2(n4225), .ZN(n2078) );
  NAND2_X1 U2783 ( .A1(n4376), .A2(REG2_REG_7__SCAN_IN), .ZN(n2190) );
  OR2_X1 U2784 ( .A1(n2234), .A2(n3858), .ZN(n2079) );
  AND4_X1 U2785 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n3574)
         );
  INV_X1 U2786 ( .A(n3574), .ZN(n3950) );
  INV_X1 U2787 ( .A(n2131), .ZN(n2130) );
  NOR2_X1 U2788 ( .A1(n3915), .A2(n2132), .ZN(n2131) );
  INV_X1 U2789 ( .A(n3885), .ZN(n3567) );
  NAND2_X1 U2790 ( .A1(n2079), .A2(n2230), .ZN(n2080) );
  INV_X1 U2791 ( .A(IR_REG_19__SCAN_IN), .ZN(n2608) );
  AND2_X1 U2792 ( .A1(n2128), .A2(n2126), .ZN(n2081) );
  AND2_X1 U2793 ( .A1(n4147), .A2(n2540), .ZN(n2082) );
  NAND2_X1 U2794 ( .A1(n2249), .A2(n3689), .ZN(n2083) );
  INV_X1 U2795 ( .A(IR_REG_31__SCAN_IN), .ZN(n2723) );
  OR2_X1 U2796 ( .A1(n2278), .A2(n2274), .ZN(n2084) );
  OR2_X1 U2797 ( .A1(n2697), .A2(n2872), .ZN(n4540) );
  INV_X2 U2798 ( .A(n4540), .ZN(n4543) );
  INV_X1 U2799 ( .A(n3897), .ZN(n3617) );
  AOI21_X1 U2800 ( .B1(n3698), .B2(n3697), .A(n2071), .ZN(n3757) );
  NAND2_X1 U2801 ( .A1(n2453), .A2(n2452), .ZN(n3220) );
  NAND2_X1 U2802 ( .A1(n2264), .A2(n2262), .ZN(n3103) );
  OR2_X1 U2803 ( .A1(n4536), .A2(n2717), .ZN(n2085) );
  AND2_X1 U2804 ( .A1(n4540), .A2(n2713), .ZN(n2086) );
  INV_X1 U2805 ( .A(n3925), .ZN(n3929) );
  INV_X1 U2806 ( .A(n4037), .ZN(n2180) );
  AND2_X1 U2807 ( .A1(n2768), .A2(n3392), .ZN(n4429) );
  INV_X1 U2808 ( .A(n3690), .ZN(n3683) );
  OR2_X1 U2809 ( .A1(n3578), .A2(n3577), .ZN(n2087) );
  AND2_X1 U2810 ( .A1(n2045), .A2(DATAI_27_), .ZN(n3708) );
  AND2_X1 U2811 ( .A1(n2092), .A2(n4245), .ZN(n2088) );
  INV_X1 U2812 ( .A(n4258), .ZN(n4100) );
  AND2_X1 U2813 ( .A1(n2046), .A2(DATAI_25_), .ZN(n4258) );
  NOR2_X1 U2814 ( .A1(n4505), .A2(n4046), .ZN(n2103) );
  AND2_X1 U2815 ( .A1(n2923), .A2(n2339), .ZN(n2880) );
  INV_X1 U2816 ( .A(n2283), .ZN(n2210) );
  OR2_X1 U2817 ( .A1(n2101), .A2(n2100), .ZN(n2089) );
  INV_X1 U2818 ( .A(n2090), .ZN(n3485) );
  INV_X1 U2819 ( .A(n2093), .ZN(n3502) );
  MUX2_X1 U2820 ( .A(n2095), .B(n2094), .S(n2351), .Z(n2867) );
  NAND2_X1 U2821 ( .A1(n4026), .A2(n4375), .ZN(n2096) );
  XNOR2_X1 U2822 ( .A(n4026), .B(n4375), .ZN(n4028) );
  NAND2_X1 U2823 ( .A1(n4475), .A2(n2099), .ZN(n2097) );
  OAI211_X1 U2824 ( .C1(n4475), .C2(n2089), .A(n2098), .B(n2097), .ZN(n4053)
         );
  NOR2_X1 U2825 ( .A1(n4475), .A2(n4045), .ZN(n4485) );
  INV_X1 U2826 ( .A(n4045), .ZN(n2102) );
  NOR2_X1 U2827 ( .A1(n2894), .A2(n2893), .ZN(n2895) );
  NOR2_X1 U2828 ( .A1(n2855), .A2(n2856), .ZN(n2894) );
  NOR2_X1 U2829 ( .A1(n2850), .A2(n2067), .ZN(n2856) );
  INV_X1 U2830 ( .A(n3737), .ZN(n2110) );
  OAI21_X1 U2831 ( .B1(n2110), .B2(n2112), .A(n2111), .ZN(n3718) );
  NAND2_X1 U2832 ( .A1(n3790), .A2(n2081), .ZN(n2122) );
  OAI211_X1 U2833 ( .C1(n3790), .C2(n2127), .A(n2123), .B(n2122), .ZN(n3714)
         );
  NAND2_X1 U2834 ( .A1(n3790), .A2(n3788), .ZN(n2133) );
  NAND2_X1 U2835 ( .A1(n2135), .A2(n3524), .ZN(n2134) );
  INV_X1 U2836 ( .A(n3055), .ZN(n2135) );
  INV_X1 U2837 ( .A(n2504), .ZN(n2144) );
  OAI21_X1 U2838 ( .B1(n2144), .B2(n2723), .A(n2145), .ZN(n2610) );
  NAND2_X1 U2839 ( .A1(n2148), .A2(n2151), .ZN(n3747) );
  NAND3_X1 U2840 ( .A1(n3604), .A2(n2149), .A3(n3797), .ZN(n2148) );
  NAND3_X1 U2841 ( .A1(n3604), .A2(n3797), .A3(n3800), .ZN(n2160) );
  NAND2_X1 U2842 ( .A1(n3463), .A2(n2164), .ZN(n2161) );
  NAND2_X1 U2843 ( .A1(n2161), .A2(n2162), .ZN(n2654) );
  NAND3_X1 U2844 ( .A1(n2172), .A2(n2718), .A3(n2085), .ZN(U3515) );
  NAND2_X1 U2845 ( .A1(n2178), .A2(n2177), .ZN(n3506) );
  NAND2_X1 U2846 ( .A1(n2638), .A2(n3325), .ZN(n3179) );
  NAND2_X1 U2847 ( .A1(n2926), .A2(n2632), .ZN(n2885) );
  NAND2_X1 U2848 ( .A1(n3506), .A2(n3251), .ZN(n2703) );
  AOI21_X1 U2849 ( .B1(n2703), .B2(n3257), .A(n2702), .ZN(n2704) );
  NAND2_X1 U2850 ( .A1(n2644), .A2(n3362), .ZN(n3397) );
  OAI21_X1 U2851 ( .B1(n4061), .B2(n2063), .A(n2216), .ZN(n2716) );
  NOR2_X1 U2852 ( .A1(n2217), .A2(n2086), .ZN(n2216) );
  NAND2_X1 U2853 ( .A1(n2184), .A2(n2183), .ZN(n4005) );
  NAND3_X1 U2854 ( .A1(n2186), .A2(n2190), .A3(n2192), .ZN(n2184) );
  OAI21_X1 U2855 ( .B1(n2819), .B2(n2189), .A(n2187), .ZN(n2191) );
  INV_X1 U2856 ( .A(n2819), .ZN(n2186) );
  INV_X1 U2857 ( .A(n2191), .ZN(n2915) );
  NAND2_X1 U2858 ( .A1(n2631), .A2(n2924), .ZN(n2923) );
  NOR2_X1 U2859 ( .A1(n2619), .A2(n2066), .ZN(n2706) );
  NAND2_X1 U2860 ( .A1(n2453), .A2(n2208), .ZN(n2207) );
  NAND3_X1 U2861 ( .A1(n2386), .A2(n2057), .A3(n2214), .ZN(n2213) );
  NOR2_X2 U2862 ( .A1(n3096), .A2(n3348), .ZN(n3095) );
  NAND2_X1 U2863 ( .A1(n2701), .A2(n2219), .ZN(n2218) );
  NAND2_X1 U2864 ( .A1(n2224), .A2(n2222), .ZN(n2221) );
  NAND2_X1 U2865 ( .A1(n3571), .A2(n3570), .ZN(n3780) );
  NAND2_X1 U2866 ( .A1(n3917), .A2(n2239), .ZN(n2238) );
  OAI211_X1 U2867 ( .C1(n3917), .C2(n2240), .A(n2238), .B(n3696), .ZN(U3217)
         );
  OR2_X1 U2868 ( .A1(n3476), .A2(n2254), .ZN(n2251) );
  NAND2_X1 U2869 ( .A1(n2251), .A2(n2252), .ZN(n4186) );
  INV_X1 U2870 ( .A(n3122), .ZN(n2265) );
  OAI21_X1 U2871 ( .B1(n3122), .B2(n2068), .A(n2257), .ZN(n2256) );
  NAND2_X1 U2872 ( .A1(n2268), .A2(n2082), .ZN(n4154) );
  NAND2_X1 U2873 ( .A1(n2680), .A2(n2679), .ZN(n2669) );
  NAND2_X1 U2874 ( .A1(n2668), .A2(n2667), .ZN(n2269) );
  NAND2_X1 U2875 ( .A1(n3558), .A2(n2270), .ZN(n3737) );
  NAND2_X1 U2876 ( .A1(n2273), .A2(n2272), .ZN(n2595) );
  OAI21_X1 U2877 ( .B1(n3771), .B2(n2084), .A(n2275), .ZN(n3663) );
  INV_X1 U2878 ( .A(IR_REG_6__SCAN_IN), .ZN(n2317) );
  CLKBUF_X1 U2879 ( .A(n2338), .Z(n2998) );
  OR2_X1 U2880 ( .A1(n2343), .A2(n2342), .ZN(n2346) );
  OR2_X1 U2881 ( .A1(n2343), .A2(n2333), .ZN(n2336) );
  NAND2_X1 U2882 ( .A1(n2595), .A2(n2594), .ZN(n2701) );
  NAND2_X1 U2883 ( .A1(n3829), .A2(n3828), .ZN(n3827) );
  NOR2_X2 U2884 ( .A1(n3095), .A2(n2052), .ZN(n3122) );
  NAND2_X1 U2885 ( .A1(n2338), .A2(n2932), .ZN(n2632) );
  BUF_X1 U2886 ( .A(n2323), .Z(n2664) );
  AND2_X1 U2887 ( .A1(n3863), .A2(n3949), .ZN(n2283) );
  INV_X1 U2888 ( .A(n3568), .ZN(n3951) );
  AND4_X1 U2889 ( .A1(n2433), .A2(n2432), .A3(n2431), .A4(n2430), .ZN(n3568)
         );
  NAND2_X1 U2890 ( .A1(n4154), .A2(n2546), .ZN(n4127) );
  OR2_X1 U2891 ( .A1(n3513), .A2(n4362), .ZN(n2284) );
  OR2_X1 U2892 ( .A1(n3513), .A2(n4305), .ZN(n2285) );
  NAND2_X1 U2893 ( .A1(n4536), .A2(n4317), .ZN(n4362) );
  NAND2_X1 U2894 ( .A1(n3600), .A2(n3599), .ZN(n3797) );
  AND2_X1 U2895 ( .A1(n3660), .A2(n3661), .ZN(n2286) );
  INV_X1 U2896 ( .A(IR_REG_25__SCAN_IN), .ZN(n2296) );
  NAND2_X1 U2897 ( .A1(n4193), .A2(n4286), .ZN(n2539) );
  INV_X1 U2898 ( .A(n3598), .ZN(n3599) );
  OR2_X1 U2899 ( .A1(n2343), .A2(n2326), .ZN(n2330) );
  INV_X1 U2900 ( .A(IR_REG_17__SCAN_IN), .ZN(n2516) );
  NOR2_X1 U2901 ( .A1(n2495), .A2(n2494), .ZN(n2508) );
  NAND2_X1 U2902 ( .A1(n2407), .A2(REG3_REG_9__SCAN_IN), .ZN(n2415) );
  INV_X1 U2903 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2457) );
  AND2_X1 U2904 ( .A1(n2508), .A2(REG3_REG_18__SCAN_IN), .ZN(n2527) );
  NOR2_X1 U2905 ( .A1(n2465), .A2(n4708), .ZN(n2472) );
  NAND2_X1 U2906 ( .A1(n2569), .A2(REG3_REG_25__SCAN_IN), .ZN(n2579) );
  OR2_X1 U2907 ( .A1(n4176), .A2(n4160), .ZN(n4131) );
  NAND2_X1 U2908 ( .A1(n2527), .A2(n2526), .ZN(n2534) );
  NAND2_X1 U2909 ( .A1(n3567), .A2(n3568), .ZN(n2440) );
  AND2_X1 U2910 ( .A1(n2405), .A2(REG3_REG_8__SCAN_IN), .ZN(n2407) );
  INV_X1 U2911 ( .A(n2882), .ZN(n3295) );
  INV_X1 U2912 ( .A(n4160), .ZN(n3648) );
  INV_X1 U2913 ( .A(n3953), .ZN(n3549) );
  INV_X1 U2914 ( .A(n4291), .ZN(n4311) );
  INV_X1 U2915 ( .A(n2550), .ZN(n2548) );
  OR2_X1 U2916 ( .A1(n2485), .A2(n4653), .ZN(n2495) );
  NAND2_X1 U2917 ( .A1(n2374), .A2(REG3_REG_5__SCAN_IN), .ZN(n2387) );
  OR2_X1 U2918 ( .A1(n2458), .A2(n2457), .ZN(n2465) );
  NAND2_X1 U2919 ( .A1(n2426), .A2(REG3_REG_11__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U2920 ( .A1(n2472), .A2(REG3_REG_15__SCAN_IN), .ZN(n2485) );
  OR2_X1 U2921 ( .A1(n2579), .A2(n3918), .ZN(n2599) );
  OR2_X1 U2922 ( .A1(n2534), .A2(n3773), .ZN(n2550) );
  INV_X1 U2923 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4708) );
  AOI21_X1 U2924 ( .B1(n3433), .B2(n2484), .A(n2483), .ZN(n3418) );
  AND2_X1 U2925 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2374) );
  AND2_X1 U2926 ( .A1(n2629), .A2(n3289), .ZN(n2865) );
  INV_X1 U2927 ( .A(n4197), .ZN(n4222) );
  INV_X1 U2928 ( .A(n4287), .ZN(n4314) );
  OR2_X1 U2929 ( .A1(n2869), .A2(n4372), .ZN(n3130) );
  INV_X1 U2930 ( .A(IR_REG_23__SCAN_IN), .ZN(n2679) );
  AND2_X1 U2931 ( .A1(n2570), .A2(n2561), .ZN(n4120) );
  INV_X1 U2932 ( .A(n3581), .ZN(n3863) );
  AND2_X1 U2933 ( .A1(n2525), .A2(n2511), .ZN(n3898) );
  AND3_X1 U2934 ( .A1(n2874), .A2(n2785), .A3(n2871), .ZN(n2861) );
  OR2_X1 U2935 ( .A1(n2599), .A2(n2596), .ZN(n4066) );
  AND4_X1 U2936 ( .A1(n2463), .A2(n2462), .A3(n2461), .A4(n2460), .ZN(n3582)
         );
  AND2_X1 U2937 ( .A1(n2747), .A2(n2745), .ZN(n2768) );
  INV_X1 U2938 ( .A(n4317), .ZN(n2985) );
  INV_X1 U2939 ( .A(n3750), .ZN(n4225) );
  INV_X1 U2940 ( .A(n3932), .ZN(n3593) );
  AND2_X1 U2941 ( .A1(n2800), .A2(n4504), .ZN(n2811) );
  AND2_X1 U2942 ( .A1(n2439), .A2(n2447), .ZN(n4023) );
  NAND2_X1 U2943 ( .A1(n2861), .A2(n2807), .ZN(n3925) );
  INV_X1 U2944 ( .A(n3685), .ZN(n4247) );
  INV_X1 U2945 ( .A(n4151), .ZN(n4269) );
  INV_X1 U2946 ( .A(n3585), .ZN(n3948) );
  INV_X1 U2947 ( .A(n3533), .ZN(n3955) );
  INV_X1 U2948 ( .A(n4513), .ZN(n4406) );
  OR2_X1 U2949 ( .A1(n3487), .A2(n2985), .ZN(n4231) );
  NAND2_X1 U2950 ( .A1(n4543), .A2(n4317), .ZN(n4305) );
  OR2_X1 U2951 ( .A1(n4067), .A2(n4362), .ZN(n2718) );
  OR2_X1 U2952 ( .A1(n2697), .A2(n2785), .ZN(n4534) );
  INV_X1 U2953 ( .A(n4022), .ZN(n4509) );
  INV_X1 U2954 ( .A(n2770), .ZN(n4378) );
  NOR2_X2 U2955 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2349)
         );
  INV_X1 U2956 ( .A(IR_REG_11__SCAN_IN), .ZN(n2437) );
  NAND3_X1 U2957 ( .A1(n2291), .A2(n2315), .A3(n2290), .ZN(n2454) );
  INV_X1 U2958 ( .A(n2454), .ZN(n2295) );
  NAND2_X1 U2959 ( .A1(n2295), .A2(n2051), .ZN(n2613) );
  NAND2_X1 U2960 ( .A1(n2660), .A2(n2297), .ZN(n2298) );
  NAND2_X1 U2961 ( .A1(n2323), .A2(n2301), .ZN(n2304) );
  INV_X1 U2962 ( .A(n2305), .ZN(n2309) );
  NAND2_X1 U2963 ( .A1(n2323), .A2(n2303), .ZN(n2622) );
  NAND2_X1 U2964 ( .A1(n3230), .A2(REG0_REG_9__SCAN_IN), .ZN(n2314) );
  INV_X1 U2965 ( .A(n2407), .ZN(n2307) );
  INV_X1 U2966 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2306) );
  NAND2_X1 U2967 ( .A1(n2307), .A2(n2306), .ZN(n2308) );
  NAND2_X1 U2968 ( .A1(n2415), .A2(n2308), .ZN(n3105) );
  INV_X1 U2969 ( .A(n3105), .ZN(n3841) );
  NAND2_X1 U2970 ( .A1(n2601), .A2(n3841), .ZN(n2313) );
  NAND2_X1 U2971 ( .A1(n2536), .A2(REG1_REG_9__SCAN_IN), .ZN(n2312) );
  NAND2_X1 U2972 ( .A1(n3229), .A2(REG2_REG_9__SCAN_IN), .ZN(n2311) );
  NAND4_X1 U2973 ( .A1(n2314), .A2(n2313), .A3(n2312), .A4(n2311), .ZN(n3953)
         );
  NOR2_X1 U2974 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2316)
         );
  NAND2_X1 U2975 ( .A1(n2315), .A2(n2316), .ZN(n2382) );
  NAND3_X1 U2976 ( .A1(n2317), .A2(n2402), .A3(n4613), .ZN(n2318) );
  NOR2_X1 U2977 ( .A1(n2401), .A2(n2318), .ZN(n2422) );
  OR2_X1 U2978 ( .A1(n2422), .A2(n2723), .ZN(n2319) );
  XNOR2_X1 U2979 ( .A(n2319), .B(IR_REG_9__SCAN_IN), .ZN(n4025) );
  NAND2_X1 U2980 ( .A1(n2664), .A2(n2320), .ZN(n2673) );
  MUX2_X2 U2981 ( .A(n2705), .B(n2706), .S(n2325), .Z(n2351) );
  MUX2_X1 U2982 ( .A(n4025), .B(DATAI_9_), .S(n2046), .Z(n3840) );
  INV_X1 U2983 ( .A(n3840), .ZN(n3548) );
  INV_X1 U2984 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2326) );
  NAND2_X1 U2985 ( .A1(n2341), .A2(REG0_REG_1__SCAN_IN), .ZN(n2329) );
  NAND2_X1 U2986 ( .A1(n2340), .A2(REG3_REG_1__SCAN_IN), .ZN(n2328) );
  NAND2_X1 U2987 ( .A1(n2344), .A2(REG2_REG_1__SCAN_IN), .ZN(n2327) );
  NAND4_X1 U2988 ( .A1(n2330), .A2(n2329), .A3(n2328), .A4(n2327), .ZN(n2332)
         );
  NAND2_X1 U2989 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2331)
         );
  MUX2_X1 U2990 ( .A(n4382), .B(DATAI_1_), .S(n2351), .Z(n2932) );
  NAND2_X1 U2991 ( .A1(n2332), .A2(n2987), .ZN(n3332) );
  INV_X1 U2992 ( .A(n2332), .ZN(n2338) );
  NAND2_X1 U2993 ( .A1(n2340), .A2(REG3_REG_0__SCAN_IN), .ZN(n2337) );
  INV_X1 U2994 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2333) );
  NAND2_X1 U2995 ( .A1(n2344), .A2(REG2_REG_0__SCAN_IN), .ZN(n2335) );
  NAND2_X1 U2996 ( .A1(n2341), .A2(REG0_REG_0__SCAN_IN), .ZN(n2334) );
  AND2_X1 U2997 ( .A1(n3962), .A2(n2931), .ZN(n2924) );
  INV_X1 U2998 ( .A(n2338), .ZN(n2808) );
  NAND2_X1 U2999 ( .A1(n2808), .A2(n2932), .ZN(n2339) );
  NAND2_X1 U3000 ( .A1(n2340), .A2(REG3_REG_2__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U3001 ( .A1(n2341), .A2(REG0_REG_2__SCAN_IN), .ZN(n2347) );
  INV_X1 U3002 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2342) );
  NAND2_X1 U3003 ( .A1(n2344), .A2(REG2_REG_2__SCAN_IN), .ZN(n2345) );
  AND4_X2 U3004 ( .A1(n2348), .A2(n2347), .A3(n2346), .A4(n2345), .ZN(n2352)
         );
  INV_X1 U3005 ( .A(n2352), .ZN(n3960) );
  MUX2_X1 U3006 ( .A(n4381), .B(DATAI_2_), .S(n2351), .Z(n2899) );
  INV_X1 U3007 ( .A(n2899), .ZN(n2997) );
  NAND2_X1 U3008 ( .A1(n3960), .A2(n2997), .ZN(n3338) );
  NAND2_X1 U3009 ( .A1(n2352), .A2(n2899), .ZN(n3335) );
  NAND2_X1 U3010 ( .A1(n2880), .A2(n2882), .ZN(n2881) );
  NAND2_X1 U3011 ( .A1(n2352), .A2(n2997), .ZN(n2353) );
  NAND2_X1 U3012 ( .A1(n2881), .A2(n2353), .ZN(n2903) );
  NAND2_X1 U3013 ( .A1(n3230), .A2(REG0_REG_3__SCAN_IN), .ZN(n2358) );
  INV_X1 U3014 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2354) );
  NAND2_X1 U3015 ( .A1(n2601), .A2(n2354), .ZN(n2357) );
  NAND2_X1 U3016 ( .A1(n2536), .A2(REG1_REG_3__SCAN_IN), .ZN(n2356) );
  NAND2_X1 U3017 ( .A1(n3229), .A2(REG2_REG_3__SCAN_IN), .ZN(n2355) );
  NOR2_X1 U3018 ( .A1(n2315), .A2(n2723), .ZN(n2359) );
  NAND2_X1 U3019 ( .A1(n2359), .A2(IR_REG_3__SCAN_IN), .ZN(n2361) );
  INV_X1 U3020 ( .A(n2359), .ZN(n2360) );
  NAND2_X1 U3021 ( .A1(n2360), .A2(n4696), .ZN(n2370) );
  MUX2_X1 U3022 ( .A(n4380), .B(DATAI_3_), .S(n2045), .Z(n2980) );
  NAND2_X1 U3023 ( .A1(n3959), .A2(n2980), .ZN(n2362) );
  NAND2_X1 U3024 ( .A1(n2903), .A2(n2362), .ZN(n2364) );
  NAND2_X1 U3025 ( .A1(n2999), .A2(n3077), .ZN(n2363) );
  NAND2_X1 U3026 ( .A1(n2364), .A2(n2363), .ZN(n2940) );
  INV_X1 U3027 ( .A(n2940), .ZN(n2372) );
  NAND2_X1 U3028 ( .A1(n3229), .A2(REG2_REG_4__SCAN_IN), .ZN(n2369) );
  NAND2_X1 U3029 ( .A1(n3230), .A2(REG0_REG_4__SCAN_IN), .ZN(n2368) );
  NOR2_X1 U3030 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2365) );
  NOR2_X1 U3031 ( .A1(n2374), .A2(n2365), .ZN(n3832) );
  NAND2_X1 U3032 ( .A1(n2601), .A2(n3832), .ZN(n2367) );
  NAND2_X1 U3033 ( .A1(n2536), .A2(REG1_REG_4__SCAN_IN), .ZN(n2366) );
  AND4_X2 U3034 ( .A1(n2369), .A2(n2368), .A3(n2367), .A4(n2366), .ZN(n3065)
         );
  NAND2_X1 U3035 ( .A1(n2370), .A2(IR_REG_31__SCAN_IN), .ZN(n2371) );
  XNOR2_X1 U3036 ( .A(n2371), .B(IR_REG_4__SCAN_IN), .ZN(n4379) );
  MUX2_X1 U3037 ( .A(n4379), .B(DATAI_4_), .S(n2046), .Z(n3831) );
  INV_X1 U3038 ( .A(n3831), .ZN(n3046) );
  NAND2_X1 U3039 ( .A1(n3958), .A2(n3046), .ZN(n3345) );
  NAND2_X1 U3040 ( .A1(n3065), .A2(n3831), .ZN(n3341) );
  NAND2_X1 U3041 ( .A1(n2372), .A2(n2938), .ZN(n2942) );
  NAND2_X1 U3042 ( .A1(n3958), .A2(n3831), .ZN(n2373) );
  NAND2_X1 U3043 ( .A1(n3230), .A2(REG0_REG_5__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U3044 ( .A1(n2536), .A2(REG1_REG_5__SCAN_IN), .ZN(n2380) );
  INV_X1 U3045 ( .A(n2374), .ZN(n2376) );
  INV_X1 U3046 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2375) );
  NAND2_X1 U3047 ( .A1(n2376), .A2(n2375), .ZN(n2377) );
  AND2_X1 U3048 ( .A1(n2377), .A2(n2387), .ZN(n3037) );
  NAND2_X1 U3049 ( .A1(n2601), .A2(n3037), .ZN(n2379) );
  NAND2_X1 U3050 ( .A1(n3229), .A2(REG2_REG_5__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U3051 ( .A1(n2382), .A2(IR_REG_31__SCAN_IN), .ZN(n2383) );
  MUX2_X1 U3052 ( .A(IR_REG_31__SCAN_IN), .B(n2383), .S(IR_REG_5__SCAN_IN), 
        .Z(n2384) );
  NAND2_X1 U3053 ( .A1(n2384), .A2(n2401), .ZN(n2770) );
  INV_X1 U3054 ( .A(DATAI_5_), .ZN(n4705) );
  MUX2_X1 U3055 ( .A(n2770), .B(n4705), .S(n2046), .Z(n3057) );
  NAND2_X1 U3056 ( .A1(n3053), .A2(n3057), .ZN(n2385) );
  INV_X1 U3057 ( .A(n3053), .ZN(n3957) );
  NAND2_X1 U3058 ( .A1(n3957), .A2(n3068), .ZN(n2386) );
  NAND2_X1 U3059 ( .A1(n3229), .A2(REG2_REG_6__SCAN_IN), .ZN(n2392) );
  NAND2_X1 U3060 ( .A1(n3230), .A2(REG0_REG_6__SCAN_IN), .ZN(n2391) );
  AND2_X1 U3061 ( .A1(n2387), .A2(n2775), .ZN(n2388) );
  NOR2_X1 U3062 ( .A1(n2395), .A2(n2388), .ZN(n3910) );
  NAND2_X1 U3063 ( .A1(n2601), .A2(n3910), .ZN(n2390) );
  NAND2_X1 U3064 ( .A1(n2536), .A2(REG1_REG_6__SCAN_IN), .ZN(n2389) );
  NAND4_X1 U3065 ( .A1(n2392), .A2(n2391), .A3(n2390), .A4(n2389), .ZN(n3956)
         );
  NAND2_X1 U3066 ( .A1(n2401), .A2(IR_REG_31__SCAN_IN), .ZN(n2393) );
  XNOR2_X1 U3067 ( .A(n2393), .B(IR_REG_6__SCAN_IN), .ZN(n4377) );
  MUX2_X1 U3068 ( .A(n4377), .B(DATAI_6_), .S(n2046), .Z(n3909) );
  NAND2_X1 U3069 ( .A1(n3527), .A2(n3526), .ZN(n2394) );
  NAND2_X1 U3070 ( .A1(n3229), .A2(REG2_REG_7__SCAN_IN), .ZN(n2400) );
  NAND2_X1 U3071 ( .A1(n3230), .A2(REG0_REG_7__SCAN_IN), .ZN(n2399) );
  NOR2_X1 U3072 ( .A1(n2395), .A2(REG3_REG_7__SCAN_IN), .ZN(n2396) );
  OR2_X1 U3073 ( .A1(n2405), .A2(n2396), .ZN(n3090) );
  INV_X1 U3074 ( .A(n3090), .ZN(n3702) );
  NAND2_X1 U3075 ( .A1(n2601), .A2(n3702), .ZN(n2398) );
  NAND2_X1 U3076 ( .A1(n2536), .A2(REG1_REG_7__SCAN_IN), .ZN(n2397) );
  OAI21_X1 U3077 ( .B1(n2401), .B2(IR_REG_6__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2403) );
  NAND2_X1 U3078 ( .A1(n2403), .A2(n2402), .ZN(n2412) );
  OR2_X1 U3079 ( .A1(n2403), .A2(n2402), .ZN(n2404) );
  MUX2_X1 U3080 ( .A(n4376), .B(DATAI_7_), .S(n2046), .Z(n3701) );
  NAND2_X1 U3081 ( .A1(n3533), .A2(n3701), .ZN(n2635) );
  NAND2_X1 U3082 ( .A1(n3955), .A2(n3532), .ZN(n3351) );
  NAND2_X1 U3083 ( .A1(n3230), .A2(REG0_REG_8__SCAN_IN), .ZN(n2411) );
  NAND2_X1 U3084 ( .A1(n2536), .A2(REG1_REG_8__SCAN_IN), .ZN(n2410) );
  NOR2_X1 U3085 ( .A1(n2405), .A2(REG3_REG_8__SCAN_IN), .ZN(n2406) );
  OR2_X1 U3086 ( .A1(n2407), .A2(n2406), .ZN(n4491) );
  INV_X1 U3087 ( .A(n4491), .ZN(n3763) );
  NAND2_X1 U3088 ( .A1(n2601), .A2(n3763), .ZN(n2409) );
  NAND2_X1 U3089 ( .A1(n3229), .A2(REG2_REG_8__SCAN_IN), .ZN(n2408) );
  NAND4_X1 U3090 ( .A1(n2411), .A2(n2410), .A3(n2409), .A4(n2408), .ZN(n3954)
         );
  NAND2_X1 U3091 ( .A1(n2412), .A2(IR_REG_31__SCAN_IN), .ZN(n2413) );
  XNOR2_X1 U3092 ( .A(n2413), .B(IR_REG_8__SCAN_IN), .ZN(n4375) );
  MUX2_X1 U3093 ( .A(n4375), .B(DATAI_8_), .S(n2046), .Z(n3762) );
  INV_X1 U3094 ( .A(n3954), .ZN(n3115) );
  INV_X1 U3095 ( .A(n3762), .ZN(n3124) );
  NAND2_X1 U3096 ( .A1(n3230), .A2(REG0_REG_10__SCAN_IN), .ZN(n2420) );
  NAND2_X1 U3097 ( .A1(n2536), .A2(REG1_REG_10__SCAN_IN), .ZN(n2419) );
  INV_X1 U3098 ( .A(n2426), .ZN(n2428) );
  INV_X1 U3099 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4664) );
  NAND2_X1 U3100 ( .A1(n2415), .A2(n4664), .ZN(n2416) );
  AND2_X1 U3101 ( .A1(n2428), .A2(n2416), .ZN(n3741) );
  NAND2_X1 U3102 ( .A1(n2601), .A2(n3741), .ZN(n2418) );
  NAND2_X1 U3103 ( .A1(n3229), .A2(REG2_REG_10__SCAN_IN), .ZN(n2417) );
  AND2_X1 U3104 ( .A1(n2422), .A2(n2421), .ZN(n2435) );
  OR2_X1 U3105 ( .A1(n2435), .A2(n2723), .ZN(n2423) );
  XNOR2_X1 U3106 ( .A(n2423), .B(IR_REG_10__SCAN_IN), .ZN(n4513) );
  INV_X1 U3107 ( .A(DATAI_10_), .ZN(n2424) );
  MUX2_X1 U3108 ( .A(n4406), .B(n2424), .S(n2046), .Z(n3559) );
  NAND2_X1 U3109 ( .A1(n3561), .A2(n3559), .ZN(n2425) );
  NAND2_X1 U3110 ( .A1(n3230), .A2(REG0_REG_11__SCAN_IN), .ZN(n2433) );
  NAND2_X1 U3111 ( .A1(n2536), .A2(REG1_REG_11__SCAN_IN), .ZN(n2432) );
  INV_X1 U3112 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2427) );
  NAND2_X1 U3113 ( .A1(n2428), .A2(n2427), .ZN(n2429) );
  AND2_X1 U3114 ( .A1(n2441), .A2(n2429), .ZN(n3886) );
  NAND2_X1 U3115 ( .A1(n2601), .A2(n3886), .ZN(n2431) );
  NAND2_X1 U3116 ( .A1(n3229), .A2(REG2_REG_11__SCAN_IN), .ZN(n2430) );
  AOI21_X1 U3117 ( .B1(n2435), .B2(n2434), .A(n2723), .ZN(n2436) );
  NAND2_X1 U3118 ( .A1(n2436), .A2(IR_REG_11__SCAN_IN), .ZN(n2439) );
  INV_X1 U3119 ( .A(n2436), .ZN(n2438) );
  NAND2_X1 U3120 ( .A1(n2438), .A2(n2437), .ZN(n2447) );
  MUX2_X1 U3121 ( .A(n4023), .B(DATAI_11_), .S(n2045), .Z(n3885) );
  NAND2_X1 U3122 ( .A1(n3568), .A2(n3885), .ZN(n3176) );
  NAND2_X1 U3123 ( .A1(n3951), .A2(n3567), .ZN(n3178) );
  NAND2_X1 U3124 ( .A1(n3176), .A2(n3178), .ZN(n3275) );
  NAND2_X1 U3125 ( .A1(n3164), .A2(n3275), .ZN(n3163) );
  NAND2_X1 U3126 ( .A1(n3163), .A2(n2440), .ZN(n3175) );
  NAND2_X1 U3127 ( .A1(n3229), .A2(REG2_REG_12__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U3128 ( .A1(n3230), .A2(REG0_REG_12__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U3129 ( .A1(n2441), .A2(n4662), .ZN(n2442) );
  AND2_X1 U3130 ( .A1(n2458), .A2(n2442), .ZN(n3783) );
  NAND2_X1 U3131 ( .A1(n2601), .A2(n3783), .ZN(n2444) );
  NAND2_X1 U3132 ( .A1(n2536), .A2(REG1_REG_12__SCAN_IN), .ZN(n2443) );
  NAND2_X1 U3133 ( .A1(n2447), .A2(IR_REG_31__SCAN_IN), .ZN(n2448) );
  XNOR2_X1 U3134 ( .A(n2448), .B(IR_REG_12__SCAN_IN), .ZN(n4033) );
  INV_X1 U3135 ( .A(DATAI_12_), .ZN(n2449) );
  MUX2_X1 U3136 ( .A(n4510), .B(n2449), .S(n2046), .Z(n3572) );
  NAND2_X1 U3137 ( .A1(n3175), .A2(n2451), .ZN(n2453) );
  NAND2_X1 U3138 ( .A1(n2454), .A2(IR_REG_31__SCAN_IN), .ZN(n2455) );
  XNOR2_X1 U3139 ( .A(n2455), .B(IR_REG_13__SCAN_IN), .ZN(n4022) );
  INV_X1 U3140 ( .A(DATAI_13_), .ZN(n2456) );
  MUX2_X1 U3141 ( .A(n4509), .B(n2456), .S(n2046), .Z(n3581) );
  NAND2_X1 U3142 ( .A1(n3229), .A2(REG2_REG_13__SCAN_IN), .ZN(n2463) );
  NAND2_X1 U3143 ( .A1(n3230), .A2(REG0_REG_13__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U3144 ( .A1(n2458), .A2(n2457), .ZN(n2459) );
  AND2_X1 U3145 ( .A1(n2465), .A2(n2459), .ZN(n3864) );
  NAND2_X1 U3146 ( .A1(n2601), .A2(n3864), .ZN(n2461) );
  NAND2_X1 U3147 ( .A1(n2536), .A2(REG1_REG_13__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U31480 ( .A1(n3230), .A2(REG0_REG_14__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U31490 ( .A1(n2536), .A2(REG1_REG_14__SCAN_IN), .ZN(n2469) );
  INV_X1 U3150 ( .A(n2472), .ZN(n2474) );
  NAND2_X1 U3151 ( .A1(n2465), .A2(n4708), .ZN(n2466) );
  NAND2_X1 U3152 ( .A1(n2601), .A2(n3723), .ZN(n2468) );
  NAND2_X1 U3153 ( .A1(n3229), .A2(REG2_REG_14__SCAN_IN), .ZN(n2467) );
  NAND2_X1 U3154 ( .A1(n2504), .A2(IR_REG_31__SCAN_IN), .ZN(n2471) );
  XNOR2_X1 U3155 ( .A(n2471), .B(IR_REG_14__SCAN_IN), .ZN(n4037) );
  MUX2_X1 U3156 ( .A(n4037), .B(DATAI_14_), .S(n2046), .Z(n3719) );
  NAND2_X1 U3157 ( .A1(n3585), .A2(n3719), .ZN(n3236) );
  NAND2_X1 U3158 ( .A1(n3948), .A2(n3583), .ZN(n3328) );
  NAND2_X1 U3159 ( .A1(n3236), .A2(n3328), .ZN(n3399) );
  NAND2_X1 U3160 ( .A1(n3398), .A2(n2073), .ZN(n3433) );
  NAND2_X1 U3161 ( .A1(n3229), .A2(REG2_REG_15__SCAN_IN), .ZN(n2479) );
  NAND2_X1 U3162 ( .A1(n3230), .A2(REG0_REG_15__SCAN_IN), .ZN(n2478) );
  INV_X1 U3163 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3164 ( .A1(n2474), .A2(n2473), .ZN(n2475) );
  AND2_X1 U3165 ( .A1(n2485), .A2(n2475), .ZN(n3935) );
  NAND2_X1 U3166 ( .A1(n2601), .A2(n3935), .ZN(n2477) );
  NAND2_X1 U3167 ( .A1(n2536), .A2(REG1_REG_15__SCAN_IN), .ZN(n2476) );
  NAND4_X1 U3168 ( .A1(n2479), .A2(n2478), .A3(n2477), .A4(n2476), .ZN(n3947)
         );
  OAI21_X1 U3169 ( .B1(n2504), .B2(IR_REG_14__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2481) );
  INV_X1 U3170 ( .A(IR_REG_15__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U3171 ( .A1(n2481), .A2(n2480), .ZN(n2491) );
  OR2_X1 U3172 ( .A1(n2481), .A2(n2480), .ZN(n2482) );
  MUX2_X1 U3173 ( .A(n4021), .B(DATAI_15_), .S(n2046), .Z(n3932) );
  NAND2_X1 U3174 ( .A1(n3947), .A2(n3932), .ZN(n2484) );
  NOR2_X1 U3175 ( .A1(n3947), .A2(n3932), .ZN(n2483) );
  NAND2_X1 U3176 ( .A1(n3229), .A2(REG2_REG_16__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U3177 ( .A1(n3230), .A2(REG0_REG_16__SCAN_IN), .ZN(n2489) );
  NAND2_X1 U3178 ( .A1(n2485), .A2(n4653), .ZN(n2486) );
  AND2_X1 U3179 ( .A1(n2495), .A2(n2486), .ZN(n3803) );
  NAND2_X1 U3180 ( .A1(n2601), .A2(n3803), .ZN(n2488) );
  NAND2_X1 U3181 ( .A1(n2536), .A2(REG1_REG_16__SCAN_IN), .ZN(n2487) );
  NAND2_X1 U3182 ( .A1(n2491), .A2(IR_REG_31__SCAN_IN), .ZN(n2492) );
  XNOR2_X1 U3183 ( .A(n2492), .B(IR_REG_16__SCAN_IN), .ZN(n4041) );
  MUX2_X1 U3184 ( .A(n4041), .B(DATAI_16_), .S(n2046), .Z(n4309) );
  NAND2_X1 U3185 ( .A1(n3602), .A2(n4309), .ZN(n3243) );
  INV_X1 U3186 ( .A(n4309), .ZN(n3601) );
  NAND2_X1 U3187 ( .A1(n3946), .A2(n3601), .ZN(n3329) );
  NAND2_X1 U3188 ( .A1(n3243), .A2(n3329), .ZN(n3420) );
  NAND2_X1 U3189 ( .A1(n3418), .A2(n3420), .ZN(n3419) );
  NAND2_X1 U3190 ( .A1(n3946), .A2(n4309), .ZN(n2493) );
  NAND2_X1 U3191 ( .A1(n3419), .A2(n2493), .ZN(n3465) );
  INV_X1 U3192 ( .A(n3465), .ZN(n2507) );
  NAND2_X1 U3193 ( .A1(n3230), .A2(REG0_REG_17__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U3194 ( .A1(n2536), .A2(REG1_REG_17__SCAN_IN), .ZN(n2499) );
  INV_X1 U3195 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2494) );
  INV_X1 U3196 ( .A(n2508), .ZN(n2510) );
  NAND2_X1 U3197 ( .A1(n2495), .A2(n2494), .ZN(n2496) );
  NAND2_X1 U3198 ( .A1(n2601), .A2(n3814), .ZN(n2498) );
  NAND2_X1 U3199 ( .A1(n3229), .A2(REG2_REG_17__SCAN_IN), .ZN(n2497) );
  NAND2_X1 U3200 ( .A1(n2502), .A2(n2501), .ZN(n2503) );
  OR2_X1 U3201 ( .A1(n2517), .A2(n2723), .ZN(n2505) );
  XNOR2_X1 U3202 ( .A(n2505), .B(IR_REG_17__SCAN_IN), .ZN(n4044) );
  MUX2_X1 U3203 ( .A(n4044), .B(DATAI_17_), .S(n2046), .Z(n3813) );
  INV_X1 U3204 ( .A(n4312), .ZN(n2646) );
  INV_X1 U3205 ( .A(n3813), .ZN(n3469) );
  OAI22_X2 U3206 ( .A1(n2507), .A2(n2506), .B1(n2646), .B2(n3469), .ZN(n3476)
         );
  INV_X1 U3207 ( .A(n2527), .ZN(n2525) );
  INV_X1 U3208 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2509) );
  NAND2_X1 U3209 ( .A1(n2510), .A2(n2509), .ZN(n2511) );
  NAND2_X1 U32100 ( .A1(n3898), .A2(n2601), .ZN(n2515) );
  NAND2_X1 U32110 ( .A1(n3230), .A2(REG0_REG_18__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U32120 ( .A1(n2536), .A2(REG1_REG_18__SCAN_IN), .ZN(n2513) );
  NAND2_X1 U32130 ( .A1(n3229), .A2(REG2_REG_18__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U32140 ( .A1(n2056), .A2(IR_REG_31__SCAN_IN), .ZN(n2518) );
  XNOR2_X1 U32150 ( .A(n2518), .B(IR_REG_18__SCAN_IN), .ZN(n4020) );
  MUX2_X1 U32160 ( .A(n4020), .B(DATAI_18_), .S(n2045), .Z(n3897) );
  NAND2_X1 U32170 ( .A1(n3619), .A2(n3897), .ZN(n4212) );
  NAND2_X1 U32180 ( .A1(n4220), .A2(n3617), .ZN(n4213) );
  NAND2_X1 U32190 ( .A1(n3619), .A2(n3617), .ZN(n2519) );
  XNOR2_X1 U32200 ( .A(n2525), .B(REG3_REG_19__SCAN_IN), .ZN(n4228) );
  NAND2_X1 U32210 ( .A1(n4228), .A2(n2601), .ZN(n2523) );
  NAND2_X1 U32220 ( .A1(n3229), .A2(REG2_REG_19__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U32230 ( .A1(n3230), .A2(REG0_REG_19__SCAN_IN), .ZN(n2521) );
  NAND2_X1 U32240 ( .A1(n2536), .A2(REG1_REG_19__SCAN_IN), .ZN(n2520) );
  NAND4_X1 U32250 ( .A1(n2523), .A2(n2522), .A3(n2521), .A4(n2520), .ZN(n3945)
         );
  MUX2_X1 U32260 ( .A(n4374), .B(DATAI_19_), .S(n2046), .Z(n3750) );
  INV_X1 U32270 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4300) );
  INV_X1 U32280 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2524) );
  INV_X1 U32290 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3852) );
  OAI21_X1 U32300 ( .B1(n2525), .B2(n2524), .A(n3852), .ZN(n2528) );
  AND2_X1 U32310 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2526) );
  NAND2_X1 U32320 ( .A1(n2528), .A2(n2534), .ZN(n4204) );
  NAND2_X1 U32330 ( .A1(n3229), .A2(REG2_REG_20__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U32340 ( .A1(n3230), .A2(REG0_REG_20__SCAN_IN), .ZN(n2529) );
  AND2_X1 U32350 ( .A1(n2530), .A2(n2529), .ZN(n2531) );
  NAND2_X1 U32360 ( .A1(n4186), .A2(n3304), .ZN(n2533) );
  INV_X1 U32370 ( .A(n4288), .ZN(n4218) );
  NAND2_X1 U32380 ( .A1(n4218), .A2(n4202), .ZN(n3305) );
  NAND2_X1 U32390 ( .A1(n2533), .A2(n3305), .ZN(n4169) );
  INV_X1 U32400 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3773) );
  NAND2_X1 U32410 ( .A1(n2534), .A2(n3773), .ZN(n2535) );
  NAND2_X1 U32420 ( .A1(n2550), .A2(n2535), .ZN(n3772) );
  AOI22_X1 U32430 ( .A1(n2536), .A2(REG1_REG_21__SCAN_IN), .B1(n3229), .B2(
        REG2_REG_21__SCAN_IN), .ZN(n2538) );
  NAND2_X1 U32440 ( .A1(n3230), .A2(REG0_REG_21__SCAN_IN), .ZN(n2537) );
  NAND2_X1 U32450 ( .A1(n2046), .A2(DATAI_21_), .ZN(n4181) );
  INV_X1 U32460 ( .A(n4181), .ZN(n4286) );
  INV_X1 U32470 ( .A(n4193), .ZN(n3873) );
  NAND2_X1 U32480 ( .A1(n3873), .A2(n4181), .ZN(n2540) );
  XNOR2_X1 U32490 ( .A(n2550), .B(REG3_REG_22__SCAN_IN), .ZN(n4162) );
  NAND2_X1 U32500 ( .A1(n4162), .A2(n2601), .ZN(n2545) );
  INV_X1 U32510 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4284) );
  NAND2_X1 U32520 ( .A1(n3230), .A2(REG0_REG_22__SCAN_IN), .ZN(n2542) );
  NAND2_X1 U32530 ( .A1(n3229), .A2(REG2_REG_22__SCAN_IN), .ZN(n2541) );
  OAI211_X1 U32540 ( .C1(n3234), .C2(n4284), .A(n2542), .B(n2541), .ZN(n2543)
         );
  INV_X1 U32550 ( .A(n2543), .ZN(n2544) );
  NAND2_X1 U32560 ( .A1(n2046), .A2(DATAI_22_), .ZN(n4160) );
  NAND2_X1 U32570 ( .A1(n4176), .A2(n4160), .ZN(n2652) );
  NAND2_X1 U32580 ( .A1(n4176), .A2(n3648), .ZN(n2546) );
  AND2_X1 U32590 ( .A1(REG3_REG_22__SCAN_IN), .A2(REG3_REG_23__SCAN_IN), .ZN(
        n2547) );
  INV_X1 U32600 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3872) );
  INV_X1 U32610 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2549) );
  OAI21_X1 U32620 ( .B1(n2550), .B2(n3872), .A(n2549), .ZN(n2551) );
  NAND2_X1 U32630 ( .A1(n2560), .A2(n2551), .ZN(n4141) );
  INV_X1 U32640 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4279) );
  NAND2_X1 U32650 ( .A1(n3229), .A2(REG2_REG_23__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32660 ( .A1(n3230), .A2(REG0_REG_23__SCAN_IN), .ZN(n2552) );
  OAI211_X1 U32670 ( .C1(n4279), .C2(n3234), .A(n2553), .B(n2552), .ZN(n2554)
         );
  INV_X1 U32680 ( .A(n2554), .ZN(n2555) );
  NAND2_X1 U32690 ( .A1(n2045), .A2(DATAI_23_), .ZN(n4138) );
  NAND2_X1 U32700 ( .A1(n4151), .A2(n4138), .ZN(n2557) );
  INV_X1 U32710 ( .A(n4138), .ZN(n2558) );
  NAND2_X1 U32720 ( .A1(n4269), .A2(n2558), .ZN(n2559) );
  INV_X1 U32730 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4648) );
  NAND2_X1 U32740 ( .A1(n2560), .A2(n4648), .ZN(n2561) );
  NAND2_X1 U32750 ( .A1(n4120), .A2(n2601), .ZN(n2566) );
  INV_X1 U32760 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4275) );
  NAND2_X1 U32770 ( .A1(n3229), .A2(REG2_REG_24__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U32780 ( .A1(n3230), .A2(REG0_REG_24__SCAN_IN), .ZN(n2562) );
  OAI211_X1 U32790 ( .C1(n4275), .C2(n3234), .A(n2563), .B(n2562), .ZN(n2564)
         );
  INV_X1 U32800 ( .A(n2564), .ZN(n2565) );
  NAND2_X1 U32810 ( .A1(n2046), .A2(DATAI_24_), .ZN(n4267) );
  NOR2_X1 U32820 ( .A1(n4134), .A2(n4267), .ZN(n2567) );
  NAND2_X1 U32830 ( .A1(n4134), .A2(n4267), .ZN(n2568) );
  INV_X1 U32840 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4595) );
  NAND2_X1 U32850 ( .A1(n2570), .A2(n4595), .ZN(n2571) );
  NAND2_X1 U32860 ( .A1(n2579), .A2(n2571), .ZN(n4104) );
  INV_X1 U32870 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4265) );
  NAND2_X1 U32880 ( .A1(n3229), .A2(REG2_REG_25__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U32890 ( .A1(n3230), .A2(REG0_REG_25__SCAN_IN), .ZN(n2572) );
  OAI211_X1 U32900 ( .C1(n4265), .C2(n3234), .A(n2573), .B(n2572), .ZN(n2574)
         );
  INV_X1 U32910 ( .A(n2574), .ZN(n2575) );
  NOR2_X1 U32920 ( .A1(n4119), .A2(n4258), .ZN(n2578) );
  NAND2_X1 U32930 ( .A1(n4119), .A2(n4258), .ZN(n2577) );
  INV_X1 U32940 ( .A(n4073), .ZN(n2586) );
  INV_X1 U32950 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3918) );
  NAND2_X1 U32960 ( .A1(n2579), .A2(n3918), .ZN(n2580) );
  NAND2_X1 U32970 ( .A1(n2599), .A2(n2580), .ZN(n4088) );
  INV_X1 U32980 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4256) );
  NAND2_X1 U32990 ( .A1(n3229), .A2(REG2_REG_26__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U33000 ( .A1(n3230), .A2(REG0_REG_26__SCAN_IN), .ZN(n2581) );
  OAI211_X1 U33010 ( .C1(n4256), .C2(n3234), .A(n2582), .B(n2581), .ZN(n2583)
         );
  INV_X1 U33020 ( .A(n2583), .ZN(n2584) );
  NAND2_X1 U33030 ( .A1(n2046), .A2(DATAI_26_), .ZN(n4085) );
  NAND2_X1 U33040 ( .A1(n4262), .A2(n4085), .ZN(n2587) );
  XNOR2_X1 U33050 ( .A(n2599), .B(REG3_REG_27__SCAN_IN), .ZN(n3711) );
  NAND2_X1 U33060 ( .A1(n3711), .A2(n2601), .ZN(n2593) );
  INV_X1 U33070 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U33080 ( .A1(n3229), .A2(REG2_REG_27__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U33090 ( .A1(n3230), .A2(REG0_REG_27__SCAN_IN), .ZN(n2588) );
  OAI211_X1 U33100 ( .C1(n2590), .C2(n3234), .A(n2589), .B(n2588), .ZN(n2591)
         );
  INV_X1 U33110 ( .A(n2591), .ZN(n2592) );
  NAND2_X1 U33120 ( .A1(n3943), .A2(n3708), .ZN(n2594) );
  NAND2_X1 U33130 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2596) );
  INV_X1 U33140 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2598) );
  INV_X1 U33150 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2597) );
  OAI21_X1 U33160 ( .B1(n2599), .B2(n2598), .A(n2597), .ZN(n2600) );
  NAND2_X1 U33170 ( .A1(n3691), .A2(n2601), .ZN(n2607) );
  INV_X1 U33180 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U33190 ( .A1(n3229), .A2(REG2_REG_28__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U33200 ( .A1(n3230), .A2(REG0_REG_28__SCAN_IN), .ZN(n2602) );
  OAI211_X1 U33210 ( .C1(n2604), .C2(n3234), .A(n2603), .B(n2602), .ZN(n2605)
         );
  INV_X1 U33220 ( .A(n2605), .ZN(n2606) );
  AND2_X1 U33230 ( .A1(n2046), .A2(DATAI_28_), .ZN(n3690) );
  NAND2_X1 U33240 ( .A1(n3685), .A2(n3690), .ZN(n3252) );
  NAND2_X1 U33250 ( .A1(n4247), .A2(n3683), .ZN(n3257) );
  NAND2_X1 U33260 ( .A1(n3252), .A2(n3257), .ZN(n3317) );
  XNOR2_X1 U33270 ( .A(n2701), .B(n3317), .ZN(n3521) );
  NAND2_X1 U33280 ( .A1(n2613), .A2(IR_REG_31__SCAN_IN), .ZN(n2614) );
  INV_X1 U33290 ( .A(n2668), .ZN(n2615) );
  NAND2_X1 U33300 ( .A1(n2615), .A2(IR_REG_31__SCAN_IN), .ZN(n2616) );
  XNOR2_X1 U33310 ( .A(n2799), .B(n4372), .ZN(n2617) );
  NAND2_X1 U33320 ( .A1(n2617), .A2(n4051), .ZN(n4200) );
  NAND2_X1 U33330 ( .A1(n2618), .A2(n4374), .ZN(n2869) );
  NAND2_X1 U33340 ( .A1(n4200), .A2(n3130), .ZN(n4527) );
  INV_X1 U33350 ( .A(n4527), .ZN(n4321) );
  NOR2_X1 U33360 ( .A1(n2619), .A2(n2723), .ZN(n2620) );
  MUX2_X1 U33370 ( .A(n2723), .B(n2620), .S(IR_REG_28__SCAN_IN), .Z(n2621) );
  INV_X1 U33380 ( .A(n2621), .ZN(n2623) );
  NAND2_X1 U33390 ( .A1(n2623), .A2(n2622), .ZN(n2858) );
  INV_X1 U33400 ( .A(n2858), .ZN(n2728) );
  AND2_X1 U33410 ( .A1(n4372), .A2(n4373), .ZN(n2790) );
  INV_X1 U33420 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U33430 ( .A1(n3229), .A2(REG2_REG_29__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U33440 ( .A1(n3230), .A2(REG0_REG_29__SCAN_IN), .ZN(n2624) );
  OAI211_X1 U33450 ( .C1(n2713), .C2(n3234), .A(n2625), .B(n2624), .ZN(n2626)
         );
  INV_X1 U33460 ( .A(n2626), .ZN(n2627) );
  OAI21_X1 U33470 ( .B1(n4066), .B2(n2628), .A(n2627), .ZN(n3942) );
  INV_X1 U33480 ( .A(n3942), .ZN(n3259) );
  NAND2_X1 U33490 ( .A1(n2858), .A2(n2790), .ZN(n4291) );
  INV_X1 U33500 ( .A(n2618), .ZN(n2730) );
  INV_X1 U33510 ( .A(n4372), .ZN(n2629) );
  INV_X1 U33520 ( .A(n4373), .ZN(n3289) );
  NAND2_X1 U3353 ( .A1(n2730), .A2(n2865), .ZN(n4244) );
  OAI22_X1 U33540 ( .A1(n3259), .A2(n4291), .B1(n3683), .B2(n4244), .ZN(n2630)
         );
  AOI21_X1 U3355 ( .B1(n4287), .B2(n3943), .A(n2630), .ZN(n2659) );
  INV_X1 U3356 ( .A(n3962), .ZN(n2988) );
  NAND2_X1 U3357 ( .A1(n2988), .A2(n2931), .ZN(n2925) );
  NAND2_X1 U3358 ( .A1(n2885), .A2(n3295), .ZN(n2884) );
  NAND2_X1 U3359 ( .A1(n2884), .A2(n3335), .ZN(n2905) );
  NAND2_X1 U3360 ( .A1(n2999), .A2(n2980), .ZN(n3340) );
  NAND2_X1 U3361 ( .A1(n3959), .A2(n3077), .ZN(n3337) );
  NAND2_X1 U3362 ( .A1(n2905), .A2(n3300), .ZN(n2904) );
  INV_X1 U3363 ( .A(n3341), .ZN(n2633) );
  AND2_X1 U3364 ( .A1(n3957), .A2(n3057), .ZN(n2951) );
  NAND2_X1 U3365 ( .A1(n3053), .A2(n3068), .ZN(n3321) );
  NAND2_X1 U3366 ( .A1(n3956), .A2(n3526), .ZN(n3343) );
  NAND2_X1 U3367 ( .A1(n3012), .A2(n3343), .ZN(n2634) );
  NAND2_X1 U3368 ( .A1(n3527), .A2(n3909), .ZN(n3347) );
  NAND2_X1 U3369 ( .A1(n2634), .A2(n3347), .ZN(n3084) );
  INV_X1 U3370 ( .A(n2635), .ZN(n2636) );
  NAND2_X1 U3371 ( .A1(n3115), .A2(n3762), .ZN(n3353) );
  NAND2_X1 U3372 ( .A1(n3954), .A2(n3124), .ZN(n3350) );
  AND2_X1 U3373 ( .A1(n3953), .A2(n3548), .ZN(n3100) );
  NAND2_X1 U3374 ( .A1(n3549), .A2(n3840), .ZN(n3354) );
  NAND2_X1 U3375 ( .A1(n3952), .A2(n3559), .ZN(n3320) );
  NAND2_X1 U3376 ( .A1(n3142), .A2(n3320), .ZN(n2638) );
  NAND2_X1 U3377 ( .A1(n3561), .A2(n3740), .ZN(n3325) );
  NAND2_X1 U3378 ( .A1(n3950), .A2(n3572), .ZN(n3212) );
  NAND2_X1 U3379 ( .A1(n3949), .A2(n3581), .ZN(n2639) );
  NAND2_X1 U3380 ( .A1(n3212), .A2(n2639), .ZN(n3358) );
  INV_X1 U3381 ( .A(n3178), .ZN(n3361) );
  NOR2_X1 U3382 ( .A1(n3358), .A2(n3361), .ZN(n2640) );
  NAND2_X1 U3383 ( .A1(n3179), .A2(n2640), .ZN(n2644) );
  NAND2_X1 U3384 ( .A1(n3574), .A2(n2450), .ZN(n3214) );
  NAND2_X1 U3385 ( .A1(n3176), .A2(n3214), .ZN(n2643) );
  INV_X1 U3386 ( .A(n3358), .ZN(n2642) );
  NOR2_X1 U3387 ( .A1(n3949), .A2(n3581), .ZN(n2641) );
  AOI21_X1 U3388 ( .B1(n2643), .B2(n2642), .A(n2641), .ZN(n3362) );
  NAND2_X1 U3389 ( .A1(n3397), .A2(n2206), .ZN(n2645) );
  NAND2_X1 U3390 ( .A1(n2645), .A2(n3236), .ZN(n3429) );
  INV_X1 U3391 ( .A(n3947), .ZN(n4315) );
  NAND2_X1 U3392 ( .A1(n4315), .A2(n3932), .ZN(n3242) );
  NAND2_X1 U3393 ( .A1(n3947), .A2(n3593), .ZN(n3327) );
  NAND2_X1 U3394 ( .A1(n3242), .A2(n3327), .ZN(n3432) );
  NAND2_X1 U3395 ( .A1(n3430), .A2(n3327), .ZN(n3425) );
  INV_X1 U3396 ( .A(n3420), .ZN(n3424) );
  NAND2_X1 U3397 ( .A1(n3425), .A2(n3424), .ZN(n3423) );
  NAND2_X1 U3398 ( .A1(n3423), .A2(n3329), .ZN(n3463) );
  NAND2_X1 U3399 ( .A1(n3945), .A2(n4225), .ZN(n3287) );
  NAND2_X1 U3400 ( .A1(n3287), .A2(n4213), .ZN(n3238) );
  NAND2_X1 U3401 ( .A1(n4288), .A2(n4202), .ZN(n3237) );
  INV_X1 U3402 ( .A(n3238), .ZN(n2648) );
  NAND2_X1 U3403 ( .A1(n2646), .A2(n3813), .ZN(n3477) );
  NAND2_X1 U3404 ( .A1(n4212), .A2(n3477), .ZN(n2647) );
  NAND2_X1 U3405 ( .A1(n2648), .A2(n2647), .ZN(n2649) );
  NAND2_X1 U3406 ( .A1(n4195), .A2(n3750), .ZN(n3288) );
  NAND2_X1 U3407 ( .A1(n2649), .A2(n3288), .ZN(n4187) );
  NOR2_X1 U3408 ( .A1(n4288), .A2(n4202), .ZN(n2650) );
  OR2_X1 U3409 ( .A1(n4187), .A2(n2650), .ZN(n2651) );
  NAND2_X1 U3410 ( .A1(n2651), .A2(n3237), .ZN(n3369) );
  OR2_X1 U3411 ( .A1(n4193), .A2(n4181), .ZN(n3278) );
  AND2_X1 U3412 ( .A1(n4131), .A2(n3278), .ZN(n3370) );
  NAND2_X1 U3413 ( .A1(n4269), .A2(n4138), .ZN(n3283) );
  AND2_X1 U3414 ( .A1(n3283), .A2(n2652), .ZN(n3375) );
  AND2_X1 U3415 ( .A1(n4193), .A2(n4181), .ZN(n4128) );
  NAND2_X1 U3416 ( .A1(n4131), .A2(n4128), .ZN(n2653) );
  AND2_X1 U3417 ( .A1(n3375), .A2(n2653), .ZN(n3248) );
  OR2_X1 U3418 ( .A1(n4269), .A2(n4138), .ZN(n3284) );
  NAND2_X1 U3419 ( .A1(n2654), .A2(n3284), .ZN(n4113) );
  NOR2_X1 U3420 ( .A1(n4259), .A2(n4267), .ZN(n3274) );
  INV_X1 U3421 ( .A(n4085), .ZN(n4080) );
  NAND2_X1 U3422 ( .A1(n4262), .A2(n4080), .ZN(n2655) );
  INV_X1 U3423 ( .A(n4119), .ZN(n4272) );
  NAND2_X1 U3424 ( .A1(n4272), .A2(n4258), .ZN(n4074) );
  NAND2_X1 U3425 ( .A1(n2655), .A2(n4074), .ZN(n3372) );
  INV_X1 U3426 ( .A(n3372), .ZN(n2656) );
  NAND2_X1 U3427 ( .A1(n4119), .A2(n4100), .ZN(n3282) );
  NAND2_X1 U3428 ( .A1(n4259), .A2(n4267), .ZN(n4093) );
  NAND2_X1 U3429 ( .A1(n3282), .A2(n4093), .ZN(n4075) );
  INV_X1 U3430 ( .A(n4262), .ZN(n3944) );
  AND2_X1 U3431 ( .A1(n3944), .A2(n4085), .ZN(n3260) );
  AOI21_X1 U3432 ( .B1(n2656), .B2(n4075), .A(n3260), .ZN(n3376) );
  XNOR2_X1 U3433 ( .A(n3943), .B(n3708), .ZN(n3508) );
  INV_X1 U3434 ( .A(n3708), .ZN(n4245) );
  OR2_X1 U3435 ( .A1(n3943), .A2(n4245), .ZN(n3251) );
  XOR2_X1 U3436 ( .A(n3317), .B(n2703), .Z(n2658) );
  NAND2_X1 U3437 ( .A1(n2730), .A2(n4373), .ZN(n3269) );
  NAND2_X1 U3438 ( .A1(n4374), .A2(n4372), .ZN(n2657) );
  NAND2_X1 U3439 ( .A1(n2658), .A2(n4197), .ZN(n3516) );
  OAI211_X1 U3440 ( .C1(n3521), .C2(n4321), .A(n2659), .B(n3516), .ZN(n2698)
         );
  AND2_X1 U3441 ( .A1(n2660), .A2(n2667), .ZN(n2661) );
  AOI21_X1 U3442 ( .B1(n2668), .B2(n2661), .A(n2723), .ZN(n2662) );
  MUX2_X1 U3443 ( .A(n2723), .B(n2662), .S(IR_REG_25__SCAN_IN), .Z(n2663) );
  INV_X1 U3444 ( .A(n2663), .ZN(n2666) );
  INV_X1 U3445 ( .A(n2664), .ZN(n2665) );
  NAND2_X1 U3446 ( .A1(n2666), .A2(n2665), .ZN(n2677) );
  NAND2_X1 U3447 ( .A1(n2677), .A2(B_REG_SCAN_IN), .ZN(n2671) );
  MUX2_X1 U3448 ( .A(n2671), .B(B_REG_SCAN_IN), .S(n2678), .Z(n2675) );
  NAND2_X1 U3449 ( .A1(n2665), .A2(IR_REG_31__SCAN_IN), .ZN(n2672) );
  MUX2_X1 U3450 ( .A(IR_REG_31__SCAN_IN), .B(n2672), .S(IR_REG_26__SCAN_IN), 
        .Z(n2674) );
  INV_X1 U3451 ( .A(D_REG_1__SCAN_IN), .ZN(n2738) );
  NAND2_X1 U3452 ( .A1(n2689), .A2(n2738), .ZN(n2871) );
  INV_X1 U3453 ( .A(n2736), .ZN(n2676) );
  NAND2_X1 U3454 ( .A1(n2677), .A2(n2676), .ZN(n2783) );
  NAND2_X1 U3455 ( .A1(n2871), .A2(n2783), .ZN(n2693) );
  XNOR2_X1 U3456 ( .A(n2680), .B(n2679), .ZN(n2743) );
  NAND2_X1 U3457 ( .A1(n2618), .A2(n4051), .ZN(n2789) );
  NAND2_X1 U34580 ( .A1(n2789), .A2(n2790), .ZN(n2795) );
  NAND2_X1 U34590 ( .A1(n2811), .A2(n2795), .ZN(n2870) );
  NOR2_X1 U3460 ( .A1(n3130), .A2(n4373), .ZN(n2812) );
  NOR2_X1 U3461 ( .A1(n2870), .A2(n2812), .ZN(n2692) );
  NOR4_X1 U3462 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2684) );
  NOR4_X1 U3463 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2683) );
  NOR4_X1 U3464 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2682) );
  NOR4_X1 U3465 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2681) );
  NAND4_X1 U3466 ( .A1(n2684), .A2(n2683), .A3(n2682), .A4(n2681), .ZN(n2691)
         );
  NOR2_X1 U34670 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .ZN(n2688) );
  NOR4_X1 U3468 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2687) );
  NOR4_X1 U34690 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2686) );
  NOR4_X1 U3470 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2685) );
  NAND4_X1 U34710 ( .A1(n2688), .A2(n2687), .A3(n2686), .A4(n2685), .ZN(n2690)
         );
  OAI21_X1 U3472 ( .B1(n2691), .B2(n2690), .A(n2689), .ZN(n2784) );
  NAND3_X1 U34730 ( .A1(n2693), .A2(n2692), .A3(n2784), .ZN(n2697) );
  OAI22_X1 U3474 ( .A1(n2732), .A2(D_REG_0__SCAN_IN), .B1(n2736), .B2(n2678), 
        .ZN(n2872) );
  MUX2_X1 U34750 ( .A(REG1_REG_28__SCAN_IN), .B(n2698), .S(n4543), .Z(n2694)
         );
  INV_X1 U3476 ( .A(n2694), .ZN(n2696) );
  NOR2_X1 U34770 ( .A1(n2934), .A2(n2899), .ZN(n2909) );
  NOR2_X1 U3478 ( .A1(n3502), .A2(n3683), .ZN(n2695) );
  NAND2_X1 U34790 ( .A1(n2696), .A2(n2285), .ZN(U3546) );
  INV_X1 U3480 ( .A(n2872), .ZN(n2785) );
  MUX2_X1 U34810 ( .A(REG0_REG_28__SCAN_IN), .B(n2698), .S(n4536), .Z(n2699)
         );
  INV_X1 U3482 ( .A(n2699), .ZN(n2700) );
  NAND2_X1 U34830 ( .A1(n2700), .A2(n2284), .ZN(U3514) );
  NAND2_X1 U3484 ( .A1(n2046), .A2(DATAI_29_), .ZN(n4063) );
  XNOR2_X1 U34850 ( .A(n3942), .B(n4063), .ZN(n3318) );
  INV_X1 U3486 ( .A(n3252), .ZN(n2702) );
  XNOR2_X1 U34870 ( .A(n2704), .B(n3318), .ZN(n2710) );
  AND2_X1 U3488 ( .A1(n2706), .A2(n2705), .ZN(n2835) );
  AOI21_X1 U34890 ( .B1(B_REG_SCAN_IN), .B2(n2835), .A(n4291), .ZN(n4056) );
  INV_X1 U3490 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2709) );
  NAND2_X1 U34910 ( .A1(n3229), .A2(REG2_REG_30__SCAN_IN), .ZN(n2708) );
  NAND2_X1 U3492 ( .A1(n3230), .A2(REG0_REG_30__SCAN_IN), .ZN(n2707) );
  OAI211_X1 U34930 ( .C1(n3234), .C2(n2709), .A(n2708), .B(n2707), .ZN(n3941)
         );
  NAND2_X1 U3494 ( .A1(n4247), .A2(n4287), .ZN(n2711) );
  OAI21_X1 U34950 ( .B1(n2714), .B2(n4063), .A(n4239), .ZN(n4067) );
  NAND2_X1 U3496 ( .A1(n2716), .A2(n2715), .ZN(U3547) );
  INV_X1 U34970 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2717) );
  INV_X1 U3498 ( .A(n4504), .ZN(n2735) );
  NOR2_X1 U34990 ( .A1(n2800), .A2(n2735), .ZN(U4043) );
  INV_X1 U3500 ( .A(DATAI_30_), .ZN(n2720) );
  NAND2_X1 U35010 ( .A1(n2305), .A2(STATE_REG_SCAN_IN), .ZN(n2719) );
  OAI21_X1 U3502 ( .B1(STATE_REG_SCAN_IN), .B2(n2720), .A(n2719), .ZN(U3322)
         );
  INV_X1 U35030 ( .A(DATAI_26_), .ZN(n2722) );
  NAND2_X1 U3504 ( .A1(n2736), .A2(STATE_REG_SCAN_IN), .ZN(n2721) );
  OAI21_X1 U35050 ( .B1(STATE_REG_SCAN_IN), .B2(n2722), .A(n2721), .ZN(U3326)
         );
  INV_X1 U35060 ( .A(DATAI_31_), .ZN(n4651) );
  OR4_X1 U35070 ( .A1(n2304), .A2(IR_REG_30__SCAN_IN), .A3(n2723), .A4(U3149), 
        .ZN(n2724) );
  OAI21_X1 U35080 ( .B1(STATE_REG_SCAN_IN), .B2(n4651), .A(n2724), .ZN(U3321)
         );
  INV_X1 U35090 ( .A(DATAI_24_), .ZN(n4665) );
  NAND2_X1 U35100 ( .A1(n2678), .A2(STATE_REG_SCAN_IN), .ZN(n2725) );
  OAI21_X1 U35110 ( .B1(STATE_REG_SCAN_IN), .B2(n4665), .A(n2725), .ZN(U3328)
         );
  INV_X1 U35120 ( .A(DATAI_27_), .ZN(n2727) );
  NAND2_X1 U35130 ( .A1(n2835), .A2(STATE_REG_SCAN_IN), .ZN(n2726) );
  OAI21_X1 U35140 ( .B1(STATE_REG_SCAN_IN), .B2(n2727), .A(n2726), .ZN(U3325)
         );
  INV_X1 U35150 ( .A(DATAI_28_), .ZN(n4592) );
  NAND2_X1 U35160 ( .A1(n2728), .A2(STATE_REG_SCAN_IN), .ZN(n2729) );
  OAI21_X1 U35170 ( .B1(STATE_REG_SCAN_IN), .B2(n4592), .A(n2729), .ZN(U3324)
         );
  INV_X1 U35180 ( .A(DATAI_20_), .ZN(n4666) );
  NAND2_X1 U35190 ( .A1(n2730), .A2(STATE_REG_SCAN_IN), .ZN(n2731) );
  OAI21_X1 U35200 ( .B1(STATE_REG_SCAN_IN), .B2(n4666), .A(n2731), .ZN(U3332)
         );
  INV_X1 U35210 ( .A(D_REG_0__SCAN_IN), .ZN(n2734) );
  NOR3_X1 U35220 ( .A1(n2736), .A2(n2735), .A3(n2678), .ZN(n2733) );
  AOI21_X1 U35230 ( .B1(n4503), .B2(n2734), .A(n2733), .ZN(U3458) );
  NOR3_X1 U35240 ( .A1(n4371), .A2(n2736), .A3(n2735), .ZN(n2737) );
  AOI21_X1 U35250 ( .B1(n4503), .B2(n2738), .A(n2737), .ZN(U3459) );
  INV_X1 U35260 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2739) );
  AND2_X1 U35270 ( .A1(n2835), .A2(n2739), .ZN(n2740) );
  NOR2_X1 U35280 ( .A1(n2858), .A2(n2740), .ZN(n2838) );
  OAI21_X1 U35290 ( .B1(REG1_REG_0__SCAN_IN), .B2(n2835), .A(n2838), .ZN(n2741) );
  MUX2_X1 U35300 ( .A(n2741), .B(n2838), .S(IR_REG_0__SCAN_IN), .Z(n2751) );
  INV_X1 U35310 ( .A(n2811), .ZN(n2797) );
  INV_X1 U35320 ( .A(n2743), .ZN(n2742) );
  NAND2_X1 U35330 ( .A1(n2742), .A2(STATE_REG_SCAN_IN), .ZN(n3395) );
  NAND2_X1 U35340 ( .A1(n2797), .A2(n3395), .ZN(n2747) );
  NAND2_X1 U35350 ( .A1(n2743), .A2(n2790), .ZN(n2744) );
  AND2_X1 U35360 ( .A1(n2046), .A2(n2744), .ZN(n2745) );
  INV_X1 U35370 ( .A(n2768), .ZN(n2750) );
  INV_X1 U35380 ( .A(n2835), .ZN(n2765) );
  NAND3_X1 U35390 ( .A1(n4484), .A2(IR_REG_0__SCAN_IN), .A3(n2333), .ZN(n2749)
         );
  INV_X1 U35400 ( .A(n2745), .ZN(n2746) );
  AOI22_X1 U35410 ( .A1(n4482), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2748) );
  OAI211_X1 U35420 ( .C1(n2751), .C2(n2750), .A(n2749), .B(n2748), .ZN(U3240)
         );
  NOR2_X1 U35430 ( .A1(n4482), .A2(n3961), .ZN(U3148) );
  XNOR2_X1 U35440 ( .A(n4381), .B(n2342), .ZN(n3985) );
  XNOR2_X1 U35450 ( .A(n4382), .B(n2326), .ZN(n3965) );
  AND2_X1 U35460 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3964) );
  NAND2_X1 U35470 ( .A1(n3965), .A2(n3964), .ZN(n3963) );
  NAND2_X1 U35480 ( .A1(n4382), .A2(REG1_REG_1__SCAN_IN), .ZN(n2752) );
  NAND2_X1 U35490 ( .A1(n3963), .A2(n2752), .ZN(n3984) );
  NAND2_X1 U35500 ( .A1(n3985), .A2(n3984), .ZN(n3983) );
  NAND2_X1 U35510 ( .A1(n4381), .A2(REG1_REG_2__SCAN_IN), .ZN(n2753) );
  NAND2_X1 U35520 ( .A1(n3983), .A2(n2753), .ZN(n2754) );
  XNOR2_X1 U35530 ( .A(n2754), .B(n2193), .ZN(n3992) );
  NAND2_X1 U35540 ( .A1(n3992), .A2(REG1_REG_3__SCAN_IN), .ZN(n3991) );
  NAND2_X1 U35550 ( .A1(n2754), .A2(n4380), .ZN(n2755) );
  NAND2_X1 U35560 ( .A1(n3991), .A2(n2755), .ZN(n2757) );
  INV_X1 U35570 ( .A(n4379), .ZN(n2844) );
  XNOR2_X1 U35580 ( .A(n2757), .B(n2844), .ZN(n2841) );
  NAND2_X1 U35590 ( .A1(n2841), .A2(REG1_REG_4__SCAN_IN), .ZN(n2840) );
  INV_X1 U35600 ( .A(n2840), .ZN(n2756) );
  XNOR2_X1 U35610 ( .A(n4378), .B(REG1_REG_5__SCAN_IN), .ZN(n2758) );
  INV_X1 U35620 ( .A(n4484), .ZN(n2921) );
  AOI211_X1 U35630 ( .C1(n2759), .C2(n2758), .A(n2777), .B(n2921), .ZN(n2773)
         );
  INV_X1 U35640 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3977) );
  INV_X1 U35650 ( .A(n4381), .ZN(n3975) );
  MUX2_X1 U35660 ( .A(REG2_REG_2__SCAN_IN), .B(n3977), .S(n4381), .Z(n2762) );
  INV_X1 U35670 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2984) );
  MUX2_X1 U35680 ( .A(REG2_REG_1__SCAN_IN), .B(n2984), .S(n4382), .Z(n3967) );
  AND2_X1 U35690 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2760) );
  NAND2_X1 U35700 ( .A1(n3967), .A2(n2760), .ZN(n3979) );
  NAND2_X1 U35710 ( .A1(n4382), .A2(REG2_REG_1__SCAN_IN), .ZN(n3978) );
  NAND2_X1 U35720 ( .A1(n3979), .A2(n3978), .ZN(n2761) );
  XNOR2_X1 U35730 ( .A(n2763), .B(n4379), .ZN(n2839) );
  INV_X1 U35740 ( .A(n2763), .ZN(n2764) );
  AOI22_X1 U35750 ( .A1(n2839), .A2(REG2_REG_4__SCAN_IN), .B1(n4379), .B2(
        n2764), .ZN(n2767) );
  INV_X1 U35760 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3064) );
  MUX2_X1 U35770 ( .A(REG2_REG_5__SCAN_IN), .B(n3064), .S(n2770), .Z(n2766) );
  NOR2_X1 U35780 ( .A1(n2767), .A2(n2766), .ZN(n2774) );
  NOR2_X1 U35790 ( .A1(n2858), .A2(n2765), .ZN(n3392) );
  INV_X1 U35800 ( .A(n4429), .ZN(n4478) );
  AOI211_X1 U35810 ( .C1(n2767), .C2(n2766), .A(n2774), .B(n4478), .ZN(n2772)
         );
  NAND2_X1 U3582 ( .A1(n2768), .A2(n2858), .ZN(n4489) );
  NOR2_X1 U3583 ( .A1(STATE_REG_SCAN_IN), .A2(n2375), .ZN(n3059) );
  AOI21_X1 U3584 ( .B1(n4482), .B2(ADDR_REG_5__SCAN_IN), .A(n3059), .ZN(n2769)
         );
  OAI21_X1 U3585 ( .B1(n4489), .B2(n2770), .A(n2769), .ZN(n2771) );
  OR3_X1 U3586 ( .A1(n2773), .A2(n2772), .A3(n2771), .ZN(U3245) );
  AOI21_X1 U3587 ( .B1(n4378), .B2(REG2_REG_5__SCAN_IN), .A(n2774), .ZN(n2817)
         );
  XNOR2_X1 U3588 ( .A(n2817), .B(n4377), .ZN(n2819) );
  XNOR2_X1 U3589 ( .A(n2819), .B(REG2_REG_6__SCAN_IN), .ZN(n2782) );
  INV_X1 U3590 ( .A(n4489), .ZN(n3990) );
  NOR2_X1 U3591 ( .A1(STATE_REG_SCAN_IN), .A2(n2775), .ZN(n3908) );
  AOI21_X1 U3592 ( .B1(n4482), .B2(ADDR_REG_6__SCAN_IN), .A(n3908), .ZN(n2776)
         );
  INV_X1 U3593 ( .A(n2776), .ZN(n2780) );
  INV_X1 U3594 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3018) );
  NOR2_X1 U3595 ( .A1(n2778), .A2(n3018), .ZN(n2823) );
  AOI211_X1 U3596 ( .C1(n2778), .C2(n3018), .A(n2921), .B(n2823), .ZN(n2779)
         );
  AOI211_X1 U3597 ( .C1(n3990), .C2(n4377), .A(n2780), .B(n2779), .ZN(n2781)
         );
  OAI21_X1 U3598 ( .B1(n2782), .B2(n4478), .A(n2781), .ZN(U3246) );
  AND2_X1 U3599 ( .A1(n2784), .A2(n2783), .ZN(n2874) );
  INV_X1 U3600 ( .A(n2861), .ZN(n2794) );
  INV_X1 U3601 ( .A(n2799), .ZN(n2786) );
  NAND2_X2 U3602 ( .A1(n2786), .A2(n2800), .ZN(n3579) );
  NAND2_X1 U3603 ( .A1(n4051), .A2(n4372), .ZN(n2849) );
  INV_X1 U3604 ( .A(n2849), .ZN(n2787) );
  AND2_X1 U3605 ( .A1(n2787), .A2(n4504), .ZN(n2788) );
  NAND2_X1 U3606 ( .A1(n2794), .A2(n3391), .ZN(n2975) );
  INV_X1 U3607 ( .A(n2975), .ZN(n2798) );
  NAND2_X1 U3608 ( .A1(n2789), .A2(n2865), .ZN(n2792) );
  INV_X1 U3609 ( .A(n2790), .ZN(n2791) );
  NAND2_X1 U3610 ( .A1(n2792), .A2(n2791), .ZN(n2805) );
  NAND2_X1 U3611 ( .A1(n2805), .A2(n4244), .ZN(n2793) );
  NAND2_X1 U3612 ( .A1(n2794), .A2(n2793), .ZN(n2796) );
  NAND2_X1 U3613 ( .A1(n2796), .A2(n2795), .ZN(n2974) );
  NOR3_X1 U3614 ( .A1(n2798), .A2(n2974), .A3(n2797), .ZN(n2902) );
  INV_X1 U3615 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2816) );
  INV_X1 U3616 ( .A(n2800), .ZN(n2973) );
  OAI22_X1 U3617 ( .A1(n2988), .A2(n3579), .B1(n3682), .B2(n2867), .ZN(n2848)
         );
  AOI21_X1 U3618 ( .B1(n2973), .B2(REG1_REG_0__SCAN_IN), .A(n2848), .ZN(n2803)
         );
  NOR2_X1 U3619 ( .A1(n2803), .A2(n2804), .ZN(n2850) );
  AOI21_X1 U3620 ( .B1(n2804), .B2(n2803), .A(n2850), .ZN(n2833) );
  INV_X1 U3621 ( .A(n2805), .ZN(n2806) );
  AND2_X1 U3622 ( .A1(n2811), .A2(n2806), .ZN(n2807) );
  NAND2_X1 U3623 ( .A1(n2833), .A2(n3929), .ZN(n2815) );
  AND2_X1 U3624 ( .A1(n3391), .A2(n2858), .ZN(n2809) );
  AND2_X1 U3625 ( .A1(n2811), .A2(n4310), .ZN(n2810) );
  NAND2_X1 U3626 ( .A1(n2861), .A2(n2810), .ZN(n2813) );
  AOI22_X1 U3627 ( .A1(n2808), .A2(n3931), .B1(n3933), .B2(n2931), .ZN(n2814)
         );
  OAI211_X1 U3628 ( .C1(n2902), .C2(n2816), .A(n2815), .B(n2814), .ZN(U3229)
         );
  INV_X1 U3629 ( .A(n2817), .ZN(n2818) );
  INV_X1 U3630 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3091) );
  MUX2_X1 U3631 ( .A(n3091), .B(REG2_REG_7__SCAN_IN), .S(n4376), .Z(n2820) );
  AOI211_X1 U3632 ( .C1(n2821), .C2(n2820), .A(n4478), .B(n2915), .ZN(n2832)
         );
  INV_X1 U3633 ( .A(n2822), .ZN(n2824) );
  INV_X1 U3634 ( .A(n4376), .ZN(n2829) );
  INV_X1 U3635 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4541) );
  AND2_X1 U3636 ( .A1(n2829), .A2(n4541), .ZN(n2912) );
  INV_X1 U3637 ( .A(n2912), .ZN(n2825) );
  NAND2_X1 U3638 ( .A1(n4376), .A2(REG1_REG_7__SCAN_IN), .ZN(n2913) );
  NAND2_X1 U3639 ( .A1(n2825), .A2(n2913), .ZN(n2827) );
  OAI21_X1 U3640 ( .B1(n2914), .B2(n2827), .A(n4484), .ZN(n2826) );
  AOI21_X1 U3641 ( .B1(n2914), .B2(n2827), .A(n2826), .ZN(n2831) );
  INV_X1 U3642 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4690) );
  NOR2_X1 U3643 ( .A1(STATE_REG_SCAN_IN), .A2(n4690), .ZN(n3700) );
  AOI21_X1 U3644 ( .B1(n4482), .B2(ADDR_REG_7__SCAN_IN), .A(n3700), .ZN(n2828)
         );
  OAI21_X1 U3645 ( .B1(n4489), .B2(n2829), .A(n2828), .ZN(n2830) );
  OR3_X1 U3646 ( .A1(n2832), .A2(n2831), .A3(n2830), .ZN(U3247) );
  INV_X1 U3647 ( .A(n2833), .ZN(n2836) );
  NAND2_X1 U3648 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3966) );
  AOI21_X1 U3649 ( .B1(n2835), .B2(n3966), .A(n2858), .ZN(n2834) );
  OAI21_X1 U3650 ( .B1(n2836), .B2(n2835), .A(n2834), .ZN(n2837) );
  OAI211_X1 U3651 ( .C1(IR_REG_0__SCAN_IN), .C2(n2838), .A(n2837), .B(n3961), 
        .ZN(n3989) );
  XOR2_X1 U3652 ( .A(REG2_REG_4__SCAN_IN), .B(n2839), .Z(n2846) );
  OAI211_X1 U3653 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2841), .A(n4484), .B(n2840), 
        .ZN(n2843) );
  AND2_X1 U3654 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3830) );
  AOI21_X1 U3655 ( .B1(n4482), .B2(ADDR_REG_4__SCAN_IN), .A(n3830), .ZN(n2842)
         );
  OAI211_X1 U3656 ( .C1(n4489), .C2(n2844), .A(n2843), .B(n2842), .ZN(n2845)
         );
  AOI21_X1 U3657 ( .B1(n4429), .B2(n2846), .A(n2845), .ZN(n2847) );
  NAND2_X1 U3658 ( .A1(n3989), .A2(n2847), .ZN(U3244) );
  INV_X1 U3659 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2986) );
  INV_X1 U3660 ( .A(n2848), .ZN(n2851) );
  NAND2_X1 U3661 ( .A1(n2932), .A2(n3529), .ZN(n2852) );
  NAND2_X1 U3662 ( .A1(n2853), .A2(n2852), .ZN(n2892) );
  OAI22_X1 U3663 ( .A1(n2998), .A2(n3579), .B1(n3682), .B2(n2987), .ZN(n2854)
         );
  INV_X2 U3664 ( .A(n3667), .ZN(n2971) );
  XNOR2_X1 U3665 ( .A(n2854), .B(n2971), .ZN(n2891) );
  XNOR2_X1 U3666 ( .A(n2892), .B(n2891), .ZN(n2855) );
  AOI211_X1 U3667 ( .C1(n2856), .C2(n2855), .A(n3925), .B(n2894), .ZN(n2857)
         );
  INV_X1 U3668 ( .A(n2857), .ZN(n2864) );
  INV_X1 U3669 ( .A(n3391), .ZN(n2859) );
  NOR2_X1 U3670 ( .A1(n2859), .A2(n2858), .ZN(n2860) );
  INV_X1 U3671 ( .A(n3931), .ZN(n3875) );
  OAI22_X1 U3672 ( .A1(n2988), .A2(n3919), .B1(n3875), .B2(n2352), .ZN(n2862)
         );
  AOI21_X1 U3673 ( .B1(n2932), .B2(n3933), .A(n2862), .ZN(n2863) );
  OAI211_X1 U3674 ( .C1(n2902), .C2(n2986), .A(n2864), .B(n2863), .ZN(U3219)
         );
  INV_X1 U3675 ( .A(n2865), .ZN(n2866) );
  NOR2_X1 U3676 ( .A1(n2867), .A2(n2866), .ZN(n4518) );
  NAND2_X1 U3677 ( .A1(n3962), .A2(n2867), .ZN(n3333) );
  AND2_X1 U3678 ( .A1(n2925), .A2(n3333), .ZN(n3279) );
  INV_X1 U3679 ( .A(n4200), .ZN(n3166) );
  NOR2_X1 U3680 ( .A1(n3166), .A2(n4197), .ZN(n2868) );
  OAI22_X1 U3681 ( .A1(n3279), .A2(n2868), .B1(n2998), .B2(n4291), .ZN(n4517)
         );
  AOI21_X1 U3682 ( .B1(n4518), .B2(n2869), .A(n4517), .ZN(n2879) );
  INV_X1 U3683 ( .A(n2870), .ZN(n2873) );
  NAND4_X1 U3684 ( .A1(n2874), .A2(n2873), .A3(n2872), .A4(n2871), .ZN(n2875)
         );
  NAND2_X2 U3685 ( .A1(n2875), .A2(n4490), .ZN(n4493) );
  INV_X1 U3686 ( .A(n4490), .ZN(n4227) );
  AOI22_X1 U3687 ( .A1(n4229), .A2(REG2_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(n4227), .ZN(n2878) );
  INV_X1 U3688 ( .A(n3279), .ZN(n4519) );
  OR2_X1 U3689 ( .A1(n2799), .A2(n4051), .ZN(n3025) );
  INV_X1 U3690 ( .A(n3025), .ZN(n2876) );
  NAND2_X1 U3691 ( .A1(n4493), .A2(n2876), .ZN(n4210) );
  INV_X1 U3692 ( .A(n4210), .ZN(n4498) );
  NAND2_X1 U3693 ( .A1(n4519), .A2(n4498), .ZN(n2877) );
  OAI211_X1 U3694 ( .C1(n2879), .C2(n4229), .A(n2878), .B(n2877), .ZN(U3290)
         );
  INV_X1 U3695 ( .A(n3130), .ZN(n4524) );
  OAI21_X1 U3696 ( .B1(n2880), .B2(n2882), .A(n2881), .ZN(n2995) );
  AOI22_X1 U3697 ( .A1(n3959), .A2(n4311), .B1(n2899), .B2(n4310), .ZN(n2883)
         );
  OAI21_X1 U3698 ( .B1(n2998), .B2(n4314), .A(n2883), .ZN(n2888) );
  OAI21_X1 U3699 ( .B1(n3295), .B2(n2885), .A(n2884), .ZN(n2886) );
  AOI22_X1 U3700 ( .A1(n2995), .A2(n3166), .B1(n4197), .B2(n2886), .ZN(n2996)
         );
  INV_X1 U3701 ( .A(n2996), .ZN(n2887) );
  AOI211_X1 U3702 ( .C1(n4524), .C2(n2995), .A(n2888), .B(n2887), .ZN(n2959)
         );
  INV_X1 U3703 ( .A(n4362), .ZN(n4332) );
  XNOR2_X1 U3704 ( .A(n2934), .B(n2997), .ZN(n3002) );
  AOI22_X1 U3705 ( .A1(n4332), .A2(n3002), .B1(REG0_REG_2__SCAN_IN), .B2(n4534), .ZN(n2889) );
  OAI21_X1 U3706 ( .B1(n2959), .B2(n4534), .A(n2889), .ZN(U3471) );
  INV_X1 U3707 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3972) );
  OAI22_X1 U3708 ( .A1(n2352), .A2(n3684), .B1(n3579), .B2(n2997), .ZN(n2965)
         );
  OAI22_X1 U3709 ( .A1(n2352), .A2(n3579), .B1(n3682), .B2(n2997), .ZN(n2890)
         );
  XNOR2_X1 U3710 ( .A(n2890), .B(n2971), .ZN(n2964) );
  XOR2_X1 U3711 ( .A(n2965), .B(n2964), .Z(n2896) );
  AND2_X1 U3712 ( .A1(n2892), .A2(n2891), .ZN(n2893) );
  OAI21_X1 U3713 ( .B1(n2896), .B2(n2895), .A(n2967), .ZN(n2897) );
  NAND2_X1 U3714 ( .A1(n2897), .A2(n3929), .ZN(n2901) );
  OAI22_X1 U3715 ( .A1(n2999), .A2(n3875), .B1(n3919), .B2(n2998), .ZN(n2898)
         );
  AOI21_X1 U3716 ( .B1(n2899), .B2(n3933), .A(n2898), .ZN(n2900) );
  OAI211_X1 U3717 ( .C1(n2902), .C2(n3972), .A(n2901), .B(n2900), .ZN(U3234)
         );
  XOR2_X1 U3718 ( .A(n2903), .B(n3300), .Z(n3080) );
  OAI22_X1 U3719 ( .A1(n3065), .A2(n4291), .B1(n4244), .B2(n3077), .ZN(n2908)
         );
  OAI21_X1 U3720 ( .B1(n3300), .B2(n2905), .A(n2904), .ZN(n2906) );
  AOI22_X1 U3721 ( .A1(n2906), .A2(n4197), .B1(n4287), .B2(n3960), .ZN(n3083)
         );
  INV_X1 U3722 ( .A(n3083), .ZN(n2907) );
  AOI211_X1 U3723 ( .C1(n4527), .C2(n3080), .A(n2908), .B(n2907), .ZN(n2961)
         );
  INV_X1 U3724 ( .A(n2909), .ZN(n2910) );
  AOI21_X1 U3725 ( .B1(n2980), .B2(n2910), .A(n2937), .ZN(n3079) );
  AOI22_X1 U3726 ( .A1(n3079), .A2(n4332), .B1(REG0_REG_3__SCAN_IN), .B2(n4534), .ZN(n2911) );
  OAI21_X1 U3727 ( .B1(n2961), .B2(n4534), .A(n2911), .ZN(U3473) );
  AOI21_X1 U3728 ( .B1(n2914), .B2(n2913), .A(n2912), .ZN(n4026) );
  XOR2_X1 U3729 ( .A(REG1_REG_8__SCAN_IN), .B(n4028), .Z(n2922) );
  INV_X1 U3730 ( .A(n4375), .ZN(n4027) );
  XNOR2_X1 U3731 ( .A(REG2_REG_8__SCAN_IN), .B(n4006), .ZN(n2916) );
  NAND2_X1 U3732 ( .A1(n4429), .A2(n2916), .ZN(n2917) );
  NAND2_X1 U3733 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3760) );
  NAND2_X1 U3734 ( .A1(n2917), .A2(n3760), .ZN(n2918) );
  AOI21_X1 U3735 ( .B1(n4482), .B2(ADDR_REG_8__SCAN_IN), .A(n2918), .ZN(n2920)
         );
  NAND2_X1 U3736 ( .A1(n3990), .A2(n4375), .ZN(n2919) );
  OAI211_X1 U3737 ( .C1(n2922), .C2(n2921), .A(n2920), .B(n2919), .ZN(U3248)
         );
  INV_X1 U3738 ( .A(n2994), .ZN(n2928) );
  OAI21_X1 U3739 ( .B1(n3297), .B2(n2171), .A(n2926), .ZN(n2927) );
  AOI22_X1 U3740 ( .A1(n2928), .A2(n3166), .B1(n2927), .B2(n4197), .ZN(n2983)
         );
  OAI22_X1 U3741 ( .A1(n2352), .A2(n4291), .B1(n4244), .B2(n2987), .ZN(n2929)
         );
  AOI21_X1 U3742 ( .B1(n4287), .B2(n3962), .A(n2929), .ZN(n2930) );
  OAI211_X1 U3743 ( .C1(n3130), .C2(n2994), .A(n2983), .B(n2930), .ZN(n3009)
         );
  NAND2_X1 U3744 ( .A1(n2932), .A2(n2931), .ZN(n2933) );
  NAND2_X1 U3745 ( .A1(n2934), .A2(n2933), .ZN(n3007) );
  OAI22_X1 U3746 ( .A1(n4305), .A2(n3007), .B1(n4543), .B2(n2326), .ZN(n2935)
         );
  AOI21_X1 U3747 ( .B1(n3009), .B2(n4543), .A(n2935), .ZN(n2936) );
  INV_X1 U3748 ( .A(n2936), .ZN(U3519) );
  OAI211_X1 U3749 ( .C1(n2937), .C2(n3046), .A(n4317), .B(n2956), .ZN(n4521)
         );
  NOR2_X1 U3750 ( .A1(n4521), .A2(n4374), .ZN(n2947) );
  XOR2_X1 U3751 ( .A(n3296), .B(n2939), .Z(n2946) );
  NAND2_X1 U3752 ( .A1(n2940), .A2(n3296), .ZN(n2941) );
  AND2_X1 U3753 ( .A1(n2942), .A2(n2941), .ZN(n4525) );
  AOI22_X1 U3754 ( .A1(n3959), .A2(n4287), .B1(n3831), .B2(n4310), .ZN(n2943)
         );
  OAI21_X1 U3755 ( .B1(n3053), .B2(n4291), .A(n2943), .ZN(n2944) );
  AOI21_X1 U3756 ( .B1(n4525), .B2(n3166), .A(n2944), .ZN(n2945) );
  OAI21_X1 U3757 ( .B1(n2946), .B2(n4222), .A(n2945), .ZN(n4522) );
  AOI211_X1 U3758 ( .C1(n4227), .C2(n3832), .A(n2947), .B(n4522), .ZN(n2949)
         );
  AOI22_X1 U3759 ( .A1(n4525), .A2(n4498), .B1(REG2_REG_4__SCAN_IN), .B2(n4229), .ZN(n2948) );
  OAI21_X1 U3760 ( .B1(n2949), .B2(n4229), .A(n2948), .ZN(U3286) );
  INV_X1 U3761 ( .A(n2951), .ZN(n3344) );
  AND2_X1 U3762 ( .A1(n3344), .A2(n3321), .ZN(n3285) );
  XNOR2_X1 U3763 ( .A(n2950), .B(n3285), .ZN(n3072) );
  XOR2_X1 U3764 ( .A(n3285), .B(n2952), .Z(n2953) );
  NAND2_X1 U3765 ( .A1(n2953), .A2(n4197), .ZN(n3074) );
  AOI22_X1 U3766 ( .A1(n3956), .A2(n4311), .B1(n4310), .B2(n3068), .ZN(n2954)
         );
  OAI211_X1 U3767 ( .C1(n3065), .C2(n4314), .A(n3074), .B(n2954), .ZN(n2955)
         );
  AOI21_X1 U3768 ( .B1(n3072), .B2(n4527), .A(n2955), .ZN(n2963) );
  AOI21_X1 U3769 ( .B1(n3068), .B2(n2956), .A(n3016), .ZN(n3062) );
  AOI22_X1 U3770 ( .A1(n3062), .A2(n4332), .B1(REG0_REG_5__SCAN_IN), .B2(n4534), .ZN(n2957) );
  OAI21_X1 U3771 ( .B1(n2963), .B2(n4534), .A(n2957), .ZN(U3477) );
  INV_X1 U3772 ( .A(n4305), .ZN(n4252) );
  AOI22_X1 U3773 ( .A1(n4252), .A2(n3002), .B1(REG1_REG_2__SCAN_IN), .B2(n4540), .ZN(n2958) );
  OAI21_X1 U3774 ( .B1(n2959), .B2(n4540), .A(n2958), .ZN(U3520) );
  AOI22_X1 U3775 ( .A1(n3079), .A2(n4252), .B1(REG1_REG_3__SCAN_IN), .B2(n4540), .ZN(n2960) );
  OAI21_X1 U3776 ( .B1(n2961), .B2(n4540), .A(n2960), .ZN(U3521) );
  AOI22_X1 U3777 ( .A1(n3062), .A2(n4252), .B1(REG1_REG_5__SCAN_IN), .B2(n4540), .ZN(n2962) );
  OAI21_X1 U3778 ( .B1(n2963), .B2(n4540), .A(n2962), .ZN(U3523) );
  OAI22_X1 U3779 ( .A1(n2999), .A2(n3684), .B1(n3657), .B2(n3077), .ZN(n3038)
         );
  NAND2_X1 U3780 ( .A1(n3959), .A2(n3529), .ZN(n2970) );
  NAND2_X1 U3781 ( .A1(n2980), .A2(n2968), .ZN(n2969) );
  NAND2_X1 U3782 ( .A1(n2970), .A2(n2969), .ZN(n2972) );
  XNOR2_X1 U3783 ( .A(n2972), .B(n2971), .ZN(n3039) );
  XOR2_X1 U3784 ( .A(n3038), .B(n3039), .Z(n3042) );
  XOR2_X1 U3785 ( .A(n3043), .B(n3042), .Z(n2982) );
  OAI22_X1 U3786 ( .A1(n2352), .A2(n3919), .B1(n3875), .B2(n3065), .ZN(n2979)
         );
  OAI21_X1 U3787 ( .B1(n2974), .B2(n2973), .A(STATE_REG_SCAN_IN), .ZN(n2977)
         );
  AND2_X1 U3788 ( .A1(n2975), .A2(n3395), .ZN(n2976) );
  MUX2_X1 U3789 ( .A(n3936), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2978) );
  AOI211_X1 U3790 ( .C1(n2980), .C2(n3933), .A(n2979), .B(n2978), .ZN(n2981)
         );
  OAI21_X1 U3791 ( .B1(n2982), .B2(n3925), .A(n2981), .ZN(U3215) );
  MUX2_X1 U3792 ( .A(n2984), .B(n2983), .S(n4493), .Z(n2993) );
  NAND2_X1 U3793 ( .A1(n4493), .A2(n4051), .ZN(n3487) );
  INV_X1 U3794 ( .A(n3007), .ZN(n2991) );
  NAND2_X1 U3795 ( .A1(n4493), .A2(n4310), .ZN(n4180) );
  OAI22_X1 U3796 ( .A1(n4180), .A2(n2987), .B1(n2986), .B2(n4490), .ZN(n2990)
         );
  INV_X1 U3797 ( .A(n4174), .ZN(n4105) );
  INV_X1 U3798 ( .A(n4175), .ZN(n4106) );
  OAI22_X1 U3799 ( .A1(n2988), .A2(n4105), .B1(n4106), .B2(n2352), .ZN(n2989)
         );
  AOI211_X1 U3800 ( .C1(n4497), .C2(n2991), .A(n2990), .B(n2989), .ZN(n2992)
         );
  OAI211_X1 U3801 ( .C1(n2994), .C2(n4210), .A(n2993), .B(n2992), .ZN(U3289)
         );
  INV_X1 U3802 ( .A(n2995), .ZN(n3005) );
  MUX2_X1 U3803 ( .A(n3977), .B(n2996), .S(n4493), .Z(n3004) );
  OAI22_X1 U3804 ( .A1(n4180), .A2(n2997), .B1(n3972), .B2(n4490), .ZN(n3001)
         );
  OAI22_X1 U3805 ( .A1(n2999), .A2(n4106), .B1(n4105), .B2(n2998), .ZN(n3000)
         );
  AOI211_X1 U3806 ( .C1(n4497), .C2(n3002), .A(n3001), .B(n3000), .ZN(n3003)
         );
  OAI211_X1 U3807 ( .C1(n3005), .C2(n4210), .A(n3004), .B(n3003), .ZN(U3288)
         );
  INV_X1 U3808 ( .A(REG0_REG_1__SCAN_IN), .ZN(n3006) );
  OAI22_X1 U3809 ( .A1(n4362), .A2(n3007), .B1(n4536), .B2(n3006), .ZN(n3008)
         );
  AOI21_X1 U3810 ( .B1(n3009), .B2(n4536), .A(n3008), .ZN(n3010) );
  INV_X1 U3811 ( .A(n3010), .ZN(U3469) );
  AND2_X1 U3812 ( .A1(n3347), .A2(n3343), .ZN(n3298) );
  XOR2_X1 U3813 ( .A(n3011), .B(n3298), .Z(n3036) );
  XNOR2_X1 U3814 ( .A(n3012), .B(n3298), .ZN(n3033) );
  AOI22_X1 U3815 ( .A1(n3955), .A2(n4311), .B1(n3909), .B2(n4310), .ZN(n3013)
         );
  OAI21_X1 U3816 ( .B1(n3053), .B2(n4314), .A(n3013), .ZN(n3014) );
  AOI21_X1 U3817 ( .B1(n3033), .B2(n4197), .A(n3014), .ZN(n3015) );
  OAI21_X1 U3818 ( .B1(n3036), .B2(n4321), .A(n3015), .ZN(n3023) );
  NOR2_X1 U3819 ( .A1(n3016), .A2(n3526), .ZN(n3017) );
  OR2_X1 U3820 ( .A1(n3089), .A2(n3017), .ZN(n3027) );
  OAI22_X1 U3821 ( .A1(n3027), .A2(n4305), .B1(n4543), .B2(n3018), .ZN(n3019)
         );
  AOI21_X1 U3822 ( .B1(n3023), .B2(n4543), .A(n3019), .ZN(n3020) );
  INV_X1 U3823 ( .A(n3020), .ZN(U3524) );
  INV_X1 U3824 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3021) );
  OAI22_X1 U3825 ( .A1(n3027), .A2(n4362), .B1(n4536), .B2(n3021), .ZN(n3022)
         );
  AOI21_X1 U3826 ( .B1(n3023), .B2(n4536), .A(n3022), .ZN(n3024) );
  INV_X1 U3827 ( .A(n3024), .ZN(U3479) );
  NAND2_X1 U3828 ( .A1(n4200), .A2(n3025), .ZN(n3026) );
  NAND2_X1 U3829 ( .A1(n4493), .A2(n3026), .ZN(n4234) );
  INV_X1 U3830 ( .A(n3027), .ZN(n3031) );
  INV_X1 U3831 ( .A(n4180), .ZN(n4101) );
  AOI22_X1 U3832 ( .A1(n4175), .A2(n3955), .B1(n4101), .B2(n3909), .ZN(n3029)
         );
  AOI22_X1 U3833 ( .A1(n4229), .A2(REG2_REG_6__SCAN_IN), .B1(n3910), .B2(n4227), .ZN(n3028) );
  OAI211_X1 U3834 ( .C1(n3053), .C2(n4105), .A(n3029), .B(n3028), .ZN(n3030)
         );
  AOI21_X1 U3835 ( .B1(n3031), .B2(n4497), .A(n3030), .ZN(n3035) );
  NAND2_X1 U3836 ( .A1(n4493), .A2(n4197), .ZN(n3409) );
  INV_X1 U3837 ( .A(n3409), .ZN(n3032) );
  NAND2_X1 U3838 ( .A1(n3033), .A2(n3032), .ZN(n3034) );
  OAI211_X1 U3839 ( .C1(n3036), .C2(n4234), .A(n3035), .B(n3034), .ZN(U3284)
         );
  INV_X1 U3840 ( .A(n3936), .ZN(n3922) );
  INV_X1 U3841 ( .A(n3037), .ZN(n3063) );
  INV_X1 U3842 ( .A(n3038), .ZN(n3041) );
  INV_X1 U3843 ( .A(n3039), .ZN(n3040) );
  AOI22_X1 U3844 ( .A1(n3043), .A2(n3042), .B1(n3041), .B2(n3040), .ZN(n3829)
         );
  OR2_X1 U3845 ( .A1(n3065), .A2(n3684), .ZN(n3045) );
  NAND2_X1 U3846 ( .A1(n3831), .A2(n3529), .ZN(n3044) );
  NAND2_X1 U3847 ( .A1(n3045), .A2(n3044), .ZN(n3048) );
  OAI22_X1 U3848 ( .A1(n3065), .A2(n3657), .B1(n3682), .B2(n3046), .ZN(n3047)
         );
  XNOR2_X1 U3849 ( .A(n3047), .B(n2971), .ZN(n3049) );
  XOR2_X1 U3850 ( .A(n3048), .B(n3049), .Z(n3828) );
  NAND2_X1 U3851 ( .A1(n3048), .A2(n3049), .ZN(n3050) );
  NAND2_X1 U3852 ( .A1(n3827), .A2(n3050), .ZN(n3056) );
  OR2_X1 U3853 ( .A1(n3053), .A2(n3684), .ZN(n3052) );
  NAND2_X1 U3854 ( .A1(n3068), .A2(n3529), .ZN(n3051) );
  NAND2_X1 U3855 ( .A1(n3052), .A2(n3051), .ZN(n3522) );
  OAI22_X1 U3856 ( .A1(n3053), .A2(n3579), .B1(n3682), .B2(n3057), .ZN(n3054)
         );
  XNOR2_X1 U3857 ( .A(n3054), .B(n2971), .ZN(n3523) );
  XOR2_X1 U3858 ( .A(n3522), .B(n3523), .Z(n3055) );
  OAI211_X1 U3859 ( .C1(n3056), .C2(n3055), .A(n3525), .B(n3929), .ZN(n3061)
         );
  INV_X1 U3860 ( .A(n3933), .ZN(n3874) );
  OAI22_X1 U3861 ( .A1(n3874), .A2(n3057), .B1(n3919), .B2(n3065), .ZN(n3058)
         );
  AOI211_X1 U3862 ( .C1(n3931), .C2(n3956), .A(n3059), .B(n3058), .ZN(n3060)
         );
  OAI211_X1 U3863 ( .C1(n3922), .C2(n3063), .A(n3061), .B(n3060), .ZN(U3224)
         );
  INV_X1 U3864 ( .A(n3062), .ZN(n3070) );
  OAI22_X1 U3865 ( .A1(n4493), .A2(n3064), .B1(n3063), .B2(n4490), .ZN(n3067)
         );
  OAI22_X1 U3866 ( .A1(n3065), .A2(n4105), .B1(n4106), .B2(n3527), .ZN(n3066)
         );
  AOI211_X1 U3867 ( .C1(n3068), .C2(n4101), .A(n3067), .B(n3066), .ZN(n3069)
         );
  OAI21_X1 U3868 ( .B1(n3070), .B2(n4231), .A(n3069), .ZN(n3071) );
  AOI21_X1 U3869 ( .B1(n3072), .B2(n4171), .A(n3071), .ZN(n3073) );
  OAI21_X1 U3870 ( .B1(n3074), .B2(n4229), .A(n3073), .ZN(U3285) );
  INV_X1 U3871 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3993) );
  OAI22_X1 U3872 ( .A1(n4493), .A2(n3993), .B1(REG3_REG_3__SCAN_IN), .B2(n4490), .ZN(n3075) );
  AOI21_X1 U3873 ( .B1(n3958), .B2(n4175), .A(n3075), .ZN(n3076) );
  OAI21_X1 U3874 ( .B1(n3077), .B2(n4180), .A(n3076), .ZN(n3078) );
  AOI21_X1 U3875 ( .B1(n4497), .B2(n3079), .A(n3078), .ZN(n3082) );
  NAND2_X1 U3876 ( .A1(n3080), .A2(n4171), .ZN(n3081) );
  OAI211_X1 U3877 ( .C1(n3083), .C2(n4229), .A(n3082), .B(n3081), .ZN(U3287)
         );
  XNOR2_X1 U3878 ( .A(n3084), .B(n3348), .ZN(n3088) );
  NAND2_X1 U3879 ( .A1(n3956), .A2(n4287), .ZN(n3086) );
  NAND2_X1 U3880 ( .A1(n3954), .A2(n4311), .ZN(n3085) );
  OAI211_X1 U3881 ( .C1(n4244), .C2(n3532), .A(n3086), .B(n3085), .ZN(n3087)
         );
  AOI21_X1 U3882 ( .B1(n3088), .B2(n4197), .A(n3087), .ZN(n4532) );
  OAI211_X1 U3883 ( .C1(n3089), .C2(n3532), .A(n4317), .B(n3131), .ZN(n4529)
         );
  INV_X1 U3884 ( .A(n4529), .ZN(n3094) );
  INV_X1 U3885 ( .A(n3487), .ZN(n3093) );
  OAI22_X1 U3886 ( .A1(n4493), .A2(n3091), .B1(n3090), .B2(n4490), .ZN(n3092)
         );
  AOI21_X1 U3887 ( .B1(n3094), .B2(n3093), .A(n3092), .ZN(n3099) );
  INV_X1 U3888 ( .A(n3095), .ZN(n3097) );
  NAND2_X1 U3889 ( .A1(n3096), .A2(n3348), .ZN(n4528) );
  NAND3_X1 U3890 ( .A1(n3097), .A2(n4171), .A3(n4528), .ZN(n3098) );
  OAI211_X1 U3891 ( .C1(n4532), .C2(n4229), .A(n3099), .B(n3098), .ZN(U3283)
         );
  INV_X1 U3892 ( .A(n3100), .ZN(n3326) );
  AND2_X1 U3893 ( .A1(n3326), .A2(n3354), .ZN(n3301) );
  XOR2_X1 U3894 ( .A(n3301), .B(n3101), .Z(n3102) );
  NAND2_X1 U3895 ( .A1(n3102), .A2(n4197), .ZN(n3114) );
  XNOR2_X1 U3896 ( .A(n3103), .B(n3301), .ZN(n3117) );
  NAND2_X1 U3897 ( .A1(n3117), .A2(n4171), .ZN(n3112) );
  NAND2_X1 U3898 ( .A1(n3133), .A2(n3840), .ZN(n3104) );
  AND2_X1 U3899 ( .A1(n3146), .A2(n3104), .ZN(n3119) );
  INV_X1 U3900 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4004) );
  OAI22_X1 U3901 ( .A1(n3105), .A2(n4490), .B1(n4004), .B2(n4493), .ZN(n3109)
         );
  NAND2_X1 U3902 ( .A1(n3952), .A2(n4175), .ZN(n3107) );
  NAND2_X1 U3903 ( .A1(n4174), .A2(n3954), .ZN(n3106) );
  OAI211_X1 U3904 ( .C1(n4180), .C2(n3548), .A(n3107), .B(n3106), .ZN(n3108)
         );
  OR2_X1 U3905 ( .A1(n3109), .A2(n3108), .ZN(n3110) );
  AOI21_X1 U3906 ( .B1(n3119), .B2(n4497), .A(n3110), .ZN(n3111) );
  OAI211_X1 U3907 ( .C1(n4229), .C2(n3114), .A(n3112), .B(n3111), .ZN(U3281)
         );
  AOI22_X1 U3908 ( .A1(n3952), .A2(n4311), .B1(n4310), .B2(n3840), .ZN(n3113)
         );
  OAI211_X1 U3909 ( .C1(n3115), .C2(n4314), .A(n3114), .B(n3113), .ZN(n3116)
         );
  AOI21_X1 U3910 ( .B1(n3117), .B2(n4527), .A(n3116), .ZN(n3121) );
  AOI22_X1 U3911 ( .A1(n3119), .A2(n4332), .B1(REG0_REG_9__SCAN_IN), .B2(n4534), .ZN(n3118) );
  OAI21_X1 U3912 ( .B1(n3121), .B2(n4534), .A(n3118), .ZN(U3485) );
  AOI22_X1 U3913 ( .A1(n3119), .A2(n4252), .B1(REG1_REG_9__SCAN_IN), .B2(n4540), .ZN(n3120) );
  OAI21_X1 U3914 ( .B1(n3121), .B2(n4540), .A(n3120), .ZN(U3527) );
  AND2_X1 U3915 ( .A1(n3353), .A2(n3350), .ZN(n3299) );
  XOR2_X1 U3916 ( .A(n3122), .B(n3299), .Z(n4499) );
  INV_X1 U3917 ( .A(n4499), .ZN(n3129) );
  XNOR2_X1 U3918 ( .A(n3123), .B(n3299), .ZN(n3127) );
  OAI22_X1 U3919 ( .A1(n3533), .A2(n4314), .B1(n3124), .B2(n4244), .ZN(n3125)
         );
  AOI21_X1 U3920 ( .B1(n4311), .B2(n3953), .A(n3125), .ZN(n3126) );
  OAI21_X1 U3921 ( .B1(n3127), .B2(n4222), .A(n3126), .ZN(n3128) );
  AOI21_X1 U3922 ( .B1(n4499), .B2(n3166), .A(n3128), .ZN(n4502) );
  OAI21_X1 U3923 ( .B1(n3130), .B2(n3129), .A(n4502), .ZN(n3139) );
  NAND2_X1 U3924 ( .A1(n3131), .A2(n3762), .ZN(n3132) );
  NAND2_X1 U3925 ( .A1(n3133), .A2(n3132), .ZN(n4495) );
  INV_X1 U3926 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3134) );
  OAI22_X1 U3927 ( .A1(n4495), .A2(n4362), .B1(n4536), .B2(n3134), .ZN(n3135)
         );
  AOI21_X1 U3928 ( .B1(n3139), .B2(n4536), .A(n3135), .ZN(n3136) );
  INV_X1 U3929 ( .A(n3136), .ZN(U3483) );
  INV_X1 U3930 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3137) );
  OAI22_X1 U3931 ( .A1(n4495), .A2(n4305), .B1(n4543), .B2(n3137), .ZN(n3138)
         );
  AOI21_X1 U3932 ( .B1(n3139), .B2(n4543), .A(n3138), .ZN(n3140) );
  INV_X1 U3933 ( .A(n3140), .ZN(U3526) );
  AND2_X1 U3934 ( .A1(n3325), .A2(n3320), .ZN(n3306) );
  XNOR2_X1 U3935 ( .A(n3141), .B(n3306), .ZN(n3161) );
  XOR2_X1 U3936 ( .A(n3306), .B(n3142), .Z(n3151) );
  OAI22_X1 U3937 ( .A1(n3568), .A2(n4291), .B1(n4244), .B2(n3559), .ZN(n3143)
         );
  AOI21_X1 U3938 ( .B1(n4287), .B2(n3953), .A(n3143), .ZN(n3144) );
  OAI21_X1 U3939 ( .B1(n3151), .B2(n4222), .A(n3144), .ZN(n3145) );
  AOI21_X1 U3940 ( .B1(n3161), .B2(n4527), .A(n3145), .ZN(n3150) );
  AND2_X1 U3941 ( .A1(n3146), .A2(n3740), .ZN(n3147) );
  NOR2_X1 U3942 ( .A1(n3169), .A2(n3147), .ZN(n3152) );
  AOI22_X1 U3943 ( .A1(n3152), .A2(n4252), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4540), .ZN(n3148) );
  OAI21_X1 U3944 ( .B1(n3150), .B2(n4540), .A(n3148), .ZN(U3528) );
  AOI22_X1 U3945 ( .A1(n3152), .A2(n4332), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4534), .ZN(n3149) );
  OAI21_X1 U3946 ( .B1(n3150), .B2(n4534), .A(n3149), .ZN(U3487) );
  NOR2_X1 U3947 ( .A1(n3151), .A2(n3409), .ZN(n3160) );
  NAND2_X1 U3948 ( .A1(n3152), .A2(n4497), .ZN(n3158) );
  INV_X1 U3949 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3154) );
  INV_X1 U3950 ( .A(n3741), .ZN(n3153) );
  OAI22_X1 U3951 ( .A1(n4493), .A2(n3154), .B1(n3153), .B2(n4490), .ZN(n3155)
         );
  AOI21_X1 U3952 ( .B1(n4174), .B2(n3953), .A(n3155), .ZN(n3157) );
  AOI22_X1 U3953 ( .A1(n4175), .A2(n3951), .B1(n4101), .B2(n3740), .ZN(n3156)
         );
  NAND3_X1 U3954 ( .A1(n3158), .A2(n3157), .A3(n3156), .ZN(n3159) );
  AOI211_X1 U3955 ( .C1(n3161), .C2(n4171), .A(n3160), .B(n3159), .ZN(n3162)
         );
  INV_X1 U3956 ( .A(n3162), .ZN(U3280) );
  XNOR2_X1 U3957 ( .A(n3179), .B(n3275), .ZN(n3168) );
  OAI21_X1 U3958 ( .B1(n3164), .B2(n3275), .A(n3163), .ZN(n3194) );
  OAI22_X1 U3959 ( .A1(n3574), .A2(n4291), .B1(n4244), .B2(n3567), .ZN(n3165)
         );
  AOI21_X1 U3960 ( .B1(n3194), .B2(n3166), .A(n3165), .ZN(n3167) );
  OAI21_X1 U3961 ( .B1(n4222), .B2(n3168), .A(n3167), .ZN(n3192) );
  INV_X1 U3962 ( .A(n3192), .ZN(n3174) );
  OAI21_X1 U3963 ( .B1(n3169), .B2(n3567), .A(n3182), .ZN(n3200) );
  AOI22_X1 U3964 ( .A1(n4229), .A2(REG2_REG_11__SCAN_IN), .B1(n3886), .B2(
        n4227), .ZN(n3171) );
  NAND2_X1 U3965 ( .A1(n3952), .A2(n4174), .ZN(n3170) );
  OAI211_X1 U3966 ( .C1(n3200), .C2(n4231), .A(n3171), .B(n3170), .ZN(n3172)
         );
  AOI21_X1 U3967 ( .B1(n3194), .B2(n4498), .A(n3172), .ZN(n3173) );
  OAI21_X1 U3968 ( .B1(n3174), .B2(n4229), .A(n3173), .ZN(U3279) );
  AND2_X1 U3969 ( .A1(n3214), .A2(n3212), .ZN(n3307) );
  XOR2_X1 U3970 ( .A(n3307), .B(n3175), .Z(n3205) );
  INV_X1 U3971 ( .A(n3176), .ZN(n3177) );
  AOI21_X1 U3972 ( .B1(n3179), .B2(n3178), .A(n3177), .ZN(n3215) );
  INV_X1 U3973 ( .A(n3307), .ZN(n3180) );
  XNOR2_X1 U3974 ( .A(n3215), .B(n3180), .ZN(n3181) );
  NAND2_X1 U3975 ( .A1(n3181), .A2(n4197), .ZN(n3203) );
  NOR2_X1 U3976 ( .A1(n3203), .A2(n4229), .ZN(n3190) );
  NAND2_X1 U3977 ( .A1(n3182), .A2(n2450), .ZN(n3183) );
  NAND2_X1 U3978 ( .A1(n3221), .A2(n3183), .ZN(n3211) );
  NAND2_X1 U3979 ( .A1(n4229), .A2(REG2_REG_12__SCAN_IN), .ZN(n3185) );
  NAND2_X1 U3980 ( .A1(n4227), .A2(n3783), .ZN(n3184) );
  OAI211_X1 U3981 ( .C1(n4180), .C2(n3572), .A(n3185), .B(n3184), .ZN(n3186)
         );
  INV_X1 U3982 ( .A(n3186), .ZN(n3188) );
  AOI22_X1 U3983 ( .A1(n4174), .A2(n3951), .B1(n3949), .B2(n4175), .ZN(n3187)
         );
  OAI211_X1 U3984 ( .C1(n3211), .C2(n4231), .A(n3188), .B(n3187), .ZN(n3189)
         );
  AOI211_X1 U3985 ( .C1(n3205), .C2(n4171), .A(n3190), .B(n3189), .ZN(n3191)
         );
  INV_X1 U3986 ( .A(n3191), .ZN(U3278) );
  INV_X1 U3987 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3195) );
  NOR2_X1 U3988 ( .A1(n3561), .A2(n4314), .ZN(n3193) );
  AOI211_X1 U3989 ( .C1(n4524), .C2(n3194), .A(n3193), .B(n3192), .ZN(n3197)
         );
  MUX2_X1 U3990 ( .A(n3195), .B(n3197), .S(n4536), .Z(n3196) );
  OAI21_X1 U3991 ( .B1(n3200), .B2(n4362), .A(n3196), .ZN(U3489) );
  INV_X1 U3992 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3198) );
  MUX2_X1 U3993 ( .A(n3198), .B(n3197), .S(n4543), .Z(n3199) );
  OAI21_X1 U3994 ( .B1(n4305), .B2(n3200), .A(n3199), .ZN(U3529) );
  INV_X1 U3995 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3206) );
  OAI22_X1 U3996 ( .A1(n3582), .A2(n4291), .B1(n4244), .B2(n3572), .ZN(n3201)
         );
  INV_X1 U3997 ( .A(n3201), .ZN(n3202) );
  OAI211_X1 U3998 ( .C1(n3568), .C2(n4314), .A(n3203), .B(n3202), .ZN(n3204)
         );
  AOI21_X1 U3999 ( .B1(n3205), .B2(n4527), .A(n3204), .ZN(n3208) );
  MUX2_X1 U4000 ( .A(n3206), .B(n3208), .S(n4543), .Z(n3207) );
  OAI21_X1 U4001 ( .B1(n4305), .B2(n3211), .A(n3207), .ZN(U3530) );
  INV_X1 U4002 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3209) );
  MUX2_X1 U4003 ( .A(n3209), .B(n3208), .S(n4536), .Z(n3210) );
  OAI21_X1 U4004 ( .B1(n3211), .B2(n4362), .A(n3210), .ZN(U3491) );
  XNOR2_X1 U4005 ( .A(n3582), .B(n3581), .ZN(n3293) );
  INV_X1 U4006 ( .A(n3212), .ZN(n3213) );
  AOI21_X1 U4007 ( .B1(n3215), .B2(n3214), .A(n3213), .ZN(n3216) );
  XOR2_X1 U4008 ( .A(n3293), .B(n3216), .Z(n3219) );
  OAI22_X1 U4009 ( .A1(n3585), .A2(n4291), .B1(n4244), .B2(n3581), .ZN(n3217)
         );
  AOI21_X1 U4010 ( .B1(n4287), .B2(n3950), .A(n3217), .ZN(n3218) );
  OAI21_X1 U4011 ( .B1(n3219), .B2(n4222), .A(n3218), .ZN(n3410) );
  INV_X1 U4012 ( .A(n3410), .ZN(n3227) );
  XOR2_X1 U4013 ( .A(n3293), .B(n3220), .Z(n3411) );
  INV_X1 U4014 ( .A(n3221), .ZN(n3223) );
  INV_X1 U4015 ( .A(n3402), .ZN(n3222) );
  OAI21_X1 U4016 ( .B1(n3223), .B2(n3581), .A(n3222), .ZN(n3417) );
  AOI22_X1 U4017 ( .A1(n4229), .A2(REG2_REG_13__SCAN_IN), .B1(n3864), .B2(
        n4227), .ZN(n3224) );
  OAI21_X1 U4018 ( .B1(n3417), .B2(n4231), .A(n3224), .ZN(n3225) );
  AOI21_X1 U4019 ( .B1(n3411), .B2(n4171), .A(n3225), .ZN(n3226) );
  OAI21_X1 U4020 ( .B1(n4229), .B2(n3227), .A(n3226), .ZN(U3277) );
  INV_X1 U4021 ( .A(n3941), .ZN(n3228) );
  AND2_X1 U4022 ( .A1(n2046), .A2(DATAI_30_), .ZN(n4242) );
  NOR2_X1 U4023 ( .A1(n3228), .A2(n4242), .ZN(n3382) );
  INV_X1 U4024 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3233) );
  NAND2_X1 U4025 ( .A1(n3229), .A2(REG2_REG_31__SCAN_IN), .ZN(n3232) );
  NAND2_X1 U4026 ( .A1(n3230), .A2(REG0_REG_31__SCAN_IN), .ZN(n3231) );
  OAI211_X1 U4027 ( .C1(n3234), .C2(n3233), .A(n3232), .B(n3231), .ZN(n4057)
         );
  INV_X1 U4028 ( .A(n4057), .ZN(n3235) );
  NOR2_X1 U4029 ( .A1(n3382), .A2(n3235), .ZN(n3272) );
  NAND2_X1 U4030 ( .A1(n2046), .A2(DATAI_31_), .ZN(n4058) );
  NAND2_X1 U4031 ( .A1(n3236), .A2(n3242), .ZN(n3364) );
  NAND2_X1 U4032 ( .A1(n3327), .A2(n3328), .ZN(n3241) );
  INV_X1 U4033 ( .A(n3329), .ZN(n3240) );
  NAND2_X1 U4034 ( .A1(n2053), .A2(n3237), .ZN(n3239) );
  OR2_X1 U4035 ( .A1(n3239), .A2(n3238), .ZN(n3331) );
  AOI211_X1 U4036 ( .C1(n3242), .C2(n3241), .A(n3240), .B(n3331), .ZN(n3363)
         );
  OAI21_X1 U4037 ( .B1(n3397), .B2(n3364), .A(n3363), .ZN(n3246) );
  INV_X1 U4038 ( .A(n3331), .ZN(n3245) );
  INV_X1 U4039 ( .A(n3243), .ZN(n3244) );
  NAND2_X1 U4040 ( .A1(n3245), .A2(n3244), .ZN(n3368) );
  NAND4_X1 U4041 ( .A1(n3246), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3249)
         );
  INV_X1 U4042 ( .A(n3274), .ZN(n3247) );
  NAND2_X1 U40430 ( .A1(n3247), .A2(n3284), .ZN(n3373) );
  AOI21_X1 U4044 ( .B1(n3249), .B2(n3248), .A(n3373), .ZN(n3250) );
  NOR2_X1 U4045 ( .A1(n3250), .A2(n4075), .ZN(n3256) );
  NAND2_X1 U4046 ( .A1(n3252), .A2(n3251), .ZN(n3261) );
  OR2_X1 U4047 ( .A1(n3942), .A2(n4063), .ZN(n3255) );
  INV_X1 U4048 ( .A(n4242), .ZN(n3266) );
  NAND2_X1 U4049 ( .A1(n4057), .A2(n4058), .ZN(n3380) );
  OAI21_X1 U4050 ( .B1(n3266), .B2(n3941), .A(n3380), .ZN(n3253) );
  INV_X1 U4051 ( .A(n3253), .ZN(n3254) );
  NAND2_X1 U4052 ( .A1(n3255), .A2(n3254), .ZN(n3262) );
  NOR4_X1 U4053 ( .A1(n3256), .A2(n3372), .A3(n3261), .A4(n3262), .ZN(n3268)
         );
  INV_X1 U4054 ( .A(n4063), .ZN(n3258) );
  OAI21_X1 U4055 ( .B1(n3259), .B2(n3258), .A(n3257), .ZN(n3377) );
  NOR2_X1 U4056 ( .A1(n3377), .A2(n3260), .ZN(n3265) );
  INV_X1 U4057 ( .A(n3261), .ZN(n3264) );
  INV_X1 U4058 ( .A(n3262), .ZN(n3263) );
  OAI21_X1 U4059 ( .B1(n3264), .B2(n3377), .A(n3263), .ZN(n3384) );
  AOI21_X1 U4060 ( .B1(n3508), .B2(n3265), .A(n3384), .ZN(n3267) );
  OAI22_X1 U4061 ( .A1(n3268), .A2(n3267), .B1(n3266), .B2(n4057), .ZN(n3271)
         );
  INV_X1 U4062 ( .A(n3269), .ZN(n3270) );
  OAI211_X1 U4063 ( .C1(n3272), .C2(n4058), .A(n3271), .B(n3270), .ZN(n3389)
         );
  INV_X1 U4064 ( .A(n4093), .ZN(n3273) );
  OR2_X1 U4065 ( .A1(n3274), .A2(n3273), .ZN(n4116) );
  INV_X1 U4066 ( .A(n3275), .ZN(n3277) );
  INV_X1 U4067 ( .A(n3432), .ZN(n3276) );
  NAND4_X1 U4068 ( .A1(n3277), .A2(n3276), .A3(n3424), .A4(n3348), .ZN(n3281)
         );
  INV_X1 U4069 ( .A(n3278), .ZN(n4129) );
  NOR2_X1 U4070 ( .A1(n4129), .A2(n4128), .ZN(n4170) );
  NAND2_X1 U4071 ( .A1(n4170), .A2(n3279), .ZN(n3280) );
  NOR3_X1 U4072 ( .A1(n4116), .A2(n3281), .A3(n3280), .ZN(n3315) );
  NAND2_X1 U4073 ( .A1(n4074), .A2(n3282), .ZN(n4097) );
  INV_X1 U4074 ( .A(n4097), .ZN(n3314) );
  NAND2_X1 U4075 ( .A1(n3284), .A2(n3283), .ZN(n4132) );
  NAND2_X1 U4076 ( .A1(n3285), .A2(n3479), .ZN(n3286) );
  NOR2_X1 U4077 ( .A1(n4132), .A2(n3286), .ZN(n3312) );
  NAND2_X1 U4078 ( .A1(n3288), .A2(n3287), .ZN(n4217) );
  INV_X1 U4079 ( .A(n4217), .ZN(n3294) );
  XNOR2_X1 U4080 ( .A(n3941), .B(n4242), .ZN(n3292) );
  NOR2_X1 U4081 ( .A1(n4057), .A2(n4058), .ZN(n3381) );
  INV_X1 U4082 ( .A(n3381), .ZN(n3290) );
  AND3_X1 U4083 ( .A1(n3290), .A2(n3289), .A3(n3380), .ZN(n3291) );
  AND4_X1 U4084 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3311)
         );
  NAND4_X1 U4085 ( .A1(n2206), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3303)
         );
  NAND4_X1 U4086 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3302)
         );
  NOR2_X1 U4087 ( .A1(n3303), .A2(n3302), .ZN(n3310) );
  NAND2_X1 U4088 ( .A1(n2053), .A2(n3477), .ZN(n3466) );
  INV_X1 U4089 ( .A(n3466), .ZN(n3308) );
  NAND2_X1 U4090 ( .A1(n3305), .A2(n3304), .ZN(n4190) );
  AND4_X1 U4091 ( .A1(n3308), .A2(n3307), .A3(n3306), .A4(n4190), .ZN(n3309)
         );
  AND4_X1 U4092 ( .A1(n3312), .A2(n3311), .A3(n3310), .A4(n3309), .ZN(n3313)
         );
  NAND4_X1 U4093 ( .A1(n3315), .A2(n4157), .A3(n3314), .A4(n3313), .ZN(n3316)
         );
  NOR2_X1 U4094 ( .A1(n3317), .A2(n3316), .ZN(n3319) );
  XNOR2_X1 U4095 ( .A(n4262), .B(n4085), .ZN(n4077) );
  NAND4_X1 U4096 ( .A1(n3319), .A2(n2226), .A3(n3508), .A4(n4077), .ZN(n3387)
         );
  INV_X1 U4097 ( .A(n3320), .ZN(n3360) );
  INV_X1 U4098 ( .A(n3351), .ZN(n3322) );
  NOR2_X1 U4099 ( .A1(n3322), .A2(n3321), .ZN(n3323) );
  NAND4_X1 U4100 ( .A1(n3323), .A2(n3326), .A3(n3350), .A4(n3343), .ZN(n3324)
         );
  NAND2_X1 U4101 ( .A1(n3325), .A2(n3324), .ZN(n3357) );
  NAND4_X1 U4102 ( .A1(n3329), .A2(n3328), .A3(n3327), .A4(n3326), .ZN(n3330)
         );
  NOR2_X1 U4103 ( .A1(n3331), .A2(n3330), .ZN(n3356) );
  OAI211_X1 U4104 ( .C1(n4373), .C2(n2171), .A(n3333), .B(n3332), .ZN(n3334)
         );
  NAND3_X1 U4105 ( .A1(n3335), .A2(n2632), .A3(n3334), .ZN(n3336) );
  NAND3_X1 U4106 ( .A1(n3338), .A2(n3337), .A3(n3336), .ZN(n3339) );
  NAND3_X1 U4107 ( .A1(n3341), .A2(n3340), .A3(n3339), .ZN(n3342) );
  NAND4_X1 U4108 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3346)
         );
  NAND3_X1 U4109 ( .A1(n3348), .A2(n3347), .A3(n3346), .ZN(n3349) );
  NAND3_X1 U4110 ( .A1(n3351), .A2(n3350), .A3(n3349), .ZN(n3352) );
  NAND3_X1 U4111 ( .A1(n3354), .A2(n3353), .A3(n3352), .ZN(n3355) );
  AOI22_X1 U4112 ( .A1(n3363), .A2(n3357), .B1(n3356), .B2(n3355), .ZN(n3359)
         );
  OR4_X1 U4113 ( .A1(n3361), .A2(n3360), .A3(n3359), .A4(n3358), .ZN(n3367) );
  INV_X1 U4114 ( .A(n3362), .ZN(n3365) );
  OAI21_X1 U4115 ( .B1(n3365), .B2(n3364), .A(n3363), .ZN(n3366) );
  AND4_X1 U4116 ( .A1(n3369), .A2(n3368), .A3(n3367), .A4(n3366), .ZN(n3371)
         );
  OAI21_X1 U4117 ( .B1(n4128), .B2(n3371), .A(n3370), .ZN(n3374) );
  AOI211_X1 U4118 ( .C1(n3375), .C2(n3374), .A(n3373), .B(n3372), .ZN(n3379)
         );
  INV_X1 U4119 ( .A(n3943), .ZN(n4083) );
  OAI21_X1 U4120 ( .B1(n4083), .B2(n3708), .A(n3376), .ZN(n3378) );
  NOR3_X1 U4121 ( .A1(n3379), .A2(n3378), .A3(n3377), .ZN(n3385) );
  OAI21_X1 U4122 ( .B1(n3382), .B2(n3381), .A(n3380), .ZN(n3383) );
  OAI21_X1 U4123 ( .B1(n3385), .B2(n3384), .A(n3383), .ZN(n3386) );
  MUX2_X1 U4124 ( .A(n3387), .B(n3386), .S(n2618), .Z(n3388) );
  NAND2_X1 U4125 ( .A1(n3389), .A2(n3388), .ZN(n3390) );
  XNOR2_X1 U4126 ( .A(n3390), .B(n4374), .ZN(n3396) );
  NAND2_X1 U4127 ( .A1(n3392), .A2(n3391), .ZN(n3393) );
  OAI211_X1 U4128 ( .C1(n4372), .C2(n3395), .A(n3393), .B(B_REG_SCAN_IN), .ZN(
        n3394) );
  OAI21_X1 U4129 ( .B1(n3396), .B2(n3395), .A(n3394), .ZN(U3239) );
  XNOR2_X1 U4130 ( .A(n3397), .B(n3399), .ZN(n3444) );
  OAI21_X1 U4131 ( .B1(n3400), .B2(n3399), .A(n3398), .ZN(n3446) );
  NAND2_X1 U4132 ( .A1(n3446), .A2(n4171), .ZN(n3408) );
  INV_X1 U4133 ( .A(n3435), .ZN(n3401) );
  OAI21_X1 U4134 ( .B1(n3402), .B2(n3583), .A(n3401), .ZN(n3452) );
  INV_X1 U4135 ( .A(n3452), .ZN(n3406) );
  AOI22_X1 U4136 ( .A1(n4101), .A2(n3719), .B1(n4175), .B2(n3947), .ZN(n3404)
         );
  AOI22_X1 U4137 ( .A1(n4229), .A2(REG2_REG_14__SCAN_IN), .B1(n3723), .B2(
        n4227), .ZN(n3403) );
  OAI211_X1 U4138 ( .C1(n3582), .C2(n4105), .A(n3404), .B(n3403), .ZN(n3405)
         );
  AOI21_X1 U4139 ( .B1(n3406), .B2(n4497), .A(n3405), .ZN(n3407) );
  OAI211_X1 U4140 ( .C1(n3444), .C2(n3409), .A(n3408), .B(n3407), .ZN(U3276)
         );
  INV_X1 U4141 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3412) );
  AOI21_X1 U4142 ( .B1(n3411), .B2(n4527), .A(n3410), .ZN(n3414) );
  MUX2_X1 U4143 ( .A(n3412), .B(n3414), .S(n4543), .Z(n3413) );
  OAI21_X1 U4144 ( .B1(n4305), .B2(n3417), .A(n3413), .ZN(U3531) );
  INV_X1 U4145 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3415) );
  MUX2_X1 U4146 ( .A(n3415), .B(n3414), .S(n4536), .Z(n3416) );
  OAI21_X1 U4147 ( .B1(n3417), .B2(n4362), .A(n3416), .ZN(U3493) );
  OAI21_X1 U4148 ( .B1(n3418), .B2(n3420), .A(n3419), .ZN(n4322) );
  AOI21_X1 U4149 ( .B1(n4309), .B2(n3434), .A(n2047), .ZN(n4318) );
  AOI22_X1 U4150 ( .A1(n4174), .A2(n3947), .B1(n4175), .B2(n4312), .ZN(n3422)
         );
  AOI22_X1 U4151 ( .A1(n4229), .A2(REG2_REG_16__SCAN_IN), .B1(n3803), .B2(
        n4227), .ZN(n3421) );
  OAI211_X1 U4152 ( .C1(n3601), .C2(n4180), .A(n3422), .B(n3421), .ZN(n3427)
         );
  OAI211_X1 U4153 ( .C1(n3425), .C2(n3424), .A(n3423), .B(n4197), .ZN(n4319)
         );
  NOR2_X1 U4154 ( .A1(n4319), .A2(n4229), .ZN(n3426) );
  AOI211_X1 U4155 ( .C1(n4318), .C2(n4497), .A(n3427), .B(n3426), .ZN(n3428)
         );
  OAI21_X1 U4156 ( .B1(n4322), .B2(n4234), .A(n3428), .ZN(U3274) );
  AOI21_X1 U4157 ( .B1(n3429), .B2(n3432), .A(n4222), .ZN(n3431) );
  NAND2_X1 U4158 ( .A1(n3431), .A2(n3430), .ZN(n3454) );
  XNOR2_X1 U4159 ( .A(n3433), .B(n3432), .ZN(n3456) );
  NAND2_X1 U4160 ( .A1(n3456), .A2(n4171), .ZN(n3441) );
  OAI21_X1 U4161 ( .B1(n3435), .B2(n3593), .A(n3434), .ZN(n3462) );
  INV_X1 U4162 ( .A(n3462), .ZN(n3439) );
  AOI22_X1 U4163 ( .A1(n4175), .A2(n3946), .B1(n3948), .B2(n4174), .ZN(n3437)
         );
  AOI22_X1 U4164 ( .A1(n4229), .A2(REG2_REG_15__SCAN_IN), .B1(n3935), .B2(
        n4227), .ZN(n3436) );
  OAI211_X1 U4165 ( .C1(n3593), .C2(n4180), .A(n3437), .B(n3436), .ZN(n3438)
         );
  AOI21_X1 U4166 ( .B1(n3439), .B2(n4497), .A(n3438), .ZN(n3440) );
  OAI211_X1 U4167 ( .C1(n4229), .C2(n3454), .A(n3441), .B(n3440), .ZN(U3275)
         );
  INV_X1 U4168 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3447) );
  OAI22_X1 U4169 ( .A1(n4315), .A2(n4291), .B1(n4244), .B2(n3583), .ZN(n3442)
         );
  AOI21_X1 U4170 ( .B1(n4287), .B2(n3949), .A(n3442), .ZN(n3443) );
  OAI21_X1 U4171 ( .B1(n3444), .B2(n4222), .A(n3443), .ZN(n3445) );
  AOI21_X1 U4172 ( .B1(n3446), .B2(n4527), .A(n3445), .ZN(n3449) );
  MUX2_X1 U4173 ( .A(n3447), .B(n3449), .S(n4543), .Z(n3448) );
  OAI21_X1 U4174 ( .B1(n4305), .B2(n3452), .A(n3448), .ZN(U3532) );
  INV_X1 U4175 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3450) );
  MUX2_X1 U4176 ( .A(n3450), .B(n3449), .S(n4536), .Z(n3451) );
  OAI21_X1 U4177 ( .B1(n3452), .B2(n4362), .A(n3451), .ZN(U3495) );
  INV_X1 U4178 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3457) );
  AOI22_X1 U4179 ( .A1(n3946), .A2(n4311), .B1(n3932), .B2(n4310), .ZN(n3453)
         );
  OAI211_X1 U4180 ( .C1(n3585), .C2(n4314), .A(n3454), .B(n3453), .ZN(n3455)
         );
  AOI21_X1 U4181 ( .B1(n3456), .B2(n4527), .A(n3455), .ZN(n3459) );
  MUX2_X1 U4182 ( .A(n3457), .B(n3459), .S(n4543), .Z(n3458) );
  OAI21_X1 U4183 ( .B1(n4305), .B2(n3462), .A(n3458), .ZN(U3533) );
  INV_X1 U4184 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3460) );
  MUX2_X1 U4185 ( .A(n3460), .B(n3459), .S(n4536), .Z(n3461) );
  OAI21_X1 U4186 ( .B1(n3462), .B2(n4362), .A(n3461), .ZN(U3497) );
  XNOR2_X1 U4187 ( .A(n3463), .B(n3466), .ZN(n3464) );
  NAND2_X1 U4188 ( .A1(n3464), .A2(n4197), .ZN(n3492) );
  XOR2_X1 U4189 ( .A(n3466), .B(n3465), .Z(n3494) );
  NAND2_X1 U4190 ( .A1(n3494), .A2(n4171), .ZN(n3473) );
  OAI21_X1 U4191 ( .B1(n2047), .B2(n3469), .A(n2090), .ZN(n3500) );
  INV_X1 U4192 ( .A(n3500), .ZN(n3471) );
  AOI22_X1 U4193 ( .A1(n4174), .A2(n3946), .B1(n4220), .B2(n4175), .ZN(n3468)
         );
  AOI22_X1 U4194 ( .A1(n4229), .A2(REG2_REG_17__SCAN_IN), .B1(n3814), .B2(
        n4227), .ZN(n3467) );
  OAI211_X1 U4195 ( .C1(n3469), .C2(n4180), .A(n3468), .B(n3467), .ZN(n3470)
         );
  AOI21_X1 U4196 ( .B1(n3471), .B2(n4497), .A(n3470), .ZN(n3472) );
  OAI211_X1 U4197 ( .C1(n4229), .C2(n3492), .A(n3473), .B(n3472), .ZN(U3273)
         );
  INV_X1 U4198 ( .A(n3474), .ZN(n3475) );
  AOI21_X1 U4199 ( .B1(n3479), .B2(n3476), .A(n3475), .ZN(n4308) );
  NAND2_X1 U4200 ( .A1(n3478), .A2(n3477), .ZN(n4215) );
  XNOR2_X1 U4201 ( .A(n4215), .B(n3479), .ZN(n3483) );
  NAND2_X1 U4202 ( .A1(n3945), .A2(n4311), .ZN(n3481) );
  NAND2_X1 U4203 ( .A1(n4312), .A2(n4287), .ZN(n3480) );
  OAI211_X1 U4204 ( .C1(n4244), .C2(n3617), .A(n3481), .B(n3480), .ZN(n3482)
         );
  AOI21_X1 U4205 ( .B1(n3483), .B2(n4197), .A(n3482), .ZN(n4307) );
  INV_X1 U4206 ( .A(n4307), .ZN(n3489) );
  INV_X1 U4207 ( .A(n4226), .ZN(n3484) );
  OAI211_X1 U4208 ( .C1(n3485), .C2(n3617), .A(n3484), .B(n4317), .ZN(n4306)
         );
  AOI22_X1 U4209 ( .A1(n4229), .A2(REG2_REG_18__SCAN_IN), .B1(n3898), .B2(
        n4227), .ZN(n3486) );
  OAI21_X1 U4210 ( .B1(n4306), .B2(n3487), .A(n3486), .ZN(n3488) );
  AOI21_X1 U4211 ( .B1(n3489), .B2(n4493), .A(n3488), .ZN(n3490) );
  OAI21_X1 U4212 ( .B1(n4308), .B2(n4234), .A(n3490), .ZN(U3272) );
  INV_X1 U4213 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4214 ( .A1(n4220), .A2(n4311), .B1(n4310), .B2(n3813), .ZN(n3491)
         );
  OAI211_X1 U4215 ( .C1(n3602), .C2(n4314), .A(n3492), .B(n3491), .ZN(n3493)
         );
  AOI21_X1 U4216 ( .B1(n3494), .B2(n4527), .A(n3493), .ZN(n3497) );
  MUX2_X1 U4217 ( .A(n3495), .B(n3497), .S(n4536), .Z(n3496) );
  OAI21_X1 U4218 ( .B1(n3500), .B2(n4362), .A(n3496), .ZN(U3501) );
  INV_X1 U4219 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3498) );
  MUX2_X1 U4220 ( .A(n3498), .B(n3497), .S(n4543), .Z(n3499) );
  OAI21_X1 U4221 ( .B1(n4305), .B2(n3500), .A(n3499), .ZN(U3535) );
  XNOR2_X1 U4222 ( .A(n3501), .B(n3508), .ZN(n4250) );
  AOI21_X1 U4223 ( .B1(n3708), .B2(n4084), .A(n3502), .ZN(n4333) );
  AOI22_X1 U4224 ( .A1(n4101), .A2(n3708), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4229), .ZN(n3503) );
  OAI21_X1 U4225 ( .B1(n4262), .B2(n4105), .A(n3503), .ZN(n3504) );
  AOI21_X1 U4226 ( .B1(n3711), .B2(n4227), .A(n3504), .ZN(n3505) );
  OAI21_X1 U4227 ( .B1(n3685), .B2(n4106), .A(n3505), .ZN(n3511) );
  OAI21_X1 U4228 ( .B1(n3508), .B2(n3507), .A(n3506), .ZN(n3509) );
  NAND2_X1 U4229 ( .A1(n3509), .A2(n4197), .ZN(n4248) );
  NOR2_X1 U4230 ( .A1(n4248), .A2(n4229), .ZN(n3510) );
  AOI211_X1 U4231 ( .C1(n4497), .C2(n4333), .A(n3511), .B(n3510), .ZN(n3512)
         );
  OAI21_X1 U4232 ( .B1(n4250), .B2(n4234), .A(n3512), .ZN(U3263) );
  INV_X1 U4233 ( .A(n3513), .ZN(n3519) );
  AOI22_X1 U4234 ( .A1(n4101), .A2(n3690), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4229), .ZN(n3515) );
  AOI22_X1 U4235 ( .A1(n3942), .A2(n4175), .B1(n3691), .B2(n4227), .ZN(n3514)
         );
  OAI211_X1 U4236 ( .C1(n4083), .C2(n4105), .A(n3515), .B(n3514), .ZN(n3518)
         );
  NOR2_X1 U4237 ( .A1(n3516), .A2(n4229), .ZN(n3517) );
  AOI211_X1 U4238 ( .C1(n4497), .C2(n3519), .A(n3518), .B(n3517), .ZN(n3520)
         );
  OAI21_X1 U4239 ( .B1(n3521), .B2(n4234), .A(n3520), .ZN(U3262) );
  NAND2_X1 U4240 ( .A1(n3522), .A2(n3523), .ZN(n3524) );
  OAI22_X1 U4241 ( .A1(n3527), .A2(n3684), .B1(n3657), .B2(n3526), .ZN(n3903)
         );
  OAI22_X1 U4242 ( .A1(n3527), .A2(n3579), .B1(n3682), .B2(n3526), .ZN(n3528)
         );
  XNOR2_X1 U4243 ( .A(n3528), .B(n2971), .ZN(n3904) );
  OR2_X1 U4244 ( .A1(n3533), .A2(n3684), .ZN(n3531) );
  NAND2_X1 U4245 ( .A1(n3701), .A2(n3529), .ZN(n3530) );
  NAND2_X1 U4246 ( .A1(n3531), .A2(n3530), .ZN(n3536) );
  OAI22_X1 U4247 ( .A1(n3533), .A2(n3657), .B1(n3682), .B2(n3532), .ZN(n3534)
         );
  XNOR2_X1 U4248 ( .A(n3534), .B(n2971), .ZN(n3535) );
  XOR2_X1 U4249 ( .A(n3536), .B(n3535), .Z(n3697) );
  NAND2_X1 U4250 ( .A1(n3954), .A2(n3529), .ZN(n3538) );
  NAND2_X1 U4251 ( .A1(n3762), .A2(n2968), .ZN(n3537) );
  NAND2_X1 U4252 ( .A1(n3538), .A2(n3537), .ZN(n3539) );
  XNOR2_X1 U4253 ( .A(n3539), .B(n2971), .ZN(n3543) );
  NAND2_X1 U4254 ( .A1(n3954), .A2(n3540), .ZN(n3542) );
  NAND2_X1 U4255 ( .A1(n3762), .A2(n3529), .ZN(n3541) );
  NAND2_X1 U4256 ( .A1(n3542), .A2(n3541), .ZN(n3544) );
  NAND2_X1 U4257 ( .A1(n3543), .A2(n3544), .ZN(n3756) );
  NAND2_X1 U4258 ( .A1(n3757), .A2(n3756), .ZN(n3547) );
  INV_X1 U4259 ( .A(n3543), .ZN(n3546) );
  INV_X1 U4260 ( .A(n3544), .ZN(n3545) );
  NAND2_X1 U4261 ( .A1(n3546), .A2(n3545), .ZN(n3755) );
  NAND2_X1 U4262 ( .A1(n3547), .A2(n3755), .ZN(n3837) );
  OAI22_X1 U4263 ( .A1(n3549), .A2(n3684), .B1(n3657), .B2(n3548), .ZN(n3554)
         );
  NAND2_X1 U4264 ( .A1(n3953), .A2(n3529), .ZN(n3551) );
  NAND2_X1 U4265 ( .A1(n3840), .A2(n2968), .ZN(n3550) );
  NAND2_X1 U4266 ( .A1(n3551), .A2(n3550), .ZN(n3552) );
  XNOR2_X1 U4267 ( .A(n3552), .B(n2971), .ZN(n3553) );
  XOR2_X1 U4268 ( .A(n3554), .B(n3553), .Z(n3838) );
  NAND2_X1 U4269 ( .A1(n3837), .A2(n3838), .ZN(n3558) );
  INV_X1 U4270 ( .A(n3553), .ZN(n3556) );
  INV_X1 U4271 ( .A(n3554), .ZN(n3555) );
  NAND2_X1 U4272 ( .A1(n3556), .A2(n3555), .ZN(n3557) );
  OAI22_X1 U4273 ( .A1(n3561), .A2(n3579), .B1(n3682), .B2(n3559), .ZN(n3560)
         );
  XNOR2_X1 U4274 ( .A(n3560), .B(n2971), .ZN(n3565) );
  OR2_X1 U4275 ( .A1(n3561), .A2(n3684), .ZN(n3563) );
  NAND2_X1 U4276 ( .A1(n3740), .A2(n3529), .ZN(n3562) );
  NAND2_X1 U4277 ( .A1(n3563), .A2(n3562), .ZN(n3564) );
  XNOR2_X1 U4278 ( .A(n3565), .B(n3564), .ZN(n3735) );
  NAND2_X1 U4279 ( .A1(n3565), .A2(n3564), .ZN(n3566) );
  OAI22_X1 U4280 ( .A1(n3568), .A2(n3684), .B1(n3657), .B2(n3567), .ZN(n3880)
         );
  OAI22_X1 U4281 ( .A1(n3568), .A2(n3579), .B1(n3682), .B2(n3567), .ZN(n3569)
         );
  XNOR2_X1 U4282 ( .A(n3569), .B(n2971), .ZN(n3881) );
  OAI22_X1 U4283 ( .A1(n3574), .A2(n3579), .B1(n3682), .B2(n3572), .ZN(n3573)
         );
  XNOR2_X1 U4284 ( .A(n3573), .B(n3667), .ZN(n3578) );
  OR2_X1 U4285 ( .A1(n3574), .A2(n3684), .ZN(n3576) );
  NAND2_X1 U4286 ( .A1(n2450), .A2(n3529), .ZN(n3575) );
  NAND2_X1 U4287 ( .A1(n3578), .A2(n3577), .ZN(n3778) );
  OAI22_X1 U4288 ( .A1(n3582), .A2(n3579), .B1(n3682), .B2(n3581), .ZN(n3580)
         );
  XOR2_X1 U4289 ( .A(n2971), .B(n3580), .Z(n3859) );
  OAI22_X1 U4290 ( .A1(n3582), .A2(n3684), .B1(n3657), .B2(n3581), .ZN(n3858)
         );
  OAI22_X1 U4291 ( .A1(n3585), .A2(n3579), .B1(n3682), .B2(n3583), .ZN(n3584)
         );
  XNOR2_X1 U4292 ( .A(n3584), .B(n2971), .ZN(n3588) );
  OR2_X1 U4293 ( .A1(n3585), .A2(n3684), .ZN(n3587) );
  NAND2_X1 U4294 ( .A1(n3719), .A2(n3529), .ZN(n3586) );
  NAND2_X1 U4295 ( .A1(n3587), .A2(n3586), .ZN(n3589) );
  NAND2_X1 U4296 ( .A1(n3588), .A2(n3589), .ZN(n3716) );
  NAND2_X1 U4297 ( .A1(n3718), .A2(n3716), .ZN(n3592) );
  INV_X1 U4298 ( .A(n3588), .ZN(n3591) );
  INV_X1 U4299 ( .A(n3589), .ZN(n3590) );
  NAND2_X1 U4300 ( .A1(n3591), .A2(n3590), .ZN(n3715) );
  NAND2_X1 U4301 ( .A1(n3592), .A2(n3715), .ZN(n3597) );
  OAI22_X1 U4302 ( .A1(n4315), .A2(n3579), .B1(n3682), .B2(n3593), .ZN(n3594)
         );
  XOR2_X1 U4303 ( .A(n2971), .B(n3594), .Z(n3598) );
  NAND2_X1 U4304 ( .A1(n3597), .A2(n3598), .ZN(n3798) );
  NAND2_X1 U4305 ( .A1(n3947), .A2(n3540), .ZN(n3596) );
  NAND2_X1 U4306 ( .A1(n3932), .A2(n3529), .ZN(n3595) );
  NAND2_X1 U4307 ( .A1(n3596), .A2(n3595), .ZN(n3927) );
  NAND2_X1 U4308 ( .A1(n3798), .A2(n3927), .ZN(n3604) );
  INV_X1 U4309 ( .A(n3597), .ZN(n3600) );
  OAI22_X1 U4310 ( .A1(n3602), .A2(n3684), .B1(n3657), .B2(n3601), .ZN(n3606)
         );
  OAI22_X1 U4311 ( .A1(n3602), .A2(n3657), .B1(n3682), .B2(n3601), .ZN(n3603)
         );
  XNOR2_X1 U4312 ( .A(n3603), .B(n2971), .ZN(n3605) );
  XOR2_X1 U4313 ( .A(n3606), .B(n3605), .Z(n3800) );
  INV_X1 U4314 ( .A(n3605), .ZN(n3608) );
  INV_X1 U4315 ( .A(n3606), .ZN(n3607) );
  NAND2_X1 U4316 ( .A1(n3608), .A2(n3607), .ZN(n3609) );
  NAND2_X1 U4317 ( .A1(n4312), .A2(n3529), .ZN(n3611) );
  NAND2_X1 U4318 ( .A1(n3813), .A2(n2968), .ZN(n3610) );
  NAND2_X1 U4319 ( .A1(n3611), .A2(n3610), .ZN(n3612) );
  XNOR2_X1 U4320 ( .A(n3612), .B(n2971), .ZN(n3809) );
  NAND2_X1 U4321 ( .A1(n4312), .A2(n3540), .ZN(n3614) );
  NAND2_X1 U4322 ( .A1(n3813), .A2(n3529), .ZN(n3613) );
  NAND2_X1 U4323 ( .A1(n3614), .A2(n3613), .ZN(n3810) );
  NOR2_X1 U4324 ( .A1(n3809), .A2(n3810), .ZN(n3615) );
  NAND2_X1 U4325 ( .A1(n3809), .A2(n3810), .ZN(n3616) );
  OAI22_X1 U4326 ( .A1(n3619), .A2(n3579), .B1(n3682), .B2(n3617), .ZN(n3618)
         );
  XNOR2_X1 U4327 ( .A(n3618), .B(n3667), .ZN(n3623) );
  OR2_X1 U4328 ( .A1(n3619), .A2(n3684), .ZN(n3621) );
  NAND2_X1 U4329 ( .A1(n3897), .A2(n3529), .ZN(n3620) );
  AND2_X1 U4330 ( .A1(n3621), .A2(n3620), .ZN(n3622) );
  NOR2_X1 U4331 ( .A1(n3623), .A2(n3622), .ZN(n3891) );
  NAND2_X1 U4332 ( .A1(n3623), .A2(n3622), .ZN(n3892) );
  OAI22_X1 U4333 ( .A1(n4195), .A2(n3684), .B1(n3657), .B2(n4225), .ZN(n3628)
         );
  NAND2_X1 U4334 ( .A1(n3945), .A2(n3529), .ZN(n3625) );
  NAND2_X1 U4335 ( .A1(n3750), .A2(n2968), .ZN(n3624) );
  NAND2_X1 U4336 ( .A1(n3625), .A2(n3624), .ZN(n3626) );
  XNOR2_X1 U4337 ( .A(n3626), .B(n2971), .ZN(n3627) );
  XOR2_X1 U4338 ( .A(n3628), .B(n3627), .Z(n3746) );
  NAND2_X1 U4339 ( .A1(n3747), .A2(n3746), .ZN(n3632) );
  NAND2_X1 U4340 ( .A1(n3632), .A2(n3631), .ZN(n3847) );
  NAND2_X1 U4341 ( .A1(n4288), .A2(n3529), .ZN(n3634) );
  NAND2_X1 U4342 ( .A1(n4192), .A2(n2968), .ZN(n3633) );
  NAND2_X1 U4343 ( .A1(n3634), .A2(n3633), .ZN(n3635) );
  XNOR2_X1 U4344 ( .A(n3635), .B(n2971), .ZN(n3638) );
  NAND2_X1 U4345 ( .A1(n4288), .A2(n3540), .ZN(n3637) );
  NAND2_X1 U4346 ( .A1(n4192), .A2(n3529), .ZN(n3636) );
  NAND2_X1 U4347 ( .A1(n3637), .A2(n3636), .ZN(n3639) );
  NAND2_X1 U4348 ( .A1(n3638), .A2(n3639), .ZN(n3848) );
  NAND2_X1 U4349 ( .A1(n3847), .A2(n3848), .ZN(n3846) );
  INV_X1 U4350 ( .A(n3638), .ZN(n3641) );
  INV_X1 U4351 ( .A(n3639), .ZN(n3640) );
  NAND2_X1 U4352 ( .A1(n3641), .A2(n3640), .ZN(n3850) );
  NAND2_X1 U4353 ( .A1(n4193), .A2(n3529), .ZN(n3643) );
  OR2_X1 U4354 ( .A1(n4181), .A2(n3682), .ZN(n3642) );
  NAND2_X1 U4355 ( .A1(n3643), .A2(n3642), .ZN(n3644) );
  XNOR2_X1 U4356 ( .A(n3644), .B(n2971), .ZN(n3769) );
  NAND2_X1 U4357 ( .A1(n4193), .A2(n3540), .ZN(n3646) );
  OR2_X1 U4358 ( .A1(n4181), .A2(n3579), .ZN(n3645) );
  NAND2_X1 U4359 ( .A1(n3646), .A2(n3645), .ZN(n3768) );
  AOI22_X1 U4360 ( .A1(n4176), .A2(n3529), .B1(n2968), .B2(n3648), .ZN(n3647)
         );
  XNOR2_X1 U4361 ( .A(n3647), .B(n2971), .ZN(n3649) );
  AOI22_X1 U4362 ( .A1(n4176), .A2(n3540), .B1(n3529), .B2(n3648), .ZN(n3650)
         );
  XNOR2_X1 U4363 ( .A(n3649), .B(n3650), .ZN(n3871) );
  INV_X1 U4364 ( .A(n3649), .ZN(n3652) );
  INV_X1 U4365 ( .A(n3650), .ZN(n3651) );
  NOR2_X1 U4366 ( .A1(n3652), .A2(n3651), .ZN(n3728) );
  OAI22_X1 U4367 ( .A1(n4151), .A2(n3579), .B1(n3682), .B2(n4138), .ZN(n3653)
         );
  XNOR2_X1 U4368 ( .A(n3653), .B(n2971), .ZN(n3656) );
  OAI22_X1 U4369 ( .A1(n4151), .A2(n3684), .B1(n3657), .B2(n4138), .ZN(n3655)
         );
  XNOR2_X1 U4370 ( .A(n3656), .B(n3655), .ZN(n3727) );
  NOR2_X1 U4371 ( .A1(n3728), .A2(n3727), .ZN(n3654) );
  NAND2_X1 U4372 ( .A1(n3656), .A2(n3655), .ZN(n3660) );
  NOR2_X1 U4373 ( .A1(n4267), .A2(n3657), .ZN(n3658) );
  AOI21_X1 U4374 ( .B1(n4259), .B2(n3540), .A(n3658), .ZN(n3661) );
  OAI22_X1 U4375 ( .A1(n4134), .A2(n3579), .B1(n3682), .B2(n4267), .ZN(n3659)
         );
  XNOR2_X1 U4376 ( .A(n3659), .B(n2971), .ZN(n3822) );
  NAND2_X1 U4377 ( .A1(n3819), .A2(n3822), .ZN(n3664) );
  INV_X1 U4378 ( .A(n3661), .ZN(n3662) );
  NAND2_X1 U4379 ( .A1(n3663), .A2(n3662), .ZN(n3820) );
  NAND2_X1 U4380 ( .A1(n3664), .A2(n3820), .ZN(n3790) );
  NAND2_X1 U4381 ( .A1(n4119), .A2(n3529), .ZN(n3666) );
  NAND2_X1 U4382 ( .A1(n4258), .A2(n2968), .ZN(n3665) );
  NAND2_X1 U4383 ( .A1(n3666), .A2(n3665), .ZN(n3668) );
  XNOR2_X1 U4384 ( .A(n3668), .B(n3667), .ZN(n3670) );
  AND2_X1 U4385 ( .A1(n4258), .A2(n3529), .ZN(n3669) );
  AOI21_X1 U4386 ( .B1(n4119), .B2(n3540), .A(n3669), .ZN(n3671) );
  NAND2_X1 U4387 ( .A1(n3670), .A2(n3671), .ZN(n3788) );
  INV_X1 U4388 ( .A(n3670), .ZN(n3673) );
  INV_X1 U4389 ( .A(n3671), .ZN(n3672) );
  NAND2_X1 U4390 ( .A1(n3673), .A2(n3672), .ZN(n3789) );
  OAI22_X1 U4391 ( .A1(n4262), .A2(n3579), .B1(n3682), .B2(n4085), .ZN(n3674)
         );
  XNOR2_X1 U4392 ( .A(n3674), .B(n2971), .ZN(n3675) );
  OAI22_X1 U4393 ( .A1(n4262), .A2(n3684), .B1(n3579), .B2(n4085), .ZN(n3676)
         );
  AND2_X1 U4394 ( .A1(n3675), .A2(n3676), .ZN(n3915) );
  INV_X1 U4395 ( .A(n3675), .ZN(n3678) );
  INV_X1 U4396 ( .A(n3676), .ZN(n3677) );
  AOI22_X1 U4397 ( .A1(n3943), .A2(n3529), .B1(n3708), .B2(n2968), .ZN(n3679)
         );
  XNOR2_X1 U4398 ( .A(n3679), .B(n2971), .ZN(n3680) );
  AOI22_X1 U4399 ( .A1(n3943), .A2(n3540), .B1(n3708), .B2(n3529), .ZN(n3681)
         );
  XNOR2_X1 U4400 ( .A(n3680), .B(n3681), .ZN(n3707) );
  OAI22_X1 U4401 ( .A1(n3685), .A2(n3579), .B1(n3682), .B2(n3683), .ZN(n3688)
         );
  OAI22_X1 U4402 ( .A1(n3685), .A2(n3684), .B1(n3579), .B2(n3683), .ZN(n3686)
         );
  XNOR2_X1 U4403 ( .A(n3686), .B(n2971), .ZN(n3687) );
  XOR2_X1 U4404 ( .A(n3688), .B(n3687), .Z(n3689) );
  NAND2_X1 U4405 ( .A1(n3942), .A2(n3931), .ZN(n3694) );
  AOI22_X1 U4406 ( .A1(n3933), .A2(n3690), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3693) );
  NAND2_X1 U4407 ( .A1(n3691), .A2(n3936), .ZN(n3692) );
  NAND3_X1 U4408 ( .A1(n3694), .A2(n3693), .A3(n3692), .ZN(n3695) );
  AOI21_X1 U4409 ( .B1(n3934), .B2(n3943), .A(n3695), .ZN(n3696) );
  XOR2_X1 U4410 ( .A(n3698), .B(n3697), .Z(n3699) );
  NAND2_X1 U4411 ( .A1(n3699), .A2(n3929), .ZN(n3706) );
  AOI21_X1 U4412 ( .B1(n3931), .B2(n3954), .A(n3700), .ZN(n3705) );
  AOI22_X1 U4413 ( .A1(n3701), .A2(n3933), .B1(n3934), .B2(n3956), .ZN(n3704)
         );
  NAND2_X1 U4414 ( .A1(n3936), .A2(n3702), .ZN(n3703) );
  NAND4_X1 U4415 ( .A1(n3706), .A2(n3705), .A3(n3704), .A4(n3703), .ZN(U3210)
         );
  AOI22_X1 U4416 ( .A1(n3933), .A2(n3708), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3709) );
  OAI21_X1 U4417 ( .B1(n4262), .B2(n3919), .A(n3709), .ZN(n3710) );
  AOI21_X1 U4418 ( .B1(n4247), .B2(n3931), .A(n3710), .ZN(n3713) );
  NAND2_X1 U4419 ( .A1(n3711), .A2(n3936), .ZN(n3712) );
  OAI211_X1 U4420 ( .C1(n3714), .C2(n3925), .A(n3713), .B(n3712), .ZN(U3211)
         );
  NAND2_X1 U4421 ( .A1(n3716), .A2(n3715), .ZN(n3717) );
  XNOR2_X1 U4422 ( .A(n3718), .B(n3717), .ZN(n3725) );
  AOI22_X1 U4423 ( .A1(n3949), .A2(n3934), .B1(n3933), .B2(n3719), .ZN(n3721)
         );
  NOR2_X1 U4424 ( .A1(n4708), .A2(STATE_REG_SCAN_IN), .ZN(n4444) );
  INV_X1 U4425 ( .A(n4444), .ZN(n3720) );
  OAI211_X1 U4426 ( .C1(n4315), .C2(n3875), .A(n3721), .B(n3720), .ZN(n3722)
         );
  AOI21_X1 U4427 ( .B1(n3723), .B2(n3936), .A(n3722), .ZN(n3724) );
  OAI21_X1 U4428 ( .B1(n3725), .B2(n3925), .A(n3724), .ZN(U3212) );
  INV_X1 U4429 ( .A(n3726), .ZN(n3869) );
  OAI21_X1 U4430 ( .B1(n3869), .B2(n3728), .A(n3727), .ZN(n3730) );
  NAND3_X1 U4431 ( .A1(n3730), .A2(n3929), .A3(n3729), .ZN(n3734) );
  INV_X1 U4432 ( .A(n4176), .ZN(n4292) );
  OAI22_X1 U4433 ( .A1(n4292), .A2(n3919), .B1(n3874), .B2(n4138), .ZN(n3732)
         );
  NOR2_X1 U4434 ( .A1(n4134), .A2(n3875), .ZN(n3731) );
  AOI211_X1 U4435 ( .C1(REG3_REG_23__SCAN_IN), .C2(U3149), .A(n3732), .B(n3731), .ZN(n3733) );
  OAI211_X1 U4436 ( .C1(n3922), .C2(n4141), .A(n3734), .B(n3733), .ZN(U3213)
         );
  AOI21_X1 U4437 ( .B1(n3736), .B2(n3735), .A(n3925), .ZN(n3738) );
  NAND2_X1 U4438 ( .A1(n3738), .A2(n3737), .ZN(n3745) );
  NAND2_X1 U4439 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4399) );
  INV_X1 U4440 ( .A(n4399), .ZN(n3739) );
  AOI21_X1 U4441 ( .B1(n3951), .B2(n3931), .A(n3739), .ZN(n3744) );
  AOI22_X1 U4442 ( .A1(n3740), .A2(n3933), .B1(n3934), .B2(n3953), .ZN(n3743)
         );
  NAND2_X1 U4443 ( .A1(n3936), .A2(n3741), .ZN(n3742) );
  NAND4_X1 U4444 ( .A1(n3745), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(U3214)
         );
  XNOR2_X1 U4445 ( .A(n3747), .B(n3746), .ZN(n3748) );
  NAND2_X1 U4446 ( .A1(n3748), .A2(n3929), .ZN(n3754) );
  NAND2_X1 U4447 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4050) );
  INV_X1 U4448 ( .A(n4050), .ZN(n3749) );
  AOI21_X1 U4449 ( .B1(n3931), .B2(n4288), .A(n3749), .ZN(n3753) );
  AOI22_X1 U4450 ( .A1(n4220), .A2(n3934), .B1(n3933), .B2(n3750), .ZN(n3752)
         );
  NAND2_X1 U4451 ( .A1(n3936), .A2(n4228), .ZN(n3751) );
  NAND4_X1 U4452 ( .A1(n3754), .A2(n3753), .A3(n3752), .A4(n3751), .ZN(U3216)
         );
  NAND2_X1 U4453 ( .A1(n3756), .A2(n3755), .ZN(n3758) );
  XOR2_X1 U4454 ( .A(n3758), .B(n3757), .Z(n3759) );
  NAND2_X1 U4455 ( .A1(n3759), .A2(n3929), .ZN(n3767) );
  INV_X1 U4456 ( .A(n3760), .ZN(n3761) );
  AOI21_X1 U4457 ( .B1(n3931), .B2(n3953), .A(n3761), .ZN(n3766) );
  AOI22_X1 U4458 ( .A1(n3955), .A2(n3934), .B1(n3933), .B2(n3762), .ZN(n3765)
         );
  NAND2_X1 U4459 ( .A1(n3936), .A2(n3763), .ZN(n3764) );
  NAND4_X1 U4460 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(U3218)
         );
  XNOR2_X1 U4461 ( .A(n3769), .B(n3768), .ZN(n3770) );
  XNOR2_X1 U4462 ( .A(n3771), .B(n3770), .ZN(n3777) );
  INV_X1 U4463 ( .A(n3772), .ZN(n4177) );
  OAI22_X1 U4464 ( .A1(n3919), .A2(n4218), .B1(STATE_REG_SCAN_IN), .B2(n3773), 
        .ZN(n3775) );
  OAI22_X1 U4465 ( .A1(n4292), .A2(n3875), .B1(n3874), .B2(n4181), .ZN(n3774)
         );
  AOI211_X1 U4466 ( .C1(n4177), .C2(n3936), .A(n3775), .B(n3774), .ZN(n3776)
         );
  OAI21_X1 U4467 ( .B1(n3777), .B2(n3925), .A(n3776), .ZN(U3220) );
  NAND2_X1 U4468 ( .A1(n2087), .A2(n3778), .ZN(n3779) );
  XNOR2_X1 U4469 ( .A(n3780), .B(n3779), .ZN(n3781) );
  NAND2_X1 U4470 ( .A1(n3781), .A2(n3929), .ZN(n3787) );
  NAND2_X1 U4471 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4420) );
  INV_X1 U4472 ( .A(n4420), .ZN(n3782) );
  AOI21_X1 U4473 ( .B1(n3949), .B2(n3931), .A(n3782), .ZN(n3786) );
  AOI22_X1 U4474 ( .A1(n3951), .A2(n3934), .B1(n3933), .B2(n2450), .ZN(n3785)
         );
  NAND2_X1 U4475 ( .A1(n3936), .A2(n3783), .ZN(n3784) );
  NAND4_X1 U4476 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(U3221)
         );
  NAND2_X1 U4477 ( .A1(n3789), .A2(n3788), .ZN(n3791) );
  XOR2_X1 U4478 ( .A(n3791), .B(n3790), .Z(n3796) );
  NOR2_X1 U4479 ( .A1(n3922), .A2(n4104), .ZN(n3794) );
  AOI22_X1 U4480 ( .A1(n4259), .A2(n3934), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3792) );
  OAI21_X1 U4481 ( .B1(n3874), .B2(n4100), .A(n3792), .ZN(n3793) );
  AOI211_X1 U4482 ( .C1(n3931), .C2(n3944), .A(n3794), .B(n3793), .ZN(n3795)
         );
  OAI21_X1 U4483 ( .B1(n3796), .B2(n3925), .A(n3795), .ZN(U3222) );
  INV_X1 U4484 ( .A(n3797), .ZN(n3799) );
  OAI21_X1 U4485 ( .B1(n3799), .B2(n3927), .A(n3798), .ZN(n3801) );
  XNOR2_X1 U4486 ( .A(n3801), .B(n3800), .ZN(n3802) );
  NAND2_X1 U4487 ( .A1(n3802), .A2(n3929), .ZN(n3807) );
  AND2_X1 U4488 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4463) );
  AOI21_X1 U4489 ( .B1(n3931), .B2(n4312), .A(n4463), .ZN(n3806) );
  AOI22_X1 U4490 ( .A1(n4309), .A2(n3933), .B1(n3934), .B2(n3947), .ZN(n3805)
         );
  NAND2_X1 U4491 ( .A1(n3936), .A2(n3803), .ZN(n3804) );
  NAND4_X1 U4492 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(U3223)
         );
  XOR2_X1 U4493 ( .A(n3810), .B(n3809), .Z(n3811) );
  XNOR2_X1 U4494 ( .A(n3808), .B(n3811), .ZN(n3812) );
  NAND2_X1 U4495 ( .A1(n3812), .A2(n3929), .ZN(n3818) );
  NOR2_X1 U4496 ( .A1(STATE_REG_SCAN_IN), .A2(n2494), .ZN(n4472) );
  AOI21_X1 U4497 ( .B1(n4220), .B2(n3931), .A(n4472), .ZN(n3817) );
  AOI22_X1 U4498 ( .A1(n3946), .A2(n3934), .B1(n3933), .B2(n3813), .ZN(n3816)
         );
  NAND2_X1 U4499 ( .A1(n3936), .A2(n3814), .ZN(n3815) );
  NAND4_X1 U4500 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(U3225)
         );
  NAND2_X1 U4501 ( .A1(n3820), .A2(n3819), .ZN(n3821) );
  XOR2_X1 U4502 ( .A(n3822), .B(n3821), .Z(n3826) );
  OAI22_X1 U4503 ( .A1(n4151), .A2(n3919), .B1(STATE_REG_SCAN_IN), .B2(n4648), 
        .ZN(n3824) );
  OAI22_X1 U4504 ( .A1(n4272), .A2(n3875), .B1(n3874), .B2(n4267), .ZN(n3823)
         );
  AOI211_X1 U4505 ( .C1(n4120), .C2(n3936), .A(n3824), .B(n3823), .ZN(n3825)
         );
  OAI21_X1 U4506 ( .B1(n3826), .B2(n3925), .A(n3825), .ZN(U3226) );
  OAI211_X1 U4507 ( .C1(n3829), .C2(n3828), .A(n3827), .B(n3929), .ZN(n3836)
         );
  AOI21_X1 U4508 ( .B1(n3957), .B2(n3931), .A(n3830), .ZN(n3835) );
  AOI22_X1 U4509 ( .A1(n3831), .A2(n3933), .B1(n3934), .B2(n3959), .ZN(n3834)
         );
  NAND2_X1 U4510 ( .A1(n3936), .A2(n3832), .ZN(n3833) );
  NAND4_X1 U4511 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(U3227)
         );
  XNOR2_X1 U4512 ( .A(n3837), .B(n3838), .ZN(n3839) );
  NAND2_X1 U4513 ( .A1(n3839), .A2(n3929), .ZN(n3845) );
  NOR2_X1 U4514 ( .A1(STATE_REG_SCAN_IN), .A2(n2306), .ZN(n4395) );
  AOI21_X1 U4515 ( .B1(n3952), .B2(n3931), .A(n4395), .ZN(n3844) );
  AOI22_X1 U4516 ( .A1(n3840), .A2(n3933), .B1(n3934), .B2(n3954), .ZN(n3843)
         );
  NAND2_X1 U4517 ( .A1(n3936), .A2(n3841), .ZN(n3842) );
  NAND4_X1 U4518 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(U3228)
         );
  INV_X1 U4519 ( .A(n3846), .ZN(n3851) );
  AOI21_X1 U4520 ( .B1(n3850), .B2(n3848), .A(n3847), .ZN(n3849) );
  AOI21_X1 U4521 ( .B1(n3851), .B2(n3850), .A(n3849), .ZN(n3857) );
  INV_X1 U4522 ( .A(n4204), .ZN(n3855) );
  OAI22_X1 U4523 ( .A1(n3874), .A2(n4202), .B1(n3919), .B2(n4195), .ZN(n3854)
         );
  OAI22_X1 U4524 ( .A1(n3873), .A2(n3875), .B1(STATE_REG_SCAN_IN), .B2(n3852), 
        .ZN(n3853) );
  AOI211_X1 U4525 ( .C1(n3855), .C2(n3936), .A(n3854), .B(n3853), .ZN(n3856)
         );
  OAI21_X1 U4526 ( .B1(n3857), .B2(n3925), .A(n3856), .ZN(U3230) );
  XNOR2_X1 U4527 ( .A(n3859), .B(n3858), .ZN(n3860) );
  XNOR2_X1 U4528 ( .A(n3861), .B(n3860), .ZN(n3862) );
  NAND2_X1 U4529 ( .A1(n3862), .A2(n3929), .ZN(n3868) );
  NOR2_X1 U4530 ( .A1(STATE_REG_SCAN_IN), .A2(n2457), .ZN(n4433) );
  AOI21_X1 U4531 ( .B1(n3948), .B2(n3931), .A(n4433), .ZN(n3867) );
  AOI22_X1 U4532 ( .A1(n3950), .A2(n3934), .B1(n3933), .B2(n3863), .ZN(n3866)
         );
  NAND2_X1 U4533 ( .A1(n3936), .A2(n3864), .ZN(n3865) );
  NAND4_X1 U4534 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(U3231)
         );
  AOI21_X1 U4535 ( .B1(n3871), .B2(n3870), .A(n3869), .ZN(n3879) );
  OAI22_X1 U4536 ( .A1(n3873), .A2(n3919), .B1(STATE_REG_SCAN_IN), .B2(n3872), 
        .ZN(n3877) );
  OAI22_X1 U4537 ( .A1(n4151), .A2(n3875), .B1(n3874), .B2(n4160), .ZN(n3876)
         );
  AOI211_X1 U4538 ( .C1(n4162), .C2(n3936), .A(n3877), .B(n3876), .ZN(n3878)
         );
  OAI21_X1 U4539 ( .B1(n3879), .B2(n3925), .A(n3878), .ZN(U3232) );
  XNOR2_X1 U4540 ( .A(n3881), .B(n3880), .ZN(n3882) );
  XNOR2_X1 U4541 ( .A(n3883), .B(n3882), .ZN(n3884) );
  NAND2_X1 U4542 ( .A1(n3884), .A2(n3929), .ZN(n3890) );
  AND2_X1 U4543 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4416) );
  AOI21_X1 U4544 ( .B1(n3950), .B2(n3931), .A(n4416), .ZN(n3889) );
  AOI22_X1 U4545 ( .A1(n3952), .A2(n3934), .B1(n3933), .B2(n3885), .ZN(n3888)
         );
  NAND2_X1 U4546 ( .A1(n3936), .A2(n3886), .ZN(n3887) );
  NAND4_X1 U4547 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(U3233)
         );
  INV_X1 U4548 ( .A(n3891), .ZN(n3893) );
  NAND2_X1 U4549 ( .A1(n3893), .A2(n3892), .ZN(n3894) );
  XNOR2_X1 U4550 ( .A(n3895), .B(n3894), .ZN(n3896) );
  NAND2_X1 U4551 ( .A1(n3896), .A2(n3929), .ZN(n3902) );
  AND2_X1 U4552 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4481) );
  AOI21_X1 U4553 ( .B1(n3931), .B2(n3945), .A(n4481), .ZN(n3901) );
  AOI22_X1 U4554 ( .A1(n3897), .A2(n3933), .B1(n3934), .B2(n4312), .ZN(n3900)
         );
  NAND2_X1 U4555 ( .A1(n3936), .A2(n3898), .ZN(n3899) );
  NAND4_X1 U4556 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(U3235)
         );
  XNOR2_X1 U4557 ( .A(n3904), .B(n3903), .ZN(n3905) );
  XNOR2_X1 U4558 ( .A(n3906), .B(n3905), .ZN(n3907) );
  NAND2_X1 U4559 ( .A1(n3907), .A2(n3929), .ZN(n3914) );
  AOI21_X1 U4560 ( .B1(n3955), .B2(n3931), .A(n3908), .ZN(n3913) );
  AOI22_X1 U4561 ( .A1(n3957), .A2(n3934), .B1(n3933), .B2(n3909), .ZN(n3912)
         );
  NAND2_X1 U4562 ( .A1(n3936), .A2(n3910), .ZN(n3911) );
  NAND4_X1 U4563 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(U3236)
         );
  NOR2_X1 U4564 ( .A1(n2074), .A2(n3915), .ZN(n3916) );
  XNOR2_X1 U4565 ( .A(n3917), .B(n3916), .ZN(n3926) );
  OAI22_X1 U4566 ( .A1(n4272), .A2(n3919), .B1(STATE_REG_SCAN_IN), .B2(n3918), 
        .ZN(n3920) );
  AOI21_X1 U4567 ( .B1(n4080), .B2(n3933), .A(n3920), .ZN(n3921) );
  OAI21_X1 U4568 ( .B1(n3922), .B2(n4088), .A(n3921), .ZN(n3923) );
  AOI21_X1 U4569 ( .B1(n3931), .B2(n3943), .A(n3923), .ZN(n3924) );
  OAI21_X1 U4570 ( .B1(n3926), .B2(n3925), .A(n3924), .ZN(U3237) );
  NAND2_X1 U4571 ( .A1(n3797), .A2(n3798), .ZN(n3928) );
  XNOR2_X1 U4572 ( .A(n3928), .B(n3927), .ZN(n3930) );
  NAND2_X1 U4573 ( .A1(n3930), .A2(n3929), .ZN(n3940) );
  AND2_X1 U4574 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4453) );
  AOI21_X1 U4575 ( .B1(n3946), .B2(n3931), .A(n4453), .ZN(n3939) );
  AOI22_X1 U4576 ( .A1(n3948), .A2(n3934), .B1(n3933), .B2(n3932), .ZN(n3938)
         );
  NAND2_X1 U4577 ( .A1(n3936), .A2(n3935), .ZN(n3937) );
  NAND4_X1 U4578 ( .A1(n3940), .A2(n3939), .A3(n3938), .A4(n3937), .ZN(U3238)
         );
  MUX2_X1 U4579 ( .A(DATAO_REG_31__SCAN_IN), .B(n4057), .S(n3961), .Z(U3581)
         );
  MUX2_X1 U4580 ( .A(DATAO_REG_30__SCAN_IN), .B(n3941), .S(n3961), .Z(U3580)
         );
  MUX2_X1 U4581 ( .A(DATAO_REG_29__SCAN_IN), .B(n3942), .S(n3961), .Z(U3579)
         );
  MUX2_X1 U4582 ( .A(DATAO_REG_28__SCAN_IN), .B(n4247), .S(n3961), .Z(U3578)
         );
  MUX2_X1 U4583 ( .A(DATAO_REG_27__SCAN_IN), .B(n3943), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4584 ( .A(DATAO_REG_26__SCAN_IN), .B(n3944), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4585 ( .A(DATAO_REG_25__SCAN_IN), .B(n4119), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4586 ( .A(DATAO_REG_24__SCAN_IN), .B(n4259), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4587 ( .A(DATAO_REG_23__SCAN_IN), .B(n4269), .S(n3961), .Z(U3573)
         );
  MUX2_X1 U4588 ( .A(DATAO_REG_22__SCAN_IN), .B(n4176), .S(n3961), .Z(U3572)
         );
  MUX2_X1 U4589 ( .A(DATAO_REG_21__SCAN_IN), .B(n4193), .S(n3961), .Z(U3571)
         );
  MUX2_X1 U4590 ( .A(DATAO_REG_20__SCAN_IN), .B(n4288), .S(n3961), .Z(U3570)
         );
  MUX2_X1 U4591 ( .A(DATAO_REG_19__SCAN_IN), .B(n3945), .S(n3961), .Z(U3569)
         );
  MUX2_X1 U4592 ( .A(DATAO_REG_18__SCAN_IN), .B(n4220), .S(n3961), .Z(U3568)
         );
  MUX2_X1 U4593 ( .A(DATAO_REG_17__SCAN_IN), .B(n4312), .S(n3961), .Z(U3567)
         );
  MUX2_X1 U4594 ( .A(DATAO_REG_16__SCAN_IN), .B(n3946), .S(n3961), .Z(U3566)
         );
  MUX2_X1 U4595 ( .A(DATAO_REG_15__SCAN_IN), .B(n3947), .S(n3961), .Z(U3565)
         );
  MUX2_X1 U4596 ( .A(DATAO_REG_14__SCAN_IN), .B(n3948), .S(n3961), .Z(U3564)
         );
  MUX2_X1 U4597 ( .A(DATAO_REG_13__SCAN_IN), .B(n3949), .S(n3961), .Z(U3563)
         );
  MUX2_X1 U4598 ( .A(DATAO_REG_12__SCAN_IN), .B(n3950), .S(n3961), .Z(U3562)
         );
  MUX2_X1 U4599 ( .A(DATAO_REG_11__SCAN_IN), .B(n3951), .S(n3961), .Z(U3561)
         );
  MUX2_X1 U4600 ( .A(DATAO_REG_10__SCAN_IN), .B(n3952), .S(n3961), .Z(U3560)
         );
  MUX2_X1 U4601 ( .A(DATAO_REG_9__SCAN_IN), .B(n3953), .S(n3961), .Z(U3559) );
  MUX2_X1 U4602 ( .A(DATAO_REG_8__SCAN_IN), .B(n3954), .S(n3961), .Z(U3558) );
  MUX2_X1 U4603 ( .A(DATAO_REG_7__SCAN_IN), .B(n3955), .S(n3961), .Z(U3557) );
  MUX2_X1 U4604 ( .A(DATAO_REG_6__SCAN_IN), .B(n3956), .S(n3961), .Z(U3556) );
  MUX2_X1 U4605 ( .A(DATAO_REG_5__SCAN_IN), .B(n3957), .S(n3961), .Z(U3555) );
  MUX2_X1 U4606 ( .A(DATAO_REG_4__SCAN_IN), .B(n3958), .S(n3961), .Z(U3554) );
  MUX2_X1 U4607 ( .A(DATAO_REG_3__SCAN_IN), .B(n3959), .S(n3961), .Z(U3553) );
  MUX2_X1 U4608 ( .A(DATAO_REG_2__SCAN_IN), .B(n3960), .S(n3961), .Z(U3552) );
  MUX2_X1 U4609 ( .A(DATAO_REG_1__SCAN_IN), .B(n2808), .S(n3961), .Z(U3551) );
  MUX2_X1 U4610 ( .A(DATAO_REG_0__SCAN_IN), .B(n3962), .S(n3961), .Z(U3550) );
  NAND2_X1 U4611 ( .A1(n3990), .A2(n4382), .ZN(n3971) );
  OAI211_X1 U4612 ( .C1(n3965), .C2(n3964), .A(n4484), .B(n3963), .ZN(n3970)
         );
  OAI211_X1 U4613 ( .C1(n2760), .C2(n3967), .A(n4429), .B(n3979), .ZN(n3969)
         );
  AOI22_X1 U4614 ( .A1(n4482), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3968) );
  NAND4_X1 U4615 ( .A1(n3971), .A2(n3970), .A3(n3969), .A4(n3968), .ZN(U3241)
         );
  NOR2_X1 U4616 ( .A1(n3972), .A2(STATE_REG_SCAN_IN), .ZN(n3973) );
  AOI21_X1 U4617 ( .B1(n4482), .B2(ADDR_REG_2__SCAN_IN), .A(n3973), .ZN(n3974)
         );
  OAI21_X1 U4618 ( .B1(n4489), .B2(n3975), .A(n3974), .ZN(n3976) );
  INV_X1 U4619 ( .A(n3976), .ZN(n3988) );
  MUX2_X1 U4620 ( .A(n3977), .B(REG2_REG_2__SCAN_IN), .S(n4381), .Z(n3980) );
  NAND3_X1 U4621 ( .A1(n3980), .A2(n3979), .A3(n3978), .ZN(n3981) );
  NAND3_X1 U4622 ( .A1(n4429), .A2(n3982), .A3(n3981), .ZN(n3987) );
  OAI211_X1 U4623 ( .C1(n3985), .C2(n3984), .A(n4484), .B(n3983), .ZN(n3986)
         );
  NAND4_X1 U4624 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(U3242)
         );
  NAND2_X1 U4625 ( .A1(n3990), .A2(n4380), .ZN(n3999) );
  OAI211_X1 U4626 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3992), .A(n4484), .B(n3991), 
        .ZN(n3998) );
  AOI22_X1 U4627 ( .A1(n4482), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3997) );
  XNOR2_X1 U4628 ( .A(n3994), .B(n3993), .ZN(n3995) );
  NAND2_X1 U4629 ( .A1(n4429), .A2(n3995), .ZN(n3996) );
  NAND4_X1 U4630 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(U3243)
         );
  INV_X1 U4631 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4000) );
  MUX2_X1 U4632 ( .A(n4000), .B(REG2_REG_19__SCAN_IN), .S(n4051), .Z(n4019) );
  INV_X1 U4633 ( .A(n4020), .ZN(n4505) );
  INV_X1 U4634 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4635 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4505), .B1(n4020), .B2(
        n4001), .ZN(n4480) );
  NOR2_X1 U4636 ( .A1(n4044), .A2(REG2_REG_17__SCAN_IN), .ZN(n4002) );
  AOI21_X1 U4637 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4044), .A(n4002), .ZN(n4470) );
  INV_X1 U4638 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4428) );
  NOR2_X1 U4639 ( .A1(n4428), .A2(n4509), .ZN(n4427) );
  NAND2_X1 U4640 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4023), .ZN(n4010) );
  INV_X1 U4641 ( .A(n4023), .ZN(n4512) );
  INV_X1 U4642 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4643 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4023), .B1(n4512), .B2(
        n4003), .ZN(n4412) );
  NAND2_X1 U4644 ( .A1(n4025), .A2(REG2_REG_9__SCAN_IN), .ZN(n4007) );
  INV_X1 U4645 ( .A(n4025), .ZN(n4516) );
  AOI22_X1 U4646 ( .A1(n4025), .A2(REG2_REG_9__SCAN_IN), .B1(n4004), .B2(n4516), .ZN(n4391) );
  INV_X1 U4647 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4492) );
  OAI22_X1 U4648 ( .A1(n4006), .A2(n4492), .B1(n4005), .B2(n4027), .ZN(n4390)
         );
  NAND2_X1 U4649 ( .A1(n4391), .A2(n4390), .ZN(n4389) );
  NAND2_X1 U4650 ( .A1(n4007), .A2(n4389), .ZN(n4008) );
  NAND2_X1 U4651 ( .A1(n4513), .A2(n4008), .ZN(n4009) );
  XNOR2_X1 U4652 ( .A(n4008), .B(n4406), .ZN(n4398) );
  NAND2_X1 U4653 ( .A1(n4033), .A2(n4011), .ZN(n4012) );
  XNOR2_X1 U4654 ( .A(n4011), .B(n4510), .ZN(n4419) );
  NOR2_X1 U4655 ( .A1(n2180), .A2(n4013), .ZN(n4014) );
  INV_X1 U4656 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4442) );
  NOR2_X1 U4657 ( .A1(n4442), .A2(n4441), .ZN(n4440) );
  NOR2_X1 U4658 ( .A1(n4014), .A2(n4440), .ZN(n4451) );
  NAND2_X1 U4659 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4021), .ZN(n4015) );
  OAI21_X1 U4660 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4021), .A(n4015), .ZN(n4450) );
  NOR2_X1 U4661 ( .A1(n4451), .A2(n4450), .ZN(n4449) );
  INV_X1 U4662 ( .A(n4041), .ZN(n4507) );
  NAND2_X1 U4663 ( .A1(n4016), .A2(n4507), .ZN(n4017) );
  INV_X1 U4664 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4459) );
  NAND2_X1 U4665 ( .A1(n4470), .A2(n4468), .ZN(n4469) );
  AOI21_X1 U4666 ( .B1(n4020), .B2(REG2_REG_18__SCAN_IN), .A(n4479), .ZN(n4018) );
  XOR2_X1 U4667 ( .A(n4019), .B(n4018), .Z(n4055) );
  INV_X1 U4668 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U4669 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4020), .B1(n4505), .B2(
        n4046), .ZN(n4486) );
  NOR2_X1 U4670 ( .A1(n4044), .A2(REG1_REG_17__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U4671 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4021), .ZN(n4040) );
  INV_X1 U4672 ( .A(n4021), .ZN(n4508) );
  AOI22_X1 U4673 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4021), .B1(n4508), .B2(
        n3457), .ZN(n4456) );
  NAND2_X1 U4674 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4022), .ZN(n4036) );
  AOI22_X1 U4675 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4022), .B1(n4509), .B2(
        n3412), .ZN(n4437) );
  NAND2_X1 U4676 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4023), .ZN(n4032) );
  AOI22_X1 U4677 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4023), .B1(n4512), .B2(
        n3198), .ZN(n4409) );
  NAND2_X1 U4678 ( .A1(n4025), .A2(REG1_REG_9__SCAN_IN), .ZN(n4029) );
  INV_X1 U4679 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4680 ( .A1(n4025), .A2(REG1_REG_9__SCAN_IN), .B1(n4024), .B2(n4516), .ZN(n4388) );
  NAND2_X1 U4681 ( .A1(n4513), .A2(n4030), .ZN(n4031) );
  XNOR2_X1 U4682 ( .A(n4030), .B(n4406), .ZN(n4403) );
  NAND2_X1 U4683 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4403), .ZN(n4402) );
  NAND2_X1 U4684 ( .A1(n4033), .A2(n4034), .ZN(n4035) );
  NAND2_X1 U4685 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4424), .ZN(n4423) );
  NAND2_X1 U4686 ( .A1(n4035), .A2(n4423), .ZN(n4436) );
  NAND2_X1 U4687 ( .A1(n4437), .A2(n4436), .ZN(n4435) );
  NAND2_X1 U4688 ( .A1(n4036), .A2(n4435), .ZN(n4038) );
  NAND2_X1 U4689 ( .A1(n4037), .A2(n4038), .ZN(n4039) );
  XNOR2_X1 U4690 ( .A(n4038), .B(n2180), .ZN(n4446) );
  NAND2_X1 U4691 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4446), .ZN(n4445) );
  NAND2_X1 U4692 ( .A1(n4039), .A2(n4445), .ZN(n4455) );
  NAND2_X1 U4693 ( .A1(n4456), .A2(n4455), .ZN(n4454) );
  NOR2_X1 U4694 ( .A1(n4041), .A2(n4042), .ZN(n4043) );
  INV_X1 U4695 ( .A(n4044), .ZN(n4506) );
  AOI22_X1 U4696 ( .A1(n4044), .A2(n3498), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4506), .ZN(n4473) );
  NOR2_X1 U4697 ( .A1(n4474), .A2(n4473), .ZN(n4475) );
  INV_X1 U4698 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4047) );
  MUX2_X1 U4699 ( .A(REG1_REG_19__SCAN_IN), .B(n4047), .S(n4051), .Z(n4048) );
  NAND2_X1 U4700 ( .A1(n4482), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4049) );
  OAI211_X1 U4701 ( .C1(n4489), .C2(n4051), .A(n4050), .B(n4049), .ZN(n4052)
         );
  AOI21_X1 U4702 ( .B1(n4053), .B2(n4484), .A(n4052), .ZN(n4054) );
  OAI21_X1 U4703 ( .B1(n4055), .B2(n4478), .A(n4054), .ZN(U3259) );
  XNOR2_X1 U4704 ( .A(n4238), .B(n4058), .ZN(n4326) );
  NAND2_X1 U4705 ( .A1(n4057), .A2(n4056), .ZN(n4240) );
  OAI21_X1 U4706 ( .B1(n4058), .B2(n4244), .A(n4240), .ZN(n4323) );
  NAND2_X1 U4707 ( .A1(n4323), .A2(n4493), .ZN(n4060) );
  NAND2_X1 U4708 ( .A1(n4229), .A2(REG2_REG_31__SCAN_IN), .ZN(n4059) );
  OAI211_X1 U4709 ( .C1(n4326), .C2(n4231), .A(n4060), .B(n4059), .ZN(U3260)
         );
  INV_X1 U4710 ( .A(n4061), .ZN(n4072) );
  INV_X1 U4711 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4062) );
  OAI22_X1 U4712 ( .A1(n4180), .A2(n4063), .B1(n4062), .B2(n4493), .ZN(n4064)
         );
  AOI21_X1 U4713 ( .B1(n4247), .B2(n4174), .A(n4064), .ZN(n4071) );
  INV_X1 U4714 ( .A(n4065), .ZN(n4069) );
  OAI22_X1 U4715 ( .A1(n4067), .A2(n4231), .B1(n4066), .B2(n4490), .ZN(n4068)
         );
  OAI21_X1 U4716 ( .B1(n4069), .B2(n4068), .A(n4493), .ZN(n4070) );
  OAI211_X1 U4717 ( .C1(n4072), .C2(n4234), .A(n4071), .B(n4070), .ZN(U3354)
         );
  XNOR2_X1 U4718 ( .A(n4073), .B(n4077), .ZN(n4255) );
  INV_X1 U4719 ( .A(n4255), .ZN(n4092) );
  INV_X1 U4720 ( .A(n4094), .ZN(n4076) );
  OAI21_X1 U4721 ( .B1(n4076), .B2(n4075), .A(n4074), .ZN(n4078) );
  XNOR2_X1 U4722 ( .A(n4078), .B(n4077), .ZN(n4079) );
  NAND2_X1 U4723 ( .A1(n4079), .A2(n4197), .ZN(n4082) );
  AOI22_X1 U4724 ( .A1(n4119), .A2(n4287), .B1(n4080), .B2(n4310), .ZN(n4081)
         );
  OAI211_X1 U4725 ( .C1(n4083), .C2(n4291), .A(n4082), .B(n4081), .ZN(n4254)
         );
  INV_X1 U4726 ( .A(n4099), .ZN(n4086) );
  OAI21_X1 U4727 ( .B1(n4086), .B2(n4085), .A(n4084), .ZN(n4338) );
  NOR2_X1 U4728 ( .A1(n4338), .A2(n4231), .ZN(n4090) );
  INV_X1 U4729 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4087) );
  OAI22_X1 U4730 ( .A1(n4088), .A2(n4490), .B1(n4087), .B2(n4493), .ZN(n4089)
         );
  AOI211_X1 U4731 ( .C1(n4254), .C2(n4493), .A(n4090), .B(n4089), .ZN(n4091)
         );
  OAI21_X1 U4732 ( .B1(n4092), .B2(n4234), .A(n4091), .ZN(U3264) );
  NAND2_X1 U4733 ( .A1(n4094), .A2(n4093), .ZN(n4095) );
  XNOR2_X1 U4734 ( .A(n4095), .B(n4097), .ZN(n4096) );
  NAND2_X1 U4735 ( .A1(n4096), .A2(n4197), .ZN(n4261) );
  XNOR2_X1 U4736 ( .A(n4098), .B(n4097), .ZN(n4264) );
  NAND2_X1 U4737 ( .A1(n4264), .A2(n4171), .ZN(n4111) );
  OAI21_X1 U4738 ( .B1(n4117), .B2(n4100), .A(n4099), .ZN(n4342) );
  INV_X1 U4739 ( .A(n4342), .ZN(n4109) );
  NAND2_X1 U4740 ( .A1(n4101), .A2(n4258), .ZN(n4103) );
  NAND2_X1 U4741 ( .A1(n4229), .A2(REG2_REG_25__SCAN_IN), .ZN(n4102) );
  OAI211_X1 U4742 ( .C1(n4104), .C2(n4490), .A(n4103), .B(n4102), .ZN(n4108)
         );
  OAI22_X1 U4743 ( .A1(n4262), .A2(n4106), .B1(n4134), .B2(n4105), .ZN(n4107)
         );
  AOI211_X1 U4744 ( .C1(n4109), .C2(n4497), .A(n4108), .B(n4107), .ZN(n4110)
         );
  OAI211_X1 U4745 ( .C1(n4229), .C2(n4261), .A(n4111), .B(n4110), .ZN(U3265)
         );
  INV_X1 U4746 ( .A(n4116), .ZN(n4112) );
  XNOR2_X1 U4747 ( .A(n4113), .B(n4112), .ZN(n4114) );
  NAND2_X1 U4748 ( .A1(n4114), .A2(n4197), .ZN(n4271) );
  XOR2_X1 U4749 ( .A(n4116), .B(n4115), .Z(n4274) );
  NAND2_X1 U4750 ( .A1(n4274), .A2(n4171), .ZN(n4126) );
  INV_X1 U4751 ( .A(n4117), .ZN(n4118) );
  OAI21_X1 U4752 ( .B1(n4140), .B2(n4267), .A(n4118), .ZN(n4346) );
  INV_X1 U4753 ( .A(n4346), .ZN(n4124) );
  AOI22_X1 U4754 ( .A1(n4119), .A2(n4175), .B1(n4174), .B2(n4269), .ZN(n4122)
         );
  AOI22_X1 U4755 ( .A1(n4120), .A2(n4227), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4229), .ZN(n4121) );
  OAI211_X1 U4756 ( .C1(n4267), .C2(n4180), .A(n4122), .B(n4121), .ZN(n4123)
         );
  AOI21_X1 U4757 ( .B1(n4124), .B2(n4497), .A(n4123), .ZN(n4125) );
  OAI211_X1 U4758 ( .C1(n4229), .C2(n4271), .A(n4126), .B(n4125), .ZN(U3266)
         );
  XOR2_X1 U4759 ( .A(n4132), .B(n4127), .Z(n4278) );
  INV_X1 U4760 ( .A(n4278), .ZN(n4146) );
  INV_X1 U4761 ( .A(n4128), .ZN(n4130) );
  AOI21_X1 U4762 ( .B1(n4167), .B2(n4130), .A(n4129), .ZN(n4148) );
  INV_X1 U4763 ( .A(n4157), .ZN(n4147) );
  OAI21_X1 U4764 ( .B1(n4148), .B2(n4147), .A(n4131), .ZN(n4133) );
  XNOR2_X1 U4765 ( .A(n4133), .B(n4132), .ZN(n4137) );
  OAI22_X1 U4766 ( .A1(n4134), .A2(n4291), .B1(n4138), .B2(n4244), .ZN(n4135)
         );
  AOI21_X1 U4767 ( .B1(n4287), .B2(n4176), .A(n4135), .ZN(n4136) );
  OAI21_X1 U4768 ( .B1(n4137), .B2(n4222), .A(n4136), .ZN(n4277) );
  NOR2_X1 U4769 ( .A1(n4158), .A2(n4138), .ZN(n4139) );
  OR2_X1 U4770 ( .A1(n4140), .A2(n4139), .ZN(n4350) );
  INV_X1 U4771 ( .A(n4141), .ZN(n4142) );
  AOI22_X1 U4772 ( .A1(n4142), .A2(n4227), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4229), .ZN(n4143) );
  OAI21_X1 U4773 ( .B1(n4350), .B2(n4231), .A(n4143), .ZN(n4144) );
  AOI21_X1 U4774 ( .B1(n4277), .B2(n4493), .A(n4144), .ZN(n4145) );
  OAI21_X1 U4775 ( .B1(n4146), .B2(n4234), .A(n4145), .ZN(U3267) );
  XNOR2_X1 U4776 ( .A(n4148), .B(n4147), .ZN(n4153) );
  NOR2_X1 U4777 ( .A1(n4160), .A2(n4244), .ZN(n4149) );
  AOI21_X1 U4778 ( .B1(n4193), .B2(n4287), .A(n4149), .ZN(n4150) );
  OAI21_X1 U4779 ( .B1(n4151), .B2(n4291), .A(n4150), .ZN(n4152) );
  AOI21_X1 U4780 ( .B1(n4153), .B2(n4197), .A(n4152), .ZN(n4282) );
  NAND2_X1 U4781 ( .A1(n4156), .A2(n4157), .ZN(n4281) );
  NAND3_X1 U4782 ( .A1(n4155), .A2(n4281), .A3(n4171), .ZN(n4166) );
  INV_X1 U4783 ( .A(n4172), .ZN(n4161) );
  INV_X1 U4784 ( .A(n4158), .ZN(n4159) );
  OAI21_X1 U4785 ( .B1(n4161), .B2(n4160), .A(n4159), .ZN(n4354) );
  AOI22_X1 U4786 ( .A1(n4162), .A2(n4227), .B1(n4229), .B2(
        REG2_REG_22__SCAN_IN), .ZN(n4163) );
  OAI21_X1 U4787 ( .B1(n4354), .B2(n4231), .A(n4163), .ZN(n4164) );
  INV_X1 U4788 ( .A(n4164), .ZN(n4165) );
  OAI211_X1 U4789 ( .C1(n4229), .C2(n4282), .A(n4166), .B(n4165), .ZN(U3268)
         );
  XNOR2_X1 U4790 ( .A(n4167), .B(n4170), .ZN(n4168) );
  NAND2_X1 U4791 ( .A1(n4168), .A2(n4197), .ZN(n4290) );
  XOR2_X1 U4792 ( .A(n4170), .B(n4169), .Z(n4294) );
  NAND2_X1 U4793 ( .A1(n4294), .A2(n4171), .ZN(n4185) );
  INV_X1 U4794 ( .A(n4201), .ZN(n4173) );
  OAI21_X1 U4795 ( .B1(n4173), .B2(n4181), .A(n4172), .ZN(n4358) );
  INV_X1 U4796 ( .A(n4358), .ZN(n4183) );
  AOI22_X1 U4797 ( .A1(n4176), .A2(n4175), .B1(n4174), .B2(n4288), .ZN(n4179)
         );
  AOI22_X1 U4798 ( .A1(REG2_REG_21__SCAN_IN), .A2(n4229), .B1(n4177), .B2(
        n4227), .ZN(n4178) );
  OAI211_X1 U4799 ( .C1(n4181), .C2(n4180), .A(n4179), .B(n4178), .ZN(n4182)
         );
  AOI21_X1 U4800 ( .B1(n4183), .B2(n4497), .A(n4182), .ZN(n4184) );
  OAI211_X1 U4801 ( .C1(n4229), .C2(n4290), .A(n4185), .B(n4184), .ZN(U3269)
         );
  XNOR2_X1 U4802 ( .A(n4186), .B(n4190), .ZN(n4297) );
  INV_X1 U4803 ( .A(n4187), .ZN(n4188) );
  NAND2_X1 U4804 ( .A1(n4189), .A2(n4188), .ZN(n4191) );
  XNOR2_X1 U4805 ( .A(n4191), .B(n4190), .ZN(n4198) );
  AOI22_X1 U4806 ( .A1(n4193), .A2(n4311), .B1(n4310), .B2(n4192), .ZN(n4194)
         );
  OAI21_X1 U4807 ( .B1(n4195), .B2(n4314), .A(n4194), .ZN(n4196) );
  AOI21_X1 U4808 ( .B1(n4198), .B2(n4197), .A(n4196), .ZN(n4199) );
  OAI21_X1 U4809 ( .B1(n4297), .B2(n4200), .A(n4199), .ZN(n4298) );
  NAND2_X1 U4810 ( .A1(n4298), .A2(n4493), .ZN(n4209) );
  INV_X1 U4811 ( .A(n4224), .ZN(n4203) );
  OAI21_X1 U4812 ( .B1(n4203), .B2(n4202), .A(n4201), .ZN(n4363) );
  INV_X1 U4813 ( .A(n4363), .ZN(n4207) );
  INV_X1 U4814 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4205) );
  OAI22_X1 U4815 ( .A1(n4493), .A2(n4205), .B1(n4204), .B2(n4490), .ZN(n4206)
         );
  AOI21_X1 U4816 ( .B1(n4207), .B2(n4497), .A(n4206), .ZN(n4208) );
  OAI211_X1 U4817 ( .C1(n4297), .C2(n4210), .A(n4209), .B(n4208), .ZN(U3270)
         );
  XNOR2_X1 U4818 ( .A(n4211), .B(n4217), .ZN(n4303) );
  INV_X1 U4819 ( .A(n4303), .ZN(n4235) );
  INV_X1 U4820 ( .A(n4212), .ZN(n4214) );
  OAI21_X1 U4821 ( .B1(n4215), .B2(n4214), .A(n4213), .ZN(n4216) );
  XOR2_X1 U4822 ( .A(n4217), .B(n4216), .Z(n4223) );
  OAI22_X1 U4823 ( .A1(n4218), .A2(n4291), .B1(n4244), .B2(n4225), .ZN(n4219)
         );
  AOI21_X1 U4824 ( .B1(n4287), .B2(n4220), .A(n4219), .ZN(n4221) );
  OAI21_X1 U4825 ( .B1(n4223), .B2(n4222), .A(n4221), .ZN(n4302) );
  OAI21_X1 U4826 ( .B1(n4226), .B2(n4225), .A(n4224), .ZN(n4367) );
  AOI22_X1 U4827 ( .A1(n4229), .A2(REG2_REG_19__SCAN_IN), .B1(n4228), .B2(
        n4227), .ZN(n4230) );
  OAI21_X1 U4828 ( .B1(n4367), .B2(n4231), .A(n4230), .ZN(n4232) );
  AOI21_X1 U4829 ( .B1(n4302), .B2(n4493), .A(n4232), .ZN(n4233) );
  OAI21_X1 U4830 ( .B1(n4235), .B2(n4234), .A(n4233), .ZN(U3271) );
  NAND2_X1 U4831 ( .A1(n4323), .A2(n4543), .ZN(n4237) );
  NAND2_X1 U4832 ( .A1(n4540), .A2(REG1_REG_31__SCAN_IN), .ZN(n4236) );
  OAI211_X1 U4833 ( .C1(n4326), .C2(n4305), .A(n4237), .B(n4236), .ZN(U3549)
         );
  AOI21_X1 U4834 ( .B1(n4242), .B2(n4239), .A(n4238), .ZN(n4383) );
  INV_X1 U4835 ( .A(n4383), .ZN(n4329) );
  INV_X1 U4836 ( .A(n4240), .ZN(n4241) );
  AOI21_X1 U4837 ( .B1(n4242), .B2(n4310), .A(n4241), .ZN(n4385) );
  MUX2_X1 U4838 ( .A(n2709), .B(n4385), .S(n4543), .Z(n4243) );
  OAI21_X1 U4839 ( .B1(n4329), .B2(n4305), .A(n4243), .ZN(U3548) );
  OAI22_X1 U4840 ( .A1(n4262), .A2(n4314), .B1(n4245), .B2(n4244), .ZN(n4246)
         );
  AOI21_X1 U4841 ( .B1(n4247), .B2(n4311), .A(n4246), .ZN(n4249) );
  OAI211_X1 U4842 ( .C1(n4250), .C2(n4321), .A(n4249), .B(n4248), .ZN(n4330)
         );
  MUX2_X1 U4843 ( .A(REG1_REG_27__SCAN_IN), .B(n4330), .S(n4543), .Z(n4251) );
  AOI21_X1 U4844 ( .B1(n4252), .B2(n4333), .A(n4251), .ZN(n4253) );
  INV_X1 U4845 ( .A(n4253), .ZN(U3545) );
  AOI21_X1 U4846 ( .B1(n4255), .B2(n4527), .A(n4254), .ZN(n4335) );
  MUX2_X1 U4847 ( .A(n4256), .B(n4335), .S(n4543), .Z(n4257) );
  OAI21_X1 U4848 ( .B1(n4305), .B2(n4338), .A(n4257), .ZN(U3544) );
  AOI22_X1 U4849 ( .A1(n4259), .A2(n4287), .B1(n4258), .B2(n4310), .ZN(n4260)
         );
  OAI211_X1 U4850 ( .C1(n4262), .C2(n4291), .A(n4261), .B(n4260), .ZN(n4263)
         );
  AOI21_X1 U4851 ( .B1(n4264), .B2(n4527), .A(n4263), .ZN(n4339) );
  MUX2_X1 U4852 ( .A(n4265), .B(n4339), .S(n4543), .Z(n4266) );
  OAI21_X1 U4853 ( .B1(n4305), .B2(n4342), .A(n4266), .ZN(U3543) );
  INV_X1 U4854 ( .A(n4267), .ZN(n4268) );
  AOI22_X1 U4855 ( .A1(n4269), .A2(n4287), .B1(n4310), .B2(n4268), .ZN(n4270)
         );
  OAI211_X1 U4856 ( .C1(n4272), .C2(n4291), .A(n4271), .B(n4270), .ZN(n4273)
         );
  AOI21_X1 U4857 ( .B1(n4274), .B2(n4527), .A(n4273), .ZN(n4343) );
  MUX2_X1 U4858 ( .A(n4275), .B(n4343), .S(n4543), .Z(n4276) );
  OAI21_X1 U4859 ( .B1(n4305), .B2(n4346), .A(n4276), .ZN(U3542) );
  AOI21_X1 U4860 ( .B1(n4278), .B2(n4527), .A(n4277), .ZN(n4347) );
  MUX2_X1 U4861 ( .A(n4279), .B(n4347), .S(n4543), .Z(n4280) );
  OAI21_X1 U4862 ( .B1(n4305), .B2(n4350), .A(n4280), .ZN(U3541) );
  NAND3_X1 U4863 ( .A1(n4155), .A2(n4281), .A3(n4527), .ZN(n4283) );
  AND2_X1 U4864 ( .A1(n4283), .A2(n4282), .ZN(n4351) );
  MUX2_X1 U4865 ( .A(n4284), .B(n4351), .S(n4543), .Z(n4285) );
  OAI21_X1 U4866 ( .B1(n4305), .B2(n4354), .A(n4285), .ZN(U3540) );
  INV_X1 U4867 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4295) );
  AOI22_X1 U4868 ( .A1(n4288), .A2(n4287), .B1(n4286), .B2(n4310), .ZN(n4289)
         );
  OAI211_X1 U4869 ( .C1(n4292), .C2(n4291), .A(n4290), .B(n4289), .ZN(n4293)
         );
  AOI21_X1 U4870 ( .B1(n4294), .B2(n4527), .A(n4293), .ZN(n4355) );
  MUX2_X1 U4871 ( .A(n4295), .B(n4355), .S(n4543), .Z(n4296) );
  OAI21_X1 U4872 ( .B1(n4305), .B2(n4358), .A(n4296), .ZN(U3539) );
  INV_X1 U4873 ( .A(n4297), .ZN(n4299) );
  AOI21_X1 U4874 ( .B1(n4524), .B2(n4299), .A(n4298), .ZN(n4359) );
  MUX2_X1 U4875 ( .A(n4300), .B(n4359), .S(n4543), .Z(n4301) );
  OAI21_X1 U4876 ( .B1(n4305), .B2(n4363), .A(n4301), .ZN(U3538) );
  AOI21_X1 U4877 ( .B1(n4303), .B2(n4527), .A(n4302), .ZN(n4364) );
  MUX2_X1 U4878 ( .A(n4047), .B(n4364), .S(n4543), .Z(n4304) );
  OAI21_X1 U4879 ( .B1(n4305), .B2(n4367), .A(n4304), .ZN(U3537) );
  OAI211_X1 U4880 ( .C1(n4308), .C2(n4321), .A(n4307), .B(n4306), .ZN(n4368)
         );
  MUX2_X1 U4881 ( .A(REG1_REG_18__SCAN_IN), .B(n4368), .S(n4543), .Z(U3536) );
  AOI22_X1 U4882 ( .A1(n4312), .A2(n4311), .B1(n4310), .B2(n4309), .ZN(n4313)
         );
  OAI21_X1 U4883 ( .B1(n4315), .B2(n4314), .A(n4313), .ZN(n4316) );
  AOI21_X1 U4884 ( .B1(n4318), .B2(n4317), .A(n4316), .ZN(n4320) );
  OAI211_X1 U4885 ( .C1(n4322), .C2(n4321), .A(n4320), .B(n4319), .ZN(n4369)
         );
  MUX2_X1 U4886 ( .A(REG1_REG_16__SCAN_IN), .B(n4369), .S(n4543), .Z(U3534) );
  NAND2_X1 U4887 ( .A1(n4323), .A2(n4536), .ZN(n4325) );
  NAND2_X1 U4888 ( .A1(n4534), .A2(REG0_REG_31__SCAN_IN), .ZN(n4324) );
  OAI211_X1 U4889 ( .C1(n4326), .C2(n4362), .A(n4325), .B(n4324), .ZN(U3517)
         );
  INV_X1 U4890 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4327) );
  MUX2_X1 U4891 ( .A(n4327), .B(n4385), .S(n4536), .Z(n4328) );
  OAI21_X1 U4892 ( .B1(n4329), .B2(n4362), .A(n4328), .ZN(U3516) );
  MUX2_X1 U4893 ( .A(REG0_REG_27__SCAN_IN), .B(n4330), .S(n4536), .Z(n4331) );
  AOI21_X1 U4894 ( .B1(n4333), .B2(n4332), .A(n4331), .ZN(n4334) );
  INV_X1 U4895 ( .A(n4334), .ZN(U3513) );
  INV_X1 U4896 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4336) );
  MUX2_X1 U4897 ( .A(n4336), .B(n4335), .S(n4536), .Z(n4337) );
  OAI21_X1 U4898 ( .B1(n4338), .B2(n4362), .A(n4337), .ZN(U3512) );
  INV_X1 U4899 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4340) );
  MUX2_X1 U4900 ( .A(n4340), .B(n4339), .S(n4536), .Z(n4341) );
  OAI21_X1 U4901 ( .B1(n4342), .B2(n4362), .A(n4341), .ZN(U3511) );
  INV_X1 U4902 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4344) );
  MUX2_X1 U4903 ( .A(n4344), .B(n4343), .S(n4536), .Z(n4345) );
  OAI21_X1 U4904 ( .B1(n4346), .B2(n4362), .A(n4345), .ZN(U3510) );
  INV_X1 U4905 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4348) );
  MUX2_X1 U4906 ( .A(n4348), .B(n4347), .S(n4536), .Z(n4349) );
  OAI21_X1 U4907 ( .B1(n4350), .B2(n4362), .A(n4349), .ZN(U3509) );
  INV_X1 U4908 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4352) );
  MUX2_X1 U4909 ( .A(n4352), .B(n4351), .S(n4536), .Z(n4353) );
  OAI21_X1 U4910 ( .B1(n4354), .B2(n4362), .A(n4353), .ZN(U3508) );
  INV_X1 U4911 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4356) );
  MUX2_X1 U4912 ( .A(n4356), .B(n4355), .S(n4536), .Z(n4357) );
  OAI21_X1 U4913 ( .B1(n4358), .B2(n4362), .A(n4357), .ZN(U3507) );
  INV_X1 U4914 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4360) );
  MUX2_X1 U4915 ( .A(n4360), .B(n4359), .S(n4536), .Z(n4361) );
  OAI21_X1 U4916 ( .B1(n4363), .B2(n4362), .A(n4361), .ZN(U3506) );
  INV_X1 U4917 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4365) );
  MUX2_X1 U4918 ( .A(n4365), .B(n4364), .S(n4536), .Z(n4366) );
  OAI21_X1 U4919 ( .B1(n4367), .B2(n4362), .A(n4366), .ZN(U3505) );
  MUX2_X1 U4920 ( .A(REG0_REG_18__SCAN_IN), .B(n4368), .S(n4536), .Z(U3503) );
  MUX2_X1 U4921 ( .A(REG0_REG_16__SCAN_IN), .B(n4369), .S(n4536), .Z(U3499) );
  MUX2_X1 U4922 ( .A(n4370), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U4923 ( .A(DATAI_25_), .B(n4371), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U4924 ( .A(DATAI_22_), .B(n4372), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4925 ( .A(n4373), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4926 ( .A(n4374), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4927 ( .A(DATAI_8_), .B(n4375), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4928 ( .A(n4376), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4929 ( .A(n4377), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4930 ( .A(n4378), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4931 ( .A(n4379), .B(DATAI_4_), .S(U3149), .Z(U3348) );
  MUX2_X1 U4932 ( .A(n4380), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4933 ( .A(n4381), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4934 ( .A(n4382), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4935 ( .A1(n4383), .A2(n4497), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4229), .ZN(n4384) );
  OAI21_X1 U4936 ( .B1(n4229), .B2(n4385), .A(n4384), .ZN(U3261) );
  OAI211_X1 U4937 ( .C1(n4388), .C2(n4387), .A(n4484), .B(n4386), .ZN(n4393)
         );
  OAI211_X1 U4938 ( .C1(n4391), .C2(n4390), .A(n4429), .B(n4389), .ZN(n4392)
         );
  OAI211_X1 U4939 ( .C1(n4489), .C2(n4516), .A(n4393), .B(n4392), .ZN(n4394)
         );
  AOI211_X1 U4940 ( .C1(n4482), .C2(ADDR_REG_9__SCAN_IN), .A(n4395), .B(n4394), 
        .ZN(n4396) );
  INV_X1 U4941 ( .A(n4396), .ZN(U3249) );
  OAI211_X1 U4942 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4398), .A(n4429), .B(n4397), .ZN(n4400) );
  NAND2_X1 U4943 ( .A1(n4400), .A2(n4399), .ZN(n4401) );
  AOI21_X1 U4944 ( .B1(n4482), .B2(ADDR_REG_10__SCAN_IN), .A(n4401), .ZN(n4405) );
  OAI211_X1 U4945 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4403), .A(n4484), .B(n4402), .ZN(n4404) );
  OAI211_X1 U4946 ( .C1(n4489), .C2(n4406), .A(n4405), .B(n4404), .ZN(U3250)
         );
  OAI211_X1 U4947 ( .C1(n4409), .C2(n4408), .A(n4484), .B(n4407), .ZN(n4414)
         );
  OAI211_X1 U4948 ( .C1(n4412), .C2(n4411), .A(n4429), .B(n4410), .ZN(n4413)
         );
  OAI211_X1 U4949 ( .C1(n4489), .C2(n4512), .A(n4414), .B(n4413), .ZN(n4415)
         );
  AOI211_X1 U4950 ( .C1(n4482), .C2(ADDR_REG_11__SCAN_IN), .A(n4416), .B(n4415), .ZN(n4417) );
  INV_X1 U4951 ( .A(n4417), .ZN(U3251) );
  OAI211_X1 U4952 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4419), .A(n4429), .B(n4418), .ZN(n4421) );
  NAND2_X1 U4953 ( .A1(n4421), .A2(n4420), .ZN(n4422) );
  AOI21_X1 U4954 ( .B1(n4482), .B2(ADDR_REG_12__SCAN_IN), .A(n4422), .ZN(n4426) );
  OAI211_X1 U4955 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4424), .A(n4484), .B(n4423), .ZN(n4425) );
  OAI211_X1 U4956 ( .C1(n4489), .C2(n4510), .A(n4426), .B(n4425), .ZN(U3252)
         );
  AOI21_X1 U4957 ( .B1(n4428), .B2(n4509), .A(n4427), .ZN(n4432) );
  OAI21_X1 U4958 ( .B1(n4432), .B2(n4431), .A(n4429), .ZN(n4430) );
  AOI21_X1 U4959 ( .B1(n4432), .B2(n4431), .A(n4430), .ZN(n4434) );
  AOI211_X1 U4960 ( .C1(n4482), .C2(ADDR_REG_13__SCAN_IN), .A(n4434), .B(n4433), .ZN(n4439) );
  OAI211_X1 U4961 ( .C1(n4437), .C2(n4436), .A(n4484), .B(n4435), .ZN(n4438)
         );
  OAI211_X1 U4962 ( .C1(n4489), .C2(n4509), .A(n4439), .B(n4438), .ZN(U3253)
         );
  AOI211_X1 U4963 ( .C1(n4442), .C2(n4441), .A(n4440), .B(n4478), .ZN(n4443)
         );
  AOI211_X1 U4964 ( .C1(n4482), .C2(ADDR_REG_14__SCAN_IN), .A(n4444), .B(n4443), .ZN(n4448) );
  OAI211_X1 U4965 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4446), .A(n4484), .B(n4445), .ZN(n4447) );
  OAI211_X1 U4966 ( .C1(n4489), .C2(n2180), .A(n4448), .B(n4447), .ZN(U3254)
         );
  AOI211_X1 U4967 ( .C1(n4451), .C2(n4450), .A(n4449), .B(n4478), .ZN(n4452)
         );
  AOI211_X1 U4968 ( .C1(n4482), .C2(ADDR_REG_15__SCAN_IN), .A(n4453), .B(n4452), .ZN(n4458) );
  OAI211_X1 U4969 ( .C1(n4456), .C2(n4455), .A(n4484), .B(n4454), .ZN(n4457)
         );
  OAI211_X1 U4970 ( .C1(n4489), .C2(n4508), .A(n4458), .B(n4457), .ZN(U3255)
         );
  AOI221_X1 U4971 ( .B1(n4461), .B2(n4460), .C1(n4459), .C2(n4460), .A(n4478), 
        .ZN(n4462) );
  AOI211_X1 U4972 ( .C1(n4482), .C2(ADDR_REG_16__SCAN_IN), .A(n4463), .B(n4462), .ZN(n4467) );
  OAI221_X1 U4973 ( .B1(n4465), .B2(REG1_REG_16__SCAN_IN), .C1(n4465), .C2(
        n4464), .A(n4484), .ZN(n4466) );
  OAI211_X1 U4974 ( .C1(n4489), .C2(n4507), .A(n4467), .B(n4466), .ZN(U3256)
         );
  AOI221_X1 U4975 ( .B1(n4470), .B2(n4469), .C1(n4468), .C2(n4469), .A(n4478), 
        .ZN(n4471) );
  AOI211_X1 U4976 ( .C1(n4482), .C2(ADDR_REG_17__SCAN_IN), .A(n4472), .B(n4471), .ZN(n4477) );
  OAI221_X1 U4977 ( .B1(n4475), .B2(n4474), .C1(n4475), .C2(n4473), .A(n4484), 
        .ZN(n4476) );
  OAI211_X1 U4978 ( .C1(n4489), .C2(n4506), .A(n4477), .B(n4476), .ZN(U3257)
         );
  OAI211_X1 U4979 ( .C1(n4486), .C2(n4485), .A(n4484), .B(n4483), .ZN(n4487)
         );
  OAI211_X1 U4980 ( .C1(n4489), .C2(n4505), .A(n4488), .B(n4487), .ZN(U3258)
         );
  OAI22_X1 U4981 ( .A1(n4493), .A2(n4492), .B1(n4491), .B2(n4490), .ZN(n4494)
         );
  INV_X1 U4982 ( .A(n4494), .ZN(n4501) );
  INV_X1 U4983 ( .A(n4495), .ZN(n4496) );
  AOI22_X1 U4984 ( .A1(n4499), .A2(n4498), .B1(n4497), .B2(n4496), .ZN(n4500)
         );
  OAI211_X1 U4985 ( .C1(n4229), .C2(n4502), .A(n4501), .B(n4500), .ZN(U3282)
         );
  AND2_X1 U4986 ( .A1(D_REG_31__SCAN_IN), .A2(n4503), .ZN(U3291) );
  AND2_X1 U4987 ( .A1(D_REG_30__SCAN_IN), .A2(n4503), .ZN(U3292) );
  AND2_X1 U4988 ( .A1(D_REG_29__SCAN_IN), .A2(n4503), .ZN(U3293) );
  AND2_X1 U4989 ( .A1(D_REG_28__SCAN_IN), .A2(n4503), .ZN(U3294) );
  AND2_X1 U4990 ( .A1(D_REG_27__SCAN_IN), .A2(n4503), .ZN(U3295) );
  AND2_X1 U4991 ( .A1(D_REG_26__SCAN_IN), .A2(n4503), .ZN(U3296) );
  AND2_X1 U4992 ( .A1(D_REG_25__SCAN_IN), .A2(n4503), .ZN(U3297) );
  AND2_X1 U4993 ( .A1(D_REG_24__SCAN_IN), .A2(n4503), .ZN(U3298) );
  AND2_X1 U4994 ( .A1(D_REG_23__SCAN_IN), .A2(n4503), .ZN(U3299) );
  AND2_X1 U4995 ( .A1(D_REG_22__SCAN_IN), .A2(n4503), .ZN(U3300) );
  AND2_X1 U4996 ( .A1(D_REG_21__SCAN_IN), .A2(n4503), .ZN(U3301) );
  AND2_X1 U4997 ( .A1(D_REG_20__SCAN_IN), .A2(n4503), .ZN(U3302) );
  AND2_X1 U4998 ( .A1(D_REG_19__SCAN_IN), .A2(n4503), .ZN(U3303) );
  AND2_X1 U4999 ( .A1(D_REG_18__SCAN_IN), .A2(n4503), .ZN(U3304) );
  AND2_X1 U5000 ( .A1(D_REG_17__SCAN_IN), .A2(n4503), .ZN(U3305) );
  AND2_X1 U5001 ( .A1(D_REG_16__SCAN_IN), .A2(n4503), .ZN(U3306) );
  AND2_X1 U5002 ( .A1(D_REG_15__SCAN_IN), .A2(n4503), .ZN(U3307) );
  AND2_X1 U5003 ( .A1(D_REG_14__SCAN_IN), .A2(n4503), .ZN(U3308) );
  AND2_X1 U5004 ( .A1(D_REG_13__SCAN_IN), .A2(n4503), .ZN(U3309) );
  AND2_X1 U5005 ( .A1(D_REG_12__SCAN_IN), .A2(n4503), .ZN(U3310) );
  AND2_X1 U5006 ( .A1(D_REG_11__SCAN_IN), .A2(n4503), .ZN(U3311) );
  AND2_X1 U5007 ( .A1(D_REG_10__SCAN_IN), .A2(n4503), .ZN(U3312) );
  AND2_X1 U5008 ( .A1(D_REG_9__SCAN_IN), .A2(n4503), .ZN(U3313) );
  AND2_X1 U5009 ( .A1(D_REG_8__SCAN_IN), .A2(n4503), .ZN(U3314) );
  AND2_X1 U5010 ( .A1(D_REG_7__SCAN_IN), .A2(n4503), .ZN(U3315) );
  AND2_X1 U5011 ( .A1(D_REG_6__SCAN_IN), .A2(n4503), .ZN(U3316) );
  AND2_X1 U5012 ( .A1(D_REG_5__SCAN_IN), .A2(n4503), .ZN(U3317) );
  AND2_X1 U5013 ( .A1(D_REG_4__SCAN_IN), .A2(n4503), .ZN(U3318) );
  AND2_X1 U5014 ( .A1(D_REG_3__SCAN_IN), .A2(n4503), .ZN(U3319) );
  AND2_X1 U5015 ( .A1(D_REG_2__SCAN_IN), .A2(n4503), .ZN(U3320) );
  INV_X1 U5016 ( .A(DATAI_23_), .ZN(n4647) );
  AOI21_X1 U5017 ( .B1(U3149), .B2(n4647), .A(n4504), .ZN(U3329) );
  INV_X1 U5018 ( .A(DATAI_18_), .ZN(n4553) );
  AOI22_X1 U5019 ( .A1(STATE_REG_SCAN_IN), .A2(n4505), .B1(n4553), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5020 ( .A(DATAI_17_), .ZN(n4706) );
  AOI22_X1 U5021 ( .A1(STATE_REG_SCAN_IN), .A2(n4506), .B1(n4706), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5022 ( .A(DATAI_16_), .ZN(n4619) );
  AOI22_X1 U5023 ( .A1(STATE_REG_SCAN_IN), .A2(n4507), .B1(n4619), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5024 ( .A(DATAI_15_), .ZN(n4654) );
  AOI22_X1 U5025 ( .A1(STATE_REG_SCAN_IN), .A2(n4508), .B1(n4654), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5026 ( .A(DATAI_14_), .ZN(n4582) );
  AOI22_X1 U5027 ( .A1(STATE_REG_SCAN_IN), .A2(n2180), .B1(n4582), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5028 ( .A1(STATE_REG_SCAN_IN), .A2(n4509), .B1(n2456), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5029 ( .A1(STATE_REG_SCAN_IN), .A2(n4510), .B1(n2449), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5030 ( .A(DATAI_11_), .ZN(n4511) );
  AOI22_X1 U5031 ( .A1(STATE_REG_SCAN_IN), .A2(n4512), .B1(n4511), .B2(U3149), 
        .ZN(U3341) );
  OAI22_X1 U5032 ( .A1(U3149), .A2(n4513), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4514) );
  INV_X1 U5033 ( .A(n4514), .ZN(U3342) );
  INV_X1 U5034 ( .A(DATAI_9_), .ZN(n4515) );
  AOI22_X1 U5035 ( .A1(STATE_REG_SCAN_IN), .A2(n4516), .B1(n4515), .B2(U3149), 
        .ZN(U3343) );
  AOI211_X1 U5036 ( .C1(n4524), .C2(n4519), .A(n4518), .B(n4517), .ZN(n4537)
         );
  INV_X1 U5037 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4520) );
  AOI22_X1 U5038 ( .A1(n4536), .A2(n4537), .B1(n4520), .B2(n4534), .ZN(U3467)
         );
  INV_X1 U5039 ( .A(n4521), .ZN(n4523) );
  AOI211_X1 U5040 ( .C1(n4525), .C2(n4524), .A(n4523), .B(n4522), .ZN(n4539)
         );
  INV_X1 U5041 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4526) );
  AOI22_X1 U5042 ( .A1(n4536), .A2(n4539), .B1(n4526), .B2(n4534), .ZN(U3475)
         );
  NAND2_X1 U5043 ( .A1(n4528), .A2(n4527), .ZN(n4530) );
  OAI21_X1 U5044 ( .B1(n3095), .B2(n4530), .A(n4529), .ZN(n4531) );
  INV_X1 U5045 ( .A(n4531), .ZN(n4533) );
  AND2_X1 U5046 ( .A1(n4533), .A2(n4532), .ZN(n4542) );
  INV_X1 U5047 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4535) );
  AOI22_X1 U5048 ( .A1(n4536), .A2(n4542), .B1(n4535), .B2(n4534), .ZN(U3481)
         );
  AOI22_X1 U5049 ( .A1(n4543), .A2(n4537), .B1(n2333), .B2(n4540), .ZN(U3518)
         );
  INV_X1 U5050 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4538) );
  AOI22_X1 U5051 ( .A1(n4543), .A2(n4539), .B1(n4538), .B2(n4540), .ZN(U3522)
         );
  AOI22_X1 U5052 ( .A1(n4543), .A2(n4542), .B1(n4541), .B2(n4540), .ZN(U3525)
         );
  INV_X1 U5053 ( .A(keyinput_g53), .ZN(n4726) );
  AOI22_X1 U5054 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(DATAI_29_), .B2(
        keyinput_f2), .ZN(n4544) );
  OAI221_X1 U5055 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(DATAI_29_), .C2(
        keyinput_f2), .A(n4544), .ZN(n4551) );
  AOI22_X1 U5056 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(REG3_REG_28__SCAN_IN), 
        .B2(keyinput_f40), .ZN(n4545) );
  OAI221_X1 U5057 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(REG3_REG_28__SCAN_IN), .C2(keyinput_f40), .A(n4545), .ZN(n4550) );
  AOI22_X1 U5058 ( .A1(DATAI_15_), .A2(keyinput_f16), .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_f44), .ZN(n4546) );
  OAI221_X1 U5059 ( .B1(DATAI_15_), .B2(keyinput_f16), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_f44), .A(n4546), .ZN(n4549) );
  AOI22_X1 U5060 ( .A1(DATAI_17_), .A2(keyinput_f14), .B1(DATAI_19_), .B2(
        keyinput_f12), .ZN(n4547) );
  OAI221_X1 U5061 ( .B1(DATAI_17_), .B2(keyinput_f14), .C1(DATAI_19_), .C2(
        keyinput_f12), .A(n4547), .ZN(n4548) );
  NOR4_X1 U5062 ( .A1(n4551), .A2(n4550), .A3(n4549), .A4(n4548), .ZN(n4579)
         );
  XOR2_X1 U5063 ( .A(U3149), .B(keyinput_f32), .Z(n4559) );
  AOI22_X1 U5064 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(n4553), .B2(
        keyinput_f13), .ZN(n4552) );
  OAI221_X1 U5065 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(n4553), .C2(
        keyinput_f13), .A(n4552), .ZN(n4558) );
  AOI22_X1 U5066 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(DATAI_27_), .B2(
        keyinput_f4), .ZN(n4554) );
  OAI221_X1 U5067 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(DATAI_27_), .C2(
        keyinput_f4), .A(n4554), .ZN(n4557) );
  AOI22_X1 U5068 ( .A1(DATAI_2_), .A2(keyinput_f29), .B1(DATAI_26_), .B2(
        keyinput_f5), .ZN(n4555) );
  OAI221_X1 U5069 ( .B1(DATAI_2_), .B2(keyinput_f29), .C1(DATAI_26_), .C2(
        keyinput_f5), .A(n4555), .ZN(n4556) );
  NOR4_X1 U5070 ( .A1(n4559), .A2(n4558), .A3(n4557), .A4(n4556), .ZN(n4578)
         );
  AOI22_X1 U5071 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_f39), .B1(
        REG3_REG_27__SCAN_IN), .B2(keyinput_f34), .ZN(n4560) );
  OAI221_X1 U5072 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_f39), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_f34), .A(n4560), .ZN(n4567) );
  AOI22_X1 U5073 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(REG3_REG_9__SCAN_IN), 
        .B2(keyinput_f51), .ZN(n4561) );
  OAI221_X1 U5074 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(REG3_REG_9__SCAN_IN), 
        .C2(keyinput_f51), .A(n4561), .ZN(n4566) );
  AOI22_X1 U5075 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_f37), .ZN(n4562) );
  OAI221_X1 U5076 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(
        REG3_REG_10__SCAN_IN), .C2(keyinput_f37), .A(n4562), .ZN(n4565) );
  AOI22_X1 U5077 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_f46), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_f60), .ZN(n4563) );
  OAI221_X1 U5078 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_f46), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_f60), .A(n4563), .ZN(n4564) );
  NOR4_X1 U5079 ( .A1(n4567), .A2(n4566), .A3(n4565), .A4(n4564), .ZN(n4577)
         );
  AOI22_X1 U5080 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_f33), .B1(
        IR_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n4568) );
  OAI221_X1 U5081 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_f33), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n4568), .ZN(n4575) );
  AOI22_X1 U5082 ( .A1(DATAI_7_), .A2(keyinput_f24), .B1(DATAI_10_), .B2(
        keyinput_f21), .ZN(n4569) );
  OAI221_X1 U5083 ( .B1(DATAI_7_), .B2(keyinput_f24), .C1(DATAI_10_), .C2(
        keyinput_f21), .A(n4569), .ZN(n4574) );
  AOI22_X1 U5084 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(IR_REG_7__SCAN_IN), 
        .B2(keyinput_f62), .ZN(n4570) );
  OAI221_X1 U5085 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(IR_REG_7__SCAN_IN), 
        .C2(keyinput_f62), .A(n4570), .ZN(n4573) );
  AOI22_X1 U5086 ( .A1(DATAI_0_), .A2(keyinput_f31), .B1(IR_REG_3__SCAN_IN), 
        .B2(keyinput_f58), .ZN(n4571) );
  OAI221_X1 U5087 ( .B1(DATAI_0_), .B2(keyinput_f31), .C1(IR_REG_3__SCAN_IN), 
        .C2(keyinput_f58), .A(n4571), .ZN(n4572) );
  NOR4_X1 U5088 ( .A1(n4575), .A2(n4574), .A3(n4573), .A4(n4572), .ZN(n4576)
         );
  NAND4_X1 U5089 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(n4629)
         );
  AOI22_X1 U5090 ( .A1(n2494), .A2(keyinput_f48), .B1(keyinput_f19), .B2(n2449), .ZN(n4580) );
  OAI221_X1 U5091 ( .B1(n2494), .B2(keyinput_f48), .C1(n2449), .C2(
        keyinput_f19), .A(n4580), .ZN(n4589) );
  INV_X1 U5092 ( .A(DATAI_25_), .ZN(n4650) );
  AOI22_X1 U5093 ( .A1(n4650), .A2(keyinput_f6), .B1(keyinput_f17), .B2(n4582), 
        .ZN(n4581) );
  OAI221_X1 U5094 ( .B1(n4650), .B2(keyinput_f6), .C1(n4582), .C2(keyinput_f17), .A(n4581), .ZN(n4588) );
  XNOR2_X1 U5095 ( .A(DATAI_21_), .B(keyinput_f10), .ZN(n4586) );
  XNOR2_X1 U5096 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_f52), .ZN(n4584) );
  XNOR2_X1 U5097 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_f35), .ZN(n4583) );
  NAND4_X1 U5098 ( .A1(n4586), .A2(n4585), .A3(n4584), .A4(n4583), .ZN(n4587)
         );
  NOR3_X1 U5099 ( .A1(n4589), .A2(n4588), .A3(n4587), .ZN(n4627) );
  INV_X1 U5100 ( .A(DATAI_6_), .ZN(n4591) );
  AOI22_X1 U5101 ( .A1(n4592), .A2(keyinput_f3), .B1(keyinput_f25), .B2(n4591), 
        .ZN(n4590) );
  OAI221_X1 U5102 ( .B1(n4592), .B2(keyinput_f3), .C1(n4591), .C2(keyinput_f25), .A(n4590), .ZN(n4601) );
  INV_X1 U5103 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4691) );
  AOI22_X1 U5104 ( .A1(n2375), .A2(keyinput_f47), .B1(n4691), .B2(keyinput_f41), .ZN(n4593) );
  OAI221_X1 U5105 ( .B1(n2375), .B2(keyinput_f47), .C1(n4691), .C2(
        keyinput_f41), .A(n4593), .ZN(n4600) );
  AOI22_X1 U5106 ( .A1(DATAI_23_), .A2(keyinput_f8), .B1(n4595), .B2(
        keyinput_f45), .ZN(n4594) );
  OAI221_X1 U5107 ( .B1(DATAI_23_), .B2(keyinput_f8), .C1(n4595), .C2(
        keyinput_f45), .A(n4594), .ZN(n4599) );
  XOR2_X1 U5108 ( .A(n4651), .B(keyinput_f0), .Z(n4597) );
  XNOR2_X1 U5109 ( .A(DATAI_3_), .B(keyinput_f28), .ZN(n4596) );
  NAND2_X1 U5110 ( .A1(n4597), .A2(n4596), .ZN(n4598) );
  NOR4_X1 U5111 ( .A1(n4601), .A2(n4600), .A3(n4599), .A4(n4598), .ZN(n4626)
         );
  INV_X1 U5112 ( .A(DATAI_4_), .ZN(n4603) );
  AOI22_X1 U5113 ( .A1(n2457), .A2(keyinput_f54), .B1(keyinput_f27), .B2(n4603), .ZN(n4602) );
  OAI221_X1 U5114 ( .B1(n2457), .B2(keyinput_f54), .C1(n4603), .C2(
        keyinput_f27), .A(n4602), .ZN(n4611) );
  INV_X1 U5115 ( .A(DATAI_8_), .ZN(n4634) );
  XNOR2_X1 U5116 ( .A(keyinput_f23), .B(n4634), .ZN(n4610) );
  XNOR2_X1 U5117 ( .A(keyinput_f18), .B(n2456), .ZN(n4609) );
  XNOR2_X1 U5118 ( .A(DATAI_11_), .B(keyinput_f20), .ZN(n4607) );
  XNOR2_X1 U5119 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_f42), .ZN(n4606) );
  XNOR2_X1 U5120 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_f57), .ZN(n4605) );
  XNOR2_X1 U5121 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_f50), .ZN(n4604) );
  NAND4_X1 U5122 ( .A1(n4607), .A2(n4606), .A3(n4605), .A4(n4604), .ZN(n4608)
         );
  NOR4_X1 U5123 ( .A1(n4611), .A2(n4610), .A3(n4609), .A4(n4608), .ZN(n4625)
         );
  AOI22_X1 U5124 ( .A1(n4613), .A2(keyinput_f63), .B1(keyinput_f49), .B2(n4648), .ZN(n4612) );
  OAI221_X1 U5125 ( .B1(n4613), .B2(keyinput_f63), .C1(n4648), .C2(
        keyinput_f49), .A(n4612), .ZN(n4623) );
  XNOR2_X1 U5126 ( .A(n4614), .B(keyinput_f59), .ZN(n4622) );
  XNOR2_X1 U5127 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_f43), .ZN(n4618) );
  XNOR2_X1 U5128 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_f38), .ZN(n4617) );
  XNOR2_X1 U5129 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_f55), .ZN(n4616) );
  XNOR2_X1 U5130 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_f36), .ZN(n4615) );
  NAND4_X1 U5131 ( .A1(n4618), .A2(n4617), .A3(n4616), .A4(n4615), .ZN(n4621)
         );
  XNOR2_X1 U5132 ( .A(keyinput_f15), .B(n4619), .ZN(n4620) );
  NOR4_X1 U5133 ( .A1(n4623), .A2(n4622), .A3(n4621), .A4(n4620), .ZN(n4624)
         );
  NAND4_X1 U5134 ( .A1(n4627), .A2(n4626), .A3(n4625), .A4(n4624), .ZN(n4628)
         );
  OAI22_X1 U5135 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput_f53), .B1(n4629), 
        .B2(n4628), .ZN(n4630) );
  AOI222_X1 U5136 ( .A1(REG3_REG_20__SCAN_IN), .A2(n4630), .B1(
        REG3_REG_20__SCAN_IN), .B2(keyinput_f53), .C1(n4630), .C2(n4726), .ZN(
        n4725) );
  AOI22_X1 U5137 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_g54), .B1(
        REG3_REG_25__SCAN_IN), .B2(keyinput_g45), .ZN(n4631) );
  OAI221_X1 U5138 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_g54), .C1(
        REG3_REG_25__SCAN_IN), .C2(keyinput_g45), .A(n4631), .ZN(n4723) );
  AOI22_X1 U5139 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_g50), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput_g40), .ZN(n4632) );
  OAI221_X1 U5140 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_g50), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput_g40), .A(n4632), .ZN(n4722) );
  AOI22_X1 U5141 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_g42), .B1(n4634), 
        .B2(keyinput_g23), .ZN(n4633) );
  OAI221_X1 U5142 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_g42), .C1(n4634), 
        .C2(keyinput_g23), .A(n4633), .ZN(n4644) );
  OAI22_X1 U5143 ( .A1(DATAI_26_), .A2(keyinput_g5), .B1(keyinput_g29), .B2(
        DATAI_2_), .ZN(n4635) );
  AOI221_X1 U5144 ( .B1(DATAI_26_), .B2(keyinput_g5), .C1(DATAI_2_), .C2(
        keyinput_g29), .A(n4635), .ZN(n4642) );
  OAI22_X1 U5145 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput_g32), .B1(DATAI_1_), 
        .B2(keyinput_g30), .ZN(n4636) );
  AOI221_X1 U5146 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput_g32), .C1(
        keyinput_g30), .C2(DATAI_1_), .A(n4636), .ZN(n4641) );
  OAI22_X1 U5147 ( .A1(DATAI_29_), .A2(keyinput_g2), .B1(keyinput_g3), .B2(
        DATAI_28_), .ZN(n4637) );
  AOI221_X1 U5148 ( .B1(DATAI_29_), .B2(keyinput_g2), .C1(DATAI_28_), .C2(
        keyinput_g3), .A(n4637), .ZN(n4640) );
  OAI22_X1 U5149 ( .A1(DATAI_22_), .A2(keyinput_g9), .B1(DATAI_30_), .B2(
        keyinput_g1), .ZN(n4638) );
  AOI221_X1 U5150 ( .B1(DATAI_22_), .B2(keyinput_g9), .C1(keyinput_g1), .C2(
        DATAI_30_), .A(n4638), .ZN(n4639) );
  NAND4_X1 U5151 ( .A1(n4642), .A2(n4641), .A3(n4640), .A4(n4639), .ZN(n4643)
         );
  AOI211_X1 U5152 ( .C1(keyinput_g4), .C2(DATAI_27_), .A(n4644), .B(n4643), 
        .ZN(n4645) );
  OAI21_X1 U5153 ( .B1(keyinput_g4), .B2(DATAI_27_), .A(n4645), .ZN(n4721) );
  AOI22_X1 U5154 ( .A1(n4648), .A2(keyinput_g49), .B1(keyinput_g8), .B2(n4647), 
        .ZN(n4646) );
  OAI221_X1 U5155 ( .B1(n4648), .B2(keyinput_g49), .C1(n4647), .C2(keyinput_g8), .A(n4646), .ZN(n4660) );
  AOI22_X1 U5156 ( .A1(n4651), .A2(keyinput_g0), .B1(n4650), .B2(keyinput_g6), 
        .ZN(n4649) );
  OAI221_X1 U5157 ( .B1(n4651), .B2(keyinput_g0), .C1(n4650), .C2(keyinput_g6), 
        .A(n4649), .ZN(n4659) );
  AOI22_X1 U5158 ( .A1(n4654), .A2(keyinput_g16), .B1(n4653), .B2(keyinput_g46), .ZN(n4652) );
  OAI221_X1 U5159 ( .B1(n4654), .B2(keyinput_g16), .C1(n4653), .C2(
        keyinput_g46), .A(n4652), .ZN(n4658) );
  XNOR2_X1 U5160 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_g57), .ZN(n4656) );
  XNOR2_X1 U5161 ( .A(DATAI_19_), .B(keyinput_g12), .ZN(n4655) );
  NAND2_X1 U5162 ( .A1(n4656), .A2(n4655), .ZN(n4657) );
  NOR4_X1 U5163 ( .A1(n4660), .A2(n4659), .A3(n4658), .A4(n4657), .ZN(n4719)
         );
  AOI22_X1 U5164 ( .A1(n4662), .A2(keyinput_g44), .B1(keyinput_g51), .B2(n2306), .ZN(n4661) );
  OAI221_X1 U5165 ( .B1(n4662), .B2(keyinput_g44), .C1(n2306), .C2(
        keyinput_g51), .A(n4661), .ZN(n4673) );
  AOI22_X1 U5166 ( .A1(n4665), .A2(keyinput_g7), .B1(n4664), .B2(keyinput_g37), 
        .ZN(n4663) );
  OAI221_X1 U5167 ( .B1(n4665), .B2(keyinput_g7), .C1(n4664), .C2(keyinput_g37), .A(n4663), .ZN(n4672) );
  XOR2_X1 U5168 ( .A(n4666), .B(keyinput_g11), .Z(n4670) );
  XNOR2_X1 U5169 ( .A(DATAI_0_), .B(keyinput_g31), .ZN(n4669) );
  XNOR2_X1 U5170 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_g55), .ZN(n4668) );
  XNOR2_X1 U5171 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_g63), .ZN(n4667) );
  NAND4_X1 U5172 ( .A1(n4670), .A2(n4669), .A3(n4668), .A4(n4667), .ZN(n4671)
         );
  NOR3_X1 U5173 ( .A1(n4673), .A2(n4672), .A3(n4671), .ZN(n4718) );
  OAI22_X1 U5174 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_g59), .B1(
        REG3_REG_5__SCAN_IN), .B2(keyinput_g47), .ZN(n4674) );
  AOI221_X1 U5175 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_g59), .C1(
        keyinput_g47), .C2(REG3_REG_5__SCAN_IN), .A(n4674), .ZN(n4680) );
  OAI22_X1 U5176 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_g34), .B1(
        keyinput_g20), .B2(DATAI_11_), .ZN(n4675) );
  AOI221_X1 U5177 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_g34), .C1(
        DATAI_11_), .C2(keyinput_g20), .A(n4675), .ZN(n4678) );
  OAI22_X1 U5178 ( .A1(IR_REG_7__SCAN_IN), .A2(keyinput_g62), .B1(DATAI_9_), 
        .B2(keyinput_g22), .ZN(n4676) );
  AOI221_X1 U5179 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_g62), .C1(
        keyinput_g22), .C2(DATAI_9_), .A(n4676), .ZN(n4677) );
  NAND4_X1 U5180 ( .A1(n4680), .A2(n4679), .A3(n4678), .A4(n4677), .ZN(n4716)
         );
  OAI22_X1 U5181 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput_g38), .B1(DATAI_10_), 
        .B2(keyinput_g21), .ZN(n4681) );
  AOI221_X1 U5182 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput_g38), .C1(
        keyinput_g21), .C2(DATAI_10_), .A(n4681), .ZN(n4688) );
  OAI22_X1 U5183 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(DATAI_18_), .B2(
        keyinput_g13), .ZN(n4682) );
  AOI221_X1 U5184 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(keyinput_g13), .C2(
        DATAI_18_), .A(n4682), .ZN(n4687) );
  OAI22_X1 U5185 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(keyinput_g25), .B2(DATAI_6_), .ZN(n4683) );
  AOI221_X1 U5186 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(DATAI_6_), 
        .C2(keyinput_g25), .A(n4683), .ZN(n4686) );
  OAI22_X1 U5187 ( .A1(DATAI_14_), .A2(keyinput_g17), .B1(keyinput_g24), .B2(
        DATAI_7_), .ZN(n4684) );
  AOI221_X1 U5188 ( .B1(DATAI_14_), .B2(keyinput_g17), .C1(DATAI_7_), .C2(
        keyinput_g24), .A(n4684), .ZN(n4685) );
  NAND4_X1 U5189 ( .A1(n4688), .A2(n4687), .A3(n4686), .A4(n4685), .ZN(n4715)
         );
  OAI22_X1 U5190 ( .A1(n4691), .A2(keyinput_g41), .B1(n4690), .B2(keyinput_g33), .ZN(n4689) );
  AOI221_X1 U5191 ( .B1(n4691), .B2(keyinput_g41), .C1(keyinput_g33), .C2(
        n4690), .A(n4689), .ZN(n4701) );
  XNOR2_X1 U5192 ( .A(DATAI_3_), .B(keyinput_g28), .ZN(n4695) );
  XNOR2_X1 U5193 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_g52), .ZN(n4694) );
  XNOR2_X1 U5194 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_g36), .ZN(n4693) );
  XNOR2_X1 U5195 ( .A(keyinput_g48), .B(REG3_REG_17__SCAN_IN), .ZN(n4692) );
  NAND4_X1 U5196 ( .A1(n4695), .A2(n4694), .A3(n4693), .A4(n4692), .ZN(n4699)
         );
  XNOR2_X1 U5197 ( .A(n4696), .B(keyinput_g58), .ZN(n4698) );
  XNOR2_X1 U5198 ( .A(keyinput_g19), .B(n2449), .ZN(n4697) );
  NOR3_X1 U5199 ( .A1(n4699), .A2(n4698), .A3(n4697), .ZN(n4700) );
  NAND2_X1 U5200 ( .A1(n4701), .A2(n4700), .ZN(n4714) );
  OAI22_X1 U5201 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_g43), .B1(DATAI_13_), .B2(keyinput_g18), .ZN(n4702) );
  AOI221_X1 U5202 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_g43), .C1(
        keyinput_g18), .C2(DATAI_13_), .A(n4702), .ZN(n4712) );
  OAI22_X1 U5203 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_g39), .B1(DATAI_16_), .B2(keyinput_g15), .ZN(n4703) );
  AOI221_X1 U5204 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_g39), .C1(
        keyinput_g15), .C2(DATAI_16_), .A(n4703), .ZN(n4711) );
  OAI22_X1 U5205 ( .A1(n4706), .A2(keyinput_g14), .B1(n4705), .B2(keyinput_g26), .ZN(n4704) );
  AOI221_X1 U5206 ( .B1(n4706), .B2(keyinput_g14), .C1(keyinput_g26), .C2(
        n4705), .A(n4704), .ZN(n4710) );
  OAI22_X1 U5207 ( .A1(n4708), .A2(keyinput_g35), .B1(keyinput_g60), .B2(
        IR_REG_5__SCAN_IN), .ZN(n4707) );
  AOI221_X1 U5208 ( .B1(n4708), .B2(keyinput_g35), .C1(IR_REG_5__SCAN_IN), 
        .C2(keyinput_g60), .A(n4707), .ZN(n4709) );
  NAND4_X1 U5209 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .ZN(n4713)
         );
  NOR4_X1 U5210 ( .A1(n4716), .A2(n4715), .A3(n4714), .A4(n4713), .ZN(n4717)
         );
  NAND3_X1 U5211 ( .A1(n4719), .A2(n4718), .A3(n4717), .ZN(n4720) );
  NOR4_X1 U5212 ( .A1(n4723), .A2(n4722), .A3(n4721), .A4(n4720), .ZN(n4724)
         );
  AOI211_X1 U5213 ( .C1(REG3_REG_20__SCAN_IN), .C2(n4726), .A(n4725), .B(n4724), .ZN(n4729) );
  AOI22_X1 U5214 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n4728) );
  XNOR2_X1 U5215 ( .A(n4729), .B(n4728), .ZN(U3352) );
endmodule

